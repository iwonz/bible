DAN|1|1|In the third year of the reign of Jehoiakim king of Judah, Nebuchadnezzar king of Babylon came to Jerusalem and besieged it.
DAN|1|2|And the Lord gave Jehoiakim king of Judah into his hand, with some of the vessels of the house of God. And he brought them to the land of Shinar, to the house of his god, and placed the vessels in the treasury of his god.
DAN|1|3|Then the king commanded Ashpenaz, his chief eunuch, to bring some of the people of Israel, both of the royal family and of the nobility,
DAN|1|4|youths without blemish, of good appearance and skillful in all wisdom, endowed with knowledge, understanding learning, and competent to stand in the king's palace, and to teach them the literature and language of the Chaldeans.
DAN|1|5|The king assigned them a daily portion of the food that the king ate, and of the wine that he drank. They were to be educated for three years, and at the end of that time they were to stand before the king.
DAN|1|6|Among these were Daniel, Hananiah, Mishael, and Azariah of the tribe of Judah.
DAN|1|7|And the chief of the eunuchs gave them names: Daniel he called Belteshazzar, Hananiah he called Shadrach, Mishael he called Meshach, and Azariah he called Abednego.
DAN|1|8|But Daniel resolved that he would not defile himself with the king's food, or with the wine that he drank. Therefore he asked the chief of the eunuchs to allow him not to defile himself.
DAN|1|9|And God gave Daniel favor and compassion in the sight of the chief of the eunuchs,
DAN|1|10|and the chief of the eunuchs said to Daniel, "I fear my lord the king, who assigned your food and your drink; for why should he see that you were in worse condition than the youths who are of your own age? So you would endanger my head with the king."
DAN|1|11|Then Daniel said to the steward whom the chief of the eunuchs had assigned over Daniel, Hananiah, Mishael, and Azariah,
DAN|1|12|"Test your servants for ten days; let us be given vegetables to eat and water to drink.
DAN|1|13|Then let our appearance and the appearance of the youths who eat the king's food be observed by you, and deal with your servants according to what you see."
DAN|1|14|So he listened to them in this matter, and tested them for ten days.
DAN|1|15|At the end of ten days it was seen that they were better in appearance and fatter in flesh than all the youths who ate the king's food.
DAN|1|16|So the steward took away their food and the wine they were to drink, and gave them vegetables.
DAN|1|17|As for these four youths, God gave them learning and skill in all literature and wisdom, and Daniel had understanding in all visions and dreams.
DAN|1|18|At the end of the time, when the king had commanded that they should be brought in, the chief of the eunuchs brought them in before Nebuchadnezzar.
DAN|1|19|And the king spoke with them, and among all of them none was found like Daniel, Hananiah, Mishael, and Azariah. Therefore they stood before the king.
DAN|1|20|And in every matter of wisdom and understanding about which the king inquired of them, he found them ten times better than all the magicians and enchanters that were in all his kingdom.
DAN|1|21|And Daniel was there until the first year of King Cyrus.
DAN|2|1|In the second year of the reign of Nebuchadnezzar, Nebuchadnezzar had dreams; his spirit was troubled, and his sleep left him.
DAN|2|2|Then the king commanded that the magicians, the enchanters, the sorcerers, and the Chaldeans be summoned to tell the king his dreams. So they came in and stood before the king.
DAN|2|3|And the king said to them, "I had a dream, and my spirit is troubled to know the dream."
DAN|2|4|Then the Chaldeans said to the king in Aramaic, "O king, live forever! Tell your servants the dream, and we will show the interpretation."
DAN|2|5|The king answered and said to the Chaldeans, "The word from me is firm: if you do not make known to me the dream and its interpretation, you shall be torn limb from limb, and your houses shall be laid in ruins.
DAN|2|6|But if you show the dream and its interpretation, you shall receive from me gifts and rewards and great honor. Therefore show me the dream and its interpretation."
DAN|2|7|They answered a second time and said, "Let the king tell his servants the dream, and we will show its interpretation."
DAN|2|8|The king answered and said, "I know with certainty that you are trying to gain time, because you see that the word from me is firm-
DAN|2|9|if you do not make the dream known to me, there is but one sentence for you. You have agreed to speak lying and corrupt words before me till the times change. Therefore tell me the dream, and I shall know that you can show me its interpretation."
DAN|2|10|The Chaldeans answered the king and said, "There is not a man on earth who can meet the king's demand, for no great and powerful king has asked such a thing of any magician or enchanter or Chaldean.
DAN|2|11|The thing that the king asks is difficult, and no one can show it to the king except the gods, whose dwelling is not with flesh."
DAN|2|12|Because of this the king was angry and very furious, and commanded that all the wise men of Babylon be destroyed.
DAN|2|13|So the decree went out, and the wise men were about to be killed; and they sought Daniel and his companions, to kill them.
DAN|2|14|Then Daniel replied with prudence and discretion to Arioch, the captain of the king's guard, who had gone out to kill the wise men of Babylon.
DAN|2|15|He declared to Arioch, the king's captain, "Why is the decree of the king so urgent?" Then Arioch made the matter known to Daniel.
DAN|2|16|And Daniel went in and requested the king to appoint him a time, that he might show the interpretation to the king.
DAN|2|17|Then Daniel went to his house and made the matter known to Hananiah, Mishael, and Azariah, his companions,
DAN|2|18|and told them to seek mercy from the God of heaven concerning this mystery, so that Daniel and his companions might not be destroyed with the rest of the wise men of Babylon.
DAN|2|19|Then the mystery was revealed to Daniel in a vision of the night. Then Daniel blessed the God of heaven.
DAN|2|20|Daniel answered and said: "Blessed be the name of God forever and ever, to whom belong wisdom and might.
DAN|2|21|He changes times and seasons; he removes kings and sets up kings; he gives wisdom to the wise and knowledge to those who have understanding;
DAN|2|22|he reveals deep and hidden things; he knows what is in the darkness, and the light dwells with him.
DAN|2|23|To you, O God of my fathers, I give thanks and praise, for you have given me wisdom and might, and have now made known to me what we asked of you, for you have made known to us the king's matter."
DAN|2|24|Therefore Daniel went in to Arioch, whom the king had appointed to destroy the wise men of Babylon. He went and said thus to him, "Do not destroy the wise men of Babylon; bring me in before the king, and I will show the king the interpretation."
DAN|2|25|Then Arioch brought in Daniel before the king in haste and said thus to him: "I have found among the exiles from Judah a man who will make known to the king the interpretation."
DAN|2|26|The king said to Daniel, whose name was Belteshazzar, "Are you able to make known to me the dream that I have seen and its interpretation?"
DAN|2|27|Daniel answered the king and said, "No wise men, enchanters, magicians, or astrologers can show to the king the mystery that the king has asked,
DAN|2|28|but there is a God in heaven who reveals mysteries, and he has made known to King Nebuchadnezzar what will be in the latter days. Your dream and the visions of your head as you lay in bed are these:
DAN|2|29|To you, O king, as you lay in bed came thoughts of what would be after this, and he who reveals mysteries made known to you what is to be.
DAN|2|30|But as for me, this mystery has been revealed to me, not because of any wisdom that I have more than all the living, but in order that the interpretation may be made known to the king, and that you may know the thoughts of your mind.
DAN|2|31|"You saw, O king, and behold, a great image. This image, mighty and of exceeding brightness, stood before you, and its appearance was frightening.
DAN|2|32|The head of this image was of fine gold, its chest and arms of silver, its middle and thighs of bronze,
DAN|2|33|its legs of iron, its feet partly of iron and partly of clay.
DAN|2|34|As you looked, a stone was cut out by no human hand, and it struck the image on its feet of iron and clay, and broke them in pieces.
DAN|2|35|Then the iron, the clay, the bronze, the silver, and the gold, all together were broken in pieces, and became like the chaff of the summer threshing floors; and the wind carried them away, so that not a trace of them could be found. But the stone that struck the image became a great mountain and filled the whole earth.
DAN|2|36|"This was the dream. Now we will tell the king its interpretation.
DAN|2|37|You, O king, the king of kings, to whom the God of heaven has given the kingdom, the power, and the might, and the glory,
DAN|2|38|and into whose hand he has given, wherever they dwell, the children of man, the beasts of the field, and the birds of the heavens, making you rule over them all- you are the head of gold.
DAN|2|39|Another kingdom inferior to you shall arise after you, and yet a third kingdom of bronze, which shall rule over all the earth.
DAN|2|40|And there shall be a fourth kingdom, strong as iron, because iron breaks to pieces and shatters all things. And like iron that crushes, it shall break and crush all these.
DAN|2|41|And as you saw the feet and toes, partly of potter's clay and partly of iron, it shall be a divided kingdom, but some of the firmness of iron shall be in it, just as you saw iron mixed with the soft clay.
DAN|2|42|And as the toes of the feet were partly iron and partly clay, so the kingdom shall be partly strong and partly brittle.
DAN|2|43|As you saw the iron mixed with soft clay, so they will mix with one another in marriage, but they will not hold together, just as iron does not mix with clay.
DAN|2|44|And in the days of those kings the God of heaven will set up a kingdom that shall never be destroyed, nor shall the kingdom be left to another people. It shall break in pieces all these kingdoms and bring them to an end, and it shall stand forever,
DAN|2|45|just as you saw that a stone was cut from a mountain by no human hand, and that it broke in pieces the iron, the bronze, the clay, the silver, and the gold. A great God has made known to the king what shall be after this. The dream is certain, and its interpretation sure."
DAN|2|46|Then King Nebuchadnezzar fell upon his face and paid homage to Daniel, and commanded that an offering and incense be offered up to him.
DAN|2|47|The king answered and said to Daniel, "Truly, your God is God of gods and Lord of kings, and a revealer of mysteries, for you have been able to reveal this mystery."
DAN|2|48|Then the king gave Daniel high honors and many great gifts, and made him ruler over the whole province of Babylon and chief prefect over all the wise men of Babylon.
DAN|2|49|Daniel made a request of the king, and he appointed Shadrach, Meshach, and Abednego over the affairs of the province of Babylon. But Daniel remained at the king's court.
DAN|3|1|King Nebuchadnezzar made an image of gold, whose height was sixty cubits and its breadth six cubits. He set it up on the plain of Dura, in the province of Babylon.
DAN|3|2|Then King Nebuchadnezzar sent to gather the satraps, the prefects, and the governors, the counselors, the treasurers, the justices, the magistrates, and all the officials of the provinces to come to the dedication of the image that King Nebuchadnezzar had set up.
DAN|3|3|Then the satraps, the prefects, and the governors, the counselors, the treasurers, the justices, the magistrates, and all the officials of the provinces gathered for the dedication of the image that King Nebuchadnezzar had set up. And they stood before the image that Nebuchadnezzar had set up.
DAN|3|4|And the herald proclaimed aloud, "You are commanded, O peoples, nations, and languages,
DAN|3|5|that when you hear the sound of the horn, pipe, lyre, trigon, harp, bagpipe, and every kind of music, you are to fall down and worship the golden image that King Nebuchadnezzar has set up.
DAN|3|6|And whoever does not fall down and worship shall immediately be cast into a burning fiery furnace."
DAN|3|7|Therefore, as soon as all the peoples heard the sound of the horn, pipe, lyre, trigon, harp, bagpipe, and every kind of music, all the peoples, nations, and languages fell down and worshiped the golden image that King Nebuchadnezzar had set up.
DAN|3|8|Therefore at that time certain Chaldeans came forward and maliciously accused the Jews.
DAN|3|9|They declared to King Nebuchadnezzar, "O king, live forever!
DAN|3|10|You, O king, have made a decree, that every man who hears the sound of the horn, pipe, lyre, trigon, harp, bagpipe, and every kind of music, shall fall down and worship the golden image.
DAN|3|11|And whoever does not fall down and worship shall be cast into a burning fiery furnace.
DAN|3|12|There are certain Jews whom you have appointed over the affairs of the province of Babylon: Shadrach, Meshach, and Abednego. These men, O king, pay no attention to you; they do not serve your gods or worship the golden image that you have set up."
DAN|3|13|Then Nebuchadnezzar in furious rage commanded that Shadrach, Meshach, and Abednego be brought. So they brought these men before the king.
DAN|3|14|Nebuchadnezzar answered and said to them, "Is it true, O Shadrach, Meshach, and Abednego, that you do not serve my gods or worship the golden image that I have set up?
DAN|3|15|Now if you are ready when you hear the sound of the horn, pipe, lyre, trigon, harp, bagpipe, and every kind of music, to fall down and worship the image that I have made, well and good. But if you do not worship, you shall immediately be cast into a burning fiery furnace. And who is the god who will deliver you out of my hands?"
DAN|3|16|Shadrach, Meshach, and Abednego answered and said to the king, "O Nebuchadnezzar, we have no need to answer you in this matter.
DAN|3|17|If this be so, our God whom we serve is able to deliver us from the burning fiery furnace, and he will deliver us out of your hand, O king.
DAN|3|18|But if not, be it known to you, O king, that we will not serve your gods or worship the golden image that you have set up."
DAN|3|19|Then Nebuchadnezzar was filled with fury, and the expression of his face was changed against Shadrach, Meshach, and Abednego. He ordered the furnace heated seven times more than it was usually heated.
DAN|3|20|And he ordered some of the mighty men of his army to bind Shadrach, Meshach, and Abednego, and to cast them into the burning fiery furnace.
DAN|3|21|Then these men were bound in their cloaks, their tunics, their hats, and their other garments, and they were thrown into the burning fiery furnace.
DAN|3|22|Because the king's order was urgent and the furnace overheated, the flame of the fire killed those men who took up Shadrach, Meshach, and Abednego.
DAN|3|23|And these three men, Shadrach, Meshach, and Abednego, fell bound into the burning fiery furnace.
DAN|3|24|Then King Nebuchadnezzar was astonished and rose up in haste. He declared to his counselors, "Did we not cast three men bound into the fire?" They answered and said to the king, "True, O king."
DAN|3|25|He answered and said, "But I see four men unbound, walking in the midst of the fire, and they are not hurt; and the appearance of the fourth is like a son of the gods."
DAN|3|26|Then Nebuchadnezzar came near to the door of the burning fiery furnace; he declared, "Shadrach, Meshach, and Abednego, servants of the Most High God, come out, and come here!" Then Shadrach, Meshach, and Abednego came out from the fire.
DAN|3|27|And the satraps, the prefects, the governors, and the king's counselors gathered together and saw that the fire had not had any power over the bodies of those men. The hair of their heads was not singed, their cloaks were not harmed, and no smell of fire had come upon them.
DAN|3|28|Nebuchadnezzar answered and said, "Blessed be the God of Shadrach, Meshach, and Abednego, who has sent his angel and delivered his servants, who trusted in him, and set aside the king's command, and yielded up their bodies rather than serve and worship any god except their own God.
DAN|3|29|Therefore I make a decree: Any people, nation, or language that speaks anything against the God of Shadrach, Meshach, and Abednego shall be torn limb from limb, and their houses laid in ruins, for there is no other god who is able to rescue in this way."
DAN|3|30|Then the king promoted Shadrach, Meshach, and Abednego in the province of Babylon.
DAN|4|1|King Nebuchadnezzar to all peo- ples, nations, and languages, that dwell in all the earth: Peace be multiplied to you!
DAN|4|2|It has seemed good to me to show the signs and wonders that the Most High God has done for me.
DAN|4|3|How great are his signs, how mighty his wonders! His kingdom is an everlasting kingdom, and his dominion endures from generation to generation.
DAN|4|4|I, Nebuchadnezzar, was at ease in my house and prospering in my palace.
DAN|4|5|I saw a dream that made me afraid. As I lay in bed the fancies and the visions of my head alarmed me.
DAN|4|6|So I made a decree that all the wise men of Babylon should be brought before me, that they might make known to me the interpretation of the dream.
DAN|4|7|Then the magicians, the enchanters, the Chaldeans, and the astrologers came in, and I told them the dream, but they could not make known to me its interpretation.
DAN|4|8|At last Daniel came in before me- he who was named Belteshazzar after the name of my god, and in whom is the spirit of the holy gods- and I told him the dream, saying,
DAN|4|9|"O Belteshazzar, chief of the magicians, because I know that the spirit of the holy gods is in you and that no mystery is too difficult for you, tell me the visions of my dream that I saw and their interpretation.
DAN|4|10|The visions of my head as I lay in bed were these: I saw, and behold, a tree in the midst of the earth, and its height was great.
DAN|4|11|The tree grew and became strong, and its top reached to heaven, and it was visible to the end of the whole earth.
DAN|4|12|Its leaves were beautiful and its fruit abundant, and in it was food for all. The beasts of the field found shade under it, and the birds of the heavens lived in its branches, and all flesh was fed from it.
DAN|4|13|"I saw in the visions of my head as I lay in bed, and behold, a watcher, a holy one, came down from heaven.
DAN|4|14|He proclaimed aloud and said thus: 'Chop down the tree and lop off its branches, strip off its leaves and scatter its fruit. Let the beasts flee from under it and the birds from its branches.
DAN|4|15|But leave the stump of its roots in the earth, bound with a band of iron and bronze, amid the tender grass of the field. Let him be wet with the dew of heaven. Let his portion be with the beasts in the grass of the earth.
DAN|4|16|Let his mind be changed from a man's, and let a beast's mind be given to him; and let seven periods of time pass over him.
DAN|4|17|The sentence is by the decree of the watchers, the decision by the word of the holy ones, to the end that the living may know that the Most High rules the kingdom of men and gives it to whom he will and sets over it the lowliest of men.'
DAN|4|18|This dream I, King Nebuchadnezzar, saw. And you, O Belteshazzar, tell me the interpretation, because all the wise men of my kingdom are not able to make known to me the interpretation, but you are able, for the spirit of the holy gods is in you."
DAN|4|19|Then Daniel, whose name was Belteshazzar, was dismayed for a while, and his thoughts alarmed him. The king answered and said, "Belteshazzar, let not the dream or the interpretation alarm you." Belteshazzar answered and said, "My lord, may the dream be for those who hate you and its interpretation for your enemies!
DAN|4|20|The tree you saw, which grew and became strong, so that its top reached to heaven, and it was visible to the end of the whole earth,
DAN|4|21|whose leaves were beautiful and its fruit abundant, and in which was food for all, under which beasts of the field found shade, and in whose branches the birds of the heavens lived-
DAN|4|22|it is you, O king, who have grown and become strong. Your greatness has grown and reaches to heaven, and your dominion to the ends of the earth.
DAN|4|23|And because the king saw a watcher, a holy one, coming down from heaven and saying, 'Chop down the tree and destroy it, but leave the stump of its roots in the earth, bound with a band of iron and bronze, in the tender grass of the field, and let him be wet with the dew of heaven, and let his portion be with the beasts of the field, till seven periods of time pass over him,'
DAN|4|24|this is the interpretation, O king: It is a decree of the Most High, which has come upon my lord the king,
DAN|4|25|that you shall be driven from among men, and your dwelling shall be with the beasts of the field. You shall be made to eat grass like an ox, and you shall be wet with the dew of heaven, and seven periods of time shall pass over you, till you know that the Most High rules the kingdom of men and gives it to whom he will.
DAN|4|26|And as it was commanded to leave the stump of the roots of the tree, your kingdom shall be confirmed for you from the time that you know that Heaven rules.
DAN|4|27|Therefore, O king, let my counsel be acceptable to you: break off your sins by practicing righteousness, and your iniquities by showing mercy to the oppressed, that there may perhaps be a lengthening of your prosperity."
DAN|4|28|All this came upon King Nebuchadnezzar.
DAN|4|29|At the end of twelve months he was walking on the roof of the royal palace of Babylon,
DAN|4|30|and the king answered and said, "Is not this great Babylon, which I have built by my mighty power as a royal residence and for the glory of my majesty?"
DAN|4|31|While the words were still in the king's mouth, there fell a voice from heaven, "O King Nebuchadnezzar, to you it is spoken: The kingdom has departed from you,
DAN|4|32|and you shall be driven from among men, and your dwelling shall be with the beasts of the field. And you shall be made to eat grass like an ox, and seven periods of time shall pass over you, until you know that the Most High rules the kingdom of men and gives it to whom he will."
DAN|4|33|Immediately the word was fulfilled against Nebuchadnezzar. He was driven from among men and ate grass like an ox, and his body was wet with the dew of heaven till his hair grew as long as eagles' feathers, and his nails were like birds' claws.
DAN|4|34|At the end of the days I, Nebuchadnezzar, lifted my eyes to heaven, and my reason returned to me, and I blessed the Most High, and praised and honored him who lives forever, for his dominion is an everlasting dominion, and his kingdom endures from generation to generation;
DAN|4|35|all the inhabitants of the earth are accounted as nothing, and he does according to his will among the host of heaven and among the inhabitants of the earth; and none can stay his hand or say to him, "What have you done?"
DAN|4|36|At the same time my reason returned to me, and for the glory of my kingdom, my majesty and splendor returned to me. My counselors and my lords sought me, and I was established in my kingdom, and still more greatness was added to me.
DAN|4|37|Now I, Nebuchadnezzar, praise and extol and honor the King of heaven, for all his works are right and his ways are just; and those who walk in pride he is able to humble.
DAN|5|1|King Belshazzar made a great feast for a thousand of his lords and drank wine in front of the thousand.
DAN|5|2|Belshazzar, when he tasted the wine, commanded that the vessels of gold and of silver that Nebuchadnezzar his father had taken out of the temple in Jerusalem be brought, that the king and his lords, his wives, and his concubines might drink from them.
DAN|5|3|Then they brought in the golden vessels that had been taken out of the temple, the house of God in Jerusalem, and the king and his lords, his wives, and his concubines drank from them.
DAN|5|4|They drank wine and praised the gods of gold and silver, bronze, iron, wood, and stone.
DAN|5|5|Immediately the fingers of a human hand appeared and wrote on the plaster of the wall of the king's palace, opposite the lampstand. And the king saw the hand as it wrote.
DAN|5|6|Then the king's color changed, and his thoughts alarmed him; his limbs gave way, and his knees knocked together.
DAN|5|7|The king called loudly to bring in the enchanters, the Chaldeans, and the astrologers. The king declared to the wise men of Babylon, "Whoever reads this writing, and shows me its interpretation, shall be clothed with purple and have a chain of gold around his neck and shall be the third ruler in the kingdom."
DAN|5|8|Then all the king's wise men came in, but they could not read the writing or make known to the king the interpretation.
DAN|5|9|Then King Belshazzar was greatly alarmed, and his color changed, and his lords were perplexed.
DAN|5|10|The queen, because of the words of the king and his lords, came into the banqueting hall, and the queen declared, "O king, live forever! Let not your thoughts alarm you or your color change.
DAN|5|11|There is a man in your kingdom in whom is the spirit of the holy gods. In the days of your father, light and understanding and wisdom like the wisdom of the gods were found in him, and King Nebuchadnezzar, your father- your father the king- made him chief of the magicians, enchanters, Chaldeans, and astrologers,
DAN|5|12|because an excellent spirit, knowledge, and understanding to interpret dreams, explain riddles, and solve problems were found in this Daniel, whom the king named Belteshazzar. Now let Daniel be called, and he will show the interpretation."
DAN|5|13|Then Daniel was brought in before the king. The king answered and said to Daniel, "You are that Daniel, one of the exiles of Judah, whom the king my father brought from Judah.
DAN|5|14|I have heard of you that the spirit of the gods is in you, and that light and understanding and excellent wisdom are found in you.
DAN|5|15|Now the wise men, the enchanters, have been brought in before me to read this writing and make known to me its interpretation, but they could not show the interpretation of the matter.
DAN|5|16|But I have heard that you can give interpretations and solve problems. Now if you can read the writing and make known to me its interpretation, you shall be clothed with purple and have a chain of gold around your neck and shall be the third ruler in the kingdom."
DAN|5|17|Then Daniel answered and said before the king, "Let your gifts be for yourself, and give your rewards to another. Nevertheless, I will read the writing to the king and make known to him the interpretation.
DAN|5|18|O king, the Most High God gave Nebuchadnezzar your father kingship and greatness and glory and majesty.
DAN|5|19|And because of the greatness that he gave him, all peoples, nations, and languages trembled and feared before him. Whom he would, he killed, and whom he would, he kept alive; whom he would, he raised up, and whom he would, he humbled.
DAN|5|20|But when his heart was lifted up and his spirit was hardened so that he dealt proudly, he was brought down from his kingly throne, and his glory was taken from him.
DAN|5|21|He was driven from among the children of mankind, and his mind was made like that of a beast, and his dwelling was with the wild donkeys. He was fed grass like an ox, and his body was wet with the dew of heaven, until he knew that the Most High God rules the kingdom of mankind and sets over it whom he will.
DAN|5|22|And you his son, Belshazzar, have not humbled your heart, though you knew all this,
DAN|5|23|but you have lifted up yourself against the Lord of heaven. And the vessels of his house have been brought in before you, and you and your lords, your wives, and your concubines have drunk wine from them. And you have praised the gods of silver and gold, of bronze, iron, wood, and stone, which do not see or hear or know, but the God in whose hand is your breath, and whose are all your ways, you have not honored.
DAN|5|24|"Then from his presence the hand was sent, and this writing was inscribed.
DAN|5|25|And this is the writing that was inscribed: MENE, MENE, TEKEL, and PARSIN.
DAN|5|26|This is the interpretation of the matter: MENE, God has numbered the days of your kingdom and brought it to an end;
DAN|5|27|TEKEL, you have been weighed in the balances and found wanting;
DAN|5|28|PERES, your kingdom is divided and given to the Medes and Persians."
DAN|5|29|Then Belshazzar gave the command, and Daniel was clothed with purple, a chain of gold was put around his neck, and a proclamation was made about him, that he should be the third ruler in the kingdom.
DAN|5|30|That very night Belshazzar the Chaldean king was killed.
DAN|5|31|And Darius the Mede received the kingdom, being about sixty-two years old.
DAN|6|1|It pleased Darius to set over the kingdom 120 satraps, to be throughout the whole kingdom;
DAN|6|2|and over them three presidents, of whom Daniel was one, to whom these satraps should give account, so that the king might suffer no loss.
DAN|6|3|Then this Daniel became distinguished above all the other presidents and satraps, because an excellent spirit was in him. And the king planned to set him over the whole kingdom.
DAN|6|4|Then the presidents and the satraps sought to find a ground for complaint against Daniel with regard to the kingdom, but they could find no ground for complaint or any fault, because he was faithful, and no error or fault was found in him.
DAN|6|5|Then these men said, "We shall not find any ground for complaint against this Daniel unless we find it in connection with the law of his God."
DAN|6|6|Then these presidents and satraps came by agreement to the king and said to him, "O King Darius, live forever!
DAN|6|7|All the presidents of the kingdom, the prefects and the satraps, the counselors and the governors are agreed that the king should establish an ordinance and enforce an injunction, that whoever makes petition to any god or man for thirty days, except to you, O king, shall be cast into the den of lions.
DAN|6|8|Now, O king, establish the injunction and sign the document, so that it cannot be changed, according to the law of the Medes and the Persians, which cannot be revoked."
DAN|6|9|Therefore King Darius signed the document and injunction.
DAN|6|10|When Daniel knew that the document had been signed, he went to his house where he had windows in his upper chamber open toward Jerusalem. He got down on his knees three times a day and prayed and gave thanks before his God, as he had done previously.
DAN|6|11|Then these men came by agreement and found Daniel making petition and plea before his God.
DAN|6|12|Then they came near and said before the king, concerning the injunction, "O king! Did you not sign an injunction, that anyone who makes petition to any god or man within thirty days except to you, O king, shall be cast into the den of lions?" The king answered and said, "The thing stands fast, according to the law of the Medes and Persians, which cannot be revoked."
DAN|6|13|Then they answered and said before the king, "Daniel, who is one of the exiles from Judah, pays no attention to you, O king, or the injunction you have signed, but makes his petition three times a day."
DAN|6|14|Then the king, when he heard these words, was much distressed and set his mind to deliver Daniel. And he labored till the sun went down to rescue him.
DAN|6|15|Then these men came by agreement to the king and said to the king, "Know, O king, that it is a law of the Medes and Persians that no injunction or ordinance that the king establishes can be changed."
DAN|6|16|Then the king commanded, and Daniel was brought and cast into the den of lions. The king declared to Daniel, "May your God, whom you serve continually, deliver you!"
DAN|6|17|And a stone was brought and laid on the mouth of the den, and the king sealed it with his own signet and with the signet of his lords, that nothing might be changed concerning Daniel.
DAN|6|18|Then the king went to his palace and spent the night fasting; no diversions were brought to him, and sleep fled from him.
DAN|6|19|Then, at break of day, the king arose and went in haste to the den of lions.
DAN|6|20|As he came near to the den where Daniel was, he cried out in a tone of anguish. The king declared to Daniel, "O Daniel, servant of the living God, has your God, whom you serve continually, been able to deliver you from the lions?"
DAN|6|21|Then Daniel said to the king, "O king, live forever!
DAN|6|22|My God sent his angel and shut the lions' mouths, and they have not harmed me, because I was found blameless before him; and also before you, O king, I have done no harm."
DAN|6|23|Then the king was exceedingly glad, and commanded that Daniel be taken up out of the den. So Daniel was taken up out of the den, and no kind of harm was found on him, because he had trusted in his God.
DAN|6|24|And the king commanded, and those men who had maliciously accused Daniel were brought and cast into the den of lions- they, their children, and their wives. And before they reached the bottom of the den, the lions overpowered them and broke all their bones in pieces.
DAN|6|25|Then King Darius wrote to all the peoples, nations, and languages that dwell in all the earth: "Peace be multiplied to you.
DAN|6|26|I make a decree, that in all my royal dominion people are to tremble and fear before the God of Daniel, for he is the living God, enduring forever; his kingdom shall never be destroyed, and his dominion shall be to the end.
DAN|6|27|He delivers and rescues; he works signs and wonders in heaven and on earth, he who has saved Daniel from the power of the lions."
DAN|6|28|So this Daniel prospered during the reign of Darius and the reign of Cyrus the Persian.
DAN|7|1|In the first year of Belshazzar king of Babylon, Daniel saw a dream and visions of his head as he lay in his bed. Then he wrote down the dream and told the sum of the matter.
DAN|7|2|Daniel declared, "I saw in my vision by night, and behold, the four winds of heaven were stirring up the great sea.
DAN|7|3|And four great beasts came up out of the sea, different from one another.
DAN|7|4|The first was like a lion and had eagles' wings. Then as I looked its wings were plucked off, and it was lifted up from the ground and made to stand on two feet like a man, and the mind of a man was given to it.
DAN|7|5|And behold, another beast, a second one, like a bear. It was raised up on one side. It had three ribs in its mouth between its teeth; and it was told, 'Arise, devour much flesh.'
DAN|7|6|After this I looked, and behold, another, like a leopard, with four wings of a bird on its back. And the beast had four heads, and dominion was given to it.
DAN|7|7|After this I saw in the night visions, and behold, a fourth beast, terrifying and dreadful and exceedingly strong. It had great iron teeth; it devoured and broke in pieces and stamped what was left with its feet. It was different from all the beasts that were before it, and it had ten horns.
DAN|7|8|I considered the horns, and behold, there came up among them another horn, a little one, before which three of the first horns were plucked up by the roots. And behold, in this horn were eyes like the eyes of a man, and a mouth speaking great things.
DAN|7|9|As I looked, thrones were placed, and the Ancient of days took his seat; his clothing was white as snow, and the hair of his head like pure wool; his throne was fiery flames; its wheels were burning fire.
DAN|7|10|A stream of fire issued and came out from before him; a thousand thousands served him, and ten thousand times ten thousand stood before him; the court sat in judgment, and the books were opened.
DAN|7|11|I looked then because of the sound of the great words that the horn was speaking. And as I looked, the beast was killed, and its body destroyed and given over to be burned with fire.
DAN|7|12|As for the rest of the beasts, their dominion was taken away, but their lives were prolonged for a season and a time.
DAN|7|13|I saw in the night visions, and behold, with the clouds of heaven there came one like a son of man, and he came to the Ancient of Days and was presented before him.
DAN|7|14|And to him was given dominion and glory and a kingdom, that all peoples, nations, and languages should serve him; his dominion is an everlasting dominion, which shall not pass away, and his kingdom one that shall not be destroyed.
DAN|7|15|"As for me, Daniel, my spirit within me was anxious, and the visions of my head alarmed me.
DAN|7|16|I approached one of those who stood there and asked him the truth concerning all this. So he told me and made known to me the interpretation of the things.
DAN|7|17|'These four great beasts are four kings who shall arise out of the earth.
DAN|7|18|But the saints of the Most High shall receive the kingdom and possess the kingdom forever, forever and ever.'
DAN|7|19|"Then I desired to know the truth about the fourth beast, which was different from all the rest, exceedingly terrifying, with its teeth of iron and claws of bronze, and which devoured and broke in pieces and stamped what was left with its feet,
DAN|7|20|and about the ten horns that were on its head, and the other horn that came up and before which three of them fell, the horn that had eyes and a mouth that spoke great things, and that seemed greater than its companions.
DAN|7|21|As I looked, this horn made war with the saints and prevailed over them,
DAN|7|22|until the Ancient of Days came, and judgment was given for the saints of the Most High, and the time came when the saints possessed the kingdom.
DAN|7|23|"Thus he said: 'As for the fourth beast, there shall be a fourth kingdom on earth, which shall be different from all the kingdoms, and it shall devour the whole earth, and trample it down, and break it to pieces.
DAN|7|24|As for the ten horns, out of this kingdom ten kings shall arise, and another shall arise after them; he shall be different from the former ones, and shall put down three kings.
DAN|7|25|He shall speak words against the Most High, and shall wear out the saints of the Most High, and shall think to change the times and the law; and they shall be given into his hand for a time, times, and half a time.
DAN|7|26|But the court shall sit in judgment, and his dominion shall be taken away, to be consumed and destroyed to the end.
DAN|7|27|And the kingdom and the dominion and the greatness of the kingdoms under the whole heaven shall be given to the people of the saints of the Most High; their kingdom shall be an everlasting kingdom, and all dominions shall serve and obey them.'
DAN|7|28|"Here is the end of the matter. As for me, Daniel, my thoughts greatly alarmed me, and my color changed, but I kept the matter in my heart."
DAN|8|1|In the third year of the reign of King Belshazzar a vision appeared to me, Daniel, after that which appeared to me at the first.
DAN|8|2|And I saw in the vision; and when I saw, I was in Susa the capital, which is in the province of Elam. And I saw in the vision, and I was at the Ulai canal.
DAN|8|3|I raised my eyes and saw, and behold, a ram standing on the bank of the canal. It had two horns, and both horns were high, but one was higher than the other, and the higher one came up last.
DAN|8|4|I saw the ram charging westward and northward and southward. No beast could stand before him, and there was no one who could rescue from his power. He did as he pleased and became great.
DAN|8|5|As I was considering, behold, a male goat came from the west across the face of the whole earth, without touching the ground. And the goat had a conspicuous horn between his eyes.
DAN|8|6|He came to the ram with the two horns, which I had seen standing on the bank of the canal, and he ran at him in his powerful wrath.
DAN|8|7|I saw him come close to the ram, and he was enraged against him and struck the ram and broke his two horns. And the ram had no power to stand before him, but he cast him down to the ground and trampled on him. And there was no one who could rescue the ram from his power.
DAN|8|8|Then the goat became exceedingly great, but when he was strong, the great horn was broken, and instead of it there came up four conspicuous horns toward the four winds of heaven.
DAN|8|9|Out of one of them came a little horn, which grew exceedingly great toward the south, toward the east, and toward the glorious land.
DAN|8|10|It grew great, even to the host of heaven. And some of the host and some of the stars it threw down to the ground and trampled on them.
DAN|8|11|It became great, even as great as the Prince of the host. And the regular burnt offering was taken away from him, and the place of his sanctuary was overthrown.
DAN|8|12|And a host will be given over to it together with the regular burnt offering because of transgression, and it will throw truth to the ground, and it will act and prosper.
DAN|8|13|Then I heard a holy one speaking, and another holy one said to the one who spoke, "For how long is the vision concerning the regular burnt offering, the transgression that makes desolate, and the giving over of the sanctuary and host to be trampled underfoot?"
DAN|8|14|And he said to me, "For 2,300 evenings and mornings. Then the sanctuary shall be restored to its rightful state."
DAN|8|15|When I, Daniel, had seen the vision, I sought to understand it. And behold, there stood before me one having the appearance of a man.
DAN|8|16|And I heard a man's voice between the banks of the Ulai, and it called, "Gabriel, make this man understand the vision."
DAN|8|17|So he came near where I stood. And when he came, I was frightened and fell on my face. But he said to me, "Understand, O son of man, that the vision is for the time of the end."
DAN|8|18|And when he had spoken to me, I fell into a deep sleep with my face to the ground. But he touched me and made me stand up.
DAN|8|19|He said, "Behold, I will make known to you what shall be at the latter end of the indignation, for it refers to the appointed time of the end.
DAN|8|20|As for the ram that you saw with the two horns, these are the kings of Media and Persia.
DAN|8|21|And the goat is the king of Greece. And the great horn between his eyes is the first king.
DAN|8|22|As for the horn that was broken, in place of which four others arose, four kingdoms shall arise from his nation, but not with his power.
DAN|8|23|And at the latter end of their kingdom, when the transgressors have reached their limit, a king of bold face, one who understands riddles, shall arise.
DAN|8|24|His power shall be great- but not by his own power; and he shall cause fearful destruction and shall succeed in what he does, and destroy mighty men and the people who are the saints.
DAN|8|25|By his cunning he shall make deceit prosper under his hand, and in his own mind he shall become great. Without warning he shall destroy many. And he shall even rise up against the Prince of princes, and he shall be broken- but by no human hand.
DAN|8|26|The vision of the evenings and the mornings that has been told is true, but seal up the vision, for it refers to many days from now."
DAN|8|27|And I, Daniel, was overcome and lay sick for some days. Then I rose and went about the king's business, but I was appalled by the vision and did not understand it.
DAN|9|1|In the first year of Darius the son of Ahasuerus, by descent a Mede, who was made king over the realm of the Chaldeans-
DAN|9|2|in the first year of his reign, I, Daniel, perceived in the books the number of years that, according to the word of the LORD to Jeremiah the prophet, must pass before the end of the desolations of Jerusalem, namely, seventy years.
DAN|9|3|Then I turned my face to the Lord God, seeking him by prayer and pleas for mercy with fasting and sackcloth and ashes.
DAN|9|4|I prayed to the LORD my God and made confession, saying, "O Lord, the great and awesome God, who keeps covenant and steadfast love with those who love him and keep his commandments,
DAN|9|5|we have sinned and done wrong and acted wickedly and rebelled, turning aside from your commandments and rules.
DAN|9|6|We have not listened to your servants the prophets, who spoke in your name to our kings, our princes, and our fathers, and to all the people of the land.
DAN|9|7|To you, O Lord, belongs righteousness, but to us open shame, as at this day, to the men of Judah, to the inhabitants of Jerusalem, and to all Israel, those who are near and those who are far away, in all the lands to which you have driven them, because of the treachery that they have committed against you.
DAN|9|8|To us, O Lord, belongs open shame, to our kings, to our princes, and to our fathers, because we have sinned against you.
DAN|9|9|To the Lord our God belong mercy and forgiveness, for we have rebelled against him
DAN|9|10|and have not obeyed the voice of the LORD our God by walking in his laws, which he set before us by his servants the prophets.
DAN|9|11|All Israel has transgressed your law and turned aside, refusing to obey your voice. And the curse and oath that are written in the Law of Moses the servant of God have been poured out upon us, because we have sinned against him.
DAN|9|12|He has confirmed his words, which he spoke against us and against our rulers who ruled us, by bringing upon us a great calamity. For under the whole heaven there has not been done anything like what has been done against Jerusalem.
DAN|9|13|As it is written in the Law of Moses, all this calamity has come upon us; yet we have not entreated the favor of the LORD our God, turning from our iniquities and gaining insight by your truth.
DAN|9|14|Therefore the LORD has kept ready the calamity and has brought it upon us, for the LORD our God is righteous in all the works that he has done, and we have not obeyed his voice.
DAN|9|15|And now, O Lord our God, who brought your people out of the land of Egypt with a mighty hand, and have made a name for yourself, as at this day, we have sinned, we have done wickedly.
DAN|9|16|"O Lord, according to all your righteous acts, let your anger and your wrath turn away from your city Jerusalem, your holy hill, because for our sins, and for the iniquities of our fathers, Jerusalem and your people have become a byword among all who are around us.
DAN|9|17|Now therefore, O our God, listen to the prayer of your servant and to his pleas for mercy, and for your own sake, O Lord, make your face to shine upon your sanctuary, which is desolate.
DAN|9|18|O my God, incline your ear and hear. Open your eyes and see our desolations, and the city that is called by your name. For we do not present our pleas before you because of our righteousness, but because of your great mercy.
DAN|9|19|O Lord, hear; O Lord, forgive. O Lord, pay attention and act. Delay not, for your own sake, O my God, because your city and your people are called by your name."
DAN|9|20|While I was speaking and praying, confessing my sin and the sin of my people Israel, and presenting my plea before the LORD my God for the holy hill of my God,
DAN|9|21|while I was speaking in prayer, the man Gabriel, whom I had seen in the vision at the first, came to me in swift flight at the time of the evening sacrifice.
DAN|9|22|He made me understand, speaking with me and saying, "O Daniel, I have now come out to give you insight and understanding.
DAN|9|23|At the beginning of your pleas for mercy a word went out, and I have come to tell it to you, for you are greatly loved. Therefore consider the word and understand the vision.
DAN|9|24|"Seventy weeks are decreed about your people and your holy city, to finish the transgression, to put an end to sin, and to atone for iniquity, to bring in everlasting righteousness, to seal both vision and prophet, and to anoint a most holy place.
DAN|9|25|Know therefore and understand that from the going out of the word to restore and build Jerusalem to the coming of an anointed one, a prince, there shall be seven weeks. Then for sixty-two weeks it shall be built again with squares and moat, but in a troubled time.
DAN|9|26|And after the sixty-two weeks, an anointed one shall be cut off and shall have nothing. And the people of the prince who is to come shall destroy the city and the sanctuary. Its end shall come with a flood, and to the end there shall be war. Desolations are decreed.
DAN|9|27|And he shall make a strong covenant with many for one week, and for half of the week he shall put an end to sacrifice and offering. And on the wing of abominations shall come one who makes desolate, until the decreed end is poured out on the desolator."
DAN|10|1|In the third year of Cyrus king of Persia a word was revealed to Daniel, who was named Belteshazzar. And the word was true, and it was a great conflict. And he understood the word and had understanding of the vision.
DAN|10|2|In those days I, Daniel, was mourning for three weeks.
DAN|10|3|I ate no delicacies, no meat or wine entered my mouth, nor did I anoint myself at all, for the full three weeks.
DAN|10|4|On the twenty-fourth day of the first month, as I was standing on the bank of the great river (that is, the Tigris)
DAN|10|5|I lifted up my eyes and looked, and behold, a man clothed in linen, with a belt of fine gold from Uphaz around his waist.
DAN|10|6|His body was like beryl, his face like the appearance of lightning, his eyes like flaming torches, his arms and legs like the gleam of burnished bronze, and the sound of his words like the sound of a multitude.
DAN|10|7|And I, Daniel, alone saw the vision, for the men who were with me did not see the vision, but a great trembling fell upon them, and they fled to hide themselves.
DAN|10|8|So I was left alone and saw this great vision, and no strength was left in me. My radiant appearance was fearfully changed, and I retained no strength.
DAN|10|9|Then I heard the sound of his words, and as I heard the sound of his words, I fell on my face in deep sleep with my face to the ground.
DAN|10|10|And behold, a hand touched me and set me trembling on my hands and knees.
DAN|10|11|And he said to me, "O Daniel, man greatly loved, understand the words that I speak to you, and stand upright, for now I have been sent to you." And when he had spoken this word to me, I stood up trembling.
DAN|10|12|Then he said to me, "Fear not, Daniel, for from the first day that you set your heart to understand and humbled yourself before your God, your words have been heard, and I have come because of your words.
DAN|10|13|The prince of the kingdom of Persia withstood me twenty-one days, but Michael, one of the chief princes, came to help me, for I was left there with the kings of Persia,
DAN|10|14|and came to make you understand what is to happen to your people in the latter days. For the vision is for days yet to come."
DAN|10|15|When he had spoken to me according to these words, I turned my face toward the ground and was mute.
DAN|10|16|And behold, one in the likeness of the children of man touched my lips. Then I opened my mouth and spoke. I said to him who stood before me, "O my lord, by reason of the vision pains have come upon me, and I retain no strength.
DAN|10|17|How can my lord's servant talk with my lord? For now no strength remains in me, and no breath is left in me."
DAN|10|18|Again one having the appearance of a man touched me and strengthened me.
DAN|10|19|And he said, "O man greatly loved, fear not, peace be with you; be strong and of good courage." And as he spoke to me, I was strengthened and said, "Let my lord speak, for you have strengthened me."
DAN|10|20|Then he said, "Do you know why I have come to you? But now I will return to fight against the prince of Persia; and when I go out, behold, the prince of Greece will come.
DAN|10|21|But I will tell you what is inscribed in the book of truth: there is none who contends by my side against these except Michael, your prince.
DAN|11|1|And as for me, in the first year of Darius the Mede, I stood up to confirm and strengthen him.
DAN|11|2|"And now I will show you the truth. Behold, three more kings shall arise in Persia, and a fourth shall be far richer than all of them. And when he has become strong through his riches, he shall stir up all against the kingdom of Greece.
DAN|11|3|Then a mighty king shall arise, who shall rule with great dominion and do as he wills.
DAN|11|4|And as soon as he has arisen, his kingdom shall be broken and divided toward the four winds of heaven, but not to his posterity, nor according to the authority with which he ruled, for his kingdom shall be plucked up and go to others besides these.
DAN|11|5|"Then the king of the south shall be strong, but one of his princes shall be stronger than he and shall rule, and his authority shall be a great authority.
DAN|11|6|After some years they shall make an alliance, and the daughter of the king of the south shall come to the king of the north to make an agreement. But she shall not retain the strength of her arm, and he and his arm shall not endure, but she shall be given up, and her attendants, he who fathered her, and he who supported her in those times.
DAN|11|7|"And from a branch from her roots one shall arise in his place. He shall come against the army and enter the fortress of the king of the north, and he shall deal with them and shall prevail.
DAN|11|8|He shall also carry off to Egypt their gods with their metal images and their precious vessels of silver and gold, and for some years he shall refrain from attacking the king of the north.
DAN|11|9|Then the latter shall come into the realm of the king of the south but shall return to his own land.
DAN|11|10|"His sons shall wage war and assemble a multitude of great forces, which shall keep coming and overflow and pass through, and again shall carry the war as far as his fortress.
DAN|11|11|Then the king of the south, moved with rage, shall come out and fight with the king of the north. And he shall raise a great multitude, but it shall be given into his hand.
DAN|11|12|And when the multitude is taken away, his heart shall be exalted, and he shall cast down tens of thousands, but he shall not prevail.
DAN|11|13|For the king of the north shall again raise a multitude, greater than the first. And after some years he shall come on with a great army and abundant supplies.
DAN|11|14|"In those times many shall rise against the king of the south, and the violent among your own people shall lift themselves up in order to fulfill the vision, but they shall fail.
DAN|11|15|Then the king of the north shall come and throw up siegeworks and take a well-fortified city. And the forces of the south shall not stand, or even his best troops, for there shall be no strength to stand.
DAN|11|16|But he who comes against him shall do as he wills, and none shall stand before him. And he shall stand in the glorious land, with destruction in his hand.
DAN|11|17|He shall set his face to come with the strength of his whole kingdom, and he shall bring terms of an agreement and perform them. He shall give him the daughter of women to destroy the kingdom, but it shall not stand or be to his advantage.
DAN|11|18|Afterward he shall turn his face to the coastlands and shall capture many of them, but a commander shall put an end to his insolence. Indeed, he shall turn his insolence back upon him.
DAN|11|19|Then he shall turn his face back toward the fortresses of his own land, but he shall stumble and fall, and shall not be found.
DAN|11|20|"Then shall arise in his place one who shall send an exactor of tribute for the glory of the kingdom. But within a few days he shall be broken, neither in anger nor in battle.
DAN|11|21|In his place shall arise a contemptible person to whom royal majesty has not been given. He shall come in without warning and obtain the kingdom by flatteries.
DAN|11|22|Armies shall be utterly swept away before him and broken, even the prince of the covenant.
DAN|11|23|And from the time that an alliance is made with him he shall act deceitfully, and he shall become strong with a small people.
DAN|11|24|Without warning he shall come into the richest parts of the province, and he shall do what neither his fathers nor his fathers' fathers have done, scattering among them plunder, spoil, and goods. He shall devise plans against strongholds, but only for a time.
DAN|11|25|And he shall stir up his power and his heart against the king of the south with a great army. And the king of the south shall wage war with an exceedingly great and mighty army, but he shall not stand, for plots shall be devised against him.
DAN|11|26|Even those who eat his food shall break him. His army shall be swept away, and many shall fall down slain.
DAN|11|27|And as for the two kings, their hearts shall be bent on doing evil. They shall speak lies at the same table, but to no avail, for the end is yet to be at the time appointed.
DAN|11|28|And he shall return to his land with great wealth, but his heart shall be set against the holy covenant. And he shall work his will and return to his own land.
DAN|11|29|"At the time appointed he shall return and come into the south, but it shall not be this time as it was before.
DAN|11|30|For ships of Kittim shall come against him, and he shall be afraid and withdraw, and shall turn back and be enraged and take action against the holy covenant. He shall turn back and pay attention to those who forsake the holy covenant.
DAN|11|31|Forces from him shall appear and profane the temple and fortress, and shall take away the regular burnt offering. And they shall set up the abomination that makes desolate.
DAN|11|32|He shall seduce with flattery those who violate the covenant, but the people who know their God shall stand firm and take action.
DAN|11|33|And the wise among the people shall make many understand, though for some days they shall stumble by sword and flame, by captivity and plunder.
DAN|11|34|When they stumble, they shall receive a little help. And many shall join themselves to them with flattery,
DAN|11|35|and some of the wise shall stumble, so that they may be refined, purified, and made white, until the time of the end, for it still awaits the appointed time.
DAN|11|36|"And the king shall do as he wills. He shall exalt himself and magnify himself above every god, and shall speak astonishing things against the God of gods. He shall prosper till the indignation is accomplished; for what is decreed shall be done.
DAN|11|37|He shall pay no attention to the gods of his fathers, or to the one beloved by women. He shall not pay attention to any other god, for he shall magnify himself above all.
DAN|11|38|He shall honor the god of fortresses instead of these. A god whom his fathers did not know he shall honor with gold and silver, with precious stones and costly gifts.
DAN|11|39|He shall deal with the strongest fortresses with the help of a foreign god. Those who acknowledge him he shall load with honor. He shall make them rulers over many and shall divide the land for a price.
DAN|11|40|"At the time of the end, the king of the south shall attack him, but the king of the north shall rush upon him like a whirlwind, with chariots and horsemen, and with many ships. And he shall come into countries and shall overflow and pass through.
DAN|11|41|He shall come into the glorious land. And tens of thousands shall fall, but these shall be delivered out of his hand: Edom and Moab and the main part of the Ammonites.
DAN|11|42|He shall stretch out his hand against the countries, and the land of Egypt shall not escape.
DAN|11|43|He shall become ruler of the treasures of gold and of silver, and all the precious things of Egypt, and the Libyans and the Cushites shall follow in his train.
DAN|11|44|But news from the east and the north shall alarm him, and he shall go out with great fury to destroy and devote many to destruction.
DAN|11|45|And he shall pitch his palatial tents between the sea and the glorious holy mountain. Yet he shall come to his end, with none to help him.
DAN|12|1|"At that time shall arise Michael, the great prince who has charge of your people. And there shall be a time of trouble, such as never has been since there was a nation till that time. But at that time your people shall be delivered, everyone whose name shall be found written in the book.
DAN|12|2|And many of those who sleep in the dust of the earth shall awake, some to everlasting life, and some to shame and everlasting contempt.
DAN|12|3|And those who are wise shall shine like the brightness of the sky above; and those who turn many to righteousness, like the stars forever and ever.
DAN|12|4|But you, Daniel, shut up the words and seal the book, until the time of the end. Many shall run to and fro, and knowledge shall increase."
DAN|12|5|Then I, Daniel, looked, and behold, two others stood, one on this bank of the stream and one on that bank of the stream.
DAN|12|6|And someone said to the man clothed in linen, who was above the waters of the stream, "How long shall it be till the end of these wonders?"
DAN|12|7|And I heard the man clothed in linen, who was above the waters of the stream; he raised his right hand and his left hand toward heaven and swore by him who lives forever that it would be for a time, times, and half a time, and that when the shattering of the power of the holy people comes to an end all these things would be finished.
DAN|12|8|I heard, but I did not understand. Then I said, "O my lord, what shall be the outcome of these things?"
DAN|12|9|He said, "Go your way, Daniel, for the words are shut up and sealed until the time of the end.
DAN|12|10|Many shall purify themselves and make themselves white and be refined, but the wicked shall act wickedly. And none of the wicked shall understand, but those who are wise shall understand.
DAN|12|11|And from the time that the regular burnt offering is taken away and the abomination that makes desolate is set up, there shall be 1,290 days.
DAN|12|12|Blessed is he who waits and arrives at the 1,335 days.
DAN|12|13|But go your way till the end. And you shall rest and shall stand in your allotted place at the end of the days."
