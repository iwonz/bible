JOSH|1|1|耶和华的仆人 摩西 死了以后，耶和华对 摩西 的助手 嫩 的儿子 约书亚 说：
JOSH|1|2|“我的仆人 摩西 死了。现在你要起来，和众百姓过这 约旦河 ，往我所要赐给 以色列 人的地去。
JOSH|1|3|凡你们脚掌所踏之地，我都照我所应许 摩西 的话赐给你们了。
JOSH|1|4|从旷野和这 黎巴嫩 ，直到 大河 ，就是 幼发拉底河 ， 赫 人的全地，又到 大海 日落的方向，都要作你们的疆土。
JOSH|1|5|你一生的日子，必无人能在你面前站立得住。我怎样与 摩西 同在，也必照样与你同在；我必不撇下你，也不丢弃你。
JOSH|1|6|你当刚强壮胆，因为你必使这百姓承受那地为业，就是我向他们列祖起誓要给他们的地。
JOSH|1|7|只要刚强，大大壮胆，谨守遵行我仆人 摩西 所吩咐你的一切律法，不可偏离左右，使你无论往哪里去， 都可以顺利。
JOSH|1|8|这律法书不可离开你的口，总要昼夜思想 ，好使你谨守遵行这书上所写的一切话。如此，你的道路就可以亨通，凡事顺利。
JOSH|1|9|我岂没有吩咐你吗？你当刚强壮胆，不要惧怕，也不要惊惶，因为你无论往哪里去，耶和华你的上帝必与你同在。”
JOSH|1|10|于是， 约书亚 吩咐百姓的官长说：
JOSH|1|11|“你们要走遍营中，吩咐百姓说：‘当预备食物， 因为三日之内你们要过这 约旦河 ，进去得耶和华－你们上帝赐给你们为业之地。’”
JOSH|1|12|约书亚 对 吕便 人、 迦得 人和 玛拿西 半支派的人说：
JOSH|1|13|“你们要记得耶和华的仆人 摩西 所吩咐你们的话说：‘耶和华－你们的上帝使你们得享安宁，必将这地赐给你们。’
JOSH|1|14|你们的妻子、孩子和牲畜可以留在 约旦河 东、 摩西 所给你们的地。但你们中间所有大能的勇士都要带着兵器，在你们的弟兄前面过去，你们要帮助他们。
JOSH|1|15|等到耶和华使你们的弟兄和你们一样得享平静，并且得着耶和华－你们上帝所赐他们为业之地的时候，你们才可以回到你们所得之地，承受为业，就是耶和华的仆人 摩西 在 约旦河 东、向日出的方向所给你们的地。”
JOSH|1|16|他们回答 约书亚 说：“凡你吩咐我们的，我们都必做；凡你差我们去的地方，我们都必去。
JOSH|1|17|我们在一切事上怎样听从 摩西 ，也必照样听从你。惟愿耶和华－你的上帝与你同在，像与 摩西 同在一样。
JOSH|1|18|无论什么人违背你的命令，不听从你所吩咐他的一切话，就必处死。你只要刚强壮胆！”
JOSH|2|1|嫩 的儿子 约书亚 从 什亭 暗中派两个人作探子，说：“你们去窥探那地和 耶利哥 。”于是二人去了，来到一个名叫 喇合 的妓女家里，在那里睡觉。
JOSH|2|2|有人告诉 耶利哥 王说：“看哪，今夜有 以色列 人到这里来窥探此地。”
JOSH|2|3|耶利哥 王派人到 喇合 那里， 说：“你要交出那来到你这里、进了你家的人，因为他们来是要窥探全地。”
JOSH|2|4|但女人已把二人藏起来，却说：“那两个人确实到我这里来过，他们从哪里来，我却不知道。
JOSH|2|5|天黑、要关城门的时候，他们就出去了。他们往哪里去我也不知道。你们赶快去追他们，就必追上。”
JOSH|2|6|其实，这女人已经领二人上了屋顶，把他们藏在她摆列在屋顶的的亚麻梗中。
JOSH|2|7|那些人就往 约旦河 的路上追赶他们，直到渡口。追赶他们的人一出去，城门就关了。
JOSH|2|8|二人还没有睡之前，女人就上屋顶，到他们那里，
JOSH|2|9|对他们说：“我知道耶和华已经把这地赐给你们了，并且我们也都惧怕你们。这地所有的居民在你们面前都融化了。
JOSH|2|10|因为我们听见你们出 埃及 的时候，耶和华怎样在你们前面使 红海 的水干了，并且你们怎样处置 约旦河 东的两个 亚摩利 王， 西宏 和 噩 ，把他们完全消灭。
JOSH|2|11|我们一听见就胆战心惊 ，人人因你们的缘故勇气全失。耶和华－你们的上帝是天上地下的上帝。
JOSH|2|12|现在我既然恩待你们，求你们指着耶和华向我起誓，你们也要恩待我的父家。请你们给我一个确实的凭据，
JOSH|2|13|要救活我的父母、兄弟、姊妹，和所有属他们的，拯救我们的性命脱离死亡。”
JOSH|2|14|那二人对她说：“我们愿意以性命来替你们死。你们若不泄漏我们这件事，当耶和华将这地赐给我们的时候，我们必以慈爱和诚信待你。”
JOSH|2|15|于是女人用绳子把二人从窗户缒下去，因为她的屋子是在城墙边上，她也住在城墙上。
JOSH|2|16|她对他们说：“你们暂且往山上去，免得追赶的人遇见你们。要在那里躲藏三天，等追赶的人回来，你们才可以走自己的路。”
JOSH|2|17|二人对她说：“你叫我们所起的誓与我们无关，
JOSH|2|18|除非，看哪，当我们来到这地的时候，你把这条朱红线绳子系在缒我们下去的窗户上，并要叫你的父母、兄弟和你父的全家都聚集在你家中。
JOSH|2|19|凡离开你家门往街上去的，他的血必归到自己头上，与我们无关；凡在你家里的，若有人下手害他，他的血就归到我们头上。
JOSH|2|20|你若泄漏我们这件事，你叫我们所起的誓 就与我们无关了。”
JOSH|2|21|女人说：“就照你们的话吧！”于是她送他们走了，就把朱红绳子系在窗户上。
JOSH|2|22|二人离开，到山上去，在那里停留三天，直等到追赶的人回去。追赶的人一路寻找，却找不着。
JOSH|2|23|二人回来，下了山，过了河，来到 嫩 的儿子 约书亚 那里，向他报告他们所遭遇的一切事。
JOSH|2|24|他们对 约书亚 说：“耶和华果然将那全地交在我们手中了，并且那地所有的居民在我们面前都融化了。”
JOSH|3|1|约书亚 清早起来，和 以色列 众人起行，离开 什亭 ，来到 约旦河 ，过河以前住在那里。
JOSH|3|2|过了三天，官长走遍营中，
JOSH|3|3|吩咐百姓说：“当你们看见 利未 家的祭司抬着耶和华－你们上帝的约柜的时候，你们就要起行离开所住的地方，跟着约柜走，
JOSH|3|4|使你们知道所当走的路，因为这条路是你们从来没有走过的。只是你们要与约柜相隔约二千肘，不可太靠近约柜。”
JOSH|3|5|约书亚 吩咐百姓说：“你们要使自己分别为圣，因为明天耶和华必在你们中间行奇事。”
JOSH|3|6|约书亚 对祭司说：“你们抬起约柜，在百姓的前面过去。”于是他们抬起约柜，走在百姓前面。
JOSH|3|7|耶和华对 约书亚 说：“从今日起，我必使你在 以色列 众人眼前被尊为大，使他们知道我怎样与 摩西 同在，也必照样与你同在。
JOSH|3|8|你要吩咐抬约柜的祭司说：‘你们到了 约旦河 的水边，要在 约旦河 中站着。’”
JOSH|3|9|约书亚 对 以色列 人说：“你们近前，到这里来，听耶和华－你们上帝的话。”
JOSH|3|10|约书亚 说：“你们因这事会知道永生的上帝在你们中间，他必从你们面前赶出 迦南 人、 赫 人、 希未 人、 比利洗 人、 革迦撒 人、 亚摩利 人、 耶布斯 人。
JOSH|3|11|看哪！全地之主的约柜必在你们的前面过去，到 约旦河 里。
JOSH|3|12|现在， 你们要从 以色列 支派中选出十二个人，每支派一人。
JOSH|3|13|当抬耶和华全地之主约柜的祭司，脚掌踏入 约旦河 水里的时候， 约旦河 的水，就是从上往下流的水，必然中断，竖立成垒。”
JOSH|3|14|百姓起行离开帐棚过 约旦河 的时候，抬约柜的祭司在百姓的前面。
JOSH|3|15|那时正是收割的日子， 约旦河 的水涨满两岸。抬约柜的人到了 约旦河 ，抬约柜的祭司脚一入水边，
JOSH|3|16|那从上往下流的水就在很远的地方，在 撒拉但 旁边的 亚当城 那里停住，竖立成垒；那往 亚拉巴海 ，就是 盐海 下流的水全然中断。于是，百姓在 耶利哥 的对面过了河。
JOSH|3|17|抬耶和华约柜的祭司在 约旦河 中的干地上稳稳站着， 以色列 众人都从干地上过去，直到全国都过了 约旦河 。
JOSH|4|1|当全国都过了 约旦河 ，耶和华对 约书亚 说：
JOSH|4|2|“你要从百姓中选出十二个人，每支派一人，
JOSH|4|3|吩咐他们说：‘你们从这里，从 约旦河 中祭司的脚稳稳站立的地方，取十二块石头 ，一起带过去，放在你们今夜住宿的地方。’”
JOSH|4|4|于是 约书亚 召集了他从 以色列 人中所选的十二个人，每支派一人。
JOSH|4|5|约书亚 对他们说：“你们要过去，到 约旦河 中，耶和华－你们上帝的约柜前面，按 以色列 人支派的数目，每人各取一块石头扛在肩上。
JOSH|4|6|这些石头在你们中间将成为记号。日后，你们的子孙问你们说：‘这些石头对你们有什么意思呢？’
JOSH|4|7|你们就对他们说：‘这是因为 约旦河 的水在耶和华的约柜前中断；约柜过 约旦河 的时候， 约旦河 的水就中断了。这些石头要作 以色列 人永远的纪念。’”
JOSH|4|8|以色列 人就照 约书亚 所吩咐的做了。他们按 以色列 人支派的数目，从 约旦河 中取了十二块石头，正如耶和华所吩咐 约书亚 的。他们把石头带过去，到他们所住宿的地方，就放在那里。
JOSH|4|9|约书亚 另外把十二块石头立在 约旦河 的中间，在抬约柜祭司的脚站立的地方；直到今日，石头还在那里。
JOSH|4|10|抬约柜的祭司站在 约旦河 的中间，直到耶和华命令 约书亚 告诉百姓的一切事办完为止，正如 摩西 所吩咐 约书亚 的一切话。 于是，百姓急速过了河。
JOSH|4|11|全体百姓都过了河之后，耶和华的约柜和祭司才过去，到百姓的前面。
JOSH|4|12|吕便 人、 迦得 人、 玛拿西 半支派的人都照 摩西 所吩咐他们的，带着兵器在 以色列 人的前面过去。
JOSH|4|13|约有四万带兵器的军队在耶和华面前过去，到 耶利哥 的平原，准备上阵。
JOSH|4|14|在那日，耶和华使 约书亚 在 以色列 众人眼前被尊为大。在他一生的年日中，百姓敬服他，像从前敬服 摩西 一样。
JOSH|4|15|耶和华对 约书亚 说：
JOSH|4|16|“你吩咐抬法柜的祭司从 约旦河 上来。”
JOSH|4|17|约书亚 就吩咐祭司说：“你们从 约旦河 上来。”
JOSH|4|18|抬耶和华约柜的祭司从 约旦河 中上来，脚掌一落干地， 约旦河 的水就流回原处，仍旧涨满两岸。
JOSH|4|19|正月初十，百姓从 约旦河 上来，就在 耶利哥 东边的 吉甲 安营。
JOSH|4|20|约书亚 把他们从 约旦河 取来的那十二块石头立在 吉甲 ，
JOSH|4|21|对 以色列 人说：“日后，你们的子孙问他们的父亲说：‘这些石头是什么意思呢？’
JOSH|4|22|你们就让你们的子孙知道，说：‘ 以色列 人曾走干地过这 约旦河 。’
JOSH|4|23|因为耶和华－你们的上帝在你们前面使 约旦河 的水干了，直到你们过来，就如耶和华－你们的上帝从前在我们前面使 红海 干了，直到我们过来一样，
JOSH|4|24|要使地上万民都知道，耶和华的手大有能力，也要使你们天天敬畏耶和华－你们的上帝。”
JOSH|5|1|约旦河 西 亚摩利 人的众王和靠海 迦南 人的众王，听见耶和华在 以色列 人前面使 约旦河 的水干了，直到他们过了河 ，众王因 以色列 人的缘故都胆战心惊，勇气全失。
JOSH|5|2|那时，耶和华对 约书亚 说：“你要造火石刀，第二次为 以色列 人行割礼。”
JOSH|5|3|约书亚 就造了火石刀，在 哈尔拉勒山 为 以色列 人行割礼。
JOSH|5|4|约书亚 行割礼的原因是这样：从 埃及 出来的众百姓，所有能打仗的男丁，出了 埃及 以后，都死在旷野的路上。
JOSH|5|5|这些从 埃及 出来的众百姓都受过割礼；但是那些出 埃及 以后，在旷野的路上所生的众百姓却没有受过割礼。
JOSH|5|6|以色列 人在旷野走了四十年，直到那从 埃及 出来，全国能打仗的人都消灭了，因为他们没有听从耶和华的话。耶和华曾向他们起誓，必不容许他们看见耶和华向他们列祖起誓要给我们的地，就是流奶与蜜之地。
JOSH|5|7|他们的子孙，就是耶和华兴起接续他们的，都没有受过割礼；因为在路上他们没有受割礼， 约书亚 就为他们行割礼。
JOSH|5|8|全国的人都受了割礼，留在营中自己的地方，直到痊愈。
JOSH|5|9|耶和华对 约书亚 说：“我今日将 埃及 的羞辱从你们身上除掉了。”因此，那地方名叫 吉甲 ，直到今日。
JOSH|5|10|以色列 人在 吉甲 安营。正月十四日晚上，他们在 耶利哥 的平原守逾越节。
JOSH|5|11|逾越节的第二日，他们吃了当地的出产，就在那一天，吃了无酵饼和烘过的谷物。
JOSH|5|12|他们吃了当地出产的第二日，吗哪就停止了。 以色列 人不再有吗哪了。那一年，他们就吃 迦南 地的出产。
JOSH|5|13|约书亚 靠近 耶利哥 的时候，举目观看，看哪，有一个人站在他对面，手里拿着拔出来的刀。 约书亚 到他那里，对他说：“你是属我们的，还是属我们敌人的呢？”
JOSH|5|14|他说：“不，我现在来是要作耶和华军队的元帅。” 约书亚 就脸伏于地下拜，说：“我主有什么话，请吩咐仆人吧！”
JOSH|5|15|耶和华军队的元帅对 约书亚 说：“把你脚上的鞋脱下来，因为你所站的地方是圣的。” 约书亚 就照着做了。
JOSH|6|1|耶利哥 的城门因 以色列 人的缘故，关得严紧，无人出入。
JOSH|6|2|耶和华对 约书亚 说：“看，我已经把 耶利哥城 和 耶利哥 王，以及大能的勇士，都交在你手中。
JOSH|6|3|你们要围绕这城，所有的士兵绕城一次，六日你都要这样做。
JOSH|6|4|七个祭司要拿七个羊角走在约柜前。到了第七日，你们要围绕这城七次，祭司也要吹角。
JOSH|6|5|羊角声拖长的时候，你们一听见角声，众百姓要大声呼喊，城墙就必倒塌，各人要往前直上。”
JOSH|6|6|嫩 的儿子 约书亚 召了祭司来，对他们说：“你们抬起约柜来，要有七个祭司拿七个羊角在耶和华的约柜前。”
JOSH|6|7|他又对百姓说：“你们向前去围绕那城，带兵器的要在耶和华的约柜前过去。”
JOSH|6|8|按照 约书亚 对百姓所说的，七个祭司拿了七个羊角在耶和华面前过去，他们吹着角，耶和华的约柜在他们后面跟着。
JOSH|6|9|带兵器的走在吹角的祭司前面，后队跟着约柜走，号角继续在吹。
JOSH|6|10|约书亚 吩咐百姓说：“你们不可呼喊，不可让人听见你们的声音，连一句话也不可出你们的口，直到我对你们说‘呼喊’的那日，你们才呼喊。”
JOSH|6|11|这样， 约书亚 使耶和华的约柜围绕那城，把城绕了一次。然后，众人回到营里，就在营里住宿。
JOSH|6|12|约书亚 清早起来，祭司又抬起耶和华的约柜。
JOSH|6|13|七个祭司拿七个羊角，走在耶和华的约柜前，他们吹着角；带兵器的走在他们前面，后队跟着耶和华的约柜走，号角继续在吹。
JOSH|6|14|第二日，他们再把城围绕一次，就回营里去。六日都是这样做。
JOSH|6|15|第七日清早黎明时，他们起来，以同样的方式围绕城七次；惟独这一日他们围绕城七次。
JOSH|6|16|到了第七次，祭司吹角的时候， 约书亚 对百姓说：“呼喊吧，因为耶和华已经把城交给你们了！
JOSH|6|17|这城和其中所有的都要永献给耶和华作当毁灭的，只有妓女 喇合 与她家中所有的可以存活，因为她隐藏了我们所派的使者。
JOSH|6|18|但你们务必谨慎，不可取那当灭的物，免得你们受诅咒，取了那当灭的物，使 以色列 全营成为诅咒而遭受灾祸。
JOSH|6|19|只有金子、银子和铜铁的器皿都要归耶和华为圣，放入耶和华的库房中。”
JOSH|6|20|于是百姓呼喊，祭司吹角。百姓一听见角声就大声呼喊，城墙随着倒塌。百姓上去进城，各人往前直上，把城夺取。
JOSH|6|21|他们把城中所有的，无论男女老少，牛羊和驴，都用刀杀尽。
JOSH|6|22|约书亚 对窥探这地的两个人说：“你们进那妓女的家，照你们向她所起的誓，将那女人和她所有的都从那里带出来。”
JOSH|6|23|两个作过探子的青年进去，把 喇合 与她的父母、兄弟，和她所有的带出来，他们把她所有的亲属都带出来，安置在 以色列 的营外。
JOSH|6|24|他们用火焚烧了那城和其中所有的，只有金子、银子和铜铁的器皿都放在耶和华殿的库房中。
JOSH|6|25|至于妓女 喇合 和她父家，以及她所有的， 约书亚 保存了他们的性命。她就住在 以色列 中，直到今日，因为她隐藏了 约书亚 派来窥探 耶利哥 的使者。
JOSH|6|26|当时， 约书亚 叫众人起誓说：“凡兴起重修这 耶利哥城 的，当在耶和华面前受诅咒。 他立根基的时候，必丧长子， 安城门的时候，必丧幼子。”
JOSH|6|27|耶和华与 约书亚 同在， 约书亚 的名声传遍全地。
JOSH|7|1|以色列 人在当灭之物上犯了罪。 犹大 支派中， 谢拉 的曾孙， 撒底 的孙子， 迦米 的儿子 亚干 取了当灭之物，耶和华的怒气就向 以色列 人发作。
JOSH|7|2|约书亚 从 耶利哥 派人往 伯特利 东边，靠近 伯．亚文 的 艾城 去，对他们说：“你们上去窥探那地。”那些人就上去窥探 艾城 。
JOSH|7|3|他们回到 约书亚 那里，对他说：“众百姓不必都上去，只要二、三千人上去就能攻取 艾城 ；不必劳动众百姓都上去，因为他们人少。”
JOSH|7|4|于是百姓中约有三千人上那里去，但他们竟在 艾城 的人面前逃跑。
JOSH|7|5|艾城 的人击杀他们约三十六人，从城门前追赶他们，直到 示巴琳 ，在下坡的地方击败他们。他们都胆战心惊，融化如水。
JOSH|7|6|约书亚 和 以色列 的长老就撕裂衣服，在耶和华的约柜前脸伏于地，直到晚上。他们把灰撒在头上。
JOSH|7|7|约书亚 说：“唉！主耶和华啊，你为什么领这百姓过 约旦河 ，把我们交在 亚摩利 人手中，使我们灭亡呢？我们不如住在 约旦河 的那边！
JOSH|7|8|主啊，求求你， 以色列 人既在仇敌面前转身逃跑，我还有什么可说的呢？
JOSH|7|9|迦南 人和这地所有的居民听见了就必围困我们，把我们的名从地上除去。那时，你为你至大的名要怎样做呢？”
JOSH|7|10|耶和华对 约书亚 说：“起来！你的脸为何这样俯伏呢？
JOSH|7|11|以色列 犯了罪，又违背了我所吩咐他们的约，又取了当灭之物。他们又偷窃，又行诡诈，又把那当灭的物与自己的器皿放在一起。
JOSH|7|12|因此， 以色列 人在仇敌面前站立不住。他们在仇敌面前转身逃跑，因为他们成了当灭的物。你们若不把当灭的物从你们中间除掉，我就不再与你们同在了。
JOSH|7|13|你起来，去叫百姓分别为圣，说：‘你们要为了明天使自己分别为圣，因为耶和华－ 以色列 的上帝这样说： 以色列 啊，在你中间有当灭的物；你们若不把你们中间当灭之物除掉，你在仇敌面前必站立不住！’
JOSH|7|14|到了早晨，你们要按着支派近前来。耶和华所选的支派，要按着宗族近前来；耶和华所选的宗族，要按着家族近前来；耶和华所选的家族，要按着男丁，一个一个近前来。
JOSH|7|15|被选的人有当灭之物在他那里，他和他所有的必被火焚烧，因为他违背了耶和华的约，又因他在 以色列 中做了愚妄的事。”
JOSH|7|16|于是， 约书亚 清早起来，召 以色列 按着支派近前来。选出来的是 犹大 支派。
JOSH|7|17|他召 犹大 的宗族近前来，选出来的是 谢拉 宗族。他召 谢拉 宗族，按着男丁 ，一个一个近前来，选出来的是 撒底 。
JOSH|7|18|他召 撒底 的家族，按着男丁，一个一个近前来，就选出 犹大 支派， 谢拉 的曾孙， 撒底 的孙子， 迦米 的儿子 亚干 。
JOSH|7|19|约书亚 对 亚干 说：“我儿，我劝你将荣耀归给耶和华－ 以色列 的上帝，在他面前认罪，把你所做的事告诉我，不可向我隐瞒。”
JOSH|7|20|亚干 回答 约书亚 说：“我实在得罪了耶和华－ 以色列 的上帝。这是我所做的：
JOSH|7|21|我在所夺取的财物中看见一件美好的 示拿 外袍，二百舍客勒银子，一条重五十舍客勒的金子。我贪爱这些物件，就拿去了。看哪，这些东西都埋在我帐棚内的地里，银子在外袍底下。”
JOSH|7|22|约书亚 就派使者跑到 亚干 的帐棚里。看哪，那件外袍藏在他的帐棚里，银子在外袍底下。
JOSH|7|23|他们从帐棚里把这些东西取出来，拿到 约书亚 和 以色列 众人 那里，倒在耶和华面前。
JOSH|7|24|约书亚 和 以色列 众人把 谢拉 的曾孙 亚干 和那银子、那件外袍、那条金子，以及 亚干 的儿女、牛、驴、羊、帐棚，和他所有的，都带着上到 亚割谷 去。
JOSH|7|25|约书亚 说：“你为什么给我们招惹灾祸呢？今日耶和华必使你遭受灾祸。”于是 以色列 众人用石头打死他，用火焚烧他们，把石头扔在其上。
JOSH|7|26|众人在 亚干 身上堆了一大堆石头，直存到今日。于是耶和华转意，不发他的烈怒。因此，那地方名叫 亚割谷 ，直到今日。
JOSH|8|1|耶和华对 约书亚 说：“不要惧怕，也不要惊惶。你起来，率领所有作战的士兵上 艾城 去。看，我已经把 艾城 的王和他的百姓、他的城，以及他的地，都交在你手里。
JOSH|8|2|你怎样处置 耶利哥 和 耶利哥 的王，也当照样处置 艾城 和 艾城 的王。只是城内所夺的财物和牲畜，你们可以取为自己的掠物。你要在城的后面设下伏兵。
JOSH|8|3|于是， 约书亚 和所有作战的士兵都起来，上 艾城 去。 约书亚 选了三万大能的勇士，夜间派遣他们前去，
JOSH|8|4|吩咐他们说：“看，你们要在城的后面埋伏，不可离城太远，各人都要准备。
JOSH|8|5|我与我所带领的众士兵要向城前进。城里的人像上一次那样出来迎击我们的时候，我们就在他们面前逃跑。
JOSH|8|6|他们会出来追赶我们，直到我们引诱他们远离那城。因为他们必说：‘这些人像上次那样在我们面前逃跑。’所以我们要在他们面前逃跑 。
JOSH|8|7|那时，你们就从埋伏的地方起来，夺取那城，因为耶和华－你们的上帝必把城交在你们的手里。
JOSH|8|8|你们夺了城以后，要放火烧城，照耶和华的话去做。看，这是我吩咐你们的。”
JOSH|8|9|于是， 约书亚 派遣他们前去。他们行军到埋伏的地方，伏在 伯特利 和 艾城 的中间，就是 艾城 的西边。这夜， 约书亚 在士兵中间过夜。
JOSH|8|10|约书亚 清早起来，点齐士兵。他和 以色列 的长老在百姓前面上 艾城 去。
JOSH|8|11|所有跟他一起作战的士兵都上去，向前逼近，来到城前，就在 艾城 北边安营。 约书亚 与 艾城 之间隔着一个山谷。
JOSH|8|12|他选了约五千人，安排他们埋伏在 伯特利 和 艾城 的中间，就是 艾城 的西边。
JOSH|8|13|于是，他们布署军队，就是城北的全军和城西的伏兵。当夜 约书亚 进入山谷之中。
JOSH|8|14|艾城 的王看见了，就和城里的人清早起来，急忙出去，他和所有的士兵到了所定的地点，在 亚拉巴 前，迎击 以色列 ，与之交战；王并不知道城的后面有伏兵。
JOSH|8|15|约书亚 和 以色列 众人在他们面前装败，往旷野的路逃跑。
JOSH|8|16|城内所有的百姓都被召来追赶他们。 艾城 的人追赶 约书亚 的时候，就被引诱远离了城。
JOSH|8|17|艾城 和 伯特利 没有一人不出来追赶 以色列 人的。他们撇下敞开的城门，去追赶 以色列 人。
JOSH|8|18|耶和华对 约书亚 说：“你向 艾城 伸出手里的标枪，因为我要把那城交在你手里。” 约书亚 就向那城伸出手里的标枪。
JOSH|8|19|他一伸手，伏兵立刻从埋伏的地方冲出来，直攻入城，夺了它，立刻放火烧城。
JOSH|8|20|艾城 的人回头，往后一看，看哪，城中烟气冲天，他们向这边或那边都无处可逃。往旷野逃跑的百姓就转身攻击那些追赶他们的人。
JOSH|8|21|约书亚 和 以色列 众人见伏兵已经夺了城，城中烟气上腾，就转身击杀 艾城 的人。
JOSH|8|22|伏兵也出城追击他们，他们就被 以色列 人前后夹攻，四面受敌。于是 以色列 人击杀他们，没有留下一个幸存者，也没有一个逃脱。
JOSH|8|23|以色列 人生擒了 艾城 的王，把他解到 约书亚 那里。
JOSH|8|24|以色列 人在田间和旷野杀尽了追赶他们的 艾城 所有的居民。他们全倒在刀下，直到灭尽。 以色列 众人就回到 艾城 ，用刀杀了城中的人。
JOSH|8|25|当日杀死的人，连男带女共有一万二千，这也是 艾城 所有的人。
JOSH|8|26|约书亚 没有收回手里所伸出来的标枪，直到他灭绝 艾城 所有的居民。
JOSH|8|27|只是牲畜和城内所夺的财物， 以色列 人都照耶和华所吩咐 约书亚 的话，取为自己的掠物。
JOSH|8|28|约书亚 焚烧 艾城 ，使城成为永远的废墟，直到今日还是荒凉。
JOSH|8|29|他把 艾城 的王挂在树上，直到晚上。日落的时候， 约书亚 吩咐人把尸首从树上取下来，丢在城门口，并在尸首上堆了一大堆石头，直存到今日。
JOSH|8|30|那时， 约书亚 在 以巴路山 上为耶和华－ 以色列 的上帝筑一座坛。
JOSH|8|31|这坛是照耶和华的仆人 摩西 吩咐 以色列 人，用没有动过铁器的整块石头所筑的，正如 摩西 律法书上所写的。他们在这坛上给耶和华奉献燔祭，又宰牲作为平安祭。
JOSH|8|32|约书亚 在那里，当着 以色列 人面前，将 摩西 所写的律法抄写在石头上。
JOSH|8|33|以色列 众人，无论是本地人或寄居的，都和他们的长老、官长和审判官，站在约柜两旁，在抬耶和华约柜的 利未 家的祭司面前，一半对着 基利心山 ，一半对着 以巴路山 ，照耶和华的仆人 摩西 先前所吩咐的，为 以色列 百姓祝福。
JOSH|8|34|随后， 约书亚 将律法上祝福和诅咒的话，照着律法书上一切所写的，宣读一遍。
JOSH|8|35|摩西 所吩咐的一切话， 约书亚 在 以色列 全会众和妇女、孩童，以及住在他们中间的外人面前，没有一句不宣读的。
JOSH|9|1|约旦河 西，住山区、低地和沿 大海 一带直到 黎巴嫩 的诸王，就是 赫 人、 亚摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人的诸王，听见这事，
JOSH|9|2|就都聚集，同心合意要与 约书亚 和 以色列 人作战。
JOSH|9|3|基遍 的居民听见 约书亚 向 耶利哥 和 艾城 所做的事，
JOSH|9|4|就设诡计，假扮使者 出去。他们拿旧布袋和破裂补过的旧皮酒袋驮在驴上，
JOSH|9|5|将补过的旧鞋穿在脚上，把旧衣服穿在身上，作食物的饼都又干又长了霉 。
JOSH|9|6|他们到 吉甲 营中 约书亚 那里，对他和 以色列 人说：“我们是从远地来的，现在求你与我们立约。”
JOSH|9|7|以色列 人对 希未 人说：“或许你是住在我附近的。若是这样，我怎能和你立约呢？”
JOSH|9|8|他们对 约书亚 说：“我们是你的仆人。” 约书亚 对他们说：“你们是什么人？是从哪里来的？”
JOSH|9|9|他们对他说：“你的仆人是因耶和华－你上帝的名从极远之地来的。我们听见他的名声，他在 埃及 所做的一切，
JOSH|9|10|以及他向 约旦河 东的两个 亚摩利 王， 希实本 王 西宏 和在 亚斯她录 的 巴珊 王 噩 所做的一切。
JOSH|9|11|我们的长老和我们当地所有的居民对我们说：‘你们手里要带着路上用的干粮去迎接 以色列 人，对他们说：我们是你们的仆人。现在求你们与我们立约。’
JOSH|9|12|我们出来要往你们这里来的那日，这从我们家里带出来的饼是热的；看哪，现在这饼又干又长了霉。
JOSH|9|13|这些皮酒袋，我们盛酒的时候还是新的；看哪，现在已经破裂了。我们这些衣服和鞋，因为路途非常遥远，也都穿旧了。”
JOSH|9|14|以色列 人收下他们的一些食物，但是没有求问耶和华的指示。
JOSH|9|15|于是 约书亚 与他们建立和好关系，与他们立约，让他们存活；会众的领袖也向他们起誓。
JOSH|9|16|以色列 人与他们立约之后，过了三天才听说他们是近邻，住在附近。
JOSH|9|17|以色列 人起行，第三天就到了他们的城镇，他们的城镇是 基遍 、 基非拉 、 比录 和 基列．耶琳 。
JOSH|9|18|因为会众的领袖已经指着耶和华－ 以色列 的上帝向他们起誓，所以 以色列 人不击杀他们。全会众就向领袖发怨言。
JOSH|9|19|众领袖对全会众说：“我们已经指着耶和华－ 以色列 的上帝向他们起誓，现在我们不能碰他们。
JOSH|9|20|我们要这样对待他们，让他们存活，免得因我们向他们所起的誓而愤怒临到我们。”
JOSH|9|21|领袖对会众说：“让他们活着吧。”于是他们照领袖所说的，为全会众作劈柴挑水的人。
JOSH|9|22|约书亚 召了他们来，对他们说：“你们为什么欺骗我们说：‘我们离你们很远’呢？其实你们就住在我们附近。
JOSH|9|23|现在你们当受诅咒！你们中间必不断有人作奴仆，为我上帝的殿作劈柴挑水的人。”
JOSH|9|24|他们回答 约书亚 说：“因为确实有人告诉你的仆人，耶和华－你的上帝曾吩咐他的仆人 摩西 ，把这全地赐给你们，并要在你们面前除灭这地所有的居民。我们因你们的缘故很怕自己丧命，就做了这事。
JOSH|9|25|现在，看哪，我们在你手中，你看怎样待我们是好的，是对的，就这样做吧！”
JOSH|9|26|于是 约书亚 就这样对待他们，他救了他们脱离 以色列 人的手， 以色列 人没有杀他们。
JOSH|9|27|那日， 约书亚 分派他们到耶和华选择的地方，为会众和耶和华的坛劈柴挑水，直到今日。
JOSH|10|1|耶路撒冷 王 亚多尼．洗德 听见 约书亚 夺了 艾城 ，彻底毁灭，处置 艾城 和 艾城 的王像处置 耶利哥 和 耶利哥 的王一样，又听见 基遍 的居民与 以色列 人立了和约，住在他们中间，
JOSH|10|2|耶路撒冷 人就很惧怕，因为 基遍 是一座大城，如京城一样，比 艾城 更大，并且城内的人都是勇士。
JOSH|10|3|耶路撒冷 王 亚多尼．洗德 派人去见 希伯仑 王 何咸 、 耶末 王 毗兰 、 拉吉 王 雅非亚 和 伊矶伦 王 底璧 ，说：
JOSH|10|4|“求你们上来帮助我，我们好攻打 基遍 ，因为它与 约书亚 和 以色列 人立了和约。”
JOSH|10|5|于是五个 亚摩利 王，就是 耶路撒冷 王、 希伯仑 王、 耶末 王、 拉吉 王和 伊矶伦 王，联合上去，率领他们所有的军队，对着 基遍 安营，要攻打 基遍 。
JOSH|10|6|基遍 人就派人到 吉甲 的营中 约书亚 那里，说：“不要袖手不顾你的仆人，求你赶快上来拯救我们，帮助我们，因为住山区 亚摩利 人的诸王已经联合来攻击我们。”
JOSH|10|7|于是 约书亚 和所有跟他一起作战的士兵，以及大能的勇士，从 吉甲 上去。
JOSH|10|8|耶和华对 约书亚 说：“不要怕他们， 因为我已将他们交在你手里，他们没有一人能在你面前站立得住。”
JOSH|10|9|约书亚 就连夜从 吉甲 上去，猛然袭击他们。
JOSH|10|10|耶和华使他们在 以色列 人面前溃乱。 约书亚 在 基遍 大大击杀他们，在 伯．和仑 的上坡路上追赶他们，击杀他们，直到 亚西加 和 玛基大 。
JOSH|10|11|他们在 以色列 人面前逃跑。正在 伯．和仑 下坡的时候，耶和华从天上降下大冰雹 在他们身上，直降到 亚西加 ，打死他们。被冰雹打死的，比 以色列 人用刀杀死的还多。
JOSH|10|12|当耶和华将 亚摩利 人交给 以色列 人的那一日， 约书亚 向耶和华说话，在 以色列 人眼前说： “太阳啊，停在 基遍 ； 月亮啊，停在 亚雅仑谷 。”
JOSH|10|13|太阳就停住，月亮就止住， 直到国民向敌人报仇。 这事岂不是写在《雅煞珥书》上吗？太阳停在天空当中，没有急速下落，约有一整天。
JOSH|10|14|在这日以前，这日以后，耶和华听人的声音，没有像这日的，这是因为耶和华为 以色列 作战。
JOSH|10|15|约书亚 和跟他一起的 以色列 众人回到 吉甲 的营中。
JOSH|10|16|那五个王逃跑，躲在 玛基大 洞里。
JOSH|10|17|有人告诉 约书亚 说：“那五个王已经找到了，都躲在 玛基大 洞里。”
JOSH|10|18|约书亚 说：“你们把几块大石头滚到洞口，派人在那里看守他们。
JOSH|10|19|你们却不可停留，要追赶你们的仇敌，从后面攻击他们，不让他们进到自己的城镇，因为耶和华－你们的上帝已经把他们交在你们手里。”
JOSH|10|20|约书亚 和 以色列 人彻底击败他们，直到把他们灭尽，只剩下少许的人逃进坚固的城。
JOSH|10|21|众百姓就安然回到 玛基大 营中 ，到 约书亚 那里。没有人敢向 以色列 人饶舌。
JOSH|10|22|约书亚 说：“打开洞口，把那五个王从洞里带出来，到我这里。”
JOSH|10|23|众人就这样做，把那五个王，就是 耶路撒冷 王、 希伯仑 王、 耶末 王、 拉吉 王和 伊矶伦 王，从洞里带出来，到 约书亚 那里。
JOSH|10|24|他们带出那五个王到 约书亚 那里的时候， 约书亚 就召了 以色列 众人来，对和他同去的军官说：“你们近前来，把脚踏在这些王的颈项上。”他们就近前来，把脚踏在这些王的颈项上。
JOSH|10|25|约书亚 对他们说：“你们不要惧怕，也不要惊惶。当刚强壮胆，因为耶和华必这样处置你们要攻打的所有仇敌。”
JOSH|10|26|随后， 约书亚 把这五个王杀死，挂在五棵树上。他们就被挂在树上，直到晚上。
JOSH|10|27|日落的时候， 约书亚 吩咐人把尸首从树上取下来，丢在他们躲过的洞里，把几块大石头放在洞口，直存到今日。
JOSH|10|28|当日， 约书亚 夺了 玛基大 ，用刀击杀城中的人和王，把城中所有人完全灭尽，没有留下一个幸存者。他处置 玛基大 王，像从前处置 耶利哥 王一样。
JOSH|10|29|约书亚 和跟他一起的 以色列 众人从 玛基大 往 立拿 去，攻打 立拿 。
JOSH|10|30|耶和华将 立拿 和 立拿 的王也交在 以色列 人手里。 约书亚 攻打这城，用刀击杀了城中所有的人，没有留下一个幸存者。他处置 立拿 王，像从前处置 耶利哥 王一样。
JOSH|10|31|约书亚 和跟他一起的 以色列 众人从 立拿 往 拉吉 去，对着 拉吉 安营，攻打这城。
JOSH|10|32|耶和华将 拉吉 交在 以色列 人的手里。第二日 约书亚 就夺了 拉吉 ，用刀击杀了城中所有的人，正如他向 立拿 一切所做的。
JOSH|10|33|那时 基色 王 何兰 上来帮助 拉吉 ， 约书亚 就把他和他的百姓都击杀了，没有留下一个幸存者。
JOSH|10|34|约书亚 和跟他一起的 以色列 众人从 拉吉 往 伊矶伦 去，对着 伊矶伦 安营，攻打这城。
JOSH|10|35|当日 约书亚 就夺了城，用刀击杀了城中的人。那日， 约书亚 把城中所有的人完全灭尽，正如他向 拉吉 一切所做的。
JOSH|10|36|约书亚 和跟他一起的 以色列 众人从 伊矶伦 上 希伯仑 去，攻打这城，
JOSH|10|37|夺了 希伯仑 ，用刀击败 希伯仑 、它的王和属它的一切城镇，以及城中所有的人；他没有留下一个幸存者，正如他向 伊矶伦 所做的，把城中所有的人完全灭尽。
JOSH|10|38|约书亚 和跟他一起的 以色列 众人回到 底璧 ，攻打这城，
JOSH|10|39|夺了 底璧 和属它的一切城镇，又擒获它的王，用刀把城中所有的人完全灭尽，没有留下一个幸存者。他处置 底璧 和它的王，像从前处置 希伯仑 ，处置 立拿 和它的王一样。
JOSH|10|40|这样， 约书亚 击败全地的人，就是山区、 尼革夫 、低地、山坡的人，和那里的众王，没有留下一个幸存者。他把凡有气息的完全灭尽，正如耶和华－ 以色列 的上帝所吩咐的。
JOSH|10|41|约书亚 从 加低斯．巴尼亚 攻到 迦萨 ，又攻打 歌珊 全地，直到 基遍 。
JOSH|10|42|约书亚 一举击败了这些王，夺了他们的地，因为耶和华－ 以色列 的上帝为 以色列 作战。
JOSH|10|43|于是 约书亚 和跟他一起的 以色列 众人回到 吉甲 的营中。
JOSH|11|1|夏琐 王 耶宾 听见了，就派人到 玛顿 王 约巴 、 伸仑 王、 押煞 王，
JOSH|11|2|和北方山区、 基尼烈 南边的 亚拉巴 、低地、西边 多珥 山冈 的诸王，
JOSH|11|3|以及东方和西方的 迦南 人、山区的 亚摩利 人、 赫 人、 比利洗 人、 耶布斯 人，和 黑门山 下 米斯巴 地的 希未 人那里。
JOSH|11|4|他们和他们的众军都出来，一大队人马，多如海边的沙，并有极多的战车战马。
JOSH|11|5|众王组成联军，来到 米伦 水边一同安营，要与 以色列 作战。
JOSH|11|6|耶和华对 约书亚 说：“你不要怕他们。明日这时，我必把他们全部交给 以色列 人杀灭。你要砍断他们马的蹄筋，用火焚烧他们的战车。”
JOSH|11|7|于是 约书亚 和所有跟他一起作战的士兵，来到 米伦 水边，突然攻击他们。
JOSH|11|8|耶和华将他们交在 以色列 人手里， 以色列 人就击杀他们，追赶他们到 西顿 大城，到 米斯利弗．玛音 ，直到东边 米斯巴 的山谷。 以色列 人击杀他们，没有留下一个幸存者。
JOSH|11|9|约书亚 照耶和华所吩咐他的去做，砍断他们马的蹄筋，用火焚烧他们的战车。
JOSH|11|10|那时， 约书亚 转回，夺了 夏琐 ，用刀杀了 夏琐 王。先前 夏琐 在这些王国中是为首的。
JOSH|11|11|以色列 人用刀击杀城中所有的人，把他们完全灭尽；凡有气息的，没有留下一个。 约书亚 又用火焚烧 夏琐 。
JOSH|11|12|约书亚 夺了这些王的一切城镇，擒获了这些王，用刀杀了他们，把他们完全灭尽，正如耶和华的仆人 摩西 所吩咐的。
JOSH|11|13|至于造在山冈上的城镇，除了 夏琐 以外， 以色列 人都没有焚烧。 约书亚 只焚烧了 夏琐 。
JOSH|11|14|从那些城镇所夺的财物和牲畜， 以色列 人都取为自己的掠物。至于所有的人，他们都用刀杀了，直到灭尽；凡有气息的，没有留下一个。
JOSH|11|15|耶和华怎样吩咐他的仆人 摩西 ， 摩西 就这样吩咐 约书亚 ， 约书亚 也照样做了。凡耶和华所吩咐 摩西 的， 约书亚 没有一件偏离不做的。
JOSH|11|16|约书亚 夺了那全地，就是山区、整个 尼革夫 、 歌珊 全地、低地、 亚拉巴 、 以色列 的山区和山下的低地，
JOSH|11|17|从上 西珥 的 哈拉山 ，直到 黑门山 下面 黎巴嫩 平原的 巴力．迦得 。他擒获了那里的众王，把他们杀死。
JOSH|11|18|约书亚 和这些王作战了很长的一段日子。
JOSH|11|19|除了 希未 人 基遍 的居民之外，没有一城与 以色列 人讲和，都是 以色列 人作战夺来的。
JOSH|11|20|因为耶和华的意思是要使他们的心刚硬，来与 以色列 人作战，好使他们全被杀灭，不蒙怜悯，反被除灭，正如耶和华所吩咐 摩西 的。
JOSH|11|21|那时 约书亚 来到，剪除了住山区、 希伯仑 、 底璧 、 亚拿伯 、整个 犹大 山区和 以色列 山区的 亚衲 族人。 约书亚 把他们和他们的城镇尽都毁灭。
JOSH|11|22|以色列 人的地中没有留下一个 亚衲 族人，只有一些还留在 迦萨 、 迦特 和 亚实突 。
JOSH|11|23|这样， 约书亚 照着耶和华所吩咐 摩西 的一切话夺了那全地，就按着 以色列 支派所得的份把地分给他们为业。于是国中太平，没有战争了。
JOSH|12|1|这些是 以色列 人在 约旦河 东，向日出的方向，从 亚嫩谷 直到 黑门山 ，以及东边 亚拉巴 的整个地区所击杀的王和所得的地：
JOSH|12|2|有住 希实本 的 亚摩利 王 西宏 ，他统治的地从 亚嫩谷 边的 亚罗珥 起，包括谷中之城和 基列 的一半，直到 亚扪 人边界的 雅博河 ，
JOSH|12|3|以及从东边的 亚拉巴 ，直到 基尼烈海 ，又向东通过 伯．耶施末 的路，直到 亚拉巴 的海，就是 盐海 ，再往南直到 毗斯迦山 斜坡的山脚。
JOSH|12|4|又有 巴珊 王 噩 ，他是 利乏音 人所剩下的，住在 亚斯她录 和 以得来 。
JOSH|12|5|他统治的地是 黑门山 、 撒迦 、 巴珊 全地，直到 基述 人和 玛迦 人的边界，以及 基列 的一半，直到 希实本 王 西宏 的边界。
JOSH|12|6|这两个王是耶和华的仆人 摩西 和 以色列 人所击杀的。耶和华的仆人 摩西 把他们的地赐给 吕便 人、 迦得 人和 玛拿西 半支派的人为业。
JOSH|12|7|这些是 约书亚 和 以色列 人在 约旦河 西所击杀的诸王，他们的地从 黎巴嫩 平原的 巴力．迦得 ，直上到 西珥 的 哈拉山 。 约书亚 按着 以色列 支派所得的份把这地分给他们为业，
JOSH|12|8|就是 赫 人、 亚摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人的地，包括山区、低地、 亚拉巴 、山坡、旷野和 尼革夫 。
JOSH|12|9|这些王是： 耶利哥 王一人， 靠近 伯特利 的 艾城 王一人，
JOSH|12|10|耶路撒冷 王一人， 希伯仑 王一人，
JOSH|12|11|耶末 王一人， 拉吉 王一人，
JOSH|12|12|伊矶伦 王一人， 基色 王一人，
JOSH|12|13|底璧 王一人， 基德 王一人，
JOSH|12|14|何珥玛 王一人， 亚拉得 王一人，
JOSH|12|15|立拿 王一人， 亚杜兰 王一人，
JOSH|12|16|玛基大 王一人， 伯特利 王一人，
JOSH|12|17|他普亚 王一人， 希弗 王一人，
JOSH|12|18|亚弗 王一人， 拉沙仑 王一人，
JOSH|12|19|玛顿 王一人， 夏琐 王一人，
JOSH|12|20|伸仑．米仑 王一人 ， 押煞 王一人，
JOSH|12|21|他纳 王一人， 米吉多 王一人，
JOSH|12|22|基低斯 王一人， 靠近 迦密 的 约念 王一人，
JOSH|12|23|多珥 山冈 的 多珥 王一人， 吉甲 的 戈印 王一人，
JOSH|12|24|得撒 王一人， 共三十一个王。
JOSH|13|1|约书亚 年纪老迈，耶和华对他说：“你年纪老迈了，还有极多剩下的未得之地。
JOSH|13|2|这是剩下的地： 非利士 人的全境和一切属于 基述 人的，
JOSH|13|3|是从 埃及 东边的 西曷河 往北，直到 以革伦 的边界，算是属 迦南 人的地，那里有 非利士 人五个领袖统治 迦萨 人、 亚实突 人、 亚实基伦 人、 迦特 人、 以革伦 人；还有属于 亚卫 人的，
JOSH|13|4|在南边；还有 迦南 人的全地，以及 西顿 人的 米亚拉 到 亚弗 ，直到 亚摩利 人的边界；
JOSH|13|5|还有 迦巴勒 人的地，以及向日出方向的 黎巴嫩 全地，从 黑门山 下的 巴力．迦得 ，直到 哈马口 ；
JOSH|13|6|从 黎巴嫩 直到 米斯利弗．玛音 ，一切山区的居民，就是所有的 西顿 人，我必在 以色列 人面前赶走他们。你只管照我所吩咐的，抽签将这地分给 以色列 人为业。
JOSH|13|7|现在你要把这地分给九个支派和 玛拿西 半个支派为业。
JOSH|13|8|吕便 、 迦得 二支派已经和 玛拿西 另外半个支派得了产业，就是耶和华的仆人 摩西 在 约旦河 东所赐给他们的：
JOSH|13|9|从 亚嫩谷 边的 亚罗珥 和谷中之城， 米底巴 的整个平原，直到 底本 ；
JOSH|13|10|还有在 希实本 作王的 亚摩利 王 西宏 的诸城，直到 亚扪 人的边界；
JOSH|13|11|还有 基列 ， 基述 人和 玛迦 人的边界，整个 黑门山 、整个 巴珊 ，直到 撒迦 ；
JOSH|13|12|还有在 亚斯她录 和 以得来 作王的 巴珊 王 噩 的整个国土， 噩 是 利乏音 人惟一存留的。 摩西 击败了这些人，把他们赶走。
JOSH|13|13|以色列 人却没有赶走 基述 人和 玛迦 人； 基述 人和 玛迦 人仍住在 以色列 中，直到今日。
JOSH|13|14|只是 利未 支派， 摩西 没有分产业给他们。他们的产业是献给耶和华－ 以色列 上帝的火祭，正如耶和华对他们说的。
JOSH|13|15|摩西 按着 吕便 支派的宗族分产业给他们。
JOSH|13|16|他们的地界是 亚嫩谷 边的 亚罗珥 和谷中之城，靠近 米底巴 的整个平原；
JOSH|13|17|还有 希实本 和属 希实本 平原的各城， 底本 、 巴末．巴力 、 伯．巴力．勉 、
JOSH|13|18|雅杂 、 基底莫 、 米法押 、
JOSH|13|19|基列亭 、 西比玛 、谷中山冈上的 细列．沙辖 、
JOSH|13|20|伯．毗珥 、 毗斯迦山 斜坡、 伯．耶施末 ；
JOSH|13|21|还有平原的各城，和 亚摩利 王 西宏 的整个国土。这 西宏 曾在 希实本 作王， 摩西 把他和 米甸 的族长 以未 、 利金 、 苏珥 、 户珥 、 利巴 击杀了；他们都是属 西宏 的领袖，曾住在这地。
JOSH|13|22|以色列 人杀了这些人时，也用刀杀了 比珥 的儿子占卜的 巴兰 。
JOSH|13|23|吕便 人的地界就是 约旦河 和靠近 约旦河 的地。以上是 吕便 人按着宗族所得为业的城镇和所属的村庄。
JOSH|13|24|摩西 按着 迦得 支派的宗族分产业给他们。
JOSH|13|25|他们的地界是 雅谢 和 基列 的各城，以及 亚扪 人之地的一半，直到 拉巴 前面的 亚罗珥 ；
JOSH|13|26|还有从 希实本 到 拉抹．米斯巴 和 比多宁 ，又从 玛哈念 到 底璧 的边界，
JOSH|13|27|和谷中的 伯．亚兰 、 伯．宁拉 、 疏割 、 撒分 ，就是 希实本 王 西宏 国土中其余的地，以及 约旦河 与靠近 约旦河 的地，直到 基尼烈海 的边缘，都在 约旦河 东。
JOSH|13|28|以上是 迦得 人按着宗族所得为业的城镇和所属的村庄。
JOSH|13|29|摩西 分产业给 玛拿西 半支派，这是按着 玛拿西 半支派的宗族分的。
JOSH|13|30|他们的地界是从 玛哈念 起，包括整个 巴珊 全地，就是 巴珊 王 噩 的整个国土，以及在 巴珊 、 睚珥 的一切城镇，共六十个；
JOSH|13|31|还有 基列 的一半，以及 巴珊 国的王 噩 的 亚斯她录 和 以得来 两座城。这些地是按着宗族分给 玛拿西 儿子 玛吉 子孙的，就是给 玛吉 一半子孙的。
JOSH|13|32|以上是 摩西 在 约旦河 东， 耶利哥 对面的 摩押 平原所分配的产业。
JOSH|13|33|只是 利未 支派， 摩西 没有把产业分给他们。耶和华－ 以色列 的上帝是他们的产业，正如耶和华对他们说的。
JOSH|14|1|这是 以色列 人在 迦南 地所得的产业，就是祭司 以利亚撒 和 嫩 的儿子 约书亚 ，以及 以色列 人各支派父系的领袖所分给他们的。
JOSH|14|2|他们照耶和华藉 摩西 所吩咐的，抽签分产业给九个半支派。
JOSH|14|3|摩西 在 约旦河 东已经分了产业给另外两个半支派。但是，他在他们中间没有分产业给 利未 人。
JOSH|14|4|因 约瑟 的子孙成了两个支派，就是 玛拿西 和 以法莲 。虽然他们没有分地给 利未 人，却给 利未 人城镇居住，以及城镇的郊外供他们牧养牲畜，安置财物。
JOSH|14|5|耶和华怎样吩咐 摩西 ， 以色列 人就照样做，把地分了。
JOSH|14|6|犹大 人来到 吉甲 ， 约书亚 那里， 基尼洗 族 耶孚尼 的儿子 迦勒 对 约书亚 说：“耶和华在 加低斯．巴尼亚 指着我和你对神人 摩西 所说的话，你都知道。
JOSH|14|7|耶和华的仆人 摩西 从 加低斯．巴尼亚 差派我窥探这地的时候，我刚四十岁。我把心里的话向他报告。
JOSH|14|8|虽然同我上去的众弟兄使百姓胆战心惊，我仍然专心跟从耶和华－我的上帝。
JOSH|14|9|那日， 摩西 起誓说：‘你脚所踏之地必要归你和你的子孙永远为业，因为你专心跟从耶和华－我的上帝。’
JOSH|14|10|现在，看哪，耶和华照他所说的使我活了这四十五年。当 以色列 人在旷野飘流的时候，耶和华曾对 摩西 说了这话。现在，看哪，我已经八十五岁了。
JOSH|14|11|现今我还很健壮，像 摩西 差派我去的那天一样；无论是战争，是出入，我现在的力量和那时的力量一样。
JOSH|14|12|请你将耶和华那日所说的这山区给我。那日你也曾听说，这里有 亚衲 族人，以及宽大坚固的城，或许耶和华会照他所说的与我同在，我就把他们赶出去。”
JOSH|14|13|于是 约书亚 为 耶孚尼 的儿子 迦勒 祝福，把 希伯仑 给他为业。
JOSH|14|14|所以 希伯仑 成了 基尼洗 族 耶孚尼 的儿子 迦勒 的产业，直到今日，因为他专心跟从耶和华－ 以色列 的上帝。
JOSH|14|15|希伯仑 从前名叫 基列．亚巴 ； 亚巴 是 亚衲 族最尊贵的人。于是国中太平，没有战争了。
JOSH|15|1|犹大 支派按着宗族抽签所得之地是在最南端，到 以东 的边界，往南直到 寻 的旷野。
JOSH|15|2|他们南边的地界是从 盐海 的顶端，就是朝南的海湾开始，
JOSH|15|3|通到 亚克拉滨 斜坡的南边，经过 寻 ，上到 加低斯．巴尼亚 的南边，又经过 希斯仑 ，上到 亚达珥 ，转到 甲加 ，
JOSH|15|4|再经过 押们 ，顺着 埃及 溪谷，这地界直通到海为止。这就是你们 南边的地界。
JOSH|15|5|东边的地界是从 盐海 到 约旦河 口。北边的地界是从 约旦河 口的海湾开始，
JOSH|15|6|这地界上到 伯．曷拉 ，经过 伯．亚拉巴 的北边，这地界上到 吕便 之子 波罕 的磐石。
JOSH|15|7|这地界是从 亚割谷 往北上到 底璧 ，直向 亚都冥 斜坡对面的 吉甲 ，就是河的南边，这地界再经过 隐．示麦 泉，直通到 隐．罗结 。
JOSH|15|8|这地界又上到 欣嫩子谷 ， 耶布斯 斜坡的南方， 耶布斯 就是 耶路撒冷 ，这地界又上到 欣嫩谷 西边对面的山顶，就是在 利乏音谷 的最北端。
JOSH|15|9|这地界又从山顶延伸到 尼弗多亚 水泉，通到 以弗仑山 的城镇，这地界又延伸到 巴拉 ， 巴拉 就是 基列．耶琳 。
JOSH|15|10|这地界又从 巴拉 往西绕到 西珥山 ，经过 耶琳山 斜坡的北边， 耶琳 就是 基撒仑 ，从那里又下到 伯．示麦 ，经过 亭拿 ，
JOSH|15|11|这地界通到 以革伦 斜坡的北边。这地界又延伸到 施基仑 ，经过 巴拉山 到 雅比聂 ，这地界直通到海为止。
JOSH|15|12|西边的地界就是 大海 和沿海一带之地。这是 犹大 人按着宗族所得之地四围的边界。
JOSH|15|13|约书亚 照耶和华所指示的，把 犹大 人中的一份土地，就是 基列．亚巴 ，分给 耶孚尼 的儿子 迦勒 。 亚巴 是 亚衲 族的祖先， 基列．亚巴 就是 希伯仑 。
JOSH|15|14|迦勒 从那里赶出 亚衲 的三族，就是 亚衲 族的 示筛 人、 亚希幔 人和 挞买 人。
JOSH|15|15|他又从那里上去，攻击 底璧 的居民，这 底璧 从前名叫 基列．西弗 。
JOSH|15|16|迦勒 说：“谁能攻打 基列．西弗 ，夺取那城，我就把我女儿 押撒 嫁给他。”
JOSH|15|17|迦勒 兄弟 基纳斯 的儿子 俄陀聂 夺取了那城， 迦勒 就把女儿 押撒 嫁给他。
JOSH|15|18|押撒 来的时候，催促丈夫向她父亲要一块田。 押撒 一下驴， 迦勒 就对她说：“你要什么？”
JOSH|15|19|她说：“求你给我福分；你既然把我安置在 尼革夫 地，求你也给我水泉。”她父亲就把上泉和下泉都赐给她。
JOSH|15|20|这是 犹大 支派按着宗族所得的产业。
JOSH|15|21|犹大 支派最南端，靠近 以东 边界的城镇，是 甲薛 、 以得 、 雅姑珥 、
JOSH|15|22|基拿 、 底摩拿 、 亚大达 、
JOSH|15|23|基低斯 、 夏琐 、 以提楠 、
JOSH|15|24|西弗 、 提鍊 、 比亚绿 、
JOSH|15|25|夏琐．哈大他 、 加略．希斯仑 ， 加略．希斯仑 就是 夏琐 ，
JOSH|15|26|亚曼 、 示玛 、 摩拉大 、
JOSH|15|27|哈萨．迦大 、 黑实门 、 伯．帕列 、
JOSH|15|28|哈萨．书亚 、 别是巴 、 比斯约他 、
JOSH|15|29|巴拉 、 以因 、 以森 、
JOSH|15|30|伊勒多腊 、 基失 、 何珥玛 、
JOSH|15|31|洗革拉 、 麦玛拿 、 三撒拿 、
JOSH|15|32|利巴勿 、 实忻 、 亚因 、 临门 ，共二十九座城，还有所属的村庄。
JOSH|15|33|在低地有 以实陶 、 琐拉 、 亚实拿 、
JOSH|15|34|撒挪亚 、 隐．干宁 、 他普亚 、 以楠 、
JOSH|15|35|耶末 、 亚杜兰 、 梭哥 、 亚西加 、
JOSH|15|36|沙拉音 、 亚底他音 、 基底拉 、 基底罗他音 ，共十四座城，还有所属的村庄。
JOSH|15|37|又有 洗楠 、 哈大沙 、 麦大．迦得 、
JOSH|15|38|底连 、 米斯巴 、 约帖 、
JOSH|15|39|拉吉 、 波斯加 、 伊矶伦 、
JOSH|15|40|迦本 、 拉幔 、 基提利 、
JOSH|15|41|基低罗 、 伯．大衮 、 拿玛 、 玛基大 ，共十六座城，还有所属的村庄。
JOSH|15|42|又有 立拿 、 以帖 、 亚珊 、
JOSH|15|43|益弗他 、 亚实拿 、 尼悉 、
JOSH|15|44|基伊拉 、 亚革悉 、 玛利沙 ，共九座城，还有所属的村庄。
JOSH|15|45|又有 以革伦 和所属的乡镇 与村庄，
JOSH|15|46|从 以革伦 直到海，一切靠近 亚实突 之地，以及所属的村庄、
JOSH|15|47|亚实突 和所属的乡镇与村庄， 迦萨 和所属的乡镇与村庄，到 埃及 溪谷，直到 大海 以及沿海一带之地。
JOSH|15|48|在山区有 沙密 、 雅提珥 、 梭哥 、
JOSH|15|49|大拿 、 基列．萨拿 ， 基列．萨拿 就是 底璧 ，
JOSH|15|50|亚拿伯 、 以实提莫 、 亚念 、
JOSH|15|51|歌珊 、 何仑 、 基罗 ，共十一座城，还有所属的村庄。
JOSH|15|52|又有 亚拉 、 度玛 、 以珊 、
JOSH|15|53|雅农 、 伯．他普亚 、 亚非加 、
JOSH|15|54|宏他 、 基列．亚巴 ， 基列．亚巴 就是 希伯仑 ， 洗珥 ，共九座城，还有所属的村庄。
JOSH|15|55|又有 玛云 、 迦密 、 西弗 、 淤他 、
JOSH|15|56|耶斯列 、 约甸 、 撒挪亚 、
JOSH|15|57|该隐 、 基比亚 、 亭拿 ，共十座城，还有所属的村庄。
JOSH|15|58|又有 哈忽 、 伯．夙 、 基突 、
JOSH|15|59|玛腊 、 伯．亚诺 、 伊勒提君 ，共六座城，还有所属的村庄。
JOSH|15|60|又有 基列．巴力 ， 基列．巴力 就是 基列．耶琳 ， 拉巴 ，共两座城，还有所属的村庄。
JOSH|15|61|在旷野有 伯．亚拉巴 、 密丁 、 西迦迦 、
JOSH|15|62|匿珊 、 盐城 、 隐．基底 ，共六座城，还有所属的村庄。
JOSH|15|63|至于住 耶路撒冷 的 耶布斯 人， 犹大 人不能把他们赶出去。于是， 耶布斯 人与 犹大 人同住在 耶路撒冷 ，直到今日。
JOSH|16|1|约瑟 的子孙抽签所得之地是从靠近 耶利哥 的 约旦河 起，以 耶利哥 东边的河水为边界，经过旷野，从 耶利哥 上去，直到 伯特利 的山区；
JOSH|16|2|从 伯特利 又到 路斯 ，经过 亚基 人的边界，直到 亚大录 ；
JOSH|16|3|又往西，下到 押利提 人的边界，到 下伯．和仑 的边界，到 基色 ，直通到海为止。
JOSH|16|4|约瑟 的儿子 玛拿西 、 以法莲 得了地业。
JOSH|16|5|以法莲 子孙的地界，按着宗族所得的如下：他们地业的东界，是从 亚大录．亚达 到 上伯．和仑 ，
JOSH|16|6|这地界直通到海。在北边，这地界是从 密米他 ，向东绕到 他纳．示罗 ，又经过 雅挪哈 的东边，
JOSH|16|7|从 雅挪哈 下到 亚大录 和 拿拉 ，再到 耶利哥 ，直到 约旦河 为止。
JOSH|16|8|这地界又从 他普亚 ，顺着 加拿河 往西延伸，直通到海为止。这就是 以法莲 支派按着宗族所得的地业。
JOSH|16|9|在 玛拿西 人地业的一切城镇和所属的村庄中，也保留一些城镇给 以法莲 的子孙。
JOSH|16|10|他们却没有赶出住在 基色 的 迦南 人。 迦南 人就住在 以法莲 人中，成为服劳役的仆人，直到今日。
JOSH|17|1|玛拿西 是 约瑟 的长子，这是他的支派抽签所得之地。 玛拿西 的长子， 基列 的父亲 玛吉 ，因为是勇士，就得了 基列 和 巴珊 。
JOSH|17|2|玛拿西 其余的子孙，就是 亚比以谢 的子孙， 希勒 的子孙， 亚斯烈 的子孙， 示剑 的子孙， 希弗 的子孙， 示米大 的子孙，都按着宗族抽签得了地。这都是 约瑟 的儿子 玛拿西 子孙中各宗族的男丁。
JOSH|17|3|玛拿西 的玄孙， 玛吉 的曾孙， 基列 的孙子， 希弗 的儿子 西罗非哈 没有儿子，只有女儿。他的女儿名叫 玛拉 、 挪阿 、 曷拉 、 密迦 、 得撒 。
JOSH|17|4|她们来到 以利亚撒 祭司和 嫩 的儿子 约书亚 以及众领袖面前，说：“耶和华曾吩咐 摩西 在我们兄弟中分产业给我们。”于是 约书亚 照耶和华的指示，在她们叔伯中，把产业分给她们。
JOSH|17|5|除了 约旦河 东的 基列 和 巴珊 地之外，还有十份的地业是属于 玛拿西 的，
JOSH|17|6|因为 玛拿西 支派的女子也在男子中分得产业。 基列 地属于 玛拿西 其余的子孙。
JOSH|17|7|玛拿西 的地界是从 亚设 起，到 示剑 前面的 密米他 ，往右 到 隐．他普亚 居民之地。
JOSH|17|8|他普亚 地归于 玛拿西 ，只是 玛拿西 边界的 他普亚城 却归于 以法莲 子孙。
JOSH|17|9|这地界从那里下到 加拿河 。河南边的城镇虽然在 玛拿西 境内，却是属于 以法莲 的。 玛拿西 的地界是在河的北边直通到海为止。
JOSH|17|10|南边属于 以法莲 ，北边属于 玛拿西 ，以海为界；北边达到 亚设 ，东边达到 以萨迦 。
JOSH|17|11|玛拿西 在 以萨迦 和 亚设 境内，有 伯．善 和所属的乡镇， 以伯莲 和所属的乡镇， 多珥 和所属乡镇的居民；还有 隐．多珥 和所属乡镇的居民， 他纳 和所属乡镇的居民， 米吉多 和所属乡镇的居民，共三个山冈 。
JOSH|17|12|只是 玛拿西 的子孙不能赶出这些城镇的居民， 迦南 人仍坚持住在那地。
JOSH|17|13|以色列 人强盛的时候，就叫 迦南 人做苦工，没有把他们全然赶走。
JOSH|17|14|约瑟 的子孙对 约书亚 说：“耶和华到如今这样赐福给我，我百姓众多，你为什么只给我抽一签，分一份的土地为业呢？”
JOSH|17|15|约书亚 对他们说：“如果你百姓众多，而 以法莲 山区太窄小，那么你可以上 比利洗 人和 利乏音 人之地的树林中，在那里开垦。”
JOSH|17|16|约瑟 的子孙说：“那山区容不下我们，而且住平原的 迦南 人，就是住 伯．善 和所属的乡镇，以及住在 耶斯列 平原的人，都有铁的战车。”
JOSH|17|17|约书亚 对 约瑟 家，就是 以法莲 和 玛拿西 人，说：“你百姓众多，并且强大，不可只有一签而已。
JOSH|17|18|那山区也要归你，虽然是树林，你可以去开垦，边缘之地也必归你。 迦南 人纵然强盛，有铁的战车，你也能把他们赶出去。”
JOSH|18|1|以色列 全会众都聚集在 示罗 ，把会幕设立在那里。那地已经被他们征服了。
JOSH|18|2|以色列 人中剩下七个支派还没有分得他们的地业。
JOSH|18|3|约书亚 对 以色列 人说：“耶和华－你们列祖的上帝所赐给你们的地，你们耽延不去得，要到几时呢？
JOSH|18|4|你们每支派要选三个人，我好派他们去，他们要起身走遍那地，按照各支派应得的地业写明，然后回到我这里来。
JOSH|18|5|他们要把地分成七份。 犹大 在南方，住在他的境内。 约瑟 家在北方，住在他们的境内。
JOSH|18|6|你们把地划成七份之后，就要把所写的带到我这里来。我要在耶和华－我们的上帝面前，为你们抽签。
JOSH|18|7|利未 人在你们中间没有分得地业，因为耶和华祭司的职分就是他们的产业。 迦得 支派、 吕便 支派和 玛拿西 半支派已经在 约旦河 东得了地业，是耶和华的仆人 摩西 给他们的。”
JOSH|18|8|那些去划地的人起来正要去的时候， 约书亚 吩咐他们说：“你们去走遍那地，把地划分以后，就回到我这里来。我要在 示罗 这里，在耶和华面前为你们抽签。”
JOSH|18|9|那些人就去了，走遍那地，按照城镇把地划成七份，写在册上，回到 示罗 营中 约书亚 那里。
JOSH|18|10|约书亚 就在 示罗 ，在耶和华面前为他们抽签。 约书亚 按照 以色列 人的支派，在那里把地分给他们。
JOSH|18|11|便雅悯 支派，按着宗族抽签所得之地，是在 犹大 子孙和 约瑟 子孙之间。
JOSH|18|12|他们北边的地界是从 约旦河 起，上到 耶利哥 斜坡的北边，再往西上到山区，直到 伯．亚文 的旷野。
JOSH|18|13|这地界从那里往南经过 路斯 ，直到 路斯 的斜坡， 路斯 就是 伯特利 ，又下到 亚他录．亚达 ，直到 下伯．和仑 南边的山。
JOSH|18|14|这地界往西延伸，又转向南，从 伯．和仑 南边对面的山，直通到 犹大 人的城 基列．巴力 ， 基列．巴力 就是 基列．耶琳 。这就是西边的地界。
JOSH|18|15|南边是从 基列．耶琳 的顶端为起点，这地界往西 通到 尼弗多亚 水泉，
JOSH|18|16|这地界又下到 欣嫩子谷 对面山的边缘，就是 利乏音谷 的北边；又下到 欣嫩谷 ，沿着 耶布斯 斜坡的南边，下到 隐．罗结 ；
JOSH|18|17|又往北转弯，通到 隐．示麦 ，直到 亚都冥 斜坡对面的 基利绿 ，又下到 吕便 之子 波罕 的磐石，
JOSH|18|18|又往北经过 亚拉巴 对面的斜坡 ，下到 亚拉巴 。
JOSH|18|19|这地界又经过 伯．曷拉 斜坡的北边，直通到 盐海 的北湾，就是 约旦河 的南端为止。这就是南边的地界。
JOSH|18|20|东边的地界是 约旦河 。这是 便雅悯 人按着宗族，照着他们四围的边界所得的地业。
JOSH|18|21|便雅悯 支派按着宗族所得的城镇就是： 耶利哥 、 伯．曷拉 、 伊麦．基悉 、
JOSH|18|22|伯．亚拉巴 、 洗玛脸 、 伯特利 、
JOSH|18|23|亚文 、 巴拉 、 俄弗拉 、
JOSH|18|24|基法．阿摩尼 、 俄弗尼 和 迦巴 ，共十二座城，以及所属的村庄；
JOSH|18|25|又有 基遍 、 拉玛 、 比录 、
JOSH|18|26|米斯巴 、 基非拉 、 摩撒 、
JOSH|18|27|利坚 、 伊利毗勒 、 他拉拉 、
JOSH|18|28|洗拉 、 以利弗 、 耶布斯 ， 耶布斯 就是 耶路撒冷 ， 基比亚 、 基列 ，共十四座城，以及所属的村庄。这是 便雅悯 人按着宗族所得的地业。
JOSH|19|1|第二签是 西缅 ，是 西缅 支派的人按着宗族抽出的，他们所得的地业是在 犹大 人地业的中间。
JOSH|19|2|他们所得为业之地是： 别是巴 ，或名 示巴 ， 摩拉大 、
JOSH|19|3|哈萨．书亚 、 巴拉 、 以森 、
JOSH|19|4|伊勒多腊 、 比土力 、 何珥玛 、
JOSH|19|5|洗革拉 、 伯．玛加博 、 哈萨．苏撒 、
JOSH|19|6|伯．利巴勿 、 沙鲁险 ，共十三座城，还有所属的村庄；
JOSH|19|7|又有 亚因 、 利门 、 以帖 、 亚珊 ，共四座城，还有所属的村庄；
JOSH|19|8|以及这些城镇周围一切的村庄，直到 巴拉．比珥 ，就是 尼革夫 的 拉玛 。这是 西缅 支派的人按着宗族所得的地业。
JOSH|19|9|西缅 人的地业取自 犹大 人的土地，因为 犹大 人所得的份过多，所以 西缅 人从 犹大 人的地业中取了地业。
JOSH|19|10|第三签是 西布伦 人按着宗族抽到的。他们地业的边界延伸到 撒立 。
JOSH|19|11|他们的地界往西，上到 玛拉拉 ，达到 大巴设 ，又达到 约念 前面的河。
JOSH|19|12|又从 撒立 往东转到向日出的方向，经过 吉斯绿．他泊 的边界，到 大比拉 ，又上到 雅非亚 。
JOSH|19|13|又从那里往东，经过 迦特．希弗 ，到 以特．加汛 ，通到 临门 ，延伸到 尼亚 。
JOSH|19|14|这地界在北边绕过 尼亚 ，到 哈拿顿 ，直通到 伊弗他．伊勒谷 ，
JOSH|19|15|包括 加他 、 拿哈拉 、 伸仑 、 以大拉 、 伯利恒 ，共十二座城，还有所属的村庄。
JOSH|19|16|这些城镇和所属的村庄是 西布伦 人按着宗族所得的地业。
JOSH|19|17|第四签是 以萨迦 ，是 以萨迦 人按着宗族抽出的。
JOSH|19|18|他们的地界是到 耶斯列 、 基苏律 、 书念 、
JOSH|19|19|哈弗连 、 示按 、 亚拿哈拉 、
JOSH|19|20|拉璧 、 基善 、 亚别 、
JOSH|19|21|利篾 、 隐．干宁 、 隐．哈大 、 伯．帕薛 。
JOSH|19|22|这地界达到 他泊 、 沙哈洗玛 、 伯．示麦 ，他们的地界直通到 约旦河 为止，共十六座城，还有所属的村庄。
JOSH|19|23|这些城镇和所属的村庄是 以萨迦 支派的人按着宗族所得的地业。
JOSH|19|24|第五签是 亚设 支派的人按着宗族抽出的。
JOSH|19|25|他们的地界是 黑甲 、 哈利 、 比田 、 押煞 、
JOSH|19|26|亚拉米勒 、 亚末 、 米沙勒 ，往西达到 迦密 ，又到 希曷．立纳 ，
JOSH|19|27|又转到向日出方向的 伯．大衮 ，达到 细步纶 ；又往北到 伊弗他．伊勒谷 ，到 伯．以墨 和 尼业 ，也通到 迦步勒 的左边 ，
JOSH|19|28|又到 义伯仑 、 利合 、 哈们 、 加拿 ，直到 西顿 大城。
JOSH|19|29|这地界转到 拉玛 ，直到坚固的 推罗城 。这地界又转到 何萨 ，靠近 亚革悉 一带的地方 ，直通到海为止。
JOSH|19|30|又有 乌玛 、 亚弗 、 利合 ，共二十二座城，还有所属的村庄。
JOSH|19|31|这些城镇和所属的村庄是 亚设 支派的人按着宗族所得的地业。
JOSH|19|32|第六签是 拿弗他利 人，是 拿弗他利 人按着宗族抽出的。
JOSH|19|33|他们的地界是从 希利弗 ，从 撒拿音 的橡树、 亚大米．尼吉 和 雅比聂 ，直到 拉共 ，直通到 约旦河 为止。
JOSH|19|34|这地界往西转到 亚斯纳．他泊 ，从那里通到 户割 ，南边达到 西布伦 ，西边达到 亚设 ，向日出的方向达到 约旦河 的 犹大 。
JOSH|19|35|坚固的城有 西丁 、 侧耳 、 哈末 、 拉甲 、 基尼烈 、
JOSH|19|36|亚大玛 、 拉玛 、 夏琐 、
JOSH|19|37|基低斯 、 以得来 、 隐．夏琐 、
JOSH|19|38|以利稳 、 密大．伊勒 、 和琏 、 伯．亚纳 、 伯．示麦 ，共十九座城，还有所属的村庄。
JOSH|19|39|这些城镇和所属的村庄是 拿弗他利 支派的人按着宗族所得的地业。
JOSH|19|40|但 支派，按着宗族，抽到第七签。
JOSH|19|41|他们地业的边界是 琐拉 、 以实陶 、 伊珥．示麦 、
JOSH|19|42|沙拉宾 、 亚雅仑 、 伊提拉 、
JOSH|19|43|以伦 、 亭拿 、 以革伦 、
JOSH|19|44|伊利提基 、 基比顿 、 巴拉 、
JOSH|19|45|伊胡得 、 比尼．比拉 、 迦特．临门 、
JOSH|19|46|美．耶昆 、 拉昆 ，以及 约帕 对面的地界。
JOSH|19|47|当 但 的子孙失去他们疆土的时候，就上去攻取 利善 ，用刀击杀城中的人，得了那城，住在城中，以他们祖先 但 的名字将 利善 改名为 但 。
JOSH|19|48|这些城镇和所属的村庄是 但 支派的人按着宗族所得的地业。
JOSH|19|49|以色列 人按着疆土完成了地业的分配，就在他们中间把地给 嫩 的儿子 约书亚 为业。
JOSH|19|50|他们照着耶和华的指示，把 约书亚 所要的城，就是 以法莲 山区的 亭拿．西拉 给了他。 约书亚 修建那城，住在城中。
JOSH|19|51|这就是 以利亚撒 祭司和 嫩 的儿子 约书亚 ，以及 以色列 人各支派父系的领袖，在 示罗 会幕的门口，耶和华面前抽签所分的地业。这样， 他们就完成了分地的事。
JOSH|20|1|耶和华吩咐 约书亚 说：
JOSH|20|2|“你吩咐 以色列 人说：‘你们要照我藉 摩西 所吩咐你们的，为自己设立逃城，
JOSH|20|3|使那无意中误杀人的，可以逃到那里。这些要作为你们逃避报血仇者的城。
JOSH|20|4|杀人者要逃到这些城中的一座，站在城门口，把他的事情陈诉给那城的长老听。他们就要接他入城，给他地方，让他住在他们中间。
JOSH|20|5|若是报血仇者追上了他，长老不可把他交在报血仇者的手里，因为他是无意中杀了邻舍的，并非过去彼此之间有仇恨。
JOSH|20|6|他要住在那城里，直到他站在会众面前受审判；等到当时的大祭司死后，杀人者才可以回到本城本家，就是他所逃出来的那城。’”
JOSH|20|7|于是， 以色列 人划分 拿弗他利 山区 加利利 的 基低斯 、 以法莲 山区的 示剑 和 犹大 山区的 基列．亚巴 ， 基列．亚巴 就是 希伯仑 。
JOSH|20|8|他们在 约旦河 的另一边，就是 耶利哥 的东边，从 吕便 支派中，在旷野的平原设立 比悉 ，从 迦得 支派中设立 基列 的 拉末 ，从 玛拿西 支派中设立 巴珊 的 哥兰 。
JOSH|20|9|这都是为 以色列 众人和在他们中间寄居的外人所指定的城镇，使凡误杀人者可以逃到那里，不至于死在报血仇者的手中，直到他站在会众面前受审判 。
JOSH|21|1|利未 人的众族长近前来到 以利亚撒 祭司和 嫩 的儿子 约书亚 ，以及 以色列 人各支派父系的领袖那里，
JOSH|21|2|在 迦南 地的 示罗 对他们说：“从前耶和华曾藉着 摩西 吩咐给我们城镇居住，以及城镇的郊外供我们牧养牲畜。”
JOSH|21|3|于是 以色列 人照耶和华的指示，从自己的地业中，把这些城镇和城镇的郊外给了 利未 人。
JOSH|21|4|哥辖 族抽了签。 利未 人中 亚伦 祭司的子孙，从 犹大 支派、 西缅 支派、 便雅悯 支派的地业中，抽签得了十三座城。
JOSH|21|5|哥辖 其余的子孙，从 以法莲 支派、 但 支派、 玛拿西 半支派宗族的地业中，抽签得了十座城。
JOSH|21|6|革顺 的子孙，从 以萨迦 支派、 亚设 支派、 拿弗他利 支派、住 巴珊 的 玛拿西 半支派宗族的地业中，抽签得了十三座城。
JOSH|21|7|米拉利 的子孙，按着宗族，从 吕便 支派、 迦得 支派、 西布伦 支派的地业中，得了十二座城。
JOSH|21|8|以色列 人照耶和华藉 摩西 所吩咐的，把这些城镇和城镇的郊外，抽签给 利未 人。
JOSH|21|9|他们从 犹大 支派和 西缅 支派的地业中，给了以下所记名字的各城，
JOSH|21|10|就是给 利未 人 哥辖 宗族的 亚伦 子孙，因为他们抽到第一签：
JOSH|21|11|把 犹大 山区的 基列．亚巴 ，就是 希伯仑 ，和四围的郊野给了他们。 亚巴 是 亚衲 族的祖先。
JOSH|21|12|但是，这城的田地和所属的村庄却给了 耶孚尼 的儿子 迦勒 为业。
JOSH|21|13|他们把 希伯仑 ，就是误杀人的逃城和城的郊外，给了 亚伦 祭司的子孙；又给了 立拿 和城的郊外、
JOSH|21|14|雅提珥 和城的郊外、 以实提莫 和城的郊外、
JOSH|21|15|何仑 和城的郊外、 底璧 和城的郊外、
JOSH|21|16|亚因 和城的郊外、 淤他 和城的郊外，以及 伯．示麦 和城的郊外，共九座城，都是从这二支派中分出来的。
JOSH|21|17|又从 便雅悯 支派的地业中给了 基遍 和城的郊外、 迦巴 和城的郊外、
JOSH|21|18|亚拿突 和城的郊外，以及 亚勒们 和城的郊外，共四座城。
JOSH|21|19|亚伦 子孙作祭司的共有十三座城，以及城的郊外。
JOSH|21|20|利未 人 哥辖 的宗族，就是 哥辖 其余的子孙，抽签所得的城是从 以法莲 支派来的。
JOSH|21|21|他们把 以法莲 山区的 示剑 ，就是误杀人的逃城和城的郊外给了 哥辖 其余的子孙；又给了 基色 和城的郊外、
JOSH|21|22|基伯先 和城的郊外，以及 伯．和仑 和城的郊外，共四座城。
JOSH|21|23|又从 但 支派的地业中给了 伊利提基 和城的郊外、 基比顿 和城的郊外、
JOSH|21|24|亚雅仑 和城的郊外，以及 迦特．临门 和城的郊外，共四座城。
JOSH|21|25|又从 玛拿西 半支派的地业中给了 他纳 和城的郊外，以及 迦特．临门 和城的郊外，共两座城。
JOSH|21|26|哥辖 其余的子孙共有十座城，以及城的郊外。
JOSH|21|27|利未 人宗族中 革顺 的子孙，从 玛拿西 半支派的地业中所得的是 巴珊 的 哥兰 ，就是误杀人的逃城和城的郊外，以及 比．施提拉 和城的郊外，共两座城。
JOSH|21|28|从 以萨迦 支派的地业中所得的是 基善 和城的郊外、 大比拉 和城的郊外、
JOSH|21|29|耶末 和城的郊外，以及 隐．干宁 和城的郊外，共四座城。
JOSH|21|30|从 亚设 支派的地业中所得的是 米沙勒 和城的郊外、 押顿 和城的郊外、
JOSH|21|31|黑甲 和城的郊外，以及 利合 和城的郊外，共四座城。
JOSH|21|32|从 拿弗他利 支派的地业中所得的是 加利利 的 基低斯 ，就是误杀人的逃城和城的郊外、 哈末．多珥 和城的郊外，以及 加珥坦 和城的郊外，共三座城。
JOSH|21|33|革顺 人按着宗族共有十三个城，以及城的郊外。
JOSH|21|34|其余的 利未 人，就是 米拉利 的子孙，按着宗族从 西布伦 支派的地业中所得的是 约念 和城的郊外、 加珥他 和城的郊外、
JOSH|21|35|丁拿 和城的郊外，以及 拿哈拉 和城的郊外，共四座城。
JOSH|21|36|从 吕便 支派的地业中所得的是 比悉 和城的郊外、 雅杂 和城的郊外、
JOSH|21|37|基底莫 和城的郊外，以及 米法押 和城的郊外，共四座城。
JOSH|21|38|从 迦得 支派的地业中所得的是 基列 的 拉末 ，就是误杀人的逃城和城的郊外、 玛哈念 和城的郊外、
JOSH|21|39|希实本 和城的郊外，以及 雅谢 和城的郊外，共四座城。
JOSH|21|40|利未 宗族其余的人，就是 米拉利 的子孙，按着宗族抽签所得的，共十二座城。
JOSH|21|41|利未 人在 以色列 人的地业中所得的城，共四十八个，还有城的郊外。
JOSH|21|42|这些城的四围都有郊野，每个城都是如此。
JOSH|21|43|这样，耶和华将从前向他们列祖起誓要给他们的全地赐给 以色列 人，他们就得了为业，住在其中。
JOSH|21|44|耶和华照着向他们列祖起誓所应许的一切，赐给他们全境安宁。他们所有的仇敌，没有一个能在他们面前站立得住。耶和华把所有仇敌都交在他们手中。
JOSH|21|45|耶和华应许赐福给 以色列 家的话，一句都没有落空，全都应验了。
JOSH|22|1|此后， 约书亚 召了 吕便 人、 迦得 人和 玛拿西 半支派的人来，
JOSH|22|2|对他们说：“耶和华的仆人 摩西 所吩咐你们的，你们都遵守了；我吩咐你们的话，你们也都听从了。
JOSH|22|3|你们这许多日子，都没有撇弃你们的弟兄，直到今日，并且遵守了耶和华你们上帝所吩咐的命令。
JOSH|22|4|如今耶和华－你们的上帝已经照着他所应许的，使你们的弟兄得享安宁。你们现在可以返回自己的帐棚，回到耶和华的仆人 摩西 在 约旦河 东所赐给你们为业之地。
JOSH|22|5|只是务要谨守遵行耶和华的仆人 摩西 所吩咐你们的诫命和律法，爱耶和华－你们的上帝，行他一切的道，守他的诫命，紧紧跟随他，尽心尽性事奉他。”
JOSH|22|6|于是 约书亚 为他们祝福，送他们回去，他们就回到自己的帐棚去了。
JOSH|22|7|摩西 在 巴珊 曾把地业分给 玛拿西 的半支派；然后 约书亚 在 约旦河 的西岸，在他们弟兄中，又把地业分给 玛拿西 的另外半支派。 约书亚 送他们回帐棚的时候，为他们祝福，
JOSH|22|8|对他们说：“你们要把许多财物，许多牲畜，和金、银、铜、铁，以及许多衣服，带回你们的帐棚去，要把你们从仇敌夺来的东西分给你们的众弟兄。”
JOSH|22|9|于是 吕便 人、 迦得 人、 玛拿西 半支派的人从 迦南 地的 示罗 起行，离开 以色列 人，回到他们已得为业的 基列 地，就是他们照耶和华藉 摩西 所吩咐而得的。
JOSH|22|10|吕便 人、 迦得 人和 玛拿西 半支派的人到了 迦南 地的 约旦河 一带地方，就在 约旦河 那里筑了一座坛，一座高大壮观的坛。
JOSH|22|11|以色列 人听见了，说：“看哪， 吕便 人、 迦得 人、 玛拿西 半支派的人在 迦南 地对面， 约旦河 一带地方， 以色列 人的境内，筑了一座坛。”
JOSH|22|12|以色列 人一听见，全会众的 以色列 人就聚集在 示罗 ，要上去攻打他们。
JOSH|22|13|以色列 人派 以利亚撒 祭司的儿子 非尼哈 ，往 基列 地，到 吕便 人、 迦得 人和 玛拿西 半支派的人那里。
JOSH|22|14|和他同去的还有十个领袖， 以色列 每个支派在父家中各派一个领袖，这些人每一个在 以色列 族系中都是父家的领袖。
JOSH|22|15|他们来到 基列 地，到 吕便 人、 迦得 人和 玛拿西 半支派的人那里，对他们说：
JOSH|22|16|“耶和华全会众这样说：‘你们今日离弃耶和华不跟从他，干犯 以色列 的上帝，悖逆耶和华，为自己筑了一座坛，你们所犯的是何等的罪！
JOSH|22|17|从前我们在 毗珥 犯的罪孽，导致瘟疫临到耶和华的会众，甚至到今日都还没有洗净，这还算小事吗？
JOSH|22|18|你们今日竟然离弃耶和华不跟从他！你们今日既然悖逆耶和华，明日他必向 以色列 全会众发怒。
JOSH|22|19|若你们认为所得为业之地不洁净，可以过来，到耶和华之地，就是耶和华的帐幕所居住之地，在我们中间得地业。你们却不可悖逆耶和华，也不可背叛我们，在耶和华－我们上帝的坛以外为自己筑坛。
JOSH|22|20|从前 谢拉 的曾孙 亚干 岂不是在那当灭的物上犯了罪，导致愤怒临到 以色列 全会众吗？死在他所犯的罪中的，不只是他一个人而已！’”
JOSH|22|21|于是 吕便 人、 迦得 人、 玛拿西 半支派的人回答 以色列 族系的领袖，说：
JOSH|22|22|“大能者上帝耶和华！大能者上帝耶和华！他已知道，愿 以色列 人也知道，我们若有悖逆的行为，或是干犯耶和华，你今日就不要让我们活着！
JOSH|22|23|若我们为自己筑坛，离弃耶和华不跟从他，或将燔祭、素祭、平安祭献在坛上，愿耶和华亲自追究。
JOSH|22|24|不是这样！我们做这事的原因是惧怕将来你们的子孙对我们的子孙说：‘你们与耶和华－ 以色列 的上帝有什么关系呢？
JOSH|22|25|因为耶和华以 约旦河 作我们和你们 吕便 人、 迦得 人的交界，所以你们在耶和华里无份。’这样，你们的子孙就使我们的子孙不再敬畏耶和华了。
JOSH|22|26|因此我们说：‘不如为自己筑一座坛，不是为献燔祭，也不是为献别样的祭，
JOSH|22|27|而是为你我之间和后代子孙之间作证据，好使我们也在耶和华面前献我们的燔祭、平安祭和别样的祭来事奉他，免得你们的子孙将来对我们的子孙说，你们在耶和华里无份。’
JOSH|22|28|所以我们说：‘将来他们若对我们，或对我们的子孙这样说，我们就可以回答说：你们看，我们列祖所筑的坛是耶和华坛的样式，这并不是为献燔祭，也不是为献别样的祭，而是作为你们和我们之间的证据。’
JOSH|22|29|除了耶和华－我们上帝帐幕前的坛以外，我们绝没有意思要为着献燔祭、素祭和别样的祭而另外筑一座坛，悖逆耶和华，今日离弃不跟从他。”
JOSH|22|30|非尼哈 祭司与会众中的领袖，就是与他同来那些 以色列 族系的领袖，听见 吕便 人、 迦得 人、 玛拿西 人所说的话，就都看为美。
JOSH|22|31|以利亚撒 祭司的儿子 非尼哈 对 吕便 人、 迦得 人、 玛拿西 人说：“今日我们知道耶和华在我们中间，因为你们没有向他犯悖逆的罪。现在你们把 以色列 人从耶和华的手中救出来了。”
JOSH|22|32|以利亚撒 祭司的儿子 非尼哈 与众领袖离开了 吕便 人和 迦得 人，从 基列 地回 迦南 地，到了 以色列 人那里，就把这事向他们回报。
JOSH|22|33|以色列 人看这事为美； 以色列 人就称颂上帝，不再说要上去攻打 吕便 人和 迦得 人，毁坏他们所住的地了。
JOSH|22|34|吕便 人和 迦得 人给这坛起了名，因为这坛在我们之间见证耶和华是上帝。
JOSH|23|1|耶和华使 以色列 人从四围所有的仇敌中得享安宁，已经有很多日子了。 约书亚 年纪老迈，
JOSH|23|2|就召了全 以色列 的众长老、领袖、审判官和官长来，对他们说：“我年纪已经老迈。
JOSH|23|3|耶和华－你们的上帝因你们的缘故向这些国家所做的一切，你们都亲眼看见了，那为你们作战的是耶和华－你们的上帝。
JOSH|23|4|看，我已经把所剩下的列国，连同从 约旦河 起到 大海 日落的方向，我所剪除的列国，都抽签分给你们各支派为业了。
JOSH|23|5|耶和华－你们的上帝必将他们从你们面前赶出去，使他们离开你们，你们就必得他们的地为业，正如耶和华－你们的上帝向你们所应许的。
JOSH|23|6|你们要大大壮胆，谨守遵行写在 摩西 律法书上的一切话，不可偏离左右。
JOSH|23|7|不可与你们中间所剩下的这些国家往来。你们不可提他们神明的名，不可指着它们起誓，不可事奉它们，也不可敬拜它们。
JOSH|23|8|只要紧紧跟随耶和华－你们的上帝，就像你们直到今日所做的。
JOSH|23|9|因为耶和华已经把又大又强的列国从你们面前赶出；直到今日，没有一人能在你们面前站立得住。
JOSH|23|10|你们一人必追赶千人，因为耶和华－你们的上帝照他向你们所应许的，为你们作战。
JOSH|23|11|你们要分外谨慎，爱耶和华－你们的上帝。
JOSH|23|12|你们若断然转离，紧紧跟随你们中间所剩下的这些国家，彼此结亲，互相往来，
JOSH|23|13|就要确实知道，耶和华－你们的上帝必不再将他们从你们面前赶出；他们却要成为你们的罗网、圈套、肋上的鞭、眼中的刺，直到你们在耶和华－你们上帝所赐的这美地上灭亡。
JOSH|23|14|“看哪，我今日要走世人必走的路了。你们要一心一意知道，耶和华－你们上帝所应许要赐给你们的一切福气，没有一件落空，都应验在你们身上了。
JOSH|23|15|耶和华－你们的上帝所应许的一切福气怎样临到你们身上，耶和华也必照样使各样灾祸临到你们身上，直到他把你们从耶和华－你们上帝所赐给你们的这美地上除灭。
JOSH|23|16|你们若违背耶和华－你们上帝吩咐你们所守的约，去事奉别神，敬拜它们，耶和华的怒气必向你们发作，使你们在他所赐给你们的美地上迅速灭亡。”
JOSH|24|1|约书亚 召集 以色列 的众支派到 示剑 ，他召了 以色列 的长老、领袖、审判官和官长来；他们都站在上帝面前。
JOSH|24|2|约书亚 对众百姓说：“耶和华－ 以色列 的上帝如此说：‘古时你们的列祖，就是 亚伯拉罕 和 拿鹤 的父亲 他拉 ，住在 大河 那边事奉别神。
JOSH|24|3|我将你们的祖宗 亚伯拉罕 从 大河 那边带出来，领他走遍 迦南 全地，又使他的子孙众多。我把 以撒 赐给他，
JOSH|24|4|我又把 雅各 和 以扫 赐给 以撒 ，将 西珥山 赐给 以扫 为业。但 雅各 和他的子孙下到 埃及 去了。
JOSH|24|5|我差遣 摩西 和 亚伦 ，照我在 埃及 中间所做的，降灾与 埃及 ，然后把你们领出来。
JOSH|24|6|我领你们的祖宗出 埃及 ，你们就到了 红海 。 埃及 人带领战车骑兵，追赶你们的祖宗到 红海 。
JOSH|24|7|你们的祖宗哀求耶和华，他就用黑暗把你们和 埃及 人隔开了，又使海水冲向 埃及 人，淹没他们。我在 埃及 所做的，你们都亲眼见过。你们在旷野住了很多日子。
JOSH|24|8|我领你们到 约旦河 东 亚摩利 人所住之地。他们与你们争战，我把他们交在你们手中，你们就得了他们的地为业。我也在你们面前灭绝他们。
JOSH|24|9|那时， 摩押 王 西拨 的儿子 巴勒 起来攻击 以色列 人，派人去召 比珥 的儿子 巴兰 来诅咒你们。
JOSH|24|10|但我不愿听 巴兰 ，所以他反而为你们连连祝福。这样，我救了你们脱离他的手。
JOSH|24|11|你们过了 约旦河 ，来到 耶利哥 。 耶利哥 人、 亚摩利 人、 比利洗 人、 迦南 人、 赫 人、 革迦撒 人、 希未 人、 耶布斯 人都与你们争战，我却把他们交在你们手里。
JOSH|24|12|我派遣瘟疫 在你们前面，将 亚摩利 人的两个王从你们面前赶出，并不是用你的刀，也不是用你的弓。
JOSH|24|13|我赐给你们的地，不是你们开垦的；我赐给你们的城镇，不是你们建造的。你们却住在其中，又得吃那不是你们栽植的葡萄园和橄榄园的果子。’
JOSH|24|14|“现在你们要敬畏耶和华，诚心诚意事奉他，除掉你们列祖在 大河 那边和在 埃及 事奉的神明，事奉耶和华。
JOSH|24|15|若你们认为事奉耶和华不好，今日就可以选择所要事奉的：是你们列祖在 大河 那边所事奉的神明，或是你们所住这地 亚摩利 人的神明呢？至于我和我家，我们必定事奉耶和华。”
JOSH|24|16|百姓回答说：“我们绝不离弃耶和华去事奉别神。
JOSH|24|17|因为耶和华－我们的上帝曾领我们和我们的祖宗从 埃及 地为奴之家出来，在我们眼前行了那些大神迹，并在我们所行的一切路上，和所经过的各民族中保护了我们。
JOSH|24|18|耶和华又把各民族和住此地的 亚摩利 人都从我们面前赶出去。所以，我们也必事奉耶和华，因为他是我们的上帝。”
JOSH|24|19|约书亚 对百姓说：“你们不能事奉耶和华，因为他是神圣的上帝，是忌邪 的上帝，必不赦免你们的过犯罪恶。
JOSH|24|20|你们若离弃耶和华去事奉外邦的神明，耶和华在降福之后，必转而降祸给你们，把你们灭绝。”
JOSH|24|21|百姓对 约书亚 说：“不，我们要事奉耶和华。”
JOSH|24|22|约书亚 对百姓说：“你们选择耶和华，要事奉他，你们自己作证吧！”他们说：“我们愿意作证。”
JOSH|24|23|“现在，你们要除掉你们中间外邦的神明，专心归向耶和华－ 以色列 的上帝。”
JOSH|24|24|百姓对 约书亚 说：“我们必事奉耶和华－我们的上帝，听从他的话。”
JOSH|24|25|那日， 约书亚 就与百姓立约，在 示剑 为他们制定律例典章。
JOSH|24|26|约书亚 把这些话写在上帝的律法书上，又拿一块大石头立在橡树下耶和华圣所的旁边。
JOSH|24|27|约书亚 对众百姓说：“看哪，这石头可以向我们作见证，因为它听见了耶和华所吩咐我们的一切话；这石头将向你们作见证，免得你们背叛你们的上帝。”
JOSH|24|28|于是 约书亚 解散百姓，各自回到自己的地业去了。
JOSH|24|29|这些事以后，耶和华的仆人， 嫩 的儿子 约书亚 死了，那时他一百一十岁。
JOSH|24|30|以色列 人把他葬在他自己地业的境内， 以法莲 山区的 亭拿．西拉 ，在 迦实山 的北边。
JOSH|24|31|约书亚 在世的日子和他死了以后，那些知道耶和华为 以色列 所做一切事的长老还在世的时候， 以色列 人事奉耶和华。
JOSH|24|32|以色列 人把从 埃及 所带来 约瑟 的骸骨安葬在 示剑 ，就是 雅各 从前用一百可锡塔 向 示剑 的父亲 哈抹 的众子所买的那块地；这块地就成了 约瑟 子孙的产业。
JOSH|24|33|亚伦 的儿子 以利亚撒 也死了，他们把他葬在他儿子 非尼哈 所得 以法莲 山区的小山上 。
