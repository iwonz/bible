3JOHN|1|1|Старец – возлюбленному Гаию, которого я люблю по истине.
3JOHN|1|2|Возлюбленный! молюсь, чтобы ты здравствовал и преуспевал во всем, как преуспевает душа твоя.
3JOHN|1|3|Ибо я весьма обрадовался, когда пришли братия и засвидетельствовали о твоей верности, как ты ходишь в истине.
3JOHN|1|4|Для меня нет большей радости, как слышать, что дети мои ходят в истине.
3JOHN|1|5|Возлюбленный! ты как верный поступаешь в том, что делаешь для братьев и для странников.
3JOHN|1|6|Они засвидетельствовали перед церковью о твоей любви. Ты хорошо поступишь, если отпустишь их, как должно ради Бога,
3JOHN|1|7|ибо они ради имени Его пошли, не взяв ничего от язычников.
3JOHN|1|8|Итак мы должны принимать таковых, чтобы сделаться споспешниками истине.
3JOHN|1|9|Я писал церкви; но любящий первенствовать у них Диотреф не принимает нас.
3JOHN|1|10|Посему, если я приду, то напомню о делах, которые он делает, понося нас злыми словами, и не довольствуясь тем, и сам не принимает братьев, и запрещает желающим, и изгоняет из церкви.
3JOHN|1|11|Возлюбленный! не подражай злу, но добру. Кто делает добро, тот от Бога; а делающий зло не видел Бога.
3JOHN|1|12|О Димитрии засвидетельствовано всеми и самою истиною; свидетельствуем также и мы, и вы знаете, что свидетельство наше истинно.
3JOHN|1|13|Многое имел я писать; но не хочу писать к тебе чернилами и тростью,
3JOHN|1|14|а надеюсь скоро увидеть тебя и поговорить устами к устам.
3JOHN|1|15|Мир тебе. Приветствуют тебя друзья; приветствуй друзей поименно. Аминь.
