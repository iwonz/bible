LEV|1|1|vocavit autem Mosen et locutus est ei Dominus de tabernaculo testimonii dicens
LEV|1|2|loquere filiis Israhel et dices ad eos homo qui obtulerit ex vobis hostiam Domino de pecoribus id est de bubus et ovibus offerens victimas
LEV|1|3|si holocaustum fuerit eius oblatio ac de armento masculum inmaculatum offeret ad ostium tabernaculi testimonii ad placandum sibi Dominum
LEV|1|4|ponetque manus super caput hostiae et acceptabilis erit atque in expiationem eius proficiens
LEV|1|5|immolabitque vitulum coram Domino et offerent filii Aaron sacerdotes sanguinem eius fundentes super altaris circuitum quod est ante ostium tabernaculi
LEV|1|6|detractaque pelle hostiae artus in frusta concident
LEV|1|7|et subicient in altari ignem strue lignorum ante conposita
LEV|1|8|et membra quae caesa sunt desuper ordinantes caput videlicet et cuncta quae adherent iecori
LEV|1|9|intestinis et pedibus lotis aqua adolebitque ea sacerdos super altare in holocaustum et suavem odorem Domino
LEV|1|10|quod si de pecoribus oblatio est de ovibus sive de capris holocaustum anniculum et absque macula offeret
LEV|1|11|immolabitque ad latus altaris quod respicit ad aquilonem coram Domino sanguinem vero illius fundent super altare filii Aaron per circuitum
LEV|1|12|dividentque membra caput et omnia quae adherent iecori et inponent super ligna quibus subiciendus est ignis
LEV|1|13|intestina vero et pedes lavabunt aqua et oblata omnia adolebit sacerdos super altare in holocaustum et odorem suavissimum Domino
LEV|1|14|sin autem de avibus holocausti oblatio fuerit Domino de turturibus et pullis columbae
LEV|1|15|offeret eam sacerdos ad altare et retorto ad collum capite ac rupto vulneris loco decurrere faciet sanguinem super crepidinem altaris
LEV|1|16|vesiculam vero gutturis et plumas proiciet propter altare ad orientalem plagam in loco in quo cineres effundi solent
LEV|1|17|confringetque ascellas eius et non secabit nec ferro dividet eam et adolebit super altare lignis igne subposito holocaustum est et oblatio suavissimi odoris Domino
LEV|2|1|anima cum obtulerit oblationem sacrificii Domino simila erit eius oblatio fundetque super eam oleum et ponet tus
LEV|2|2|ac deferet ad filios Aaron sacerdotes quorum unus tollet pugillum plenum similae et olei ac totum tus et ponet memoriale super altare in odorem suavissimum Domino
LEV|2|3|quod autem reliquum fuerit de sacrificio erit Aaron et filiorum eius sanctum sanctorum de oblationibus Domini
LEV|2|4|cum autem obtuleris sacrificium coctum in clibano de simila panes scilicet absque fermento conspersos oleo et lagana azyma oleo lita
LEV|2|5|si oblatio tua fuerit de sartagine similae conspersae oleo et absque fermento
LEV|2|6|divides eam minutatim et fundes supra oleum
LEV|2|7|sin autem de craticula sacrificium aeque simila oleo conspergetur
LEV|2|8|quam offeres Domino tradens manibus sacerdotis
LEV|2|9|qui cum obtulerit eam tollet memoriale de sacrificio et adolebit super altare in odorem suavitatis Domino
LEV|2|10|quicquid autem reliquum est erit Aaron et filiorum eius sanctum sanctorum de oblationibus Domini
LEV|2|11|omnis oblatio quae offertur Domino absque fermento fiet nec quicquam fermenti ac mellis adolebitur in sacrificio Domini
LEV|2|12|primitias tantum eorum offeretis et munera super altare vero non ponentur in odorem suavitatis
LEV|2|13|quicquid obtuleris sacrificii sale condies nec auferes sal foederis Dei tui de sacrificio tuo in omni oblatione offeres sal
LEV|2|14|sin autem obtuleris munus primarum frugum tuarum Domino de spicis adhuc virentibus torres eas igni et confringes in morem farris et sic offeres primitias tuas Domino
LEV|2|15|fundens supra oleum et tus inponens quia oblatio Domini est
LEV|2|16|de qua adolebit sacerdos in memoriam muneris partem farris fracti et olei ac totum tus
LEV|3|1|quod si hostia pacificorum fuerit eius oblatio et de bubus voluerit offerre marem sive feminam inmaculata offeret coram Domino
LEV|3|2|ponetque manum super caput victimae suae quae immolabitur in introitu tabernaculi fundentque filii Aaron sacerdotes sanguinem per circuitum altaris
LEV|3|3|et offerent de hostia pacificorum in oblationem Domini adipem qui operit vitalia et quicquid pinguedinis intrinsecus est
LEV|3|4|duos renes cum adipe quo teguntur ilia et reticulum iecoris cum renunculis
LEV|3|5|adolebuntque ea super altare in holocaustum lignis igne subposito in oblationem suavissimi odoris Domino
LEV|3|6|si vero de ovibus fuerit eius oblatio et pacificorum hostia sive masculum sive feminam obtulerit inmaculata erunt
LEV|3|7|si agnum obtulerit coram Domino
LEV|3|8|ponet manum super caput victimae suae quae immolabitur in vestibulo tabernaculi testimonii fundentque filii Aaron sanguinem eius per altaris circuitum
LEV|3|9|et offerent de pacificorum hostia sacrificium Domino adipem et caudam totam
LEV|3|10|cum renibus et pinguedinem quae operit ventrem atque universa vitalia et utrumque renunculum cum adipe qui est iuxta ilia reticulumque iecoris cum renunculis
LEV|3|11|et adolebit ea sacerdos super altare in pabulum ignis et oblationis Domini
LEV|3|12|si capra fuerit eius oblatio et obtulerit eam Domino
LEV|3|13|ponet manum suam super caput eius immolabitque eam in introitu tabernaculi testimonii et fundent filii Aaron sanguinem eius per altaris circuitum
LEV|3|14|tollentque ex ea in pastum ignis dominici adipem qui operit ventrem et qui tegit universa vitalia
LEV|3|15|duos renunculos cum reticulo qui est super eos iuxta ilia et arvinam iecoris cum renunculis
LEV|3|16|adolebitque ea sacerdos super altare in alimoniam ignis et suavissimi odoris omnis adeps Domini erit
LEV|3|17|iure perpetuo in generationibus et cunctis habitaculis vestris nec adipes nec sanguinem omnino comedetis
LEV|4|1|locutusque est Dominus ad Mosen dicens
LEV|4|2|loquere filiis Israhel anima cum peccaverit per ignorantiam et de universis mandatis Domini quae praecepit ut non fierent quippiam fecerit
LEV|4|3|si sacerdos qui est unctus peccaverit delinquere faciens populum offeret pro peccato suo vitulum inmaculatum Domino
LEV|4|4|et adducet illum ad ostium tabernaculi testimonii coram Domino ponetque manum super caput eius et immolabit eum Domino
LEV|4|5|hauriet quoque de sanguine vituli inferens illud in tabernaculum testimonii
LEV|4|6|cumque intinxerit digitum in sanguinem asperget eo septies coram Domino contra velum sanctuarii
LEV|4|7|ponetque de eodem sanguine super cornua altaris thymiamatis gratissimi Domino quod est in tabernaculo testimonii omnem autem reliquum sanguinem fundet in basim altaris holocausti in introitu tabernaculi
LEV|4|8|et adipem vituli auferet pro peccato tam eum qui operit vitalia quam omnia quae intrinsecus sunt
LEV|4|9|duos renunculos et reticulum quod est super eos iuxta ilia et adipem iecoris cum renunculis
LEV|4|10|sicut aufertur de vitulo hostiae pacificorum et adolebit ea super altare holocausti
LEV|4|11|pellem vero et omnes carnes cum capite et pedibus et intestinis et fimo
LEV|4|12|et reliquo corpore efferet extra castra in locum mundum ubi cineres effundi solent incendetque ea super lignorum struem quae in loco effusorum cinerum cremabuntur
LEV|4|13|quod si omnis turba Israhel ignoraverit et per inperitiam fecerit quod contra mandatum Domini est
LEV|4|14|et postea intellexerit peccatum suum offeret vitulum pro peccato adducetque eum ad ostium tabernaculi
LEV|4|15|et ponent seniores populi manus super caput eius coram Domino immolatoque vitulo in conspectu Domini
LEV|4|16|inferet sacerdos qui unctus est de sanguine eius in tabernaculum testimonii
LEV|4|17|tincto digito aspergens septies contra velum
LEV|4|18|ponetque de eodem sanguine in cornibus altaris quod est coram Domino in tabernaculo testimonii reliquum autem sanguinem fundet iuxta basim altaris holocaustorum quod est in ostio tabernaculi testimonii
LEV|4|19|omnemque eius adipem tollet et adolebit super altare
LEV|4|20|sic faciens et de hoc vitulo quomodo fecit et prius et rogante pro eis sacerdote propitius erit Dominus
LEV|4|21|ipsum autem vitulum efferet extra castra atque conburet sicut et priorem vitulum quia pro peccato est multitudinis
LEV|4|22|si peccaverit princeps et fecerit unum e pluribus per ignorantiam quod Domini lege prohibetur
LEV|4|23|et postea intellexerit peccatum suum offeret hostiam Domino hircum de capris inmaculatum
LEV|4|24|ponetque manum suam super caput eius cumque immolaverit eum in loco ubi solet mactari holocaustum coram Domino quia pro peccato est
LEV|4|25|tinguet sacerdos digitum in sanguine hostiae pro peccato tangens cornua altaris holocausti et reliquum fundens ad basim eius
LEV|4|26|adipem vero adolebit supra sicut in victimis pacificorum fieri solet rogabitque pro eo et pro peccato eius ac dimittetur ei
LEV|4|27|quod si peccaverit anima per ignorantiam de populo terrae ut faciat quicquam ex his quae Domini lege prohibentur atque delinquat
LEV|4|28|et cognoverit peccatum suum offeret capram inmaculatam
LEV|4|29|ponetque manum super caput hostiae quae pro peccato est et immolabit eam in loco holocausti
LEV|4|30|tolletque sacerdos de sanguine in digito suo et tangens cornua altaris holocausti reliquum fundet ad basim eius
LEV|4|31|omnem autem auferens adipem sicut auferri solet de victimis pacificorum adolebit super altare in odorem suavitatis Domino rogabitque pro eo et dimittetur ei
LEV|4|32|sin autem de pecoribus obtulerit victimam pro peccato ovem scilicet inmaculatam
LEV|4|33|ponet manum super caput eius et immolabit eam in loco ubi solent holocaustorum caedi hostiae
LEV|4|34|sumetque sacerdos de sanguine eius digito suo et tangens cornua altaris holocausti reliquum fundet ad basim eius
LEV|4|35|omnem quoque auferens adipem sicut auferri solet adeps arietis qui immolatur pro pacificis et cremabit super altare in incensum Domini rogabitque pro eo et pro peccato eius et dimittetur illi
LEV|5|1|si peccaverit anima et audierit vocem iurantis testisque fuerit quod aut ipse vidit aut conscius est nisi indicaverit portabit iniquitatem suam
LEV|5|2|anima quae tetigerit aliquid inmundum sive quod occisum a bestia est aut per se mortuum vel quodlibet aliud reptile et oblita fuerit inmunditiae suae rea est et deliquit
LEV|5|3|et si tetigerit quicquam de inmunditia hominis iuxta omnem inpuritatem qua pollui solet oblitaque cognoverit postea subiacebit delicto
LEV|5|4|anima quae iuraverit et protulerit labiis suis ut vel male quid faceret vel bene et id ipsum iuramento et sermone firmaverit oblitaque postea intellexerit delictum suum
LEV|5|5|agat paenitentiam pro peccato
LEV|5|6|et offerat agnam de gregibus sive capram orabitque pro eo sacerdos et pro peccato eius
LEV|5|7|sin autem non potuerit offerre pecus offerat duos turtures vel duos pullos columbarum Domino unum pro peccato et alterum in holocaustum
LEV|5|8|dabitque eos sacerdoti qui primum offerens pro peccato retorquebit caput eius ad pinnulas ita ut collo hereat et non penitus abrumpatur
LEV|5|9|et asperget de sanguine eius parietem altaris quicquid autem reliquum fuerit faciet destillare ad fundamentum eius quia pro peccato est
LEV|5|10|alterum vero adolebit holocaustum ut fieri solet rogabitque pro eo sacerdos et pro peccato eius et dimittetur ei
LEV|5|11|quod si non quiverit manus eius offerre duos turtures vel duos pullos columbae offeret pro peccato similam partem oephi decimam non mittet in eam oleum nec turis aliquid inponet quia pro peccato est
LEV|5|12|tradetque eam sacerdoti qui plenum ex toto pugillum hauriens cremabit super altare in monumentum eius qui obtulit
LEV|5|13|rogans pro illo et expians reliquam vero partem ipse habebit in munere
LEV|5|14|locutus est Dominus ad Mosen dicens
LEV|5|15|anima si praevaricans caerimonias per errorem in his quae Domino sunt sanctificata peccaverit offeret pro delicto suo arietem inmaculatum de gregibus qui emi potest duobus siclis iuxta pondus sanctuarii
LEV|5|16|ipsumque quod intulit damni restituet et quintam partem ponet supra tradens sacerdoti qui rogabit pro eo offerens arietem et dimittetur ei
LEV|5|17|anima si peccaverit per ignorantiam feceritque unum ex his quae Domini lege prohibentur et peccati rea intellexerit iniquitatem suam
LEV|5|18|offeret arietem inmaculatum de gregibus sacerdoti iuxta mensuram aestimationemque peccati qui orabit pro eo quod nesciens fecerit et dimittetur ei
LEV|5|19|quia per errorem deliquit in Dominum
LEV|6|1|locutus est Dominus ad Mosen dicens
LEV|6|2|anima quae peccaverit et contempto Domino negaverit depositum proximo suo quod fidei eius creditum fuerat vel vi aliquid extorserit aut calumniam fecerit
LEV|6|3|sive rem perditam invenerit et infitians insuper peierarit et quodlibet aliud ex pluribus fecerit in quibus peccare solent homines
LEV|6|4|convicta delicti reddet
LEV|6|5|omnia quae per fraudem voluit obtinere integra et quintam insuper partem domino cui damnum intulerat
LEV|6|6|pro peccato autem suo offeret arietem inmaculatum de grege et dabit eum sacerdoti iuxta aestimationem mensuramque delicti
LEV|6|7|qui rogabit pro eo coram Domino et dimittetur illi pro singulis quae faciendo peccaverit
LEV|6|8|locutus est Dominus ad Mosen dicens
LEV|6|9|praecipe Aaron et filiis eius haec est lex holocausti cremabitur in altari tota nocte usque mane ignis ex eodem altari erit
LEV|6|10|vestietur sacerdos tunica et feminalibus lineis tolletque cineres quos vorans ignis exusit et ponens iuxta altare
LEV|6|11|spoliabitur prioribus vestimentis indutusque aliis efferet eos extra castra et in loco mundissimo usque ad favillam consumi faciet
LEV|6|12|ignis autem in altari semper ardebit quem nutriet sacerdos subiciens ligna mane per singulos dies et inposito holocausto desuper adolebit adipes pacificorum
LEV|6|13|ignis est iste perpetuus qui numquam deficiet in altari
LEV|6|14|haec est lex sacrificii et libamentorum quae offerent filii Aaron coram Domino et coram altari
LEV|6|15|tollet sacerdos pugillum similae quae conspersa est oleo et totum tus quod super similam positum est adolebitque illud in altari in monumentum odoris suavissimi Domino
LEV|6|16|reliquam autem partem similae comedet Aaron cum filiis suis absque fermento et comedet in loco sancto atrii tabernaculi
LEV|6|17|ideo autem non fermentabitur quia pars eius in Domini offertur incensum sanctum sanctorum erit sicut pro peccato atque delicto
LEV|6|18|mares tantum stirpis Aaron comedent illud legitimum ac sempiternum est in generationibus vestris de sacrificiis Domini omnis qui tetigerit illa sanctificabitur
LEV|6|19|et locutus est Dominus ad Mosen dicens
LEV|6|20|haec est oblatio Aaron et filiorum eius quam offerre debent Domino in die unctionis suae decimam partem oephi offerent similae in sacrificio sempiterno medium eius mane et medium vespere
LEV|6|21|quae in sartagine oleo conspersa frigetur offeret autem eam calidam in odorem suavissimum Domino
LEV|6|22|sacerdos qui patri iure successerit et tota cremabitur in altari
LEV|6|23|omne enim sacrificium sacerdotum igne consumetur nec quisquam comedet ex eo
LEV|6|24|locutus est Dominus ad Mosen dicens
LEV|6|25|loquere Aaron et filiis eius ista est lex hostiae pro peccato in loco ubi offertur holocaustum immolabitur coram Domino sanctum sanctorum est
LEV|6|26|sacerdos qui offert comedet eam in loco sancto in atrio tabernaculi
LEV|6|27|quicquid tetigerit carnes eius sanctificabitur si de sanguine illius vestis fuerit aspersa lavabitur in loco sancto
LEV|6|28|vas autem fictile in quo cocta est confringetur quod si vas aeneum fuerit defricabitur et lavabitur aqua
LEV|6|29|omnis masculus de genere sacerdotali vescetur carnibus eius quia sanctum sanctorum est
LEV|6|30|hostia enim quae caeditur pro peccato cuius sanguis infertur in tabernaculum testimonii ad expiandum in sanctuario non comedetur sed conburetur igni
LEV|7|1|haec quoque est lex hostiae pro delicto sancta sanctorum est
LEV|7|2|idcirco ubi immolatur holocaustum mactabitur et victima pro delicto sanguis eius per gyrum fundetur altaris
LEV|7|3|offerent ex ea caudam et adipem qui operit vitalia
LEV|7|4|duos renunculos et pinguedinem quae iuxta ilia est reticulumque iecoris cum renunculis
LEV|7|5|et adolebit ea sacerdos super altare incensum est Domini pro delicto
LEV|7|6|omnis masculus de sacerdotali genere in loco sancto vescetur his carnibus quia sanctum sanctorum est
LEV|7|7|sicut pro peccato offertur hostia ita et pro delicto utriusque hostiae lex una erit ad sacerdotem qui eam obtulerit pertinebit
LEV|7|8|sacerdos qui offert holocausti victimam habebit pellem eius
LEV|7|9|et omne sacrificium similae quod coquitur in clibano et quicquid in craticula vel in sartagine praeparatur eius erit sacerdotis a quo offertur
LEV|7|10|sive oleo conspersa sive arida fuerit cunctis filiis Aaron aequa mensura per singulos dividetur
LEV|7|11|haec est lex hostiae pacificorum quae offertur Domino
LEV|7|12|si pro gratiarum actione fuerit oblatio offerent panes absque fermento conspersos oleo et lagana azyma uncta oleo coctamque similam et collyridas olei admixtione conspersas
LEV|7|13|panes quoque fermentatos cum hostia gratiarum quae immolatur pro pacificis
LEV|7|14|ex quibus unus pro primitiis offeretur Domino et erit sacerdotis qui fundet hostiae sanguinem
LEV|7|15|cuius carnes eadem comedentur die nec remanebit ex eis quicquam usque mane
LEV|7|16|si voto vel sponte quisquam obtulerit hostiam eadem similiter edetur die sed et si quid in crastinum remanserit vesci licitum est
LEV|7|17|quicquid autem tertius invenerit dies ignis absumet
LEV|7|18|si quis de carnibus victimae pacificorum die tertio comederit irrita fiet oblatio nec proderit offerenti quin potius quaecumque anima tali se edulio contaminarit praevaricationis rea erit
LEV|7|19|caro quae aliquid tetigerit inmundum non comedetur sed conburetur igni qui fuerit mundus vescetur ea
LEV|7|20|anima polluta quae ederit de carnibus hostiae pacificorum quae oblata est Domino peribit de populis suis
LEV|7|21|et quae tetigerit inmunditiam hominis vel iumenti sive omnis rei quae polluere potest et comederit de huiuscemodi carnibus interibit de populis suis
LEV|7|22|locutusque est Dominus ad Mosen dicens
LEV|7|23|loquere filiis Israhel adipem bovis et ovis et caprae non comedetis
LEV|7|24|adipem cadaveris morticini et eius animalis quod a bestia captum est habebitis in usus varios
LEV|7|25|si quis adipem qui offerri debet in incensum Domini comederit peribit de populo suo
LEV|7|26|sanguinem quoque omnis animalis non sumetis in cibo tam de avibus quam de pecoribus
LEV|7|27|omnis anima quae ederit sanguinem peribit de populis suis
LEV|7|28|locutus est Dominus ad Mosen dicens
LEV|7|29|loquere filiis Israhel qui offert victimam pacificorum Domino offerat simul et sacrificium id est libamenta eius
LEV|7|30|tenebit manibus adipem hostiae et pectusculum cumque ambo oblata Domino consecrarit tradet sacerdoti
LEV|7|31|qui adolebit adipem super altare pectusculum autem erit Aaron et filiorum eius
LEV|7|32|armus quoque dexter de pacificorum hostiis cedet in primitias sacerdotis
LEV|7|33|qui obtulerit sanguinem et adipem filiorum Aaron ipse habebit et armum dextrum in portione sua
LEV|7|34|pectusculum enim elationis et armum separationis tuli a filiis Israhel de hostiis eorum pacificis et dedi Aaron sacerdoti ac filiis eius lege perpetua ab omni populo Israhel
LEV|7|35|haec est unctio Aaron et filiorum eius in caerimoniis Domini die qua obtulit eos Moses ut sacerdotio fungerentur
LEV|7|36|et quae praecepit dari eis Dominus a filiis Israhel religione perpetua in generationibus suis
LEV|7|37|ista est lex holocausti et sacrificii pro peccato atque delicto et pro consecratione et pacificorum victimis
LEV|7|38|quas constituit Dominus Mosi in monte Sinai quando mandavit filiis Israhel ut offerrent oblationes suas Domino in deserto Sinai
LEV|8|1|locutusque est Dominus ad Mosen dicens
LEV|8|2|tolle Aaron cum filiis suis vestes eorum et unctionis oleum vitulum pro peccato duos arietes canistrum cum azymis
LEV|8|3|et congregabis omnem coetum ad ostium tabernaculi
LEV|8|4|fecit Moses ut Dominus imperarat congregataque omni turba ante fores
LEV|8|5|ait iste est sermo quem iussit Dominus fieri
LEV|8|6|statimque obtulit Aaron et filios eius cumque lavisset eos
LEV|8|7|vestivit pontificem subucula linea accingens eum balteo et induens tunica hyacinthina et desuper umerale inposuit
LEV|8|8|quod adstringens cingulo aptavit rationali in quo erat doctrina et veritas
LEV|8|9|cidarim quoque texit caput et super eam contra frontem posuit lamminam auream consecratam in sanctificationem sicut praeceperat ei Dominus
LEV|8|10|tulit et unctionis oleum quo levit tabernaculum cum omni supellectili sua
LEV|8|11|cumque sanctificans aspersisset altare septem vicibus unxit illud et omnia vasa eius labrumque cum basi sua sanctificavit oleo
LEV|8|12|quod fundens super caput Aaron unxit eum et consecravit
LEV|8|13|filios quoque eius oblatos vestivit tunicis lineis et cinxit balteo inposuitque mitras ut iusserat Dominus
LEV|8|14|obtulit et vitulum pro peccato cumque super caput eius posuissent Aaron et filii eius manus suas
LEV|8|15|immolavit eum hauriens sanguinem et tincto digito tetigit cornua altaris per gyrum quo expiato et sanctificato fudit reliquum sanguinem ad fundamenta eius
LEV|8|16|adipem autem qui erat super vitalia et reticulum iecoris duosque renunculos cum arvinulis suis adolevit super altare
LEV|8|17|vitulum cum pelle carnibus et fimo cremans extra castra sicut praeceperat Dominus
LEV|8|18|obtulit et arietem in holocaustum super cuius caput cum inposuissent Aaron et filii eius manus suas
LEV|8|19|immolavit eum et fudit sanguinem eius per altaris circuitum
LEV|8|20|ipsumque arietem in frusta concidens caput eius et artus et adipem adolevit igni
LEV|8|21|lotis prius intestinis et pedibus totumque simul arietem incendit super altare eo quod esset holocaustum suavissimi odoris Domino sicut praeceperat ei
LEV|8|22|obtulit et arietem secundum in consecrationem sacerdotum posueruntque super caput illius Aaron et filii eius manus suas
LEV|8|23|quem cum immolasset Moses sumens de sanguine tetigit extremum auriculae dextrae Aaron et pollicem manus eius dextrae similiter et pedis
LEV|8|24|obtulit et filios Aaron cumque de sanguine arietis immolati tetigisset extremum auriculae singulorum dextrae et pollices manus ac pedis dextri reliquum fudit super altare per circuitum
LEV|8|25|adipem vero et caudam omnemque pinguedinem quae operit intestina reticulumque iecoris et duos renes cum adipibus suis et armo dextro separavit
LEV|8|26|tollens autem de canistro azymorum quod erat coram Domino panem absque fermento et collyridam conspersam oleo laganumque posuit super adipes et armum dextrum
LEV|8|27|tradens simul omnia Aaron et filiis eius qui postquam levaverunt ea coram Domino
LEV|8|28|rursum suscepta de manibus eorum adolevit super altare holocausti eo quod consecrationis esset oblatio in odorem suavitatis sacrificii Domini
LEV|8|29|tulit et pectusculum elevans illud coram Domino de ariete consecrationis in partem suam sicut praeceperat ei Dominus
LEV|8|30|adsumensque unguentum et sanguinem qui erat in altari aspersit super Aaron et vestimenta eius et super filios illius ac vestes eorum
LEV|8|31|cumque sanctificasset eos in vestitu suo praecepit eis dicens coquite carnes ante fores tabernaculi et ibi comedite eas panes quoque consecrationis edite qui positi sunt in canistro sicut praecepit mihi dicens Aaron et filii eius comedent eos
LEV|8|32|quicquid autem reliquum fuerit de carne et panibus ignis absumet
LEV|8|33|de ostio quoque tabernaculi non exibitis septem diebus usque ad diem quo conplebitur tempus consecrationis vestrae septem enim diebus finitur consecratio
LEV|8|34|sicut et inpraesentiarum factum est ut ritus sacrificii conpleretur
LEV|8|35|die ac nocte manebitis in tabernaculo observantes custodias Domini ne moriamini sic enim mihi praeceptum est
LEV|8|36|feceruntque Aaron et filii eius cuncta quae locutus est Dominus per manum Mosi
LEV|9|1|facto autem octavo die vocavit Moses Aaron et filios eius ac maiores natu Israhel dixitque ad Aaron
LEV|9|2|tolle de armento vitulum pro peccato et arietem in holocaustum utrumque inmaculatos et offer illos coram Domino
LEV|9|3|et ad filios Israhel loqueris tollite hircum pro peccato et vitulum atque agnum anniculos et sine macula in holocaustum
LEV|9|4|bovem et arietem pro pacificis et immolate eos coram Domino in sacrificio singulorum similam oleo conspersam offerentes hodie enim Dominus apparebit vobis
LEV|9|5|tulerunt ergo cuncta quae iusserat Moses ad ostium tabernaculi ubi cum omnis staret multitudo
LEV|9|6|ait Moses iste est sermo quem praecepit Dominus facite et apparebit vobis gloria eius
LEV|9|7|dixit et ad Aaron accede ad altare et immola pro peccato tuo offer holocaustum et deprecare pro te et pro populo cumque mactaveris hostiam populi ora pro eo sicut praecepit Dominus
LEV|9|8|statimque Aaron accedens ad altare immolavit vitulum pro peccato suo
LEV|9|9|cuius sanguinem obtulerunt ei filii sui in quo tinguens digitum tetigit cornua altaris et fudit residuum ad basim eius
LEV|9|10|adipemque et renunculos ac reticulum iecoris quae sunt pro peccato adolevit super altare sicut praeceperat Dominus Mosi
LEV|9|11|carnes vero et pellem eius extra castra conbusit igni
LEV|9|12|immolavit et holocausti victimam obtuleruntque ei filii sui sanguinem eius quem fudit per altaris circuitum
LEV|9|13|ipsam etiam hostiam in frusta concisam cum capite et membris singulis obtulerunt quae omnia super altare cremavit igni
LEV|9|14|lotis prius aqua intestinis et pedibus
LEV|9|15|et pro peccato populi offerens mactavit hircum expiatoque altari
LEV|9|16|fecit holocaustum
LEV|9|17|addens in sacrificio libamenta quae pariter offeruntur et adolens ea super altare absque caerimoniis holocausti matutini
LEV|9|18|immolavit et bovem atque arietem hostias pacificas populi obtuleruntque ei filii sui sanguinem quem fudit super altare in circuitu
LEV|9|19|adipes autem bovis et caudam arietis renunculosque cum adipibus suis et reticulum iecoris
LEV|9|20|posuerunt super pectora cumque cremati essent adipes in altari
LEV|9|21|pectora eorum et armos dextros separavit Aaron elevans coram Domino sicut praeceperat Moses
LEV|9|22|et tendens manum contra populum benedixit eis sicque conpletis hostiis pro peccato et holocaustis et pacificis descendit
LEV|9|23|ingressi autem Moses et Aaron tabernaculum testimonii et deinceps egressi benedixerunt populo apparuitque gloria Domini omni multitudini
LEV|9|24|et ecce egressus ignis a Domino devoravit holocaustum et adipes qui erant super altare quod cum vidissent turbae laudaverunt Dominum ruentes in facies suas
LEV|10|1|arreptisque Nadab et Abiu filii Aaron turibulis posuerunt ignem et incensum desuper offerentes coram Domino ignem alienum quod eis praeceptum non erat
LEV|10|2|egressusque ignis a Domino devoravit eos et mortui sunt coram Domino
LEV|10|3|dixitque Moses ad Aaron hoc est quod locutus est Dominus sanctificabor in his qui adpropinquant mihi et in conspectu omnis populi glorificabor quod audiens tacuit Aaron
LEV|10|4|vocatis autem Moses Misahel et Elsaphan filios Ozihel patrui Aaron ait ad eos ite et colligite fratres vestros de conspectu sanctuarii et asportate extra castra
LEV|10|5|confestimque pergentes tulerunt eos sicut iacebant vestitos lineis tunicis et eiecerunt foras ut sibi fuerat imperatum
LEV|10|6|locutus est Moses ad Aaron et ad Eleazar atque Ithamar filios eius capita vestra nolite nudare et vestimenta nolite scindere ne forte moriamini et super omnem coetum oriatur indignatio fratres vestri et omnis domus Israhel plangant incendium quod Dominus suscitavit
LEV|10|7|vos autem non egredimini fores tabernaculi alioquin peribitis oleum quippe sanctae unctionis est super vos qui fecerunt omnia iuxta praeceptum Mosi
LEV|10|8|dixit quoque Dominus ad Aaron
LEV|10|9|vinum et omne quod inebriare potest non bibetis tu et filii tui quando intratis tabernaculum testimonii ne moriamini quia praeceptum est sempiternum in generationes vestras
LEV|10|10|et ut habeatis scientiam discernendi inter sanctum et profanum inter pollutum et mundum
LEV|10|11|doceatisque filios Israhel omnia legitima mea quae locutus est Dominus ad eos per manum Mosi
LEV|10|12|locutusque est Moses ad Aaron et ad Eleazar atque Ithamar filios eius qui residui erant tollite sacrificium quod remansit de oblatione Domini et comedite illud absque fermento iuxta altare quia sanctum sanctorum est
LEV|10|13|comedetis autem in loco sancto quod datum est tibi et filiis tuis de oblationibus Domini sicut praeceptum est mihi
LEV|10|14|pectusculum quoque quod oblatum est et armum qui separatus est edetis in loco mundissimo tu et filii tui ac filiae tuae tecum tibi enim ac liberis tuis reposita sunt de hostiis salutaribus filiorum Israhel
LEV|10|15|eo quod armum et pectus et adipes qui cremantur in altari elevaverint coram Domino et pertineant ad te et ad filios tuos lege perpetua sicut praecepit Dominus
LEV|10|16|inter haec hircum qui oblatus fuerat pro peccato cum quaereret Moses exustum repperit iratusque contra Eleazar et Ithamar filios Aaron qui remanserant ait
LEV|10|17|cur non comedistis hostiam pro peccato in loco sancto quae sancta sanctorum est et data vobis ut portetis iniquitatem multitudinis et rogetis pro ea in conspectu Domini
LEV|10|18|praesertim cum de sanguine illius non sit inlatum intra sancta et comedere eam debueritis in sanctuario sicut praeceptum est mihi
LEV|10|19|respondit Aaron oblata est hodie victima pro peccato et holocaustum coram Domino mihi autem accidit quod vides quomodo potui comedere eam aut placere Domino in caerimoniis mente lugubri
LEV|10|20|quod cum audisset Moses recepit satisfactionem
LEV|11|1|locutus est Dominus ad Mosen et Aaron dicens
LEV|11|2|dicite filiis Israhel haec sunt animalia quae comedere debetis de cunctis animantibus terrae
LEV|11|3|omne quod habet divisam ungulam et ruminat in pecoribus comedetis
LEV|11|4|quicquid autem ruminat quidem et habet ungulam sed non dividit eam sicut camelus et cetera non comedetis illud et inter inmunda reputabitis
LEV|11|5|chyrogryllius qui ruminat ungulamque non dividit inmundus est
LEV|11|6|lepus quoque nam et ipse ruminat sed ungulam non dividit
LEV|11|7|et sus qui cum ungulam dividat non ruminat
LEV|11|8|horum carnibus non vescemini nec cadavera contingetis quia inmunda sunt vobis
LEV|11|9|haec sunt quae gignuntur in aquis et vesci licitum est omne quod habet pinnulas et squamas tam in mari quam in fluminibus et stagnis comedetis
LEV|11|10|quicquid autem pinnulas et squamas non habet eorum quae in aquis moventur et vivunt abominabile vobis
LEV|11|11|et execrandum erit carnes eorum non comedetis et morticina vitabitis
LEV|11|12|cuncta quae non habent pinnulas et squamas in aquis polluta erunt
LEV|11|13|haec sunt quae de avibus comedere non debetis et vitanda sunt vobis aquilam et grypem et alietum
LEV|11|14|milvum ac vulturem iuxta genus suum
LEV|11|15|et omne corvini generis in similitudinem suam
LEV|11|16|strutionem et noctuam et larum et accipitrem iuxta genus suum
LEV|11|17|bubonem et mergulum et ibin
LEV|11|18|cycnum et onocrotalum et porphirionem
LEV|11|19|erodionem et charadrion iuxta genus suum opupam quoque et vespertilionem
LEV|11|20|omne de volucribus quod graditur super quattuor pedes abominabile erit vobis
LEV|11|21|quicquid autem ambulat quidem super quattuor pedes sed habet longiora retro crura per quae salit super terram
LEV|11|22|comedere debetis ut est brucus in genere suo et attacus atque ophiomachus ac lucusta singula iuxta genus suum
LEV|11|23|quicquid autem ex volucribus quattuor tantum habet pedes execrabile erit vobis
LEV|11|24|et quicumque morticina eorum tetigerit polluetur et erit inmundus usque ad vesperum
LEV|11|25|et si necesse fuerit ut portet quippiam horum mortuum lavabit vestimenta sua et inmundus erit usque ad solis occasum
LEV|11|26|omne animal quod habet quidem ungulam sed non dividit eam nec ruminat inmundum erit et quicquid tetigerit illud contaminabitur
LEV|11|27|quod ambulat super manus ex cunctis animantibus quae incedunt quadrupedia inmundum erit qui tetigerit morticina eorum polluetur usque ad vesperum
LEV|11|28|et qui portaverit huiuscemodi cadavera lavabit vestimenta sua et inmundus erit usque ad vesperum quia omnia haec inmunda sunt vobis
LEV|11|29|hoc quoque inter polluta reputabitur de his quae moventur in terra mustela et mus et corcodillus singula iuxta genus suum
LEV|11|30|migale et cameleon et stelio ac lacerta et talpa
LEV|11|31|omnia haec inmunda sunt qui tetigerit morticina eorum inmundus erit usque ad vesperum
LEV|11|32|et super quod ceciderit quicquam de morticinis eorum polluetur tam vas ligneum et vestimentum quam pelles et cilicia et in quocumque fit opus tinguentur aqua et polluta erunt usque ad vesperum et sic postea mundabuntur
LEV|11|33|vas autem fictile in quo horum quicquam intro ceciderit polluetur et idcirco frangendum est
LEV|11|34|omnis cibus quem comeditis si fusa fuerit super eum aqua inmundus erit et omne liquens quod bibitur de universo vase inmundum erit
LEV|11|35|et quicquid de morticinis istiusmodi ceciderit super illud inmundum erit sive clibani sive cytropodes destruentur et inmundi erunt
LEV|11|36|fontes vero et cisternae et omnis aquarum congregatio munda erit qui morticinum eorum tetigerit polluetur
LEV|11|37|si ceciderint super sementem non polluent eam
LEV|11|38|sin autem quispiam aqua sementem perfuderit et postea morticinis tacta fuerit ilico polluetur
LEV|11|39|si mortuum fuerit animal quod licet vobis comedere qui cadaver eius tetigerit inmundus erit usque ad vesperum
LEV|11|40|et qui comederit ex eo quippiam sive portaverit lavabit vestimenta sua et inmundus erit usque ad vesperum
LEV|11|41|omne quod reptat super terram abominabile erit nec adsumetur in cibum
LEV|11|42|quicquid super pectus quadrupes graditur et multos habet pedes sive per humum trahitur non comedetis quia abominabile est
LEV|11|43|nolite contaminare animas vestras nec tangatis quicquam eorum ne inmundi sitis
LEV|11|44|ego enim sum Dominus Deus vester sancti estote quoniam et ego sanctus sum ne polluatis animas vestras in omni reptili quod movetur super terram
LEV|11|45|ego sum Dominus qui eduxi vos de terra Aegypti ut essem vobis in Deum sancti eritis quia et ego sanctus sum
LEV|11|46|ista est lex animantium et volucrum et omnis animae viventis quae movetur in aqua et reptat in terra
LEV|11|47|ut differentias noveritis mundi et inmundi et sciatis quid comedere et quid respuere debeatis
LEV|12|1|locutus est Dominus ad Mosen dicens
LEV|12|2|loquere filiis Israhel et dices ad eos mulier si suscepto semine pepererit masculum inmunda erit septem diebus iuxta dies separationis menstruae
LEV|12|3|et die octavo circumcidetur infantulus
LEV|12|4|ipsa vero triginta tribus diebus manebit in sanguine purificationis suae omne sanctum non tanget nec ingredietur sanctuarium donec impleantur dies purificationis eius
LEV|12|5|sin autem feminam pepererit inmunda erit duabus ebdomadibus iuxta ritum fluxus menstrui et sexaginta ac sex diebus manebit in sanguine purificationis suae
LEV|12|6|cumque expleti fuerint dies purificationis eius pro filio sive pro filia deferet agnum anniculum in holocaustum et pullum columbae sive turturem pro peccato ad ostium tabernaculi testimonii et tradet sacerdoti
LEV|12|7|qui offeret illa coram Domino et rogabit pro ea et sic mundabitur a profluvio sanguinis sui ista est lex parientis masculum ac feminam
LEV|12|8|quod si non invenerit manus eius nec potuerit offerre agnum sumet duos turtures vel duos pullos columbae unum in holocaustum et alterum pro peccato orabitque pro ea sacerdos et sic mundabitur
LEV|13|1|locutus est Dominus ad Mosen et Aaron dicens
LEV|13|2|homo in cuius carne et cute ortus fuerit diversus color sive pustula aut quasi lucens quippiam id est plaga leprae adducetur ad Aaron sacerdotem vel ad unum quemlibet filiorum eius
LEV|13|3|qui cum viderit lepram in cute et pilos in album mutatos colorem ipsamque speciem leprae humiliorem cute et carne reliqua plaga leprae est et ad arbitrium eius separabitur
LEV|13|4|sin autem lucens candor fuerit in cute nec humilior carne reliqua et pili coloris pristini recludet eum sacerdos septem diebus
LEV|13|5|et considerabit die septimo et siquidem lepra ultra non creverit nec transierit in cute priores terminos rursum includet eum septem diebus aliis
LEV|13|6|et die septimo contemplabitur si obscurior fuerit lepra et non creverit in cute mundabit eum quia scabies est lavabitque homo vestimenta sua et mundus erit
LEV|13|7|quod si postquam a sacerdote visus est et redditus munditiae iterum lepra creverit adducetur ad eum
LEV|13|8|et inmunditiae condemnabitur
LEV|13|9|plaga leprae si fuerit in homine adducetur ad sacerdotem
LEV|13|10|et videbit eum cumque color albus in cute fuerit et capillorum mutarit aspectum ipsa quoque caro viva apparuerit
LEV|13|11|lepra vetustissima iudicabitur atque inolita cuti contaminabit itaque eum sacerdos et non recludet quia perspicue inmunditia est
LEV|13|12|sin autem effloruerit discurrens lepra in cute et operuerit omnem carnem a capite usque ad pedes quicquid sub aspectu oculorum cadit
LEV|13|13|considerabit eum sacerdos et teneri lepra mundissima iudicabit eo quod omnis in candorem versa sit et idcirco homo mundus erit
LEV|13|14|quando vero caro vivens in eo apparuerit
LEV|13|15|tunc sacerdotis iudicio polluetur et inter inmundos reputabitur caro enim viva si lepra aspergatur inmunda est
LEV|13|16|quod si rursum versa fuerit in alborem et totum hominem operuerit
LEV|13|17|considerabit eum sacerdos et mundum esse decernet
LEV|13|18|caro et cutis in qua ulcus natum est et sanatum
LEV|13|19|et in loco ulceris cicatrix apparuerit alba sive subrufa adducetur homo ad sacerdotem
LEV|13|20|qui cum viderit locum leprae humiliorem carne reliqua et pilos versos in candorem contaminabit eum plaga enim leprae orta est in ulcere
LEV|13|21|quod si pilus coloris est pristini et cicatrix subobscura et vicina carne non est humilior recludet eum septem diebus
LEV|13|22|et siquidem creverit adiudicabit eum leprae
LEV|13|23|sin autem steterit in loco suo ulceris est cicatrix et homo mundus erit
LEV|13|24|caro et cutis quam ignis exuserit et sanata albam sive rufam habuerit cicatricem
LEV|13|25|considerabit eam sacerdos et ecce versa est in alborem et locus eius reliqua cute humilior contaminabit eum quia plaga leprae in cicatrice orta est
LEV|13|26|quod si pilorum color non fuerit inmutatus nec humilior plaga carne reliqua et ipsa leprae species fuerit subobscura recludet eum septem diebus
LEV|13|27|et die septimo contemplabitur si creverit in cute lepra contaminabit eum
LEV|13|28|sin autem in loco suo candor steterit non satis clarus plaga conbustionis est et idcirco mundabitur quia cicatrix est conbusturae
LEV|13|29|vir sive mulier in cuius capite vel barba germinarit lepra videbit eos sacerdos
LEV|13|30|et siquidem humilior fuerit locus carne reliqua et capillus flavus solitoque subtilior contaminabit eos quia lepra capitis ac barbae est
LEV|13|31|sin autem viderit et locum maculae aequalem vicinae carni et capillum nigrum recludet eos septem diebus
LEV|13|32|et die septimo intuebitur si non creverit macula et capillus sui coloris est et locus plagae carni reliquae aequalis
LEV|13|33|radetur homo absque loco maculae et includetur septem diebus aliis
LEV|13|34|si die septimo visa fuerit stetisse plaga in loco suo nec humilior carne reliqua mundabit eum lotisque vestibus mundus erit
LEV|13|35|sin autem post emundationem rursus creverit macula in cute
LEV|13|36|non quaeret amplius utrum capillus in flavum colorem sit commutatus quia aperte inmundus est
LEV|13|37|porro si steterit macula et capilli nigri fuerint noverit hominem esse sanatum et confidenter eum pronuntiet mundum
LEV|13|38|vir et mulier in cuius cute candor apparuerit
LEV|13|39|intuebitur eos sacerdos si deprehenderit subobscurum alborem lucere in cute sciat non esse lepram sed maculam coloris candidi et hominem mundum
LEV|13|40|vir de cuius capite capilli fluunt calvus ac mundus est
LEV|13|41|et si a fronte ceciderint pili recalvaster et mundus est
LEV|13|42|sin autem in calvitio sive in recalvatione albus vel rufus color fuerit exortus
LEV|13|43|et hoc sacerdos viderit condemnabit eum haut dubiae leprae quae orta est in calvitio
LEV|13|44|quicumque ergo maculatus fuerit lepra et separatus ad arbitrium sacerdotis
LEV|13|45|habebit vestimenta dissuta caput nudum os veste contectum contaminatum ac sordidum se clamabit
LEV|13|46|omni tempore quo leprosus est et inmundus solus habitabit extra castra
LEV|13|47|vestis lanea sive linea quae lepram habuerit
LEV|13|48|in stamine atque subtemine aut certe pellis vel quicquid ex pelle confectum est
LEV|13|49|si alba aut rufa macula fuerit infecta lepra reputabitur ostendeturque sacerdoti
LEV|13|50|qui consideratam recludet septem diebus
LEV|13|51|et die septimo rursus aspiciens si crevisse deprehenderit lepra perseverans est pollutum iudicabit vestimentum et omne in quo fuerit inventa
LEV|13|52|et idcirco conburetur flammis
LEV|13|53|quod si eam viderit non crevisse
LEV|13|54|praecipiet et lavabunt id in quo lepra est recludetque illud septem diebus aliis
LEV|13|55|et cum viderit faciem quidem pristinam non reversam nec tamen crevisse lepram inmundum iudicabit et igne conburet eo quod infusa sit in superficie vestimenti vel per totum lepra
LEV|13|56|sin autem obscurior fuerit locus leprae postquam vestis est lota abrumpet eum et a solido dividet
LEV|13|57|quod si ultra apparuerit in his locis quae prius inmaculata erant lepra volatilis et vaga debet igne conburi
LEV|13|58|si cessaverit lavabit ea quae pura sunt secundo et munda erunt
LEV|13|59|ista est lex leprae vestimenti lanei et linei staminis atque subteminis omnisque supellectilis pelliciae quomodo mundari debeat vel contaminari
LEV|14|1|locutusque est Dominus ad Mosen dicens
LEV|14|2|hic est ritus leprosi quando mundandus est adducetur ad sacerdotem
LEV|14|3|qui egressus e castris cum invenerit lepram esse mundatam
LEV|14|4|praecipiet ei qui purificatur ut offerat pro se duos passeres vivos quos vesci licitum est et lignum cedrinum vermiculumque et hysopum
LEV|14|5|et unum e passeribus immolari iubebit in vase fictili super aquas viventes
LEV|14|6|alium autem vivum cum ligno cedrino et cocco et hysopo tinguet in sanguine passeris immolati
LEV|14|7|quo asperget illum qui mundandus est septies ut iure purgetur et dimittet passerem vivum ut in agrum avolet
LEV|14|8|cumque laverit homo vestimenta sua radet omnes pilos corporis et lavabitur aqua purificatusque ingredietur castra ita dumtaxat ut maneat extra tabernaculum suum septem diebus
LEV|14|9|et die septimo radat capillos capitis barbamque et supercilia ac totius corporis pilos et lotis rursum vestibus et corpore
LEV|14|10|die octavo adsumet duos agnos inmaculatos et ovem anniculam absque macula et tres decimas similae in sacrificium quae conspersa sit oleo et seorsum olei sextarium
LEV|14|11|cumque sacerdos purificans hominem statuerit eum et haec omnia coram Domino in ostio tabernaculi testimonii
LEV|14|12|tollet agnum et offeret eum pro delicto oleique sextarium et oblatis ante Dominum omnibus
LEV|14|13|immolabit agnum ubi immolari solet hostia pro peccato et holocaustum id est in loco sancto sicut enim pro peccato ita et pro delicto ad sacerdotem pertinet hostia sancta sanctorum est
LEV|14|14|adsumensque sacerdos de sanguine hostiae quae immolata est pro delicto ponet super extremum auriculae dextrae eius qui mundatur et super pollices manus dextrae et pedis
LEV|14|15|et de olei sextario mittet in manum suam sinistram
LEV|14|16|tinguetque digitum dextrum in eo et asperget septies contra Dominum
LEV|14|17|quod autem reliquum est olei in leva manu fundet super extremum auriculae dextrae eius qui mundatur et super pollices manus ac pedis dextri et super sanguinem qui fusus est pro delicto
LEV|14|18|et super caput eius
LEV|14|19|rogabitque pro eo coram Domino et faciet sacrificium pro peccato tunc immolabit holocaustum
LEV|14|20|et ponet illud in altari cum libamentis suis et homo rite mundabitur
LEV|14|21|quod si pauper est et non potest manus eius invenire quae dicta sunt adsumet agnum pro delicto ad oblationem ut roget pro eo sacerdos decimamque partem similae conspersae oleo in sacrificium et olei sextarium
LEV|14|22|duosque turtures sive duos pullos columbae quorum sit unus pro peccato et alter in holocaustum
LEV|14|23|offeretque ea die octavo purificationis suae sacerdoti ad ostium tabernaculi testimonii coram Domino
LEV|14|24|qui suscipiens agnum pro delicto et sextarium olei levabit simul
LEV|14|25|immolatoque agno de sanguine eius ponet super extremum auriculae dextrae illius qui mundatur et super pollices manus eius ac pedis dextri
LEV|14|26|olei vero partem mittet in manum suam sinistram
LEV|14|27|in quo tinguens digitum dextrae manus asperget septies contra Dominum
LEV|14|28|tangetque extremum dextrae auriculae illius qui mundatur et pollices manus ac pedis dextri in loco sanguinis qui effusus est pro delicto
LEV|14|29|reliquam autem partem olei quae est in sinistra manu mittet super caput purificati ut placet pro eo Dominum
LEV|14|30|et turturem sive pullum columbae offeret
LEV|14|31|unum pro delicto et alterum in holocaustum cum libamentis suis
LEV|14|32|hoc est sacrificium leprosi qui habere non potest omnia in emundationem sui
LEV|14|33|locutus est Dominus ad Mosen et Aaron dicens
LEV|14|34|cum ingressi fueritis terram Chanaan quam ego dabo vobis in possessionem si fuerit plaga leprae in aedibus
LEV|14|35|ibit cuius est domus nuntians sacerdoti et dicet quasi plaga leprae videtur mihi esse in domo mea
LEV|14|36|at ille praecipiet ut efferant universa de domo priusquam ingrediatur eam et videat utrum lepra sit ne inmunda fiant omnia quae in domo sunt intrabitque postea ut consideret domus lepram
LEV|14|37|et cum viderit in parietibus illius quasi valliculas pallore sive rubore deformes et humiliores superficie reliqua
LEV|14|38|egredietur ostium domus et statim claudet eam septem diebus
LEV|14|39|reversusque die septimo considerabit eam si invenerit crevisse lepram
LEV|14|40|iubebit erui lapides in quibus lepra est et proici eos extra civitatem in loco inmundo
LEV|14|41|domum autem ipsam radi intrinsecus per circuitum et spargi pulverem rasurae extra urbem in loco inmundo
LEV|14|42|lapidesque alios reponi pro his qui ablati fuerint et luto alio liniri domum
LEV|14|43|sin autem postquam eruti sunt lapides et pulvis elatus et alia terra lita
LEV|14|44|ingressus sacerdos viderit reversam lepram et parietes aspersos maculis lepra est perseverans et inmunda domus
LEV|14|45|quam statim destruent et lapides eius ac ligna atque universum pulverem proicient extra oppidum in loco inmundo
LEV|14|46|qui intraverit domum quando clausa est inmundus erit usque ad vesperum
LEV|14|47|et qui dormierit in ea et comederit quippiam lavabit vestimenta sua
LEV|14|48|quod si introiens sacerdos viderit lepram non crevisse in domo postquam denuo lita est purificabit eam reddita sanitate
LEV|14|49|et in purificationem eius sumet duos passeres lignumque cedrinum et vermiculum atque hysopum
LEV|14|50|et immolato uno passere in vase fictili super aquas vivas
LEV|14|51|tollet lignum cedrinum et hysopum et coccum et passerem vivum et intinguet omnia in sanguine passeris immolati atque in aquis viventibus et asperget domum septies
LEV|14|52|purificabitque eam tam in sanguine passeris quam in aquis viventibus et in passere vivo lignoque cedrino et hysopo atque vermiculo
LEV|14|53|cumque dimiserit passerem avolare in agrum libere orabit pro domo et iure mundabitur
LEV|14|54|ista est lex omnis leprae et percussurae
LEV|14|55|leprae vestium et domorum
LEV|14|56|cicatricis et erumpentium papularum lucentis maculae et in varias species coloribus inmutatis
LEV|14|57|ut possit sciri quo tempore mundum quid vel inmundum sit
LEV|15|1|locutusque est Dominus ad Mosen et Aaron dicens
LEV|15|2|loquimini filiis Israhel et dicite eis vir qui patitur fluxum seminis inmundus erit
LEV|15|3|et tunc iudicabitur huic vitio subiacere cum per momenta singula adheserit carni illius atque concreverit foedus humor
LEV|15|4|omne stratum in quo dormierit inmundum erit et ubicumque sederit
LEV|15|5|si quis hominum tetigerit lectum eius lavabit vestimenta sua et ipse lotus aqua inmundus erit usque ad vesperum
LEV|15|6|si sederit ubi ille sederat et ipse lavabit vestimenta sua et lotus aqua inmundus erit usque ad vesperum
LEV|15|7|qui tetigerit carnem eius lavabit vestimenta sua et ipse lotus aqua inmundus erit usque ad vesperum
LEV|15|8|si salivam huiuscemodi homo iecerit super eum qui mundus est lavabit vestem suam et lotus aqua inmundus erit usque ad vesperum
LEV|15|9|sagma super quo sederit inmundum erit
LEV|15|10|et quicquid sub eo fuerit qui fluxum seminis patitur pollutum erit usque ad vesperum qui portaverit horum aliquid lavabit vestem suam et ipse lotus aqua inmundus erit usque ad vesperum
LEV|15|11|omnis quem tetigerit qui talis est non lotis ante manibus lavabit vestimenta sua et lotus aqua inmundus erit usque ad vesperum
LEV|15|12|vas fictile quod tetigerit confringetur vas autem ligneum lavabitur aqua
LEV|15|13|si sanatus fuerit qui huiuscemodi sustinet passionem numerabit septem dies post emundationem sui et lotis vestibus ac toto corpore in aquis viventibus erit mundus
LEV|15|14|die autem octavo sumet duos turtures aut duos pullos columbae et veniet in conspectu Domini ad ostium tabernaculi testimonii dabitque eos sacerdoti
LEV|15|15|qui faciet unum pro peccato et alterum in holocaustum rogabitque pro eo coram Domino ut emundetur a fluxu seminis sui
LEV|15|16|vir de quo egreditur semen coitus lavabit aqua omne corpus suum et inmundus erit usque ad vesperum
LEV|15|17|vestem et pellem quam habuerit lavabit aqua et inmunda erit usque ad vesperum
LEV|15|18|mulier cum qua coierit lavabitur aqua et inmunda erit usque ad vesperum
LEV|15|19|mulier quae redeunte mense patitur fluxum sanguinis septem diebus separabitur
LEV|15|20|omnis qui tetigerit eam inmundus erit usque ad vesperum
LEV|15|21|et in quo dormierit vel sederit diebus separationis suae polluetur
LEV|15|22|qui tetigerit lectum eius lavabit vestimenta sua et ipse lotus aqua inmundus erit usque ad vesperum
LEV|15|23|omne vas super quo illa sederit quisquis adtigerit lavabit vestimenta sua et lotus aqua pollutus erit usque ad vesperum
LEV|15|24|si coierit cum ea vir tempore sanguinis menstrualis inmundus erit septem diebus et omne stratum in quo dormierit polluetur
LEV|15|25|mulier quae patitur multis diebus fluxum sanguinis non in tempore menstruali vel quae post menstruum sanguinem fluere non cessat quamdiu huic subiacet passioni inmunda erit quasi sit in tempore menstruo
LEV|15|26|omne stratum in quo dormierit et vas in quo sederit pollutum erit
LEV|15|27|quicumque tetigerit eam lavabit vestimenta sua et ipse lotus aqua inmundus erit usque ad vesperum
LEV|15|28|si steterit sanguis et fluere cessarit numerabit septem dies purificationis suae
LEV|15|29|et octavo die offeret pro se sacerdoti duos turtures vel duos pullos columbae ad ostium tabernaculi testimonii
LEV|15|30|qui unum faciet pro peccato et alterum in holocaustum rogabitque pro ea coram Domino et pro fluxu inmunditiae eius
LEV|15|31|docebitis ergo filios Israhel ut caveant inmunditiam et non moriantur in sordibus suis cum polluerint tabernaculum meum quod est inter eos
LEV|15|32|ista est lex eius qui patitur fluxum seminis et qui polluitur coitu
LEV|15|33|et quae menstruis temporibus separatur vel quae iugi fluit sanguine et hominis qui dormierit cum ea
LEV|16|1|locutusque est Dominus ad Mosen post mortem duum filiorum Aaron quando offerentes ignem alienum interfecti sunt
LEV|16|2|et praecepit ei dicens loquere ad Aaron fratrem tuum ne omni tempore ingrediatur sanctuarium quod est intra velum coram propitiatorio quo tegitur arca ut non moriatur quia in nube apparebo super oraculum
LEV|16|3|nisi haec ante fecerit vitulum offeret pro peccato et arietem in holocaustum
LEV|16|4|tunica linea vestietur feminalibus lineis verecunda celabit accingetur zona linea cidarim lineam inponet capiti haec enim vestimenta sunt sancta quibus cunctis cum lotus fuerit induetur
LEV|16|5|suscipietque ab universa multitudine filiorum Israhel duos hircos pro peccato et unum arietem in holocaustum
LEV|16|6|cumque obtulerit vitulum et oraverit pro se et pro domo sua
LEV|16|7|duos hircos stare faciet coram Domino in ostio tabernaculi testimonii
LEV|16|8|mittens super utrumque sortem unam Domino et alteram capro emissario
LEV|16|9|cuius sors exierit Domino offeret illum pro peccato
LEV|16|10|cuius autem in caprum emissarium statuet eum vivum coram Domino ut fundat preces super eo et emittat illum in solitudinem
LEV|16|11|his rite celebratis offeret vitulum et rogans pro se et pro domo sua immolabit eum
LEV|16|12|adsumptoque turibulo quod de prunis altaris impleverit et hauriens manu conpositum thymiama in incensum ultra velum intrabit in sancta
LEV|16|13|ut positis super ignem aromatibus nebula eorum et vapor operiat oraculum quod est super testimonium et non moriatur
LEV|16|14|tollet quoque de sanguine vituli et asperget digito septies contra propitiatorium ad orientem
LEV|16|15|cumque mactaverit hircum pro peccato populi inferet sanguinem eius intra velum sicut praeceptum est de sanguine vituli ut aspergat e regione oraculi
LEV|16|16|et expiet sanctuarium ab inmunditiis filiorum Israhel et a praevaricationibus eorum cunctisque peccatis iuxta hunc ritum faciet tabernaculo testimonii quod fixum est inter eos in medio sordium habitationis eorum
LEV|16|17|nullus hominum sit in tabernaculo quando pontifex ingreditur sanctuarium ut roget pro se et pro domo sua et pro universo coetu Israhel donec egrediatur
LEV|16|18|cum autem exierit ad altare quod coram Domino est oret pro se et sumptum sanguinem vituli atque hirci fundat super cornua eius per gyrum
LEV|16|19|aspergensque digito septies expiet et sanctificet illud ab inmunditiis filiorum Israhel
LEV|16|20|postquam emundarit sanctuarium et tabernaculum et altare tunc offerat hircum viventem
LEV|16|21|et posita utraque manu super caput eius confiteatur omnes iniquitates filiorum Israhel et universa delicta atque peccata eorum quae inprecans capiti eius emittet illum per hominem paratum in desertum
LEV|16|22|cumque portaverit hircus omnes iniquitates eorum in terram solitariam et dimissus fuerit in deserto
LEV|16|23|revertetur Aaron in tabernaculum testimonii et depositis vestibus quibus prius indutus erat cum intraret sanctuarium relictisque ibi
LEV|16|24|lavabit carnem suam in loco sancto indueturque vestimentis suis et postquam egressus obtulerit holocaustum suum ac plebis rogabit tam pro se quam pro populo
LEV|16|25|et adipem qui oblatus est pro peccatis adolebit super altare
LEV|16|26|ille vero qui dimiserit caprum emissarium lavabit vestimenta sua et corpus aqua et sic ingredietur in castra
LEV|16|27|vitulum autem et hircum qui pro peccato fuerant immolati et quorum sanguis inlatus est ut in sanctuario expiatio conpleretur asportabunt foras castra et conburent igni tam pelles quam carnes eorum et fimum
LEV|16|28|et quicumque conbuserit ea lavabit vestimenta sua et carnem aqua et sic ingredietur in castra
LEV|16|29|eritque hoc vobis legitimum sempiternum mense septimo decima die mensis adfligetis animas vestras nullumque facietis opus sive indigena sive advena qui peregrinatur inter vos
LEV|16|30|in hac die expiatio erit vestri atque mundatio ab omnibus peccatis vestris coram Domino mundabimini
LEV|16|31|sabbatum enim requietionis est et adfligetis animas vestras religione perpetua
LEV|16|32|expiabit autem sacerdos qui unctus fuerit et cuius initiatae manus ut sacerdotio fungatur pro patre suo indueturque stola linea et vestibus sanctis
LEV|16|33|et expiabit sanctuarium et tabernaculum testimonii atque altare sacerdotes quoque et universum populum
LEV|16|34|eritque hoc vobis legitimum sempiternum ut oretis pro filiis Israhel et pro cunctis peccatis eorum semel in anno fecit igitur sicut praeceperat Dominus Mosi
LEV|17|1|et locutus est Dominus ad Mosen dicens
LEV|17|2|loquere Aaron et filiis eius et cunctis filiis Israhel et dices ad eos iste est sermo quem mandavit Dominus dicens
LEV|17|3|homo quilibet de domo Israhel si occiderit bovem aut ovem sive capram in castris vel extra castra
LEV|17|4|et non obtulerit ad ostium tabernaculi oblationem Domino sanguinis reus erit quasi sanguinem fuderit sic peribit de medio populi sui
LEV|17|5|ideo offerre debent sacerdoti filii Israhel hostias suas quas occidunt in agro ut sanctificentur Domino ante ostium tabernaculi testimonii et immolent eas hostias pacificas Domino
LEV|17|6|fundetque sacerdos sanguinem super altare Domini ad ostium tabernaculi testimonii et adolebit adipem in odorem suavitatis Domino
LEV|17|7|et nequaquam ultra immolabunt hostias suas daemonibus cum quibus fornicati sunt legitimum sempiternum erit illis et posteris eorum
LEV|17|8|et ad ipsos dices homo de domo Israhel et de advenis qui peregrinantur apud vos qui obtulerit holocaustum sive victimam
LEV|17|9|et ad ostium tabernaculi testimonii non adduxerit eam ut offeratur Domino interibit de populo suo
LEV|17|10|homo quilibet de domo Israhel et de advenis qui peregrinantur inter eos si comederit sanguinem obfirmabo faciem meam contra animam illius et disperdam eam de populo suo
LEV|17|11|quia anima carnis in sanguine est et ego dedi illum vobis ut super altare in eo expietis pro animabus vestris et sanguis pro animae piaculo sit
LEV|17|12|idcirco dixi filiis Israhel omnis anima ex vobis non comedet sanguinem nec ex advenis qui peregrinantur inter vos
LEV|17|13|homo quicumque de filiis Israhel et de advenis qui peregrinantur apud vos si venatione atque aucupio ceperit feram vel avem quibus vesci licitum est fundat sanguinem eius et operiat illum terra
LEV|17|14|anima enim omnis carnis in sanguine est unde dixi filiis Israhel sanguinem universae carnis non comedetis quia anima carnis in sanguine est et quicumque comederit illum interibit
LEV|17|15|anima quae comederit morticinum vel captum a bestia tam de indigenis quam de advenis lavabit vestes suas et semet ipsum aqua et contaminatus erit usque ad vesperum et hoc ordine mundus fiet
LEV|17|16|quod si non laverit vestimenta sua nec corpus portabit iniquitatem suam
LEV|18|1|locutusque est Dominus ad Mosen dicens
LEV|18|2|loquere filiis Israhel et dices ad eos ego Dominus Deus vester
LEV|18|3|iuxta consuetudinem terrae Aegypti in qua habitastis non facietis et iuxta morem regionis Chanaan ad quam ego introducturus sum vos non agetis nec in legitimis eorum ambulabitis
LEV|18|4|facietis iudicia mea et praecepta servabitis et ambulabitis in eis ego Dominus Deus vester
LEV|18|5|custodite leges meas atque iudicia quae faciens homo vivet in eis ego Dominus
LEV|18|6|omnis homo ad proximam sanguinis sui non accedet ut revelet turpitudinem eius ego Dominus
LEV|18|7|turpitudinem patris et turpitudinem matris tuae non discoperies mater tua est non revelabis turpitudinem eius
LEV|18|8|turpitudinem uxoris patris tui non discoperies turpitudo enim patris tui est
LEV|18|9|turpitudinem sororis tuae ex patre sive ex matre quae domi vel foris genita est non revelabis
LEV|18|10|turpitudinem filiae filii tui vel neptis ex filia non revelabis quia turpitudo tua est
LEV|18|11|turpitudinem filiae uxoris patris tui quam peperit patri tuo et est soror tua non revelabis
LEV|18|12|turpitudinem sororis patris tui non discoperies quia caro est patris tui
LEV|18|13|turpitudinem sororis matris tuae non revelabis eo quod caro sit matris tuae
LEV|18|14|turpitudinem patrui tui non revelabis nec accedes ad uxorem eius quae tibi adfinitate coniungitur
LEV|18|15|turpitudinem nurus tuae non revelabis quia uxor filii tui est nec discoperies ignominiam eius
LEV|18|16|turpitudinem uxoris fratris tui non revelabis quia turpitudo fratris tui est
LEV|18|17|turpitudinem uxoris tuae et filiae eius non revelabis filiam filii eius et filiam filiae illius non sumes ut reveles ignominiam eius quia caro illius sunt et talis coitus incestus est
LEV|18|18|sororem uxoris tuae in pelicatum illius non accipies nec revelabis turpitudinem eius adhuc illa vivente
LEV|18|19|ad mulierem quae patitur menstrua non accedes nec revelabis foeditatem eius
LEV|18|20|cum uxore proximi tui non coibis nec seminis commixtione maculaberis
LEV|18|21|de semine tuo non dabis ut consecretur idolo Moloch nec pollues nomen Dei tui ego Dominus
LEV|18|22|cum masculo non commisceberis coitu femineo quia abominatio est
LEV|18|23|cum omni pecore non coibis nec maculaberis cum eo mulier non subcumbet iumento nec miscebitur ei quia scelus est
LEV|18|24|ne polluamini in omnibus his quibus contaminatae sunt universae gentes quas ego eiciam ante conspectum vestrum
LEV|18|25|et quibus polluta est terra cuius ego scelera visitabo ut evomat habitatores suos
LEV|18|26|custodite legitima mea atque iudicia et non faciat ex omnibus abominationibus istis tam indigena quam colonus qui peregrinatur apud vos
LEV|18|27|omnes enim execrationes istas fecerunt accolae terrae qui fuerunt ante vos et polluerunt eam
LEV|18|28|cavete ergo ne et vos similiter evomat cum paria feceritis sicut evomuit gentem quae fuit ante vos
LEV|18|29|omnis anima quae fecerit de abominationibus his quippiam peribit de medio populi sui
LEV|18|30|custodite mandata mea nolite facere quae fecerunt hii qui fuerunt ante vos et ne polluamini in eis ego Dominus Deus vester
LEV|19|1|locutus est Dominus ad Mosen dicens
LEV|19|2|loquere ad omnem coetum filiorum Israhel et dices ad eos sancti estote quia ego sanctus sum Dominus Deus vester
LEV|19|3|unusquisque matrem et patrem suum timeat sabbata mea custodite ego Dominus Deus vester
LEV|19|4|nolite converti ad idola nec deos conflatiles faciatis vobis ego Dominus Deus vester
LEV|19|5|si immolaveritis hostiam pacificorum Domino ut sit placabilis
LEV|19|6|eo die quo fuerit immolata comedetis eam et die altero quicquid autem residuum fuerit in diem tertium igne conburetis
LEV|19|7|si quis post biduum comederit ex ea profanus erit et impietatis reus
LEV|19|8|portabit iniquitatem suam quia sanctum Domini polluit et peribit anima illa de populo suo
LEV|19|9|cum messueris segetes terrae tuae non tondebis usque ad solum superficiem terrae nec remanentes spicas colliges
LEV|19|10|neque in vinea tua racemos et grana decidentia congregabis sed pauperibus et peregrinis carpenda dimittes ego Dominus Deus vester
LEV|19|11|non facietis furtum non mentiemini nec decipiet unusquisque proximum suum
LEV|19|12|non peierabis in nomine meo nec pollues nomen Dei tui ego Dominus
LEV|19|13|non facies calumniam proximo tuo nec vi opprimes eum non morabitur opus mercennarii apud te usque mane
LEV|19|14|non maledices surdo nec coram caeco pones offendiculum sed timebis Deum tuum quia ego sum Dominus
LEV|19|15|non facies quod iniquum est nec iniuste iudicabis nec consideres personam pauperis nec honores vultum potentis iuste iudica proximo tuo
LEV|19|16|non eris criminator et susurro in populis non stabis contra sanguinem proximi tui ego Dominus
LEV|19|17|ne oderis fratrem tuum in corde tuo sed publice argue eum ne habeas super illo peccatum
LEV|19|18|non quaeres ultionem nec memor eris iniuriae civium tuorum diliges amicum tuum sicut temet ipsum ego Dominus
LEV|19|19|leges meas custodite iumenta tua non facies coire cum alterius generis animantibus agrum non seres diverso semine veste quae ex duobus texta est non indueris
LEV|19|20|homo si dormierit cum muliere coitu seminis quae sit ancilla etiam nubilis et tamen pretio non redempta nec libertate donata vapulabunt ambo et non morientur quia non fuit libera
LEV|19|21|pro delicto autem suo offeret Domino ad ostium tabernaculi testimonii arietem
LEV|19|22|orabitque pro eo sacerdos et pro delicto eius coram Domino et repropitiabitur ei dimitteturque peccatum
LEV|19|23|quando ingressi fueritis terram et plantaveritis in ea ligna pomifera auferetis praeputia eorum poma quae germinant inmunda erunt vobis nec edetis ex eis
LEV|19|24|quarto anno omnis fructus eorum sanctificabitur laudabilis Domino
LEV|19|25|quinto autem anno comedetis fructus congregantes poma quae proferunt ego Dominus Deus vester
LEV|19|26|non comedetis cum sanguine non augurabimini nec observabitis somnia
LEV|19|27|neque in rotundum adtondebitis comam nec radatis barbam
LEV|19|28|et super mortuo non incidetis carnem vestram neque figuras aliquas et stigmata facietis vobis ego Dominus
LEV|19|29|ne prostituas filiam tuam et contaminetur terra et impleatur piaculo
LEV|19|30|sabbata mea custodite et sanctuarium meum metuite ego Dominus
LEV|19|31|ne declinetis ad magos nec ab ariolis aliquid sciscitemini ut polluamini per eos ego Dominus Deus vester
LEV|19|32|coram cano capite consurge et honora personam senis et time Deum tuum ego sum Dominus
LEV|19|33|si habitaverit advena in terra vestra et moratus fuerit inter vos ne exprobretis ei
LEV|19|34|sed sit inter vos quasi indigena et diligetis eum quasi vosmet ipsos fuistis enim et vos advenae in terra Aegypti ego Dominus Deus vester
LEV|19|35|nolite facere iniquum aliquid in iudicio in regula in pondere in mensura
LEV|19|36|statera iusta et aequa sint pondera iustus modius aequusque sextarius ego Dominus Deus vester qui eduxi vos de terra Aegypti
LEV|19|37|custodite omnia praecepta mea et universa iudicia et facite ea ego Dominus
LEV|20|1|locutusque est Dominus ad Mosen dicens
LEV|20|2|haec loqueris filiis Israhel homo de filiis Israhel et de advenis qui habitant in Israhel si quis dederit de semine suo idolo Moloch morte moriatur populus terrae lapidabit eum
LEV|20|3|et ego ponam faciem meam contra illum succidamque eum de medio populi sui eo quod dederit de semine suo Moloch et contaminaverit sanctuarium meum ac polluerit nomen sanctum meum
LEV|20|4|quod si neglegens populus terrae et quasi parvipendens imperium meum dimiserit hominem qui dederit de semine suo Moloch nec voluerit eum occidere
LEV|20|5|ponam faciem meam super hominem illum et cognationem eius succidamque et ipsum et omnes qui consenserunt ei ut fornicarentur cum Moloch de medio populi sui
LEV|20|6|anima quae declinaverit ad magos et ariolos et fornicata fuerit cum eis ponam faciem meam contra eam et interficiam illam de medio populi sui
LEV|20|7|sanctificamini et estote sancti quia ego Dominus Deus vester
LEV|20|8|custodite praecepta mea et facite ea ego Dominus qui sanctifico vos
LEV|20|9|qui maledixerit patri suo et matri morte moriatur patri matrique maledixit sanguis eius sit super eum
LEV|20|10|si moechatus quis fuerit cum uxore alterius et adulterium perpetrarit cum coniuge proximi sui morte moriantur et moechus et adultera
LEV|20|11|qui dormierit cum noverca sua et revelaverit ignominiam patris sui morte moriantur ambo sanguis eorum sit super eos
LEV|20|12|si quis dormierit cum nuru sua uterque moriantur quia scelus operati sunt sanguis eorum sit super eos
LEV|20|13|qui dormierit cum masculo coitu femineo uterque operati sunt nefas morte moriantur sit sanguis eorum super eos
LEV|20|14|qui supra uxorem filiam duxerit matrem eius scelus operatus est vivus ardebit cum eis nec permanebit tantum nefas in medio vestri
LEV|20|15|qui cum iumento et pecore coierit morte moriatur pecus quoque occidite
LEV|20|16|mulier quae subcubuerit cuilibet iumento simul interficietur cum eo sanguis eorum sit super eos
LEV|20|17|qui acceperit sororem suam filiam patris sui vel filiam matris suae et viderit turpitudinem eius illaque conspexerit fratris ignominiam nefariam rem operati sunt occidentur in conspectu populi sui eo quod turpitudinem suam mutuo revelarint et portabunt iniquitatem suam
LEV|20|18|qui coierit cum muliere in fluxu menstruo et revelaverit turpitudinem eius ipsaque aperuerit fontem sanguinis sui interficientur ambo de medio populi sui
LEV|20|19|turpitudinem materterae tuae et amitae tuae non discoperies qui hoc fecerit ignominiam carnis suae nudavit portabunt ambo iniquitatem suam
LEV|20|20|qui coierit cum uxore patrui vel avunculi sui et revelaverit ignominiam cognationis suae portabunt ambo peccatum suum absque liberis morientur
LEV|20|21|qui duxerit uxorem fratris sui rem facit inlicitam turpitudinem fratris sui revelavit absque filiis erunt
LEV|20|22|custodite leges meas atque iudicia et facite ea ne et vos evomat terra quam intraturi estis et habitaturi
LEV|20|23|nolite ambulare in legitimis nationum quas ego expulsurus sum ante vos omnia enim haec fecerunt et abominatus sum eos
LEV|20|24|vobis autem loquor possidete terram eorum quam dabo vobis in hereditatem terram fluentem lacte et melle ego Dominus Deus vester qui separavi vos a ceteris populis
LEV|20|25|separate ergo et vos iumentum mundum ab inmundo et avem mundam ab inmunda ne polluatis animas vestras in pecore et in avibus et cunctis quae moventur in terra et quae vobis ostendi esse polluta
LEV|20|26|eritis sancti mihi quia sanctus ego sum Dominus et separavi vos a ceteris populis ut essetis mei
LEV|20|27|vir sive mulier in quibus pythonicus vel divinationis fuerit spiritus morte moriantur lapidibus obruent eos sanguis eorum sit super illos
LEV|21|1|dixit quoque Dominus ad Mosen loquere ad sacerdotes filios Aaron et dices eis ne contaminetur sacerdos in mortibus civium suorum
LEV|21|2|nisi tantum in consanguineis ac propinquis id est super matre et patre et filio ac filia fratre quoque
LEV|21|3|et sorore virgine quae non est nupta viro
LEV|21|4|sed nec in principe populi sui contaminabitur
LEV|21|5|non radent caput nec barbam neque in carnibus suis facient incisuras
LEV|21|6|sancti erunt Deo suo et non polluent nomen eius incensum enim Domini et panes Dei sui offerunt et ideo sancti erunt
LEV|21|7|scortum et vile prostibulum non ducet uxorem nec eam quae repudiata est a marito quia consecratus est Deo suo
LEV|21|8|et panes propositionis offert sit ergo sanctus quia et ego sanctus sum Dominus qui sanctifico vos
LEV|21|9|sacerdotis filia si deprehensa fuerit in stupro et violaverit nomen patris sui flammis exuretur
LEV|21|10|pontifex id est sacerdos maximus inter fratres suos super cuius caput fusum est unctionis oleum et cuius manus in sacerdotio consecratae sunt vestitusque est sanctis vestibus caput suum non discoperiet vestimenta non scindet
LEV|21|11|et ad omnem mortuum non ingredietur omnino super patre quoque suo et matre non contaminabitur
LEV|21|12|nec egredietur de sanctis ne polluat sanctuarium Domini quia oleum sanctae unctionis Dei sui super eum est ego Dominus
LEV|21|13|virginem ducet uxorem
LEV|21|14|viduam et repudiatam et sordidam atque meretricem non accipiet sed puellam de populo suo
LEV|21|15|ne commisceat stirpem generis sui vulgo gentis suae quia ego Dominus qui sanctifico eum
LEV|21|16|locutusque est Dominus ad Mosen dicens
LEV|21|17|loquere ad Aaron homo de semine tuo per familias qui habuerit maculam non offeret panes Deo suo
LEV|21|18|nec accedet ad ministerium eius si caecus fuerit si claudus si vel parvo vel grandi et torto naso
LEV|21|19|si fracto pede si manu
LEV|21|20|si gibbus si lippus si albuginem habens in oculo si iugem scabiem si inpetiginem in corpore vel hirniosus
LEV|21|21|omnis qui habuerit maculam de semine Aaron sacerdotis non accedet offerre hostias Domino nec panes Deo suo
LEV|21|22|vescetur tamen panibus qui offeruntur in sanctuario
LEV|21|23|ita dumtaxat ut intra velum non ingrediatur nec accedat ad altare quia maculam habet et contaminare non debet sanctuarium meum ego Dominus qui sanctifico eos
LEV|21|24|locutus est ergo Moses ad Aaron et filios eius et ad omnem Israhel cuncta quae sibi fuerant imperata
LEV|22|1|locutus quoque est Dominus ad Mosen dicens
LEV|22|2|loquere ad Aaron et ad filios eius ut caveant ab his quae consecrata sunt filiorum Israhel et non contaminent nomen sanctificatorum mihi quae ipsi offerunt ego Dominus
LEV|22|3|dic ad eos et ad posteros eorum omnis homo qui accesserit de stirpe vestra ad ea quae consecrata sunt et quae obtulerunt filii Israhel Domino in quo est inmunditia peribit coram Domino ego sum Dominus
LEV|22|4|homo de semine Aaron qui fuerit leprosus aut patiens fluxum seminis non vescetur de his quae sanctificata sunt mihi donec sanetur qui tetigerit inmundum super mortuo et ex quo egreditur semen quasi coitus
LEV|22|5|et qui tangit reptile et quodlibet inmundum cuius tactus est sordidus
LEV|22|6|inmundus erit usque ad vesperum et non vescetur his quae sanctificata sunt sed cum laverit carnem suam aqua
LEV|22|7|et occubuerit sol tunc mundatus vescetur de sanctificatis quia cibus illius est
LEV|22|8|morticinum et captum a bestia non comedent nec polluentur in eis ego sum Dominus
LEV|22|9|custodient praecepta mea ut non subiaceant peccato et moriantur in sanctuario cum polluerint illud ego Dominus qui sanctifico eos
LEV|22|10|omnis alienigena non comedet de sanctificatis inquilinus sacerdotis et mercennarius non vescentur ex eis
LEV|22|11|quem autem sacerdos emerit et qui vernaculus domus eius fuerit hii comedent ex eis
LEV|22|12|si filia sacerdotis cuilibet ex populo nupta fuerit de his quae sanctificata sunt et de primitiis non vescetur
LEV|22|13|sin autem vidua vel repudiata et absque liberis reversa fuerit ad domum patris sui sicut puella consuerat aletur cibis patris sui omnis alienigena comedendi ex eis non habet potestatem
LEV|22|14|qui comederit de sanctificatis per ignorantiam addet quintam partem cum eo quod comedit et dabit sacerdoti in sanctuarium
LEV|22|15|nec contaminabunt sanctificata filiorum Israhel quae offerunt Domino
LEV|22|16|ne forte sustineant iniquitatem delicti sui cum sanctificata comederint ego Dominus qui sanctifico eos
LEV|22|17|locutus est Dominus ad Mosen dicens
LEV|22|18|loquere ad Aaron et filios eius et ad omnes filios Israhel dicesque ad eos homo de domo Israhel et de advenis qui habitant apud vos qui obtulerit oblationem suam vel vota solvens vel sponte offerens quicquid illud obtulerit in holocaustum Domini
LEV|22|19|ut offeratur per vos masculus inmaculatus erit ex bubus et ex ovibus et ex capris
LEV|22|20|si maculam habuerit non offeretis neque erit acceptabile
LEV|22|21|homo qui obtulerit victimam pacificorum Domino vel vota solvens vel sponte offerens tam de bubus quam de ovibus inmaculatum offeret ut acceptabile sit omnis macula non erit in eo
LEV|22|22|si caecum fuerit si fractum si cicatricem habens si papulas aut scabiem vel inpetiginem non offeretis ea Domino neque adolebitis ex eis super altare Domini
LEV|22|23|bovem et ovem aure et cauda amputatis voluntarie offerre potes votum autem ex his solvi non potest
LEV|22|24|omne animal quod vel contritis vel tunsis vel sectis ablatisque testiculis est non offeretis Domino et in terra vestra hoc omnino ne faciatis
LEV|22|25|de manu alienigenae non offeretis panes Deo vestro et quicquid aliud dare voluerint quia corrupta et maculata sunt omnia non suscipietis ea
LEV|22|26|locutusque est Dominus ad Mosen dicens
LEV|22|27|bos ovis et capra cum genita fuerint septem diebus erunt sub ubere matris suae die autem octavo et deinceps offerri poterunt Domino
LEV|22|28|sive illa bos sive ovis non immolabuntur una die cum fetibus suis
LEV|22|29|si immolaveritis hostiam pro gratiarum actione Domino ut possit esse placabilis
LEV|22|30|eodem die comedetis eam non remanebit quicquam in mane alterius diei ego Dominus
LEV|22|31|custodite mandata mea et facite ea ego Dominus
LEV|22|32|ne polluatis nomen meum sanctum ut sanctificer in medio filiorum Israhel ego Dominus qui sanctifico vos
LEV|22|33|et eduxi de terra Aegypti ut essem vobis in Deum ego Dominus
LEV|23|1|locutus est Dominus ad Mosen dicens
LEV|23|2|loquere filiis Israhel et dices ad eos hae sunt feriae Domini quas vocabitis sanctas
LEV|23|3|sex diebus facietis opus dies septimus quia sabbati requies est vocabitur sanctus omne opus non facietis in eo sabbatum Domini est in cunctis habitationibus vestris
LEV|23|4|hae sunt ergo feriae Domini sanctae quas celebrare debetis temporibus suis
LEV|23|5|mense primo quartadecima die mensis ad vesperum phase Domini est
LEV|23|6|et quintadecima die mensis huius sollemnitas azymorum Domini est septem diebus azyma comedetis
LEV|23|7|dies primus erit vobis celeberrimus sanctusque omne opus servile non facietis in eo
LEV|23|8|sed offeretis sacrificium in igne Domino septem diebus dies autem septimus erit celebrior et sanctior nullumque servile opus fiet in eo
LEV|23|9|locutusque est Dominus ad Mosen dicens
LEV|23|10|loquere filiis Israhel et dices ad eos cum ingressi fueritis terram quam ego dabo vobis et messueritis segetem feretis manipulos spicarum primitias messis vestrae ad sacerdotem
LEV|23|11|qui elevabit fasciculum coram Domino ut acceptabile sit pro vobis altero die sabbati et sanctificabit illum
LEV|23|12|atque in eodem die quo manipulus consecratur caedetur agnus inmaculatus anniculus in holocaustum Domini
LEV|23|13|et libamenta offerentur cum eo duae decimae similae conspersae oleo in incensum Domini odoremque suavissimum liba quoque vini quarta pars hin
LEV|23|14|panem et pulentam et pultes non comedetis ex segete usque ad diem qua offeratis ex ea Deo vestro praeceptum est sempiternum in generationibus cunctisque habitaculis vestris
LEV|23|15|numerabitis ergo ab altero die sabbati in quo obtulistis manipulum primitiarum septem ebdomadas plenas
LEV|23|16|usque ad alteram diem expletionis ebdomadae septimae id est quinquaginta dies et sic offeretis sacrificium novum Domino
LEV|23|17|ex omnibus habitaculis vestris panes primitiarum duos de duabus decimis similae fermentatae quos coquetis in primitias Domini
LEV|23|18|offeretisque cum panibus septem agnos inmaculatos anniculos et vitulum de armento unum et arietes duos et erunt in holocausto cum libamentis suis in odorem suavissimum Domino
LEV|23|19|facietis et hircum pro peccato duosque agnos anniculos hostias pacificorum
LEV|23|20|cumque elevaverit eos sacerdos cum panibus primitiarum coram Domino cedent in usum eius
LEV|23|21|et vocabitis hunc diem celeberrimum atque sanctissimum omne opus servile non facietis in eo legitimum sempiternum erit in cunctis habitaculis et generationibus vestris
LEV|23|22|postquam autem messueritis segetem terrae vestrae non secabitis eam usque ad solum nec remanentes spicas colligetis sed pauperibus et peregrinis dimittetis eas ego Dominus Deus vester
LEV|23|23|locutusque est Dominus ad Mosen dicens
LEV|23|24|loquere filiis Israhel mense septimo prima die mensis erit vobis sabbatum memorabile clangentibus tubis et vocabitur sanctum
LEV|23|25|omne opus servile non facietis in eo et offeretis holocaustum Domino
LEV|23|26|locutusque est Dominus ad Mosen dicens
LEV|23|27|decimo die mensis huius septimi dies expiationum erit celeberrimus et vocabitur sanctus adfligetisque animas vestras in eo et offeretis holocaustum Domino
LEV|23|28|omne opus non facietis in tempore diei huius quia dies propitiationis est ut propitietur vobis Dominus Deus vester
LEV|23|29|omnis anima quae adflicta non fuerit die hoc peribit de populis suis
LEV|23|30|et quae operis quippiam fecerit delebo eam de populo suo
LEV|23|31|nihil ergo operis facietis in eo legitimum sempiternum erit vobis in cunctis generationibus et habitationibus vestris
LEV|23|32|sabbatum requietionis est adfligetis animas vestras die nono mensis a vespero usque ad vesperum celebrabitis sabbata vestra
LEV|23|33|et locutus est Dominus ad Mosen dicens
LEV|23|34|loquere filiis Israhel a quintodecimo die mensis huius septimi erunt feriae tabernaculorum septem diebus Domino
LEV|23|35|dies primus vocabitur celeberrimus atque sanctissimus omne opus servile non facietis
LEV|23|36|et septem diebus offeretis holocausta Domino dies quoque octavus erit celeberrimus atque sanctissimus et offeretis holocaustum Domino est enim coetus atque collectae omne opus servile non facietis in eo
LEV|23|37|hae sunt feriae Domini quas vocabitis celeberrimas et sanctissimas offeretisque in eis oblationes Domino holocausta et libamenta iuxta ritum uniuscuiusque diei
LEV|23|38|exceptis sabbatis Domini donisque vestris et quae offertis ex voto vel quae sponte tribuitis Domino
LEV|23|39|a quintodecimo ergo die mensis septimi quando congregaveritis omnes fructus terrae vestrae celebrabitis ferias Domini septem diebus die primo et die octavo erit sabbatum id est requies
LEV|23|40|sumetisque vobis die primo fructus arboris pulcherrimae spatulasque palmarum et ramos ligni densarum frondium et salices de torrente et laetabimini coram Domino Deo vestro
LEV|23|41|celebrabitisque sollemnitatem eius septem diebus per annum legitimum sempiternum erit in generationibus vestris mense septimo festa celebrabitis
LEV|23|42|et habitabitis in umbraculis septem diebus omnis qui de genere est Israhel manebit in tabernaculis
LEV|23|43|ut discant posteri vestri quod in tabernaculis habitare fecerim filios Israhel cum educerem eos de terra Aegypti ego Dominus Deus vester
LEV|23|44|locutusque est Moses super sollemnitatibus Domini ad filios Israhel
LEV|24|1|et locutus est Dominus ad Mosen dicens
LEV|24|2|praecipe filiis Israhel ut adferant tibi oleum de olivis purissimum ac lucidum ad concinnandas lucernas iugiter
LEV|24|3|extra velum testimonii in tabernaculo foederis ponetque eas Aaron a vespere usque in mane coram Domino cultu rituque perpetuo in generationibus vestris
LEV|24|4|super candelabro mundissimo ponentur semper in conspectu Domini
LEV|24|5|accipies quoque similam et coques ex ea duodecim panes qui singuli habebunt duas decimas
LEV|24|6|quorum senos altrinsecus super mensam purissimam coram Domino statues
LEV|24|7|et pones super eos tus lucidissimum ut sit panis in monumentum oblationis Domini
LEV|24|8|per singula sabbata mutabuntur coram Domino suscepti a filiis Israhel foedere sempiterno
LEV|24|9|eruntque Aaron et filiorum eius ut comedant eos in loco sancto quia sanctum sanctorum est de sacrificiis Domini iure perpetuo
LEV|24|10|ecce autem egressus filius mulieris israhelitis quem pepererat de viro aegyptio inter filios Israhel iurgatus est in castris cum viro israhelite
LEV|24|11|cumque blasphemasset nomen et maledixisset ei adductus est ad Mosen vocabatur autem mater eius Salumith filia Dabri de tribu Dan
LEV|24|12|miseruntque eum in carcerem donec nossent quid iuberet Dominus
LEV|24|13|qui locutus est ad Mosen
LEV|24|14|dicens educ blasphemum extra castra et ponant omnes qui audierunt manus suas super caput eius et lapidet eum populus universus
LEV|24|15|et ad filios Israhel loqueris homo qui maledixerit Deo suo portabit peccatum suum
LEV|24|16|et qui blasphemaverit nomen Domini morte moriatur lapidibus opprimet eum omnis multitudo sive ille civis seu peregrinus fuerit qui blasphemaverit nomen Domini morte moriatur
LEV|24|17|qui percusserit et occiderit hominem morte moriatur
LEV|24|18|qui percusserit animal reddat vicarium id est animam pro anima
LEV|24|19|qui inrogaverit maculam cuilibet civium suorum sicut fecit fiet ei
LEV|24|20|fracturam pro fractura oculum pro oculo dentem pro dente restituet qualem inflixerit maculam talem sustinere cogetur
LEV|24|21|qui percusserit iumentum reddet aliud qui percusserit hominem punietur
LEV|24|22|aequum iudicium sit inter vos sive peregrinus sive civis peccaverit quia ego sum Dominus Deus vester
LEV|24|23|locutusque est Moses ad filios Israhel et eduxerunt eum qui blasphemaverat extra castra ac lapidibus oppresserunt feceruntque filii Israhel sicut praeceperat Dominus Mosi
LEV|25|1|locutusque est Dominus ad Mosen in monte Sinai dicens
LEV|25|2|loquere filiis Israhel et dices ad eos quando ingressi fueritis terram quam ego dabo vobis sabbatizet sabbatum Domini
LEV|25|3|sex annis seres agrum tuum et sex annis putabis vineam tuam colligesque fructus eius
LEV|25|4|septimo autem anno sabbatum erit terrae requietionis Domini agrum non seres et vineam non putabis
LEV|25|5|quae sponte gignit humus non metes et uvas primitiarum tuarum non colliges quasi vindemiam annus enim requietionis terrae est
LEV|25|6|sed erunt vobis in cibum tibi et servo tuo ancillae et mercennario tuo et advenae qui peregrinantur apud te
LEV|25|7|iumentis tuis et pecoribus omnia quae nascuntur praebebunt cibum
LEV|25|8|numerabis quoque tibi septem ebdomades annorum id est septem septies quae simul faciunt annos quadraginta novem
LEV|25|9|et clanges bucina mense septimo decima die mensis propitiationis tempore in universa terra vestra
LEV|25|10|sanctificabisque annum quinquagesimum et vocabis remissionem cunctis habitatoribus terrae tuae ipse est enim iobeleus revertetur homo ad possessionem suam et unusquisque rediet ad familiam pristinam
LEV|25|11|quia iobeleus est et quinquagesimus annus non seretis neque metetis sponte in agro nascentia et primitias vindemiae non colligetis
LEV|25|12|ob sanctificationem iobelei sed statim ablata comedetis
LEV|25|13|anno iobelei redient omnes ad possessiones suas
LEV|25|14|quando vendes quippiam civi tuo vel emes ab eo ne contristes fratrem tuum sed iuxta numerum annorum iobelei emes ab eo
LEV|25|15|et iuxta supputationem frugum vendet tibi
LEV|25|16|quanto plus anni remanserint post iobeleum tanto crescet et pretium et quanto minus temporis numeraveris tanto minoris et emptio constabit tempus enim frugum vendet tibi
LEV|25|17|nolite adfligere contribules vestros sed timeat unusquisque Deum suum quia ego Dominus Deus vester
LEV|25|18|facite praecepta mea et iudicia custodite et implete ea ut habitare possitis in terra absque ullo pavore
LEV|25|19|et gignat vobis humus fructus suos quibus vescamini usque ad saturitatem nullius impetum formidantes
LEV|25|20|quod si dixeritis quid comedemus anno septimo si non seruerimus neque collegerimus fruges nostras
LEV|25|21|dabo benedictionem meam vobis anno sexto et faciet fructus trium annorum
LEV|25|22|seretisque anno octavo et comedetis veteres fruges usque ad nonum annum donec nova nascantur edetis vetera
LEV|25|23|terra quoque non veniet in perpetuum quia mea est et vos advenae et coloni mei estis
LEV|25|24|unde cuncta regio possessionis vestrae sub redemptionis condicione vendetur
LEV|25|25|si adtenuatus frater tuus vendiderit possessiunculam suam et voluerit propinquus eius potest redimere quod ille vendiderat
LEV|25|26|sin autem non habuerit proximum et ipse pretium ad redimendum potuerit invenire
LEV|25|27|conputabuntur fructus ex eo tempore quo vendidit et quod reliquum est reddet emptori sicque recipiet possessionem suam
LEV|25|28|quod si non invenerit manus eius ut reddat pretium habebit emptor quod emerat usque ad annum iobeleum in ipso enim omnis venditio redit ad dominum et ad possessorem pristinum
LEV|25|29|qui vendiderit domum intra urbis muros habebit licentiam redimendi donec unus impleatur annus
LEV|25|30|si non redemerit et anni circulus fuerit evolutus emptor possidebit eam et posteri eius in perpetuum et redimi non poterit etiam in iobeleo
LEV|25|31|sin autem in villa fuerit domus quae muros non habet agrorum iure vendetur si ante redempta non fuerit in iobeleo revertetur ad dominum
LEV|25|32|aedes Levitarum quae in urbibus sunt semper possunt redimi
LEV|25|33|si redemptae non fuerint in iobeleo revertentur ad dominos quia domus urbium leviticarum pro possessionibus sunt inter filios Israhel
LEV|25|34|suburbana autem eorum non venient quia possessio sempiterna est
LEV|25|35|si adtenuatus fuerit frater tuus et infirmus manu et susceperis eum quasi advenam et peregrinum et vixerit tecum
LEV|25|36|ne accipias usuras ab eo nec amplius quam dedisti time Deum tuum ut vivere possit frater tuus apud te
LEV|25|37|pecuniam tuam non dabis ei ad usuram et frugum superabundantiam non exiges
LEV|25|38|ego Dominus Deus vester qui eduxi vos de terra Aegypti ut darem vobis terram Chanaan et essem vester Deus
LEV|25|39|si paupertate conpulsus vendiderit se tibi frater tuus non eum opprimes servitute famulorum
LEV|25|40|sed quasi mercennarius et colonus erit usque ad annum iobeleum operabitur apud te
LEV|25|41|et postea egredietur cum liberis suis et revertetur ad cognationem et ad possessionem patrum suorum
LEV|25|42|mei enim servi sunt et ego eduxi eos de terra Aegypti non venient condicione servorum
LEV|25|43|ne adfligas eum per potentiam sed metuito Deum tuum
LEV|25|44|servus et ancilla sint vobis de nationibus quae in circuitu vestro sunt
LEV|25|45|et de advenis qui peregrinantur apud vos vel qui ex his nati fuerint in terra vestra hos habebitis famulos
LEV|25|46|et hereditario iure transmittetis ad posteros ac possidebitis in aeternum fratres autem vestros filios Israhel ne opprimatis per potentiam
LEV|25|47|si invaluerit apud vos manus advenae atque peregrini et adtenuatus frater tuus vendiderit se ei aut cuiquam de stirpe eius
LEV|25|48|post venditionem potest redimi qui voluerit ex fratribus suis redimet eum
LEV|25|49|et patruus et patruelis et consanguineus et adfinis sin autem et ipse potuerit redimet se
LEV|25|50|supputatis dumtaxat annis a tempore venditionis suae usque ad annum iobeleum et pecunia qua venditus fuerat iuxta annorum numerum et rationem mercennarii supputata
LEV|25|51|si plures fuerint anni qui remanent usque ad iobeleum secundum hos reddet et pretium
LEV|25|52|si pauci ponet rationem cum eo iuxta annorum numerum et reddet emptori quod reliquum est annorum
LEV|25|53|quibus ante servivit mercedibus inputatis non adfliget eum violenter in conspectu tuo
LEV|25|54|quod si per haec redimi non potuerit anno iobeleo egredietur cum liberis suis
LEV|25|55|mei sunt enim servi filii Israhel quos eduxi de terra Aegypti
LEV|26|1|ego Dominus Deus vester non facietis vobis idolum et sculptile nec titulos erigetis nec insignem lapidem ponetis in terra vestra ut adoretis eum ego enim sum Dominus Deus vester
LEV|26|2|custodite sabbata mea et pavete ad sanctuarium meum ego Dominus
LEV|26|3|si in praeceptis meis ambulaveritis et mandata mea custodieritis et feceritis ea dabo vobis pluvias temporibus suis
LEV|26|4|et terra gignet germen suum et pomis arbores replebuntur
LEV|26|5|adprehendet messium tritura vindemiam et vindemia occupabit sementem et comedetis panem vestrum in saturitatem et absque pavore habitabitis in terra vestra
LEV|26|6|dabo pacem in finibus vestris dormietis et non erit qui exterreat auferam malas bestias et gladius non transibit terminos vestros
LEV|26|7|persequemini inimicos vestros et corruent coram vobis
LEV|26|8|persequentur quinque de vestris centum alienos et centum ex vobis decem milia cadent inimici vestri in conspectu vestro gladio
LEV|26|9|respiciam vos et crescere faciam multiplicabimini et firmabo pactum meum vobiscum
LEV|26|10|comedetis vetustissima veterum et vetera novis supervenientibus proicietis
LEV|26|11|ponam tabernaculum meum in medio vestri et non abiciet vos anima mea
LEV|26|12|ambulabo inter vos et ero vester Deus vosque eritis populus meus
LEV|26|13|ego Dominus Deus vester qui eduxi vos de terra Aegyptiorum ne serviretis eis et qui confregi catenas cervicum vestrarum ut incederetis erecti
LEV|26|14|quod si non audieritis me nec feceritis omnia mandata mea
LEV|26|15|si spreveritis leges meas et iudicia mea contempseritis ut non faciatis ea quae a me constituta sunt et ad irritum perducatis pactum meum
LEV|26|16|ego quoque haec faciam vobis visitabo vos velociter in egestate et ardore qui conficiat oculos vestros et consumat animas frustra seretis sementem quae ab hostibus devorabitur
LEV|26|17|ponam faciem meam contra vos et corruetis coram hostibus vestris et subiciemini his qui oderunt vos fugietis nemine persequente
LEV|26|18|sin autem nec sic oboedieritis mihi addam correptiones vestras septuplum propter peccata vestra
LEV|26|19|et conteram superbiam duritiae vestrae daboque caelum vobis desuper sicut ferrum et terram aeneam
LEV|26|20|consumetur in cassum labor vester non proferet terra germen nec arbores poma praebebunt
LEV|26|21|si ambulaveritis ex adverso mihi nec volueritis audire me addam plagas vestras usque in septuplum propter peccata vestra
LEV|26|22|emittamque in vos bestias agri quae consumant et vos et pecora vestra et ad paucitatem cuncta redigant desertaeque fiant viae vestrae
LEV|26|23|quod si nec sic volueritis recipere disciplinam sed ambulaveritis ex adverso mihi
LEV|26|24|ego quoque contra vos adversus incedam et percutiam vos septies propter peccata vestra
LEV|26|25|inducamque super vos gladium ultorem foederis mei cumque confugeritis in urbes mittam pestilentiam in medio vestri et trademini hostium manibus
LEV|26|26|postquam confregero baculum panis vestri ita ut decem mulieres in uno clibano coquant panes et reddant eos ad pondus et comedetis et non saturabimini
LEV|26|27|sin autem nec per haec audieritis me sed ambulaveritis contra me
LEV|26|28|et ego incedam adversum vos in furore contrario et corripiam vos septem plagis propter peccata vestra
LEV|26|29|ita ut comedatis carnes filiorum et filiarum vestrarum
LEV|26|30|destruam excelsa vestra et simulacra confringam cadetis inter ruinas idolorum vestrorum et abominabitur vos anima mea
LEV|26|31|in tantum ut urbes vestras redigam in solitudinem et deserta faciam sanctuaria vestra nec recipiam ultra odorem suavissimum
LEV|26|32|disperdamque terram vestram et stupebunt super ea inimici vestri cum habitatores illius fuerint
LEV|26|33|vos autem dispergam in gentes et evaginabo post vos gladium eritque terra vestra deserta et civitates dirutae
LEV|26|34|tunc placebunt terrae sabbata sua cunctis diebus solitudinis suae quando fueritis
LEV|26|35|in terra hostili sabbatizabit et requiescet in sabbatis solitudinis suae eo quod non requieverit in sabbatis vestris quando habitabatis in ea
LEV|26|36|et qui de vobis remanserint dabo pavorem in cordibus eorum in regionibus hostium terrebit eos sonitus folii volantis et ita fugient quasi gladium cadent nullo sequente
LEV|26|37|et corruent singuli super fratres suos quasi bella fugientes nemo vestrum inimicis audebit resistere
LEV|26|38|peribitis inter gentes et hostilis vos terra consumet
LEV|26|39|quod si et de his aliqui remanserint tabescent in iniquitatibus suis in terra inimicorum suorum et propter peccata patrum suorum et sua adfligentur
LEV|26|40|donec confiteantur iniquitates suas et maiorum suorum quibus praevaricati sunt in me et ambulaverunt ex adverso mihi
LEV|26|41|ambulabo igitur et ego contra eos et inducam illos in terram hostilem donec erubescat incircumcisa mens eorum tunc orabunt pro impietatibus suis
LEV|26|42|et recordabor foederis mei quod pepigi cum Iacob et Isaac et Abraham terrae quoque memor ero
LEV|26|43|quae cum relicta fuerit ab eis conplacebit sibi in sabbatis suis patiens solitudinem propter illos ipsi vero rogabunt pro peccatis suis eo quod abiecerint iudicia mea et leges meas despexerint
LEV|26|44|et tamen etiam cum essent in terra hostili non penitus abieci eos neque sic despexi ut consumerentur et irritum facerem pactum meum cum eis ego enim sum Dominus Deus eorum
LEV|26|45|et recordabor foederis mei pristini quando eduxi eos de terra Aegypti in conspectu gentium ut essem Deus eorum ego Dominus Deus haec sunt praecepta atque iudicia et leges quas dedit Dominus inter se et inter filios Israhel in monte Sinai per manum Mosi
LEV|26|46|
LEV|27|1|locutusque est Dominus ad Mosen dicens
LEV|27|2|loquere filiis Israhel et dices ad eos homo qui votum fecerit et spoponderit Deo animam suam sub aestimatione dabit pretium
LEV|27|3|si fuerit masculus a vicesimo usque ad sexagesimum annum dabit quinquaginta siclos argenti ad mensuram sanctuarii
LEV|27|4|si mulier triginta
LEV|27|5|a quinto autem anno usque ad vicesimum masculus dabit viginti siclos femina decem
LEV|27|6|ab uno mense usque ad annum quintum pro masculo dabuntur quinque sicli pro femina tres
LEV|27|7|sexagenarius et ultra masculus dabit quindecim siclos femina decem
LEV|27|8|si pauper fuerit et aestimationem reddere non valebit stabit coram sacerdote et quantum ille aestimaverit et viderit eum posse reddere tantum dabit
LEV|27|9|animal autem quod immolari potest Domino si quis voverit sanctum erit
LEV|27|10|et mutari non poterit id est nec melius malo nec peius bono quod si mutaverit et ipsum quod mutatum est et illud pro quo mutatum est consecratum erit Domino
LEV|27|11|animal inmundum quod immolari Domino non potest si quis voverit adducetur ante sacerdotem
LEV|27|12|qui diiudicans utrum bonum an malum sit statuet pretium
LEV|27|13|quod si dare voluerit is qui offert addet supra aestimationis quintam partem
LEV|27|14|homo si voverit domum suam et sanctificaverit Domino considerabit eam sacerdos utrum bona an mala sit et iuxta pretium quod ab eo fuerit constitutum venundabitur
LEV|27|15|sin autem ille qui voverat voluerit redimere eam dabit quintam partem aestimationis supra et habebit domum
LEV|27|16|quod si agrum possessionis suae voverit et consecraverit Domino iuxta mensuram sementis aestimabitur pretium si triginta modiis hordei seritur terra quinquaginta siclis veniet argenti
LEV|27|17|si statim ab anno incipientis iobelei voverit agrum quanto valere potest tanto aestimabitur
LEV|27|18|sin autem post aliquantum temporis supputabit sacerdos pecuniam iuxta annorum qui reliqui sunt numerum usque ad iobeleum et detrahetur ex pretio
LEV|27|19|quod si voluerit redimere agrum ille qui voverat addet quintam partem aestimatae pecuniae et possidebit eum
LEV|27|20|sin autem noluerit redimere sed alteri cuilibet fuerit venundatus ultra eum qui voverat redimere non poterit
LEV|27|21|quia cum iobelei venerit dies sanctificatus erit Domino et possessio consecrata ad ius pertinet sacerdotum
LEV|27|22|si ager emptus et non de possessione maiorum sanctificatus fuerit Domino
LEV|27|23|supputabit sacerdos iuxta annorum numerum usque ad iobeleum pretium et dabit ille qui voverat eum Domino
LEV|27|24|in iobeleo autem revertetur ad priorem dominum qui vendiderat eum et habuerat in sortem possessionis suae
LEV|27|25|omnis aestimatio siclo sanctuarii ponderabitur siclus viginti obolos habet
LEV|27|26|primogenita quae ad Dominum pertinent nemo sanctificare poterit et vovere sive bos sive ovis fuerit Domini sunt
LEV|27|27|quod si inmundum est animal redimet qui obtulit iuxta aestimationem tuam et addet quintam partem pretii si redimere noluerit vendetur alteri quantocumque a te fuerit aestimatum
LEV|27|28|omne quod Domino consecratur sive homo fuerit sive animal sive ager non veniet nec redimi poterit quicquid semel fuerit consecratum sanctum sanctorum erit Domino
LEV|27|29|et omnis consecratio quae offertur ab homine non redimetur sed morte morietur
LEV|27|30|omnes decimae terrae sive de frugibus sive de pomis arborum Domini sunt et illi sanctificantur
LEV|27|31|si quis autem voluerit redimere decimas suas addet quintam partem earum
LEV|27|32|omnium decimarum boves et oves et caprae quae sub pastoris virga transeunt quicquid decimum venerit sanctificabitur Domino
LEV|27|33|non eligetur nec bonum nec malum nec altero commutabitur si quis mutaverit et quod mutatum est et pro quo mutatum est sanctificabitur Domino et non redimetur
LEV|27|34|haec sunt praecepta quae mandavit Dominus Mosi ad filios Israhel in monte Sinai
