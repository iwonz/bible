REV|1|1|apocalypsis Iesu Christi quam dedit illi Deus palam facere servis suis quae oportet fieri cito et significavit mittens per angelum suum servo suo Iohanni
REV|1|2|qui testimonium perhibuit verbo Dei et testimonium Iesu Christi quaecumque vidit
REV|1|3|beatus qui legit et qui audiunt verba prophetiae et servant ea quae in ea scripta sunt tempus enim prope est
REV|1|4|Iohannes septem ecclesiis quae sunt in Asia gratia vobis et pax ab eo qui est et qui erat et qui venturus est et a septem spiritibus qui in conspectu throni eius sunt
REV|1|5|et ab Iesu Christo qui est testis fidelis primogenitus mortuorum et princeps regum terrae qui dilexit nos et lavit nos a peccatis nostris in sanguine suo
REV|1|6|et fecit nostrum regnum sacerdotes Deo et Patri suo ipsi gloria et imperium in saecula saeculorum amen
REV|1|7|ecce venit cum nubibus et videbit eum omnis oculus et qui eum pupugerunt et plangent se super eum omnes tribus terrae etiam amen
REV|1|8|ego sum Alpha et Omega principium et finis dicit Dominus Deus qui est et qui erat et qui venturus est Omnipotens
REV|1|9|ego Iohannes frater vester et particeps in tribulatione et regno et patientia in Iesu fui in insula quae appellatur Patmos propter verbum Dei et testimonium Iesu
REV|1|10|fui in spiritu in dominica die et audivi post me vocem magnam tamquam tubae
REV|1|11|dicentis quod vides scribe in libro et mitte septem ecclesiis Ephesum et Zmyrnam et Pergamum et Thyatiram et Sardis et Philadelphiam et Laodiciam
REV|1|12|et conversus sum ut viderem vocem quae loquebatur mecum et conversus vidi septem candelabra aurea
REV|1|13|et in medio septem candelabrorum similem Filio hominis vestitum podere et praecinctum ad mamillas zonam auream
REV|1|14|caput autem eius et capilli erant candidi tamquam lana alba tamquam nix et oculi eius velut flamma ignis
REV|1|15|et pedes eius similes orichalco sicut in camino ardenti et vox illius tamquam vox aquarum multarum
REV|1|16|et habebat in dextera sua stellas septem et de ore eius gladius utraque parte acutus exiebat et facies eius sicut sol lucet in virtute sua
REV|1|17|et cum vidissem eum cecidi ad pedes eius tamquam mortuus et posuit dexteram suam super me dicens noli timere ego sum primus et novissimus
REV|1|18|et vivus et fui mortuus et ecce sum vivens in saecula saeculorum et habeo claves mortis et inferni
REV|1|19|scribe ergo quae vidisti et quae sunt et quae oportet fieri post haec
REV|1|20|sacramentum septem stellarum quas vidisti in dextera mea et septem candelabra aurea septem stellae angeli sunt septem ecclesiarum et candelabra septem septem ecclesiae sunt
REV|2|1|angelo Ephesi ecclesiae scribe haec dicit qui tenet septem stellas in dextera sua qui ambulat in medio septem candelabrorum aureorum
REV|2|2|scio opera tua et laborem et patientiam tuam et quia non potes sustinere malos et temptasti eos qui se dicunt apostolos et non sunt et invenisti eos mendaces
REV|2|3|et patientiam habes et sustinuisti propter nomen meum et non defecisti
REV|2|4|sed habeo adversus te quod caritatem tuam primam reliquisti
REV|2|5|memor esto itaque unde excideris et age paenitentiam et prima opera fac sin autem venio tibi et movebo candelabrum tuum de loco suo nisi paenitentiam egeris
REV|2|6|sed hoc habes quia odisti facta Nicolaitarum quae et ego odi
REV|2|7|qui habet aurem audiat quid Spiritus dicat ecclesiis vincenti dabo ei edere de ligno vitae quod est in paradiso Dei mei
REV|2|8|et angelo Zmyrnae ecclesiae scribe haec dicit primus et novissimus qui fuit mortuus et vivit
REV|2|9|scio tribulationem tuam et paupertatem tuam sed dives es et blasphemaris ab his qui se dicunt Iudaeos esse et non sunt sed sunt synagoga Satanae
REV|2|10|nihil horum timeas quae passurus es ecce missurus est diabolus ex vobis in carcerem ut temptemini et habebitis tribulationem diebus decem esto fidelis usque ad mortem et dabo tibi coronam vitae
REV|2|11|qui habet aurem audiat quid Spiritus dicat ecclesiis qui vicerit non laedetur a morte secunda
REV|2|12|et angelo Pergami ecclesiae scribe haec dicit qui habet rompheam utraque parte acutam
REV|2|13|scio ubi habitas ubi sedes est Satanae et tenes nomen meum et non negasti fidem meam et in diebus Antipas testis meus fidelis qui occisus est apud vos ubi Satanas habitat
REV|2|14|sed habeo adversus te pauca quia habes illic tenentes doctrinam Balaam qui docebat Balac mittere scandalum coram filiis Israhel edere et fornicari
REV|2|15|ita habes et tu tenentes doctrinam Nicolaitarum
REV|2|16|similiter paenitentiam age si quo minus venio tibi cito et pugnabo cum illis in gladio oris mei
REV|2|17|qui habet aurem audiat quid Spiritus dicat ecclesiis vincenti dabo ei manna absconditum et dabo illi calculum candidum et in calculo nomen novum scriptum quod nemo scit nisi qui accipit
REV|2|18|et angelo Thyatirae ecclesiae scribe haec dicit Filius Dei qui habet oculos ut flammam ignis et pedes eius similes orichalco
REV|2|19|novi opera tua et caritatem et fidem et ministerium et patientiam tuam et opera tua novissima plura prioribus
REV|2|20|sed habeo adversus te quia permittis mulierem Hiezabel quae se dicit propheten docere et seducere servos meos fornicari et manducare de idolothytis
REV|2|21|et dedi illi tempus ut paenitentiam ageret et non vult paeniteri a fornicatione sua
REV|2|22|ecce mitto eam in lectum et qui moechantur cum ea in tribulationem maximam nisi paenitentiam egerint ab operibus eius
REV|2|23|et filios eius interficiam in morte et scient omnes ecclesiae quia ego sum scrutans renes et corda et dabo unicuique vestrum secundum opera vestra
REV|2|24|vobis autem dico ceteris qui Thyatirae estis quicumque non habent doctrinam hanc qui non cognoverunt altitudines Satanae quemadmodum dicunt non mittam super vos aliud pondus
REV|2|25|tamen id quod habetis tenete donec veniam
REV|2|26|et qui vicerit et qui custodierit usque in finem opera mea dabo illi potestatem super gentes
REV|2|27|et reget illas in virga ferrea tamquam vas figuli confringentur
REV|2|28|sicut et ego accepi a Patre meo et dabo illi stellam matutinam
REV|2|29|qui habet aurem audiat quid Spiritus dicat ecclesiis
REV|3|1|et angelo ecclesiae Sardis scribe haec dicit qui habet septem spiritus Dei et septem stellas scio opera tua quia nomen habes quod vivas et mortuus es
REV|3|2|esto vigilans et confirma cetera quae moritura erant non enim invenio opera tua plena coram Deo meo
REV|3|3|in mente ergo habe qualiter acceperis et audieris et serva et paenitentiam age si ergo non vigilaveris veniam tamquam fur et nescies qua hora veniam ad te
REV|3|4|sed habes pauca nomina in Sardis qui non inquinaverunt vestimenta sua et ambulabunt mecum in albis quia digni sunt
REV|3|5|qui vicerit sic vestietur vestimentis albis et non delebo nomen eius de libro vitae et confitebor nomen eius coram Patre meo et coram angelis eius
REV|3|6|qui habet aurem audiat quid Spiritus dicat ecclesiis
REV|3|7|et angelo Philadelphiae ecclesiae scribe haec dicit sanctus et verus qui habet clavem David qui aperit et nemo cludit et cludit et nemo aperit
REV|3|8|scio opera tua ecce dedi coram te ostium apertum quod nemo potest cludere quia modicam habes virtutem et servasti verbum meum et non negasti nomen meum
REV|3|9|ecce dabo de synagoga Satanae qui dicunt se Iudaeos esse et non sunt sed mentiuntur ecce faciam illos ut veniant et adorent ante pedes tuos et scient quia ego dilexi te
REV|3|10|quoniam servasti verbum patientiae meae et ego te servabo ab hora temptationis quae ventura est in orbem universum temptare habitantes in terra
REV|3|11|venio cito tene quod habes ut nemo accipiat coronam tuam
REV|3|12|qui vicerit faciam illum columnam in templo Dei mei et foras non egredietur amplius et scribam super eum nomen Dei mei et nomen civitatis Dei mei novae Hierusalem quae descendit de caelo a Deo meo et nomen meum novum
REV|3|13|qui habet aurem audiat quid Spiritus dicat ecclesiis
REV|3|14|et angelo Laodiciae ecclesiae scribe haec dicit Amen testis fidelis et verus qui est principium creaturae Dei
REV|3|15|scio opera tua quia neque frigidus es neque calidus utinam frigidus esses aut calidus
REV|3|16|sed quia tepidus es et nec frigidus nec calidus incipiam te evomere ex ore meo
REV|3|17|quia dicis quod dives sum et locupletatus et nullius egeo et nescis quia tu es miser et miserabilis et pauper et caecus et nudus
REV|3|18|suadeo tibi emere a me aurum ignitum probatum ut locuples fias et vestimentis albis induaris et non appareat confusio nuditatis tuae et collyrio inungue oculos tuos ut videas
REV|3|19|ego quos amo arguo et castigo aemulare ergo et paenitentiam age
REV|3|20|ecce sto ad ostium et pulso si quis audierit vocem meam et aperuerit ianuam introibo ad illum et cenabo cum illo et ipse mecum
REV|3|21|qui vicerit dabo ei sedere mecum in throno meo sicut et ego vici et sedi cum Patre meo in throno eius
REV|3|22|qui habet aurem audiat quid Spiritus dicat ecclesiis
REV|4|1|post haec vidi et ecce ostium apertum in caelo et vox prima quam audivi tamquam tubae loquentis mecum dicens ascende huc et ostendam tibi quae oportet fieri post haec
REV|4|2|statim fui in spiritu et ecce sedis posita erat in caelo et supra sedem sedens
REV|4|3|et qui sedebat similis erat aspectui lapidis iaspidis et sardini et iris erat in circuitu sedis similis visioni zmaragdinae
REV|4|4|et in circuitu sedis sedilia viginti quattuor et super thronos viginti quattuor seniores sedentes circumamictos vestimentis albis et in capitibus eorum coronas aureas
REV|4|5|et de throno procedunt fulgura et voces et tonitrua et septem lampades ardentes ante thronum quae sunt septem spiritus Dei
REV|4|6|et in conspectu sedis tamquam mare vitreum simile cristallo et in medio sedis et in circuitu sedis quattuor animalia plena oculis ante et retro
REV|4|7|et animal primum simile leoni et secundum animal simile vitulo et tertium animal habens faciem quasi hominis et quartum animal simile aquilae volanti
REV|4|8|et quattuor animalia singula eorum habebant alas senas et in circuitu et intus plena sunt oculis et requiem non habent die et nocte dicentia sanctus sanctus sanctus Dominus Deus omnipotens qui erat et qui est et qui venturus est
REV|4|9|et cum darent illa animalia gloriam et honorem et benedictionem sedenti super thronum viventi in saecula saeculorum
REV|4|10|procident viginti quattuor seniores ante sedentem in throno et adorabunt viventem in saecula saeculorum et mittent coronas suas ante thronum dicentes
REV|4|11|dignus es Domine et Deus noster accipere gloriam et honorem et virtutem quia tu creasti omnia et propter voluntatem tuam erant et creata sunt
REV|5|1|et vidi in dextera sedentis super thronum librum scriptum intus et foris signatum sigillis septem
REV|5|2|et vidi angelum fortem praedicantem voce magna quis est dignus aperire librum et solvere signacula eius
REV|5|3|et nemo poterat in caelo neque in terra neque subtus terram aperire librum neque respicere illum
REV|5|4|et ego flebam multum quoniam nemo dignus inventus est aperire librum nec videre eum
REV|5|5|et unus de senioribus dicit mihi ne fleveris ecce vicit leo de tribu Iuda radix David aperire librum et septem signacula eius
REV|5|6|et vidi et ecce in medio throni et quattuor animalium et in medio seniorum agnum stantem tamquam occisum habentem cornua septem et oculos septem qui sunt spiritus Dei missi in omnem terram
REV|5|7|et venit et accepit de dextera sedentis de throno
REV|5|8|et cum aperuisset librum quattuor animalia et viginti quattuor seniores ceciderunt coram agno habentes singuli citharas et fialas aureas plenas odoramentorum quae sunt orationes sanctorum
REV|5|9|et cantant novum canticum dicentes dignus es accipere librum et aperire signacula eius quoniam occisus es et redemisti nos Deo in sanguine tuo ex omni tribu et lingua et populo et natione
REV|5|10|et fecisti eos Deo nostro regnum et sacerdotes et regnabunt super terram
REV|5|11|et vidi et audivi vocem angelorum multorum in circuitu throni et animalium et seniorum et erat numerus eorum milia milium
REV|5|12|dicentium voce magna dignus est agnus qui occisus est accipere virtutem et divinitatem et sapientiam et fortitudinem et honorem et gloriam et benedictionem
REV|5|13|et omnem creaturam quae in caelo est et super terram et sub terram et quae sunt in mari et quae in ea omnes audivi dicentes sedenti in throno et agno benedictio et honor et gloria et potestas in saecula saeculorum
REV|5|14|et quattuor animalia dicebant amen et seniores ceciderunt et adoraverunt
REV|6|1|et vidi quod aperuisset agnus unum de septem signaculis et audivi unum de quattuor animalibus dicentem tamquam vocem tonitrui veni
REV|6|2|et vidi et ecce equus albus et qui sedebat super illum habebat arcum et data est ei corona et exivit vincens ut vinceret
REV|6|3|et cum aperuisset sigillum secundum audivi secundum animal dicens veni
REV|6|4|et exivit alius equus rufus et qui sedebat super illum datum est ei ut sumeret pacem de terra et ut invicem se interficiant et datus est illi gladius magnus
REV|6|5|et cum aperuisset sigillum tertium audivi tertium animal dicens veni et vidi et ecce equus niger et qui sedebat super eum habebat stateram in manu sua
REV|6|6|et audivi tamquam vocem in medio quattuor animalium dicentem bilibris tritici denario et tres bilibres hordei denario et vinum et oleum ne laeseris
REV|6|7|et cum aperuisset sigillum quartum audivi vocem quarti animalis dicentis veni et vidi
REV|6|8|et ecce equus pallidus et qui sedebat desuper nomen illi Mors et inferus sequebatur eum et data est illi potestas super quattuor partes terrae interficere gladio fame et morte et bestiis terrae
REV|6|9|et cum aperuisset quintum sigillum vidi subtus altare animas interfectorum propter verbum Dei et propter testimonium quod habebant
REV|6|10|et clamabant voce magna dicentes usquequo Domine sanctus et verus non iudicas et vindicas sanguinem nostrum de his qui habitant in terra
REV|6|11|et datae sunt illis singulae stolae albae et dictum est illis ut requiescerent tempus adhuc modicum donec impleantur conservi eorum et fratres eorum qui interficiendi sunt sicut et illi
REV|6|12|et vidi cum aperuisset sigillum sextum et terraemotus factus est magnus et sol factus est niger tamquam saccus cilicinus et luna tota facta est sicut sanguis
REV|6|13|et stellae caeli ceciderunt super terram sicut ficus mittit grossos suos cum vento magno movetur
REV|6|14|et caelum recessit sicut liber involutus et omnis mons et insulae de locis suis motae sunt
REV|6|15|et reges terrae et principes et tribuni et divites et fortes et omnis servus et liber absconderunt se in speluncis et petris montium
REV|6|16|et dicunt montibus et petris cadite super nos et abscondite nos a facie sedentis super thronum et ab ira agni
REV|6|17|quoniam venit dies magnus irae ipsorum et quis poterit stare
REV|7|1|post haec vidi quattuor angelos stantes super quattuor angulos terrae tenentes quattuor ventos terrae ne flaret ventus super terram neque super mare neque in ullam arborem
REV|7|2|et vidi alterum angelum ascendentem ab ortu solis habentem signum Dei vivi et clamavit voce magna quattuor angelis quibus datum est nocere terrae et mari
REV|7|3|dicens nolite nocere terrae neque mari neque arboribus quoadusque signemus servos Dei nostri in frontibus eorum
REV|7|4|et audivi numerum signatorum centum quadraginta quattuor milia signati ex omni tribu filiorum Israhel
REV|7|5|ex tribu Iuda duodecim milia signati ex tribu Ruben duodecim milia ex tribu Gad duodecim milia
REV|7|6|ex tribu Aser duodecim milia ex tribu Nepthalim duodecim milia ex tribu Manasse duodecim milia
REV|7|7|ex tribu Symeon duodecim milia ex tribu Levi duodecim milia ex tribu Issachar duodecim milia
REV|7|8|ex tribu Zabulon duodecim milia ex tribu Ioseph duodecim milia ex tribu Beniamin duodecim milia signati
REV|7|9|post haec vidi turbam magnam quam dinumerare nemo poterat ex omnibus gentibus et tribubus et populis et linguis stantes ante thronum et in conspectu agni amicti stolas albas et palmae in manibus eorum
REV|7|10|et clamabant voce magna dicentes salus Deo nostro qui sedet super thronum et agno
REV|7|11|et omnes angeli stabant in circuitu throni et seniorum et quattuor animalium et ceciderunt in conspectu throni in facies suas et adoraverunt Deum
REV|7|12|dicentes amen benedictio et claritas et sapientia et gratiarum actio et honor et virtus et fortitudo Deo nostro in saecula saeculorum amen
REV|7|13|et respondit unus de senioribus dicens mihi hii qui amicti sunt stolis albis qui sunt et unde venerunt
REV|7|14|et dixi illi domine mi tu scis et dixit mihi hii sunt qui veniunt de tribulatione magna et laverunt stolas suas et dealbaverunt eas in sanguine agni
REV|7|15|ideo sunt ante thronum Dei et serviunt ei die ac nocte in templo eius et qui sedet in throno habitabit super illos
REV|7|16|non esurient neque sitient amplius neque cadet super illos sol neque ullus aestus
REV|7|17|quoniam agnus qui in medio throni est reget illos et deducet eos ad vitae fontes aquarum et absterget Deus omnem lacrimam ex oculis eorum
REV|8|1|et cum aperuisset sigillum septimum factum est silentium in caelo quasi media hora
REV|8|2|et vidi septem angelos stantes in conspectu Dei et datae sunt illis septem tubae
REV|8|3|et alius angelus venit et stetit ante altare habens turibulum aureum et data sunt illi incensa multa ut daret orationibus sanctorum omnium super altare aureum quod est ante thronum
REV|8|4|et ascendit fumus incensorum de orationibus sanctorum de manu angeli coram Deo
REV|8|5|et accepit angelus turibulum et implevit illud de igne altaris et misit in terram et facta sunt tonitrua et voces et fulgora et terraemotus
REV|8|6|et septem angeli qui habebant septem tubas paraverunt se ut tuba canerent
REV|8|7|et primus tuba cecinit et facta est grando et ignis mixta in sanguine et missum est in terram et tertia pars terrae conbusta est et tertia pars arborum conbusta est et omne faenum viride conbustum est
REV|8|8|et secundus angelus tuba cecinit et tamquam mons magnus igne ardens missus est in mare et facta est tertia pars maris sanguis
REV|8|9|et mortua est tertia pars creaturae quae habent animas et tertia pars navium interiit
REV|8|10|et tertius angelus tuba cecinit et cecidit de caelo stella magna ardens tamquam facula et cecidit in tertiam partem fluminum et in fontes aquarum
REV|8|11|et nomen stellae dicitur Absinthius et facta est tertia pars aquarum in absinthium et multi hominum mortui sunt de aquis quia amarae factae sunt
REV|8|12|et quartus angelus tuba cecinit et percussa est tertia pars solis et tertia pars lunae et tertia pars stellarum ut obscuraretur tertia pars eorum et diei non luceret pars tertia et nox similiter
REV|8|13|et vidi et audivi vocem unius aquilae volantis per medium caelum dicentis voce magna vae vae vae habitantibus in terra de ceteris vocibus tubae trium angelorum qui erant tuba canituri
REV|9|1|et quintus angelus tuba cecinit et vidi stellam de caelo cecidisse in terram et data est illi clavis putei abyssi
REV|9|2|et aperuit puteum abyssi et ascendit fumus putei sicut fumus fornacis magnae et obscuratus est sol et aer de fumo putei
REV|9|3|et de fumo exierunt lucustae in terram et data est illis potestas sicut habent potestatem scorpiones terrae
REV|9|4|et praeceptum est illis ne laederent faenum terrae neque omne viride neque omnem arborem nisi tantum homines qui non habent signum Dei in frontibus
REV|9|5|et datum est illis ne occiderent eos sed ut cruciarentur mensibus quinque et cruciatus eorum ut cruciatus scorpii cum percutit hominem
REV|9|6|et in diebus illis quaerent homines mortem et non invenient eam et desiderabunt mori et fugiet mors ab ipsis
REV|9|7|et similitudines lucustarum similes equis paratis in proelium et super capita earum tamquam coronae similes auro et facies earum sicut facies hominum
REV|9|8|et habebant capillos sicut capillos mulierum et dentes earum sicut leonum erant
REV|9|9|et habebant loricas sicut loricas ferreas et vox alarum earum sicut vox curruum equorum multorum currentium in bellum
REV|9|10|et habebant caudas similes scorpionum et aculei in caudis earum potestas earum nocere hominibus mensibus quinque
REV|9|11|et habebant super se regem angelum abyssi cui nomen hebraice Abaddon graece autem Apollyon et latine habet nomen Exterminans
REV|9|12|vae unum abiit ecce veniunt adhuc duo vae post haec
REV|9|13|et sextus angelus tuba cecinit et audivi vocem unum ex cornibus altaris aurei quod est ante oculos Dei
REV|9|14|dicentem sexto angelo qui habebat tubam solve quattuor angelos qui alligati sunt in flumine magno Eufrate
REV|9|15|et soluti sunt quattuor angeli qui parati erant in horam et diem et mensem et annum ut occiderent tertiam partem hominum
REV|9|16|et numerus equestris exercitus vicies milies dena milia audivi numerum eorum
REV|9|17|et ita vidi equos in visione et qui sedebant super eos habentes loricas igneas et hyacinthinas et sulphureas et capita equorum erant tamquam capita leonum et de ore ipsorum procedit ignis et fumus et sulphur
REV|9|18|ab his tribus plagis occisa est tertia pars hominum de igne et fumo et sulphure qui procedebat ex ore ipsorum
REV|9|19|potestas enim equorum in ore eorum est et in caudis eorum nam caudae illorum similes serpentibus habentes capita et in his nocent
REV|9|20|et ceteri homines qui non sunt occisi in his plagis neque paenitentiam egerunt de operibus manuum suarum ut non adorarent daemonia et simulacra aurea et argentea et aerea et lapidea et lignea quae neque videre possunt neque audire neque ambulare
REV|9|21|et non egerunt paenitentiam ab homicidiis suis neque a veneficiis suis neque a fornicatione sua neque a furtis suis
REV|10|1|et vidi alium angelum fortem descendentem de caelo amictum nube et iris in capite eius et facies eius erat ut sol et pedes eius tamquam columna ignis
REV|10|2|et habebat in manu sua libellum apertum et posuit pedem suum dextrum supra mare sinistrum autem super terram
REV|10|3|et clamavit voce magna quemadmodum cum leo rugit et cum clamasset locuta sunt septem tonitrua voces suas
REV|10|4|et cum locuta fuissent septem tonitrua scripturus eram et audivi vocem de caelo dicentem signa quae locuta sunt septem tonitrua et noli ea scribere
REV|10|5|et angelum quem vidi stantem supra mare et supra terram levavit manum suam ad caelum
REV|10|6|et iuravit per viventem in saecula saeculorum qui creavit caelum et ea quae in illo sunt et terram et ea quae in ea sunt et mare et quae in eo sunt quia tempus amplius non erit
REV|10|7|sed in diebus vocis septimi angeli cum coeperit tuba canere et consummabitur mysterium Dei sicut evangelizavit per servos suos prophetas
REV|10|8|et vox quam audivi de caelo iterum loquentem mecum et dicentem vade accipe librum apertum de manu angeli stantis supra mare et supra terram
REV|10|9|et abii ad angelum dicens ei ut daret mihi librum et dicit mihi accipe et devora illum et faciet amaricare ventrem tuum sed in ore tuo erit dulce tamquam mel
REV|10|10|et accepi librum de manu angeli et devoravi eum et erat in ore meo tamquam mel dulce et cum devorassem eum amaricatus est venter meus
REV|10|11|et dicunt mihi oportet te iterum prophetare populis et gentibus et linguis et regibus multis
REV|11|1|et datus est mihi calamus similis virgae dicens surge et metire templum Dei et altare et adorantes in eo
REV|11|2|atrium autem quod est foris templum eice foras et ne metieris eum quoniam datum est gentibus et civitatem sanctam calcabunt mensibus quadraginta duobus
REV|11|3|et dabo duobus testibus meis et prophetabunt diebus mille ducentis sexaginta amicti saccos
REV|11|4|hii sunt duo olivae et duo candelabra in conspectu Domini terrae stantes
REV|11|5|et si quis eos voluerit nocere ignis exiet de ore illorum et devorabit inimicos eorum et si quis voluerit eos laedere sic oportet eum occidi
REV|11|6|hii habent potestatem cludendi caelum ne pluat diebus prophetiae ipsorum et potestatem habent super aquas convertendi eas in sanguinem et percutere terram omni plaga quotienscumque voluerint
REV|11|7|et cum finierint testimonium suum bestia quae ascendit de abysso faciet adversus illos bellum et vincet eos et occidet illos
REV|11|8|et corpora eorum in plateis civitatis magnae quae vocatur spiritaliter Sodoma et Aegyptus ubi et Dominus eorum crucifixus est
REV|11|9|et videbunt de populis et tribubus et linguis et gentibus corpora eorum per tres dies et dimidium et corpora eorum non sinunt poni in monumentis
REV|11|10|et inhabitantes terram gaudebunt super illis et iucundabuntur et munera mittent invicem quoniam hii duo prophetae cruciaverunt eos qui inhabitant super terram
REV|11|11|et post dies tres et dimidium spiritus vitae a Deo intravit in eos et steterunt super pedes suos et timor magnus cecidit super eos qui viderunt eos
REV|11|12|et audierunt vocem magnam de caelo dicentem illis ascendite huc et ascenderunt in caelum in nube et viderunt illos inimici eorum
REV|11|13|et in illa hora factus est terraemotus magnus et decima pars civitatis cecidit et occisi sunt in terraemotu nomina hominum septem milia et reliqui in timore sunt missi et dederunt gloriam Deo caeli
REV|11|14|vae secundum abiit ecce vae tertium veniet cito
REV|11|15|et septimus angelus tuba cecinit et factae sunt voces magnae in caelo dicentes factum est regnum huius mundi Domini nostri et Christi eius et regnabit in saecula saeculorum
REV|11|16|et viginti quattuor seniores qui in conspectu Dei sedent in sedibus suis ceciderunt in facies suas et adoraverunt Deum
REV|11|17|dicentes gratias agimus tibi Domine Deus omnipotens qui es et qui eras quia accepisti virtutem tuam magnam et regnasti
REV|11|18|et iratae sunt gentes et advenit ira tua et tempus mortuorum iudicari et reddere mercedem servis tuis prophetis et sanctis et timentibus nomen tuum pusillis et magnis et exterminandi eos qui corruperunt terram
REV|11|19|et apertum est templum Dei in caelo et visa est arca testamenti eius in templo eius et facta sunt fulgora et voces et terraemotus et grando magna
REV|12|1|et signum magnum paruit in caelo mulier amicta sole et luna sub pedibus eius et in capite eius corona stellarum duodecim
REV|12|2|et in utero habens et clamat parturiens et cruciatur ut pariat
REV|12|3|et visum est aliud signum in caelo et ecce draco magnus rufus habens capita septem et cornua decem et in capitibus suis septem diademata
REV|12|4|et cauda eius trahebat tertiam partem stellarum caeli et misit eas in terram et draco stetit ante mulierem quae erat paritura ut cum peperisset filium eius devoraret
REV|12|5|et peperit filium masculum qui recturus erit omnes gentes in virga ferrea et raptus est filius eius ad Deum et ad thronum eius
REV|12|6|et mulier fugit in solitudinem ubi habet locum paratum a Deo ut ibi pascant illam diebus mille ducentis sexaginta
REV|12|7|et factum est proelium in caelo Michahel et angeli eius proeliabantur cum dracone et draco pugnabat et angeli eius
REV|12|8|et non valuerunt neque locus inventus est eorum amplius in caelo
REV|12|9|et proiectus est draco ille magnus serpens antiquus qui vocatur Diabolus et Satanas qui seducit universum orbem proiectus est in terram et angeli eius cum illo missi sunt
REV|12|10|et audivi vocem magnam in caelo dicentem nunc facta est salus et virtus et regnum Dei nostri et potestas Christi eius quia proiectus est accusator fratrum nostrorum qui accusabat illos ante conspectum Dei nostri die ac nocte
REV|12|11|et ipsi vicerunt illum propter sanguinem agni et propter verbum testimonii sui et non dilexerunt animam suam usque ad mortem
REV|12|12|propterea laetamini caeli et qui habitatis in eis vae terrae et mari quia descendit diabolus ad vos habens iram magnam sciens quod modicum tempus habet
REV|12|13|et postquam vidit draco quod proiectus est in terram persecutus est mulierem quae peperit masculum
REV|12|14|et datae sunt mulieri duae alae aquilae magnae ut volaret in desertum in locum suum ubi alitur per tempus et tempora et dimidium temporis a facie serpentis
REV|12|15|et misit serpens ex ore suo post mulierem aquam tamquam flumen ut eam faceret trahi a flumine
REV|12|16|et adiuvit terra mulierem et aperuit terra os suum et absorbuit flumen quod misit draco de ore suo
REV|12|17|et iratus est draco in mulierem et abiit facere proelium cum reliquis de semine eius qui custodiunt mandata Dei et habent testimonium Iesu
REV|12|18|et stetit super harenam maris
REV|13|1|et vidi de mare bestiam ascendentem habentem capita septem et cornua decem et super cornua eius decem diademata et super capita eius nomina blasphemiae
REV|13|2|et bestiam quam vidi similis erat pardo et pedes eius sicut ursi et os eius sicut os leonis et dedit illi draco virtutem suam et potestatem magnam
REV|13|3|et unum de capitibus suis quasi occisum in mortem et plaga mortis eius curata est et admirata est universa terra post bestiam
REV|13|4|et adoraverunt draconem quia dedit potestatem bestiae et adoraverunt bestiam dicentes quis similis bestiae et quis poterit pugnare cum ea
REV|13|5|et datum est ei os loquens magna et blasphemiae et data est illi potestas facere menses quadraginta duo
REV|13|6|et aperuit os suum in blasphemias ad Deum blasphemare nomen eius et tabernaculum eius et eos qui in caelo habitant
REV|13|7|et datum est illi bellum facere cum sanctis et vincere illos et data est ei potestas in omnem tribum et populum et linguam et gentem
REV|13|8|et adorabunt eum omnes qui inhabitant terram quorum non sunt scripta nomina in libro vitae agni qui occisus est ab origine mundi
REV|13|9|si quis habet aurem audiat
REV|13|10|qui in captivitatem in captivitatem vadit qui in gladio occiderit oportet eum gladio occidi hic est patientia et fides sanctorum
REV|13|11|et vidi aliam bestiam ascendentem de terra et habebat cornua duo similia agni et loquebatur sicut draco
REV|13|12|et potestatem prioris bestiae omnem faciebat in conspectu eius et facit terram et inhabitantes in eam adorare bestiam primam cuius curata est plaga mortis
REV|13|13|et fecit signa magna ut etiam ignem faceret de caelo descendere in terram in conspectu hominum
REV|13|14|et seducit habitantes terram propter signa quae data sunt illi facere in conspectu bestiae dicens habitantibus in terra ut faciant imaginem bestiae quae habet plagam gladii et vixit
REV|13|15|et datum est illi ut daret spiritum imagini bestiae ut et loquatur imago bestiae et faciat quicumque non adoraverint imaginem bestiae occidantur
REV|13|16|et faciet omnes pusillos et magnos et divites et pauperes et liberos et servos habere caracter in dextera manu aut in frontibus suis
REV|13|17|et ne quis possit emere aut vendere nisi qui habet caracter nomen bestiae aut numerum nominis eius
REV|13|18|hic sapientia est qui habet intellectum conputet numerum bestiae numerus enim hominis est et numerus eius est sescenti sexaginta sex
REV|14|1|et vidi et ecce agnus stabat supra montem Sion et cum illo centum quadraginta quattuor milia habentes nomen eius et nomen Patris eius scriptum in frontibus suis
REV|14|2|et audivi vocem de caelo tamquam vocem aquarum multarum et tamquam vocem tonitrui magni et vocem quam audivi sicut citharoedorum citharizantium in citharis suis
REV|14|3|et cantabant quasi canticum novum ante sedem et ante quattuor animalia et seniores et nemo poterat discere canticum nisi illa centum quadraginta quattuor milia qui empti sunt de terra
REV|14|4|hii sunt qui cum mulieribus non sunt coinquinati virgines enim sunt hii qui sequuntur agnum quocumque abierit hii empti sunt ex hominibus primitiae Deo et agno
REV|14|5|et in ore ipsorum non est inventum mendacium sine macula sunt
REV|14|6|et vidi alterum angelum volantem per medium caelum habentem evangelium aeternum ut evangelizaret sedentibus super terram et super omnem gentem et tribum et linguam et populum
REV|14|7|dicens magna voce timete Deum et date illi honorem quia venit hora iudicii eius et adorate eum qui fecit caelum et terram et mare et fontes aquarum
REV|14|8|et alius angelus secutus est dicens cecidit cecidit Babylon illa magna quae a vino irae fornicationis suae potionavit omnes gentes
REV|14|9|et alius angelus tertius secutus est illos dicens voce magna si quis adoraverit bestiam et imaginem eius et acceperit caracterem in fronte sua aut in manu sua
REV|14|10|et hic bibet de vino irae Dei qui mixtus est mero in calice irae ipsius et cruciabitur igne et sulphure in conspectu angelorum sanctorum et ante conspectum agni
REV|14|11|et fumus tormentorum eorum in saecula saeculorum ascendit nec habent requiem die ac nocte qui adoraverunt bestiam et imaginem eius et si quis acceperit caracterem nominis eius
REV|14|12|hic patientia sanctorum est qui custodiunt mandata Dei et fidem Iesu
REV|14|13|et audivi vocem de caelo dicentem scribe beati mortui qui in Domino moriuntur amodo iam dicit Spiritus ut requiescant a laboribus suis opera enim illorum sequuntur illos
REV|14|14|et vidi et ecce nubem candidam et supra nubem sedentem similem Filio hominis habentem in capite suo coronam auream et in manu sua falcem acutam
REV|14|15|et alter angelus exivit de templo clamans voce magna ad sedentem super nubem mitte falcem tuam et mete quia venit hora ut metatur quoniam aruit messis terrae
REV|14|16|et misit qui sedebat supra nubem falcem suam in terram et messa est terra
REV|14|17|et alius angelus exivit de templo quod est in caelo habens et ipse falcem acutam
REV|14|18|et alius angelus de altari qui habet potestatem supra ignem et clamavit voce magna qui habebat falcem acutam dicens mitte falcem tuam acutam et vindemia botros vineae terrae quoniam maturae sunt uvae eius
REV|14|19|et misit angelus falcem suam in terram et vindemiavit vineam terrae et misit in lacum irae Dei magnum
REV|14|20|et calcatus est lacus extra civitatem et exivit sanguis de lacu usque ad frenos equorum per stadia mille sescenta
REV|15|1|et vidi aliud signum in caelo magnum et mirabile angelos septem habentes plagas septem novissimas quoniam in illis consummata est ira Dei
REV|15|2|et vidi tamquam mare vitreum mixtum igne et eos qui vicerunt bestiam et imaginem illius et numerum nominis eius stantes supra mare vitreum habentes citharas Dei
REV|15|3|et cantant canticum Mosi servi Dei et canticum agni dicentes magna et mirabilia opera tua Domine Deus omnipotens iustae et verae viae tuae rex saeculorum
REV|15|4|quis non timebit Domine et magnificabit nomen tuum quia solus pius quoniam omnes gentes venient et adorabunt in conspectu tuo quoniam iudicia tua manifestata sunt
REV|15|5|et post haec vidi et ecce apertum est templum tabernaculi testimonii in caelo
REV|15|6|et exierunt septem angeli habentes septem plagas de templo vestiti lapide mundo candido et praecincti circa pectora zonis aureis
REV|15|7|et unus ex quattuor animalibus dedit septem angelis septem fialas aureas plenas iracundiae Dei viventis in saecula saeculorum
REV|15|8|et impletum est templum fumo a maiestate Dei et de virtute eius et nemo poterat introire in templum donec consummarentur septem plagae septem angelorum
REV|16|1|et audivi vocem magnam de templo dicentem septem angelis ite et effundite septem fialas irae Dei in terram
REV|16|2|et abiit primus et effudit fialam suam in terram et factum est vulnus saevum ac pessimum in homines qui habent caracterem bestiae et eos qui adoraverunt imaginem eius
REV|16|3|et secundus effudit fialam suam in mare et factus est sanguis tamquam mortui et omnis anima vivens mortua est in mari
REV|16|4|et tertius effudit fialam suam super flumina et super fontes aquarum et factus est sanguis
REV|16|5|et audivi angelum aquarum dicentem iustus es qui es et qui eras sanctus quia haec iudicasti
REV|16|6|quia sanguinem sanctorum et prophetarum fuderunt et sanguinem eis dedisti bibere digni sunt
REV|16|7|et audivi altare dicens etiam Domine Deus omnipotens vera et iusta iudicia tua
REV|16|8|et quartus effudit fialam suam in solem et datum est illi aestu adficere homines et igni
REV|16|9|et aestuaverunt homines aestu magno et blasphemaverunt nomen Dei habentis potestatem super has plagas neque egerunt paenitentiam ut darent illi gloriam
REV|16|10|et quintus effudit fialam suam super sedem bestiae et factum est regnum eius tenebrosum et conmanducaverunt linguas suas prae dolore
REV|16|11|et blasphemaverunt Deum caeli prae doloribus et vulneribus suis et non egerunt paenitentiam ex operibus suis
REV|16|12|et sextus effudit fialam suam in flumen illud magnum Eufraten et siccavit aquam eius ut praepararetur via regibus ab ortu solis
REV|16|13|et vidi de ore draconis et de ore bestiae et de ore pseudoprophetae spiritus tres inmundos in modum ranarum
REV|16|14|sunt enim spiritus daemoniorum facientes signa et procedunt ad reges totius terrae congregare illos in proelium ad diem magnum Dei omnipotentis
REV|16|15|ecce venio sicut fur beatus qui vigilat et custodit vestimenta sua ne nudus ambulet et videant turpitudinem eius
REV|16|16|et congregavit illos in locum qui vocatur hebraice Hermagedon
REV|16|17|et septimus effudit fialam suam in aerem et exivit vox magna de templo a throno dicens factum est
REV|16|18|et facta sunt fulgora et voces et tonitrua et terraemotus factus est magnus qualis numquam fuit ex quo homines fuerunt super terram talis terraemotus sic magnus
REV|16|19|et facta est civitas magna in tres partes et civitates gentium ceciderunt et Babylon magna venit in memoriam ante Deum dare ei calicem vini indignationis irae eius
REV|16|20|et omnis insula fugit et montes non sunt inventi
REV|16|21|et grando magna sicut talentum descendit de caelo in homines et blasphemaverunt homines Deum propter plagam grandinis quoniam magna facta est vehementer
REV|17|1|et venit unus de septem angelis qui habebant septem fialas et locutus est mecum dicens veni ostendam tibi damnationem meretricis magnae quae sedet super aquas multas
REV|17|2|cum qua fornicati sunt reges terrae et inebriati sunt qui inhabitant terram de vino prostitutionis eius
REV|17|3|et abstulit me in desertum in spiritu et vidi mulierem sedentem super bestiam coccineam plenam nominibus blasphemiae habentem capita septem et cornua decem
REV|17|4|et mulier erat circumdata purpura et coccino et inaurata auro et lapide pretioso et margaritis habens poculum aureum in manu sua plenum abominationum et inmunditia fornicationis eius
REV|17|5|et in fronte eius nomen scriptum mysterium Babylon magna mater fornicationum et abominationum terrae
REV|17|6|et vidi mulierem ebriam de sanguine sanctorum et de sanguine martyrum Iesu et miratus sum cum vidissem illam admiratione magna
REV|17|7|et dixit mihi angelus quare miraris ego tibi dicam sacramentum mulieris et bestiae quae portat eam quae habet capita septem et decem cornua
REV|17|8|bestiam quam vidisti fuit et non est et ascensura est de abysso et in interitum ibit et mirabuntur inhabitantes terram quorum non sunt scripta nomina in libro vitae a constitutione mundi videntes bestiam quia erat et non est
REV|17|9|et hic est sensus qui habet sapientiam septem capita septem montes sunt super quos mulier sedet et reges septem sunt
REV|17|10|quinque ceciderunt unus est alius nondum venit et cum venerit oportet illum breve tempus manere
REV|17|11|et bestia quae erat et non est et ipsa octava est et de septem est et in interitum vadit
REV|17|12|et decem cornua quae vidisti decem reges sunt qui regnum nondum acceperunt sed potestatem tamquam reges una hora accipiunt post bestiam
REV|17|13|hii unum consilium habent et virtutem et potestatem suam bestiae tradunt
REV|17|14|hii cum agno pugnabunt et agnus vincet illos quoniam Dominus dominorum est et rex regum et qui cum illo sunt vocati et electi et fideles
REV|17|15|et dixit mihi aquas quas vidisti ubi meretrix sedet populi sunt et gentes et linguae
REV|17|16|et decem cornua quae vidisti et bestiam hii odient fornicariam et desolatam facient illam et nudam et carnes eius manducabunt et ipsam igni concremabunt
REV|17|17|Deus enim dedit in corda eorum ut faciant quod illi placitum est ut dent regnum suum bestiae donec consummentur verba Dei
REV|17|18|et mulier quam vidisti est civitas magna quae habet regnum super reges terrae
REV|18|1|et post haec vidi alium angelum descendentem de caelo habentem potestatem magnam et terra inluminata est a gloria eius
REV|18|2|et exclamavit in forti voce dicens cecidit cecidit Babylon magna et facta est habitatio daemoniorum et custodia omnis spiritus inmundi et custodia omnis volucris inmundae
REV|18|3|quia de ira fornicationis eius biberunt omnes gentes et reges terrae cum illa fornicati sunt et mercatores terrae de virtute deliciarum eius divites facti sunt
REV|18|4|et audivi aliam vocem de caelo dicentem exite de illa populus meus ut ne participes sitis delictorum eius et de plagis eius non accipiatis
REV|18|5|quoniam pervenerunt peccata eius usque ad caelum et recordatus est Deus iniquitatum eius
REV|18|6|reddite illi sicut ipsa reddidit et duplicate duplicia secundum opera eius in poculo quo miscuit miscite illi duplum
REV|18|7|quantum glorificavit se et in deliciis fuit tantum date illi tormentum et luctum quia in corde suo dicit sedeo regina et vidua non sum et luctum non videbo
REV|18|8|ideo in una die venient plagae eius mors et luctus et fames et igni conburetur quia fortis est Deus qui iudicavit illam
REV|18|9|et flebunt et plangent se super illam reges terrae qui cum illa fornicati sunt et in deliciis vixerunt cum viderint fumum incendii eius
REV|18|10|longe stantes propter timorem tormentorum eius dicentes vae vae civitas illa magna Babylon civitas illa fortis quoniam una hora venit iudicium tuum
REV|18|11|et negotiatores terrae flebunt et lugebunt super illam quoniam merces eorum nemo emet amplius
REV|18|12|mercem auri et argenti et lapidis pretiosi et margaritis et byssi et purpurae et serici et cocci et omne lignum thyinum et omnia vasa eboris et omnia vasa de lapide pretioso et aeramento et ferro et marmore
REV|18|13|et cinnamomum et amomum et odoramentorum et unguenti et turis et vini et olei et similae et tritici et iumentorum et ovium et equorum et raedarum et mancipiorum et animarum hominum
REV|18|14|et poma tua desiderii animae discessit a te et omnia pinguia et clara perierunt a te et amplius illa iam non invenient
REV|18|15|mercatores horum qui divites facti sunt ab ea longe stabunt propter timorem tormentorum eius flentes ac lugentes
REV|18|16|et dicentes vae vae civitas illa magna quae amicta erat byssino et purpura et cocco et deaurata est auro et lapide pretioso et margaritis
REV|18|17|quoniam una hora destitutae sunt tantae divitiae et omnis gubernator et omnis qui in locum navigat et nautae et qui maria operantur longe steterunt
REV|18|18|et clamaverunt videntes locum incendii eius dicentes quae similis civitati huic magnae
REV|18|19|et miserunt pulverem super capita sua et clamaverunt flentes et lugentes dicentes vae vae civitas magna in qua divites facti sunt omnes qui habent naves in mari de pretiis eius quoniam una hora desolata est
REV|18|20|exulta super eam caelum et sancti et apostoli et prophetae quoniam iudicavit Deus iudicium vestrum de illa
REV|18|21|et sustulit unus angelus fortis lapidem quasi molarem magnum et misit in mare dicens hoc impetu mittetur Babylon magna illa civitas et ultra iam non invenietur
REV|18|22|et vox citharoedorum et musicorum et tibia canentium et tuba non audietur in te amplius et omnis artifex omnis artis non invenietur in te amplius et vox molae non audietur in te amplius
REV|18|23|et lux lucernae non lucebit tibi amplius et vox sponsi et sponsae non audietur adhuc in te quia mercatores tui erant principes terrae quia in veneficiis tuis erraverunt omnes gentes
REV|18|24|et in ea sanguis prophetarum et sanctorum inventus est et omnium qui interfecti sunt in terra
REV|19|1|post haec audivi quasi vocem magnam turbarum multarum in caelo dicentium alleluia salus et gloria et virtus Deo nostro est
REV|19|2|quia vera et iusta iudicia sunt eius quia iudicavit de meretrice magna quae corrupit terram in prostitutione sua et vindicavit sanguinem servorum suorum de manibus eius
REV|19|3|et iterum dixerunt alleluia et fumus eius ascendit in saecula saeculorum
REV|19|4|et ceciderunt seniores viginti quattuor et quattuor animalia et adoraverunt Deum sedentem super thronum dicentes amen alleluia
REV|19|5|et vox de throno exivit dicens laudem dicite Deo nostro omnes servi eius et qui timetis eum pusilli et magni
REV|19|6|et audivi quasi vocem turbae magnae et sicut vocem aquarum multarum et sicut vocem tonitruum magnorum dicentium alleluia quoniam regnavit Dominus Deus noster omnipotens
REV|19|7|gaudeamus et exultemus et demus gloriam ei quia venerunt nuptiae agni et uxor eius praeparavit se
REV|19|8|et datum est illi ut cooperiat se byssinum splendens candidum byssinum enim iustificationes sunt sanctorum
REV|19|9|et dicit mihi scribe beati qui ad cenam nuptiarum agni vocati sunt et dicit mihi haec verba vera Dei sunt
REV|19|10|et cecidi ante pedes eius ut adorarem eum et dicit mihi vide ne feceris conservus tuus sum et fratrum tuorum habentium testimonium Iesu Deum adora testimonium enim Iesu est spiritus prophetiae
REV|19|11|et vidi caelum apertum et ecce equus albus et qui sedebat super eum vocabatur Fidelis et Verax vocatur et iustitia iudicat et pugnat
REV|19|12|oculi autem eius sicut flamma ignis et in capite eius diademata multa habens nomen scriptum quod nemo novit nisi ipse
REV|19|13|et vestitus erat vestem aspersam sanguine et vocatur nomen eius Verbum Dei
REV|19|14|et exercitus qui sunt in caelo sequebantur eum in equis albis vestiti byssinum album mundum
REV|19|15|et de ore ipsius procedit gladius acutus ut in ipso percutiat gentes et ipse reget eos in virga ferrea et ipse calcat torcular vini furoris irae Dei omnipotentis
REV|19|16|et habet in vestimento et in femore suo scriptum rex regum et Dominus dominantium
REV|19|17|et vidi unum angelum stantem in sole et clamavit voce magna dicens omnibus avibus quae volabant per medium caeli venite congregamini ad cenam magnam Dei
REV|19|18|ut manducetis carnes regum et carnes tribunorum et carnes fortium et carnes equorum et sedentium in ipsis et carnes omnium liberorum ac servorum et pusillorum ac magnorum
REV|19|19|et vidi bestiam et reges terrae et exercitus eorum congregatos ad faciendum proelium cum illo qui sedebat in equo et cum exercitu eius
REV|19|20|et adprehensa est bestia et cum illo pseudopropheta qui fecit signa coram ipso quibus seduxit eos qui acceperunt caracterem bestiae qui et adorant imaginem eius vivi missi sunt hii duo in stagnum ignis ardentis sulphure
REV|19|21|et ceteri occisi sunt in gladio sedentis super equum qui procedit de ore ipsius et omnes aves saturatae sunt carnibus eorum
REV|20|1|et vidi angelum descendentem de caelo habentem clavem abyssi et catenam magnam in manu sua
REV|20|2|et adprehendit draconem serpentem antiquum qui est diabolus et Satanas et ligavit eum per annos mille
REV|20|3|et misit eum in abyssum et clusit et signavit super illum ut non seducat amplius gentes donec consummentur mille anni post haec oportet illum solvi modico tempore
REV|20|4|et vidi sedes et sederunt super eas et iudicium datum est illis et animas decollatorum propter testimonium Iesu et propter verbum Dei et qui non adoraverunt bestiam neque imaginem eius nec acceperunt caracterem in frontibus aut in manibus suis et vixerunt et regnaverunt cum Christo mille annis
REV|20|5|ceteri mortuorum non vixerunt donec consummentur mille anni haec est resurrectio prima
REV|20|6|beatus et sanctus qui habet partem in resurrectione prima in his secunda mors non habet potestatem sed erunt sacerdotes Dei et Christi et regnabunt cum illo mille annis
REV|20|7|et cum consummati fuerint mille anni solvetur Satanas de carcere suo et exibit et seducet gentes quae sunt super quattuor angulos terrae Gog et Magog et congregabit eos in proelium quorum numerus est sicut harena maris
REV|20|8|et ascenderunt super latitudinem terrae et circumierunt castra sanctorum et civitatem dilectam
REV|20|9|et descendit ignis a Deo de caelo et devoravit eos et diabolus qui seducebat eos missus est in stagnum ignis et sulphuris ubi et bestia
REV|20|10|et pseudoprophetes et cruciabuntur die ac nocte in saecula saeculorum
REV|20|11|et vidi thronum magnum candidum et sedentem super eum a cuius aspectu fugit terra et caelum et locus non est inventus ab eis
REV|20|12|et vidi mortuos magnos et pusillos stantes in conspectu throni et libri aperti sunt et alius liber apertus est qui est vitae et iudicati sunt mortui ex his quae scripta erant in libris secundum opera ipsorum
REV|20|13|et dedit mare mortuos qui in eo erant et mors et inferus dederunt mortuos qui in ipsis erant et iudicatum est de singulis secundum opera ipsorum
REV|20|14|et inferus et mors missi sunt in stagnum ignis haec mors secunda est stagnum ignis
REV|20|15|et qui non est inventus in libro vitae scriptus missus est in stagnum ignis
REV|21|1|et vidi caelum novum et terram novam primum enim caelum et prima terra abiit et mare iam non est
REV|21|2|et civitatem sanctam Hierusalem novam vidi descendentem de caelo a Deo paratam sicut sponsam ornatam viro suo
REV|21|3|et audivi vocem magnam de throno dicentem ecce tabernaculum Dei cum hominibus et habitabit cum eis et ipsi populus eius erunt et ipse Deus cum eis erit eorum Deus
REV|21|4|et absterget Deus omnem lacrimam ab oculis eorum et mors ultra non erit neque luctus neque clamor neque dolor erit ultra quae prima abierunt
REV|21|5|et dixit qui sedebat in throno ecce nova facio omnia et dicit scribe quia haec verba fidelissima sunt et vera
REV|21|6|et dixit mihi factum est ego sum Alpha et Omega initium et finis ego sitienti dabo de fonte aquae vivae gratis
REV|21|7|qui vicerit possidebit haec et ero illi Deus et ille erit mihi filius
REV|21|8|timidis autem et incredulis et execratis et homicidis et fornicatoribus et veneficis et idolatris et omnibus mendacibus pars illorum erit in stagno ardenti igne et sulphure quod est mors secunda
REV|21|9|et venit unus de septem angelis habentibus fialas plenas septem plagis novissimis et locutus est mecum dicens veni ostendam tibi sponsam uxorem agni
REV|21|10|et sustulit me in spiritu in montem magnum et altum et ostendit mihi civitatem sanctam Hierusalem descendentem de caelo a Deo
REV|21|11|habentem claritatem Dei lumen eius simile lapidi pretioso tamquam lapidi iaspidis sicut cristallum
REV|21|12|et habebat murum magnum et altum habens portas duodecim et in portis angelos duodecim et nomina inscripta quae sunt nomina duodecim tribuum filiorum Israhel
REV|21|13|ab oriente portae tres et ab aquilone portae tres et ab austro portae tres et ab occasu portae tres
REV|21|14|et murus civitatis habens fundamenta duodecim et in ipsis duodecim nomina duodecim apostolorum agni
REV|21|15|et qui loquebatur mecum habebat mensuram harundinem auream ut metiretur civitatem et portas eius et murum
REV|21|16|et civitas in quadro posita est et longitudo eius tanta est quanta et latitudo et mensus est civitatem de harundine per stadia duodecim milia longitudo et latitudo et altitudo eius aequalia sunt
REV|21|17|et mensus est murus eius centum quadraginta quattuor cubitorum mensura hominis quae est angeli
REV|21|18|et erat structura muri eius ex lapide iaspide ipsa vero civitas auro mundo simile vitro mundo
REV|21|19|fundamenta muri civitatis omni lapide pretioso ornata fundamentum primum iaspis secundus sapphyrus tertius carcedonius quartus zmaragdus
REV|21|20|quintus sardonix sextus sardinus septimus chrysolitus octavus berillus nonus topazius decimus chrysoprassus undecimus hyacinthus duodecimus amethistus
REV|21|21|et duodecim portae duodecim margaritae sunt per singulas et singulae portae erant ex singulis margaritis et platea civitatis aurum mundum tamquam vitrum perlucidum
REV|21|22|et templum non vidi in ea Dominus enim Deus omnipotens templum illius est et agnus
REV|21|23|et civitas non eget sole neque luna ut luceant in ea nam claritas Dei inluminavit eam et lucerna eius est agnus
REV|21|24|et ambulabunt gentes per lumen eius et reges terrae adferent gloriam suam et honorem in illam
REV|21|25|et portae eius non cludentur per diem nox enim non erit illic
REV|21|26|et adferent gloriam et honorem gentium in illam
REV|21|27|nec intrabit in ea aliquid coinquinatum et faciens abominationem et mendacium nisi qui scripti sunt in libro vitae agni
REV|22|1|et ostendit mihi fluvium aquae vitae splendidum tamquam cristallum procedentem de sede Dei et agni
REV|22|2|in medio plateae eius et ex utraque parte fluminis lignum vitae adferens fructus duodecim per menses singula reddentia fructum suum et folia ligni ad sanitatem gentium
REV|22|3|et omne maledictum non erit amplius et sedes Dei et agni in illa erunt et servi eius servient illi
REV|22|4|et videbunt faciem eius et nomen eius in frontibus eorum
REV|22|5|et nox ultra non erit et non egebunt lumine lucernae neque lumine solis quoniam Dominus Deus inluminat illos et regnabunt in saecula saeculorum
REV|22|6|et dixit mihi haec verba fidelissima et vera sunt et Dominus Deus spirituum prophetarum misit angelum suum ostendere servis suis quae oportet fieri cito
REV|22|7|et ecce venio velociter beatus qui custodit verba prophetiae libri huius
REV|22|8|et ego Iohannes qui audivi et vidi haec et postquam audissem et vidissem cecidi ut adorarem ante pedes angeli qui mihi haec ostendebat
REV|22|9|et dicit mihi vide ne feceris conservus tuus sum et fratrum tuorum prophetarum et eorum qui servant verba libri huius Deum adora
REV|22|10|et dicit mihi ne signaveris verba prophetiae libri huius tempus enim prope est
REV|22|11|qui nocet noceat adhuc et qui in sordibus est sordescat adhuc et iustus iustitiam faciat adhuc et sanctus sanctificetur adhuc
REV|22|12|ecce venio cito et merces mea mecum est reddere unicuique secundum opera sua
REV|22|13|ego Alpha et Omega primus et novissimus principium et finis
REV|22|14|beati qui lavant stolas suas ut sit potestas eorum in ligno vitae et portis intrent in civitatem
REV|22|15|foris canes et venefici et inpudici et homicidae et idolis servientes et omnis qui amat et facit mendacium
REV|22|16|ego Iesus misi angelum meum testificari vobis haec in ecclesiis ego sum radix et genus David stella splendida et matutina
REV|22|17|et Spiritus et sponsa dicunt veni et qui audit dicat veni et qui sitit veniat qui vult accipiat aquam vitae gratis
REV|22|18|contestor ego omni audienti verba prophetiae libri huius si quis adposuerit ad haec adponet Deus super illum plagas scriptas in libro isto
REV|22|19|et si quis deminuerit de verbis libri prophetiae huius auferet Deus partem eius de ligno vitae et de civitate sancta et de his quae scripta sunt in libro isto
REV|22|20|dicit qui testimonium perhibet istorum etiam venio cito amen veni Domine Iesu
REV|22|21|gratia Domini nostri Iesu Christi cum omnibus
