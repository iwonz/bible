ISA|1|1|visio Isaiae filii Amos quam vidit super Iudam et Hierusalem in diebus Oziae Ioatham Ahaz Ezechiae regum Iuda
ISA|1|2|audite caeli et auribus percipe terra quoniam Dominus locutus est filios enutrivi et exaltavi ipsi autem spreverunt me
ISA|1|3|cognovit bos possessorem suum et asinus praesepe domini sui Israhel non cognovit populus meus non intellexit
ISA|1|4|vae genti peccatrici populo gravi iniquitate semini nequam filiis sceleratis dereliquerunt Dominum blasphemaverunt Sanctum Israhel abalienati sunt retrorsum
ISA|1|5|super quo percutiam vos ultra addentes praevaricationem omne caput languidum et omne cor maerens
ISA|1|6|a planta pedis usque ad verticem non est in eo sanitas vulnus et livor et plaga tumens non est circumligata nec curata medicamine neque fota oleo
ISA|1|7|terra vestra deserta civitates vestrae succensae igni regionem vestram coram vobis alieni devorant et desolabitur sicut in vastitate hostili
ISA|1|8|et derelinquetur filia Sion ut umbraculum in vinea et sicut tugurium in cucumerario sicut civitas quae vastatur
ISA|1|9|nisi Dominus exercituum reliquisset nobis semen quasi Sodoma fuissemus et quasi Gomorra similes essemus
ISA|1|10|audite verbum Domini principes Sodomorum percipite auribus legem Dei nostri populus Gomorrae
ISA|1|11|quo mihi multitudinem victimarum vestrarum dicit Dominus plenus sum holocausta arietum et adipem pinguium et sanguinem vitulorum et agnorum et hircorum nolui
ISA|1|12|cum veneritis ante conspectum meum quis quaesivit haec de manibus vestris ut ambularetis in atriis meis
ISA|1|13|ne adferatis ultra sacrificium frustra incensum abominatio est mihi neomeniam et sabbatum et festivitates alias non feram iniqui sunt coetus vestri
ISA|1|14|kalendas vestras et sollemnitates vestras odivit anima mea facta sunt mihi molesta laboravi sustinens
ISA|1|15|et cum extenderitis manus vestras avertam oculos meos a vobis et cum multiplicaveritis orationem non audiam manus vestrae sanguine plenae sunt
ISA|1|16|lavamini mundi estote auferte malum cogitationum vestrarum ab oculis meis quiescite agere perverse
ISA|1|17|discite benefacere quaerite iudicium subvenite oppresso iudicate pupillo defendite viduam
ISA|1|18|et venite et arguite me dicit Dominus si fuerint peccata vestra ut coccinum quasi nix dealbabuntur et si fuerint rubra quasi vermiculus velut lana erunt
ISA|1|19|si volueritis et audieritis bona terrae comedetis
ISA|1|20|quod si nolueritis et me provocaveritis ad iracundiam gladius devorabit vos quia os Domini locutum est
ISA|1|21|quomodo facta est meretrix civitas fidelis plena iudicii iustitia habitavit in ea nunc autem homicidae
ISA|1|22|argentum tuum versum est in scoriam vinum tuum mixtum est aqua
ISA|1|23|principes tui infideles socii furum omnes diligunt munera sequuntur retributiones pupillo non iudicant et causa viduae non ingreditur ad eos
ISA|1|24|propter hoc ait Dominus exercituum Fortis Israhel heu consolabor super hostibus meis et vindicabor de inimicis meis
ISA|1|25|et convertam manum meam ad te et excoquam ad purum scoriam tuam et auferam omne stagnum tuum
ISA|1|26|et restituam iudices tuos ut fuerunt prius et consiliarios tuos sicut antiquitus post haec vocaberis civitas iusti urbs fidelis
ISA|1|27|Sion in iudicio redimetur et reducent eam in iustitia
ISA|1|28|et conteret scelestos et peccatores simul et qui dereliquerunt Dominum consumentur
ISA|1|29|confundentur enim ab idolis quibus sacrificaverunt et erubescetis super hortis quos elegeratis
ISA|1|30|cum fueritis velut quercus defluentibus foliis et velut hortus absque aqua
ISA|1|31|et erit fortitudo vestra ut favilla stuppae et opus vestrum quasi scintilla et succendetur utrumque simul et non erit qui extinguat
ISA|2|1|verbum quod vidit Isaias filius Amos super Iudam et Hierusalem
ISA|2|2|et erit in novissimis diebus praeparatus mons domus Domini in vertice montium et elevabitur super colles et fluent ad eum omnes gentes
ISA|2|3|et ibunt populi multi et dicent venite et ascendamus ad montem Domini et ad domum Dei Iacob et docebit nos vias suas et ambulabimus in semitis eius quia de Sion exibit lex et verbum Domini de Hierusalem
ISA|2|4|et iudicabit gentes et arguet populos multos et conflabunt gladios suos in vomeres et lanceas suas in falces non levabit gens contra gentem gladium nec exercebuntur ultra ad proelium
ISA|2|5|domus Iacob venite et ambulemus in lumine Domini
ISA|2|6|proiecisti enim populum tuum domum Iacob quia repleti sunt ut olim et augures habuerunt ut Philisthim et pueris alienis adheserunt
ISA|2|7|repleta est terra argento et auro et non est finis thesaurorum eius
ISA|2|8|et repleta est terra eius equis et innumerabiles quadrigae eius et repleta est terra eius idolis opus manuum suarum adoraverunt quod fecerunt digiti eorum
ISA|2|9|et incurvavit se homo et humiliatus est vir ne ergo dimittas eis
ISA|2|10|ingredere in petram abscondere fossa humo a facie timoris Domini et a gloria maiestatis eius
ISA|2|11|oculi sublimis hominis humiliati sunt et incurvabitur altitudo virorum exaltabitur autem Dominus solus in die illa
ISA|2|12|quia dies Domini exercituum super omnem superbum et excelsum et super omnem arrogantem et humiliabitur
ISA|2|13|et super omnes cedros Libani sublimes et erectas et super omnes quercus Basan
ISA|2|14|et super omnes montes excelsos et super omnes colles elevatos
ISA|2|15|et super omnem turrem excelsam et super omnem murum munitum
ISA|2|16|et super omnes naves Tharsis et super omne quod visu pulchrum est
ISA|2|17|et incurvabitur sublimitas hominum et humiliabitur altitudo virorum et elevabitur Dominus solus in die illa
ISA|2|18|et idola penitus conterentur
ISA|2|19|et introibunt in speluncas petrarum et in voragines terrae a facie formidinis Domini et a gloria maiestatis eius cum surrexerit percutere terram
ISA|2|20|in die illa proiciet homo idola argenti sui et simulacra auri sui quae fecerat sibi ut adoraret talpas et vespertiliones
ISA|2|21|et ingredietur fissuras petrarum et cavernas saxorum a facie formidinis Domini et a gloria maiestatis eius cum surrexerit percutere terram
ISA|2|22|quiescite ergo ab homine cuius spiritus in naribus eius quia excelsus reputatus est ipse
ISA|3|1|ecce enim Dominator Deus exercituum auferet ab Hierusalem et ab Iuda validum et fortem omne robur panis et omne robur aquae
ISA|3|2|fortem et virum bellatorem iudicem et prophetam et ariolum et senem
ISA|3|3|principem super quinquaginta et honorabilem vultu et consiliarium sapientem de architectis et prudentem eloquii mystici
ISA|3|4|et dabo pueros principes eorum et effeminati dominabuntur eis
ISA|3|5|et inruet populus vir ad virum unusquisque ad proximum suum tumultuabitur puer contra senem et ignobilis contra nobilem
ISA|3|6|adprehendet enim vir fratrem suum domesticum patris sui vestimentum tibi est princeps esto noster ruina autem haec sub manu tua
ISA|3|7|respondebit in die illa dicens non sum medicus et in domo mea non est panis neque vestimentum nolite constituere me principem populi
ISA|3|8|ruit enim Hierusalem et Iudas concidit quia lingua eorum et adinventiones eorum contra Dominum ut provocarent oculos maiestatis eius
ISA|3|9|agnitio vultus eorum respondit eis et peccatum suum quasi Sodomae praedicaverunt nec absconderunt vae animae eorum quoniam reddita sunt eis mala
ISA|3|10|dicite iusto quoniam bene quoniam fructum adinventionum suarum comedet
ISA|3|11|vae impio in malum retributio enim manuum eius fiet ei
ISA|3|12|populum meum exactores sui spoliaverunt et mulieres dominatae sunt eius popule meus qui beatum te dicunt ipsi te decipiunt et viam gressuum tuorum dissipant
ISA|3|13|stat ad iudicandum Dominus et stat ad iudicandos populos
ISA|3|14|Dominus ad iudicium veniet cum senibus populi sui et principibus eius vos enim depasti estis vineam meam et rapina pauperis in domo vestra
ISA|3|15|quare adteritis populum meum et facies pauperum commolitis dicit Dominus Deus exercituum
ISA|3|16|et dixit Dominus pro eo quod elevatae sunt filiae Sion et ambulaverunt extento collo et nutibus oculorum ibant et plaudebant ambulabant et in pedibus suis conposito gradu incedebant
ISA|3|17|decalvabit Dominus verticem filiarum Sion et Dominus crinem earum nudabit
ISA|3|18|in die illa auferet Dominus ornatum calciamentorum et lunulas
ISA|3|19|et torques et monilia et armillas et mitras
ISA|3|20|discriminalia et periscelidas et murenulas et olfactoriola et inaures
ISA|3|21|et anulos et gemmas in fronte pendentes
ISA|3|22|et mutatoria et pallia et linteamina et acus
ISA|3|23|et specula et sindones et vittas et theristra
ISA|3|24|et erit pro suavi odore fetor et pro zona funiculus et pro crispanti crine calvitium et pro fascia pectorali cilicium
ISA|3|25|pulcherrimi quoque viri tui gladio cadent et fortes tui in proelio
ISA|3|26|et maerebunt atque lugebunt portae eius et desolata in terra sedebit
ISA|4|1|et adprehendent septem mulieres virum unum in die illa dicentes panem nostrum comedemus et vestimentis nostris operiemur tantummodo vocetur nomen tuum super nos aufer obprobrium nostrum
ISA|4|2|in die illa erit germen Domini in magnificentia et in gloria et fructus terrae sublimis et exultatio his qui salvati fuerint de Israhel
ISA|4|3|et erit omnis qui relictus fuerit in Sion et residuus in Hierusalem sanctus vocabitur omnis qui scriptus est in vita in Hierusalem
ISA|4|4|si abluerit Dominus sordem filiarum Sion et sanguinem Hierusalem laverit de medio eius spiritu iudicii et spiritu ardoris
ISA|4|5|et creabit Dominus super omnem locum montis Sion et ubi invocatus est nubem per diem et fumum et splendorem ignis flammantis in nocte super omnem enim gloriam protectio
ISA|4|6|et tabernaculum erit in umbraculum diei ab aestu et in securitatem et absconsionem a turbine et a pluvia
ISA|5|1|cantabo dilecto meo canticum patruelis mei vineae suae vinea facta est dilecto meo in cornu filio olei
ISA|5|2|et sepivit eam et lapides elegit ex illa et plantavit eam electam et aedificavit turrem in medio eius et torcular extruxit in ea et expectavit ut faceret uvas et fecit labruscas
ISA|5|3|nunc ergo habitator Hierusalem et vir Iuda iudicate inter me et inter vineam meam
ISA|5|4|quid est quod debui ultra facere vineae meae et non feci ei an quod expectavi ut faceret uvas et fecit labruscas
ISA|5|5|et nunc ostendam vobis quid ego faciam vineae meae auferam sepem eius et erit in direptionem diruam maceriam eius et erit in conculcationem
ISA|5|6|et ponam eam desertam non putabitur et non fodietur et ascendent vepres et spinae et nubibus mandabo ne pluant super eam imbrem
ISA|5|7|vinea enim Domini exercituum domus Israhel et vir Iuda germen delectabile eius et expectavi ut faceret iudicium et ecce iniquitas et iustitiam et ecce clamor
ISA|5|8|vae qui coniungitis domum ad domum et agrum agro copulatis usque ad terminum loci numquid habitabitis soli vos in medio terrae
ISA|5|9|in auribus meis sunt haec Domini exercituum nisi domus multae desertae fuerint grandes et pulchrae absque habitatore
ISA|5|10|decem enim iuga vinearum facient lagunculam unam et triginta modii sementis facient modios tres
ISA|5|11|vae qui consurgitis mane ad ebrietatem sectandam et potandum usque ad vesperam ut vino aestuetis
ISA|5|12|cithara et lyra et tympanum et tibia et vinum in conviviis vestris et opus Domini non respicitis nec opera manuum eius consideratis
ISA|5|13|propterea captivus ductus est populus meus quia non habuit scientiam et nobiles eius interierunt fame et multitudo eius siti exaruit
ISA|5|14|propterea dilatavit infernus animam suam et aperuit os suum absque ullo termino et descendent fortes eius et populus eius et sublimes gloriosique eius ad eum
ISA|5|15|et incurvabitur homo et humiliabitur vir et oculi sublimium deprimentur
ISA|5|16|et exaltabitur Dominus exercituum in iudicio et Deus sanctus sanctificabitur in iustitia
ISA|5|17|et pascentur agni iuxta ordinem suum et deserta in ubertatem versa advenae comedent
ISA|5|18|vae qui trahitis iniquitatem in funiculis vanitatis et quasi vinculum plaustri peccatum
ISA|5|19|qui dicitis festinet et cito veniat opus eius ut videamus et adpropiet et veniat consilium Sancti Israhel et sciemus illud
ISA|5|20|vae qui dicitis malum bonum et bonum malum ponentes tenebras lucem et lucem tenebras ponentes amarum in dulce et dulce in amarum
ISA|5|21|vae qui sapientes estis in oculis vestris et coram vobismet ipsis prudentes
ISA|5|22|vae qui potentes estis ad bibendum vinum et viri fortes ad miscendam ebrietatem
ISA|5|23|qui iustificatis impium pro muneribus et iustitiam iusti aufertis ab eo
ISA|5|24|propter hoc sicut devorat stipulam lingua ignis et calor flammae exurit sic radix eorum quasi favilla erit et germen eorum ut pulvis ascendet abiecerunt enim legem Domini exercituum et eloquium Sancti Israhel blasphemaverunt
ISA|5|25|ideo iratus est furor Domini in populo suo et extendit manum suam super eum et percussit eum et conturbati sunt montes et facta sunt morticina eorum quasi stercus in medio platearum in omnibus his non est aversus furor eius sed adhuc manus eius extenta
ISA|5|26|et levabit signum nationibus procul et sibilabit ad eum de finibus terrae et ecce festinus velociter veniet
ISA|5|27|non est deficiens neque laborans in eo non dormitabit neque dormiet neque solvetur cingulum renum eius nec rumpetur corrigia calciamenti eius
ISA|5|28|sagittae eius acutae et omnes arcus eius extenti ungulae equorum eius ut silex et rotae eius quasi impetus tempestatis
ISA|5|29|rugitus eius ut leonis rugiet ut catuli leonum et frendet et tenebit praedam et amplexabitur et non erit qui eruat
ISA|5|30|et sonabit super eum in die illa sicut sonitus maris aspiciemus in terram et ecce tenebrae tribulationis et lux obtenebrata est in caligine eius
ISA|6|1|in anno quo mortuus est rex Ozias vidi Dominum sedentem super solium excelsum et elevatum et ea quae sub eo erant implebant templum
ISA|6|2|seraphin stabant super illud sex alae uni et sex alae alteri duabus velabant faciem eius et duabus velabant pedes eius et duabus volabant
ISA|6|3|et clamabant alter ad alterum et dicebant sanctus sanctus sanctus Dominus exercituum plena est omnis terra gloria eius
ISA|6|4|et commota sunt superliminaria cardinum a voce clamantis et domus impleta est fumo
ISA|6|5|et dixi vae mihi quia tacui quia vir pollutus labiis ego sum et in medio populi polluta labia habentis ego habito et Regem Dominum exercituum vidi oculis meis
ISA|6|6|et volavit ad me unus de seraphin et in manu eius calculus quem forcipe tulerat de altari
ISA|6|7|et tetigit os meum et dixit ecce tetigit hoc labia tua et auferetur iniquitas tua et peccatum tuum mundabitur
ISA|6|8|et audivi vocem Domini dicentis quem mittam et quis ibit nobis et dixi ecce ego sum mitte me
ISA|6|9|et dixit vade et dices populo huic audite audientes et nolite intellegere et videte visionem et nolite cognoscere
ISA|6|10|excaeca cor populi huius et aures eius adgrava et oculos eius claude ne forte videat oculis suis et auribus suis audiat et corde suo intellegat et convertatur et sanem eum
ISA|6|11|et dixi usquequo Domine et dixit donec desolentur civitates absque habitatore et domus sine homine et terra relinquetur deserta
ISA|6|12|et longe faciet Dominus homines et multiplicabitur quae derelicta fuerat in medio terrae
ISA|6|13|et adhuc in ea decimatio et convertetur et erit in ostensionem sicut terebinthus et sicuti quercus quae expandit ramos suos semen sanctum erit id quod steterit in ea
ISA|7|1|et factum est in diebus Ahaz filii Ioatham filii Oziae regis Iuda ascendit Rasin rex Syriae et Phacee filius Romeliae rex Israhel in Hierusalem ad proeliandum contra eam et non potuerunt debellare eam
ISA|7|2|et nuntiaverunt domui David dicentes requievit Syria super Ephraim et commotum est cor eius et cor populi eius sicut moventur ligna silvarum a facie venti
ISA|7|3|et dixit Dominus ad Isaiam egredere in occursum Ahaz tu et qui derelictus est Iasub filius tuus ad extremum aquaeductus piscinae superioris in via agri Fullonis
ISA|7|4|et dices ad eum vide ut sileas noli timere et cor tuum ne formidet a duobus caudis titionum fumigantium istorum in ira furoris Rasin et Syriae et filii Romeliae
ISA|7|5|eo quod consilium inierit contra te Syria malum Ephraim et filius Romeliae dicentes
ISA|7|6|ascendamus ad Iudam et suscitemus eum et avellamus eum ad nos et ponamus regem in medio eius filium Tabeel
ISA|7|7|haec dicit Dominus Deus non stabit et non erit istud
ISA|7|8|sed caput Syriae Damascus et caput Damasci Rasin et adhuc sexaginta et quinque anni et desinet Ephraim esse populus
ISA|7|9|et caput Ephraim Samaria et caput Samariae filius Romeliae si non credideritis non permanebitis
ISA|7|10|et adiecit Dominus loqui ad Ahaz dicens
ISA|7|11|pete tibi signum a Domino Deo tuo in profundum inferni sive in excelsum supra
ISA|7|12|et dixit Ahaz non petam et non temptabo Dominum
ISA|7|13|et dixit audite ergo domus David numquid parum vobis est molestos esse hominibus quia molesti estis et Deo meo
ISA|7|14|propter hoc dabit Dominus ipse vobis signum ecce virgo concipiet et pariet filium et vocabitis nomen eius Emmanuhel
ISA|7|15|butyrum et mel comedet ut sciat reprobare malum et eligere bonum
ISA|7|16|quia antequam sciat puer reprobare malum et eligere bonum derelinquetur terra quam tu detestaris a facie duum regum suorum
ISA|7|17|adducet Dominus super te et super populum tuum et super domum patris tui dies qui non venerunt a diebus separationis Ephraim a Iuda cum rege Assyriorum
ISA|7|18|et erit in die illa sibilabit Dominus muscae quae est in extremo fluminum Aegypti et api quae est in terra Assur
ISA|7|19|et venient et requiescent omnes in torrentibus vallium et cavernis petrarum et in omnibus frutectis et in universis foraminibus
ISA|7|20|in die illa radet Dominus in novacula conducta in his qui trans Flumen sunt in rege Assyriorum caput et pilos pedum et barbam universam
ISA|7|21|et erit in die illa nutriet homo vaccam boum et duas oves
ISA|7|22|et prae ubertate lactis comedet butyrum butyrum enim et mel manducabit omnis qui relictus fuerit in medio terrae
ISA|7|23|et erit in die illa omnis locus ubi fuerint mille vites mille argenteis et in spinas et in vepres erunt
ISA|7|24|cum sagittis et arcu ingredientur illuc vepres enim et spinae erunt in universa terra
ISA|7|25|et omnes montes qui in sarculo sarientur non veniet illuc terror spinarum et veprium et erit in pascua bovis et in conculcationem pecoris
ISA|8|1|et dixit Dominus ad me sume tibi librum grandem et scribe in eo stilo hominis Velociter spolia detrahe Cito praedare
ISA|8|2|et adhibui mihi testes fideles Uriam sacerdotem et Zacchariam filium Barachiae
ISA|8|3|et accessi ad prophetissam et concepit et peperit filium et dixit Dominus ad me voca nomen eius Adcelera spolia detrahere Festina praedari
ISA|8|4|quia antequam sciat puer vocare patrem suum et matrem suam auferetur fortitudo Damasci et spolia Samariae coram rege Assyriorum
ISA|8|5|et adiecit Dominus loqui ad me adhuc dicens
ISA|8|6|pro eo quod abiecit populus iste aquas Siloae quae vadunt cum silentio et adsumpsit magis Rasin et filium Romeliae
ISA|8|7|propter hoc ecce Dominus adducet super eos aquas Fluminis fortes et multas regem Assyriorum et omnem gloriam eius et ascendet super omnes rivos eius et fluet super universas ripas eius
ISA|8|8|et ibit per Iudam inundans et transiens usque ad collum veniet et erit extensio alarum eius implens latitudinem terrae tuae o Emmanuhel
ISA|8|9|congregamini populi et vincimini et audite universae procul terrae confortamini et vincimini accingite vos et vincimini
ISA|8|10|inite consilium et dissipabitur loquimini verbum et non fiet quia nobiscum Deus
ISA|8|11|haec enim ait Dominus ad me sicut in forti manu erudivit me ne irem in via populi huius dicens
ISA|8|12|non dicatis coniuratio omnia enim quae loquitur populus iste coniuratio est et timorem eius ne timeatis neque paveatis
ISA|8|13|Dominum exercituum ipsum sanctificate ipse pavor vester et ipse terror vester
ISA|8|14|et erit vobis in sanctificationem in lapidem autem offensionis et in petram scandali duabus domibus Israhel in laqueum et in ruinam habitantibus Hierusalem
ISA|8|15|et offendent ex eis plurimi et cadent et conterentur et inretientur et capientur
ISA|8|16|liga testimonium signa legem in discipulis meis
ISA|8|17|et expectabo Dominum qui abscondit faciem suam a domo Iacob et praestolabor eum
ISA|8|18|ecce ego et pueri quos mihi dedit Dominus in signum et in portentum Israhelis a Domino exercituum qui habitat in monte Sion
ISA|8|19|et cum dixerint ad vos quaerite a pythonibus et a divinis qui stridunt in incantationibus suis numquid non populus a Deo suo requirit pro vivis a mortuis
ISA|8|20|ad legem magis et ad testimonium quod si non dixerint iuxta verbum hoc non erit eis matutina lux
ISA|8|21|et transibit per eam corruet et esuriet et cum esurierit irascetur et maledicet regi suo et Deo suo et suspiciet sursum
ISA|8|22|et ad terram intuebitur et ecce tribulatio et tenebrae dissolutio angustia et caligo persequens et non poterit avolare de angustia sua
ISA|9|1|primo tempore adleviata est terra Zabulon et terra Nepthalim et novissimo adgravata est via maris trans Iordanem Galileae gentium
ISA|9|2|populus qui ambulabat in tenebris vidit lucem magnam habitantibus in regione umbrae mortis lux orta est eis
ISA|9|3|multiplicasti gentem non magnificasti laetitiam laetabuntur coram te sicut laetantur in messe sicut exultant quando dividunt spolia
ISA|9|4|iugum enim oneris eius et virgam umeri eius et sceptrum exactoris eius superasti sicut in die Madian
ISA|9|5|quia omnis violenta praedatio cum tumultu et vestimentum mixtum sanguine erit in conbustionem et cibus ignis
ISA|9|6|parvulus enim natus est nobis filius datus est nobis et factus est principatus super umerum eius et vocabitur nomen eius Admirabilis consiliarius Deus fortis Pater futuri saeculi Princeps pacis
ISA|9|7|multiplicabitur eius imperium et pacis non erit finis super solium David et super regnum eius ut confirmet illud et corroboret in iudicio et iustitia amodo et usque in sempiternum zelus Domini exercituum faciet hoc
ISA|9|8|verbum misit Dominus in Iacob et cecidit in Israhel
ISA|9|9|et sciet populus omnis Ephraim et habitantes Samariam in superbia et magnitudine cordis dicentes
ISA|9|10|lateres ceciderunt sed quadris lapidibus aedificabimus sycomoros succiderunt sed cedros inmutabimus
ISA|9|11|et elevabit Dominus hostes Rasin super eum et inimicos eius in tumultum vertet
ISA|9|12|Syriam ab oriente et Philisthim ab occidente et devorabunt Israhel toto ore in omnibus his non est aversus furor eius sed adhuc manus eius extenta
ISA|9|13|et populus non est reversus ad percutientem se et Dominum exercituum non inquisierunt
ISA|9|14|et disperdet Dominus ab Israhel caput et caudam incurvantem et refrenantem die una
ISA|9|15|longevus et honorabilis ipse est caput et propheta docens mendacium ipse cauda est
ISA|9|16|et erunt qui beatificant populum istum seducentes et qui beatificantur praecipitati
ISA|9|17|propter hoc super adulescentulis eius non laetabitur Dominus et pupillorum eius et viduarum non miserebitur quia omnis hypocrita est et nequam et universum os locutum est stultitiam in omnibus his non est aversus furor eius sed adhuc manus eius extenta
ISA|9|18|succensa est enim quasi ignis impietas veprem et spinam vorabit et succendetur in densitate saltus et convolvetur superbia fumi
ISA|9|19|in ira Domini exercituum conturbata est terra et erit populus quasi esca ignis vir fratri suo non parcet
ISA|9|20|et declinabit ad dexteram et esuriet et comedet ad sinistram et non saturabitur unusquisque carnem brachii sui vorabit Manasses Ephraim et Ephraim Manassen simul ipsi contra Iudam
ISA|9|21|in omnibus his non est aversus furor eius sed adhuc manus eius extenta
ISA|10|1|vae qui condunt leges iniquas et scribentes iniustitiam scripserunt
ISA|10|2|ut opprimerent in iudicio pauperes et vim facerent causae humilium populi mei ut essent viduae praeda eorum et pupillos diriperent
ISA|10|3|quid facietis in die visitationis et calamitatis de longe venientis ad cuius fugietis auxilium et ubi derelinquetis gloriam vestram
ISA|10|4|ne incurvemini sub vinculo et cum interfectis cadatis super omnibus his non est aversus furor eius sed adhuc manus eius extenta
ISA|10|5|vae Assur virga furoris mei et baculus ipse in manu eorum indignatio mea
ISA|10|6|ad gentem fallacem mittam eum et contra populum furoris mei mandabo illi ut auferat spolia et diripiat praedam et ponat illum in conculcationem quasi lutum platearum
ISA|10|7|ipse autem non sic arbitrabitur et cor eius non ita aestimabit sed ad conterendum erit cor eius et ad internicionem gentium non paucarum
ISA|10|8|dicet enim
ISA|10|9|numquid non principes mei simul reges sunt numquid non ut Charchamis sic Chalanno et ut Arfad sic Emath numquid non ut Damascus sic Samaria
ISA|10|10|quomodo invenit manus mea regna idoli sic et simulacra eorum de Hierusalem et de Samaria
ISA|10|11|numquid non sicut feci Samariae et idolis eius sic faciam Hierusalem et simulacris eius
ISA|10|12|et erit cum impleverit Dominus cuncta opera sua in monte Sion et in Hierusalem visitabo super fructum magnifici cordis regis Assur et super gloriam altitudinis oculorum eius
ISA|10|13|dixit enim in fortitudine manus meae feci et in sapientia mea intellexi et abstuli terminos populorum et principes eorum depraedatus sum et detraxi quasi potens in sublime residentes
ISA|10|14|et invenit quasi nidum manus mea fortitudinem populorum et sicut colliguntur ova quae derelicta sunt sic universam terram ego congregavi et non fuit qui moveret pinnam et aperiret os et ganniret
ISA|10|15|numquid gloriabitur securis contra eum qui secat in ea aut exaltabitur serra contra eum a quo trahitur quomodo si elevetur virga contra levantem se et exaltetur baculus qui utique lignum est
ISA|10|16|propter hoc mittet Dominator Deus exercituum in pinguibus eius tenuitatem et subtus gloriam eius succensa ardebit quasi conbustio ignis
ISA|10|17|et erit lumen Israhel in igne et Sanctus eius in flamma et succendetur et devorabitur spina eius et vepres in die una
ISA|10|18|et gloria saltus eius et Carmeli eius ab anima usque ad carnem consumetur et erit terrore profugus
ISA|10|19|et reliquiae ligni saltus eius pro paucitate numerabuntur et puer scribet eos
ISA|10|20|et erit in die illa non adiciet residuum Israhel et hii qui fugerint de domo Iacob inniti super eo qui percutit eos sed innitetur super Dominum Sanctum Israhel in veritate
ISA|10|21|reliquiae convertentur reliquiae inquam Iacob ad Deum fortem
ISA|10|22|si enim fuerit populus tuus Israhel quasi harena maris reliquiae convertentur ex eo consummatio adbreviata inundabit iustitiam
ISA|10|23|consummationem enim et adbreviationem Dominus Deus exercituum faciet in medio omnis terrae
ISA|10|24|propter hoc haec dicit Dominus Deus exercituum noli timere populus meus habitator Sion ab Assur in virga percutiet te et baculum suum levabit super te in via Aegypti
ISA|10|25|adhuc enim paululum modicumque et consummabitur indignatio et furor meus super scelus eorum
ISA|10|26|et suscitabit super eum Dominus exercituum flagellum iuxta plagam Madian in petra Oreb et virgam suam super mare et levabit eam in via Aegypti
ISA|10|27|et erit in die illa auferetur onus eius de umero tuo et iugum eius de collo tuo et conputrescet iugum a facie olei
ISA|10|28|veniet in Aiath transibit in Magron apud Machmas commendabit vasa sua
ISA|10|29|transierunt cursim Gabee sedes nostra obstipuit Rama Gabaath Saulis fugit
ISA|10|30|hinni voce tua filia Gallim adtende Laisa paupercula Anathoth
ISA|10|31|migravit Medemena habitatores Gebim confortamini
ISA|10|32|adhuc dies est ut in Nob stetur agitabit manum suam super montem filiae Sion collem Hierusalem
ISA|10|33|ecce Dominator Dominus exercituum confringet lagunculam in terrore et excelsi statura succidentur et sublimes humiliabuntur
ISA|10|34|et subvertentur condensa saltus ferro et Libanus cum excelsis cadet
ISA|11|1|et egredietur virga de radice Iesse et flos de radice eius ascendet
ISA|11|2|et requiescet super eum spiritus Domini spiritus sapientiae et intellectus spiritus consilii et fortitudinis spiritus scientiae et pietatis
ISA|11|3|et replebit eum spiritus timoris Domini non secundum visionem oculorum iudicabit neque secundum auditum aurium arguet
ISA|11|4|sed iudicabit in iustitia pauperes et arguet in aequitate pro mansuetis terrae et percutiet terram virga oris sui et spiritu labiorum suorum interficiet impium
ISA|11|5|et erit iustitia cingulum lumborum eius et fides cinctorium renis eius
ISA|11|6|habitabit lupus cum agno et pardus cum hedo accubabit vitulus et leo et ovis simul morabuntur et puer parvulus minabit eos
ISA|11|7|vitulus et ursus pascentur simul requiescent catuli eorum et leo quasi bos comedet paleas
ISA|11|8|et delectabitur infans ab ubere super foramine aspidis et in caverna reguli qui ablactatus fuerit manum suam mittet
ISA|11|9|non nocebunt et non occident in universo monte sancto meo quia repleta est terra scientia Domini sicut aquae maris operientes
ISA|11|10|in die illa radix Iesse qui stat in signum populorum ipsum gentes deprecabuntur et erit sepulchrum eius gloriosum
ISA|11|11|et erit in die illa adiciet Dominus secundo manum suam ad possidendum residuum populi sui quod relinquetur ab Assyriis et ab Aegypto et a Fetros et ab Aethiopia et ab Aelam et a Sennaar et ab Emath et ab insulis maris
ISA|11|12|et levabit signum in nationes et congregabit profugos Israhel et dispersos Iuda colliget a quattuor plagis terrae
ISA|11|13|et auferetur zelus Ephraim et hostes Iuda peribunt Ephraim non aemulabitur Iudam et Iudas non pugnabit contra Ephraim
ISA|11|14|et volabunt in umeros Philisthim per mare simul praedabuntur filios orientis Idumea et Moab praeceptum manus eorum et filii Ammon oboedientes erunt
ISA|11|15|et desolabit Dominus linguam maris Aegypti et levabit manum suam super Flumen in fortitudine spiritus sui et percutiet eum in septem rivis ita ut transeant per eum calciati
ISA|11|16|et erit via residuo populo meo qui relinquetur ab Assyriis sicut fuit Israhel in die qua ascendit de terra Aegypti
ISA|12|1|et dices in illa die confitebor tibi Domine quoniam iratus es mihi conversus est furor tuus et consolatus es me
ISA|12|2|ecce Deus salvator meus fiducialiter agam et non timebo quia fortitudo mea et laus mea Dominus Deus et factus est mihi in salutem
ISA|12|3|haurietis aquas in gaudio de fontibus salvatoris
ISA|12|4|et dicetis in illa die confitemini Domino et invocate nomen eius notas facite in populis adinventiones eius mementote quoniam excelsum est nomen eius
ISA|12|5|cantate Domino quoniam magnifice fecit adnuntiate hoc in universa terra
ISA|12|6|exulta et lauda habitatio Sion quia magnus in medio tui Sanctus Israhel
ISA|13|1|onus Babylonis quod vidit Isaias filius Amos
ISA|13|2|super montem caligosum levate signum exaltate vocem levate manum et ingrediantur portas duces
ISA|13|3|ego mandavi sanctificatis meis et vocavi fortes meos in ira mea exultantes in gloria mea
ISA|13|4|vox multitudinis in montibus quasi populorum frequentium vox sonitus regum gentium congregatarum Dominus exercituum praecepit militiae belli
ISA|13|5|venientibus de terra procul a summitate caeli Dominus et vasa furoris eius ut disperdat omnem terram
ISA|13|6|ululate quia prope est dies Domini quasi vastitas a Domino veniet
ISA|13|7|propter hoc omnes manus dissolventur et omne cor hominis tabescet
ISA|13|8|et conteretur tortiones et dolores tenebunt quasi parturiens dolebunt unusquisque ad proximum suum stupebit facies conbustae vultus eorum
ISA|13|9|ecce dies Domini venit crudelis et indignationis plenus et irae furorisque ad ponendam terram in solitudine et peccatores eius conterendos de ea
ISA|13|10|quoniam stellae caeli et splendor earum non expandent lumen suum obtenebratus est sol in ortu suo et luna non splendebit in lumine suo
ISA|13|11|et visitabo super orbis mala et contra impios iniquitatem eorum et quiescere faciam superbiam infidelium et arrogantiam fortium humiliabo
ISA|13|12|pretiosior erit vir auro et homo mundo obrizo
ISA|13|13|super hoc caelum turbabo et movebitur terra de loco suo propter indignationem Domini exercituum et propter diem irae furoris eius
ISA|13|14|et erit quasi dammula fugiens et quasi ovis et non erit qui congreget unusquisque ad populum suum convertetur et singuli ad terram suam fugient
ISA|13|15|omnis qui inventus fuerit occidetur et omnis qui supervenerit cadet in gladio
ISA|13|16|infantes eorum adlident in oculis eorum diripientur domus eorum et uxores eorum violabuntur
ISA|13|17|ecce ego suscitabo super eos Medos qui argentum non quaerant nec aurum velint
ISA|13|18|sed sagittis parvulos interficiant et lactantibus uteri non misereantur et super filios non parcat oculus eorum
ISA|13|19|et erit Babylon illa gloriosa in regnis inclita in superbia Chaldeorum sicut subvertit Deus Sodomam et Gomorram
ISA|13|20|non habitabitur usque in finem et non fundabitur usque ad generationem et generationem nec ponet ibi tentoria Arabs nec pastores requiescent ibi
ISA|13|21|sed requiescent ibi bestiae et replebuntur domus eorum draconibus et habitabunt ibi strutiones et pilosi saltabunt ibi
ISA|13|22|et respondebunt ibi ululae in aedibus eius et sirenae in delubris voluptatis
ISA|14|1|prope est ut veniat tempus eius et dies eius non elongabuntur miserebitur enim Dominus Iacob et eliget adhuc de Israhel et requiescere eos faciet super humum suam adiungetur advena ad eos et adherebit domui Iacob
ISA|14|2|et tenebunt eos populi et adducent eos in locum suum et possidebit eos domus Israhel super terram Domini in servos et ancillas et erunt capientes eos qui se ceperant et subicient exactores suos
ISA|14|3|et erit in die illa cum requiem dederit tibi Deus a labore tuo et a concussione tua et a servitute dura qua ante servisti
ISA|14|4|sumes parabolam istam contra regem Babylonis et dices quomodo cessavit exactor quievit tributum
ISA|14|5|contrivit Dominus baculum impiorum virgam dominantium
ISA|14|6|caedentem populos in indignatione plaga insanabili subicientem in furore gentes persequentem crudeliter
ISA|14|7|conquievit et siluit omnis terra gavisa est et exultavit
ISA|14|8|abietes quoque laetatae sunt super te et cedri Libani ex quo dormisti non ascendit qui succidat nos
ISA|14|9|infernus subter conturbatus est in occursum adventus tui suscitavit tibi gigantas omnes principes terrae surrexerunt de soliis suis omnes principes nationum
ISA|14|10|universi respondebunt et dicent tibi et tu vulneratus es sicut nos nostri similis effectus es
ISA|14|11|detracta est ad inferos superbia tua concidit cadaver tuum subter te sternetur tinea et operimentum tuum erunt vermes
ISA|14|12|quomodo cecidisti de caelo lucifer qui mane oriebaris corruisti in terram qui vulnerabas gentes
ISA|14|13|qui dicebas in corde tuo in caelum conscendam super astra Dei exaltabo solium meum sedebo in monte testamenti in lateribus aquilonis
ISA|14|14|ascendam super altitudinem nubium ero similis Altissimo
ISA|14|15|verumtamen ad infernum detraheris in profundum laci
ISA|14|16|qui te viderint ad te inclinabuntur teque prospicient numquid iste est vir qui conturbavit terram qui concussit regna
ISA|14|17|qui posuit orbem desertum et urbes eius destruxit vinctis eius non aperuit carcerem
ISA|14|18|omnes reges gentium universi dormierunt in gloria vir in domo sua
ISA|14|19|tu autem proiectus es de sepulchro tuo quasi stirps inutilis pollutus et obvolutus qui interfecti sunt gladio et descenderunt ad fundamenta laci quasi cadaver putridum
ISA|14|20|non habebis consortium neque cum eis in sepultura tu enim terram disperdisti tu populum occidisti non vocabitur in aeternum semen pessimorum
ISA|14|21|praeparate filios eius occisioni in iniquitate patrum eorum non consurgent nec hereditabunt terram neque implebunt faciem orbis civitatum
ISA|14|22|et consurgam super eos dicit Dominus exercituum et perdam Babylonis nomen et reliquias et germen et progeniem ait Dominus
ISA|14|23|et ponam eam in possessionem ericii et in paludes aquarum et scopabo eam in scopa terens dicit Dominus exercituum
ISA|14|24|iuravit Dominus exercituum dicens si non ut putavi ita erit et quomodo mente tractavi
ISA|14|25|sic eveniet ut conteram Assyrium in terra mea et in montibus meis conculcem eum et auferetur ab eis iugum eius et onus illius ab umero eorum tolletur
ISA|14|26|hoc consilium quod cogitavi super omnem terram et haec est manus extenta super universas gentes
ISA|14|27|Dominus enim exercituum decrevit et quis poterit infirmare et manus eius extenta et quis avertet eam
ISA|14|28|in anno quo mortuus est rex Ahaz factum est onus istud
ISA|14|29|ne laeteris Philisthea omnis tu quoniam comminuta est virga percussoris tui de radice enim colubri egredietur regulus et semen eius absorbens volucrem
ISA|14|30|et pascentur primogeniti pauperum et pauperes fiducialiter requiescent et interire faciam in fame radicem tuam et reliquias tuas interficiam
ISA|14|31|ulula porta clama civitas prostrata est Philisthea omnis ab aquilone enim fumus venit et non est qui effugiat agmen eius
ISA|14|32|et quid respondebitur nuntiis gentis quia Dominus fundavit Sion et in ipsa sperabunt pauperes populi eius
ISA|15|1|onus Moab quia nocte vastata est Ar Moab conticuit quia nocte vastatus est murus Moab conticuit
ISA|15|2|ascendit domus et Dibon ad excelsa in planctum super Nabo et super Medaba Moab ululabit in cunctis capitibus eius calvitium omnis barba radetur
ISA|15|3|in triviis eius accincti sunt sacco super tecta eius et in plateis eius omnis ululat descendit in fletum
ISA|15|4|clamavit Esebon et Eleale usque Iasa audita est vox eorum super hoc expediti Moab ululabunt anima eius ululabit sibi
ISA|15|5|cor meum ad Moab clamabit vectes eius usque ad Segor vitulam conternantem per ascensum enim Luith flens ascendet et in via Oronaim clamorem contritionis levabunt
ISA|15|6|aquae enim Nemrim desertae erunt quia aruit herba defecit germen viror omnis interiit
ISA|15|7|secundum magnitudinem operis et visitatio eorum ad torrentem salicum ducent eos
ISA|15|8|quoniam circumiit clamor terminum Moab usque ad Gallim ululatus eius et usque ad puteum Helim clamor eius
ISA|15|9|quia aquae Dibon repletae sunt sanguine ponam enim super Dibon additamenta his qui fugerint de Moab leonem et reliquiis terrae
ISA|16|1|emitte agnum dominatorem terrae de Petra deserti ad montem filiae Sion
ISA|16|2|et erit sicut avis fugiens et pulli de nido avolantes sic erunt filiae Moab in transcensu Arnon
ISA|16|3|ini consilium coge concilium pone quasi noctem umbram tuam in meridie absconde fugientes et vagos ne prodas
ISA|16|4|habitabunt apud te profugi mei Moab esto latibulum eorum a facie vastatoris finitus est enim pulvis consummatus est miser defecit qui conculcabat terram
ISA|16|5|et praeparabitur in misericordia solium et sedebit super eum in veritate in tabernaculo David iudicans et quaerens iudicium et velociter reddens quod iustum est
ISA|16|6|audivimus superbiam Moab superbus est valde superbia eius et arrogantia eius et indignatio eius plus quam fortitudo eius
ISA|16|7|idcirco ululabit Moab ad Moab universus ululabit his qui laetantur super muro cocti lateris loquimini plagas suas
ISA|16|8|quoniam suburbana Esebon deserta sunt et vinea Sabama domini gentium exciderunt flagella eius usque ad Iazer pervenerunt erraverunt in deserto propagines eius relictae sunt transierunt mare
ISA|16|9|super hoc plorabo in fletu Iazer vineam Sabama inebriabo te lacrima mea Esebon et Eleale quoniam super vindemiam tuam et super messem tuam vox calcantium inruit
ISA|16|10|et auferetur laetitia et exultatio de Carmelo et in vineis non exultabit neque iubilabit vinum in torculari non calcabit qui calcare consueverat vocem calcantium abstuli
ISA|16|11|super hoc venter meus ad Moab quasi cithara sonabit et viscera mea ad murum cocti lateris
ISA|16|12|et erit cum apparuerit quod laboravit Moab super excelsis suis ingredietur ad sancta sua ut obsecret et non valebit
ISA|16|13|hoc verbum quod locutus est Dominus ad Moab ex tunc
ISA|16|14|et nunc locutus est Dominus dicens in tribus annis quasi anni mercennarii auferetur gloria Moab super omni populo multo et relinquetur parvus et modicus nequaquam multus
ISA|17|1|onus Damasci ecce Damascus desinet esse civitas et erit sicut acervus lapidum in ruina
ISA|17|2|derelictae civitates Aroer gregibus erunt et requiescent ibi et non erit qui exterreat
ISA|17|3|et cessabit adiutorium ab Ephraim et regnum a Damasco et reliquiae Syriae sicut gloria filiorum Israhel erunt dicit Dominus exercituum
ISA|17|4|et erit in die illa adtenuabitur gloria Iacob et pingue carnis eius marcescet
ISA|17|5|et erit sicut congregans in messe quod restiterit et brachium eius spicas leget et erit sicut quaerens spicas in valle Rafaim
ISA|17|6|et relinquetur in eo sicut racemus et sicut excussio oleae duarum aut trium olivarum in summitate rami sive quattuor aut quinque in cacuminibus eius fructus eius dicit Dominus Deus Israhel
ISA|17|7|in die illa inclinabitur homo ad factorem suum et oculi eius ad Sanctum Israhel respicient
ISA|17|8|et non inclinabitur ad altaria quae fecerunt manus eius et quae operati sunt digiti eius non respiciet lucos et delubra
ISA|17|9|in die illa erunt civitates fortitudinis eius derelictae sicut aratra et segetes quae derelictae sunt a facie filiorum Israhel et erit deserta
ISA|17|10|quia oblita es Dei salvatoris tui et Fortis adiutoris tui non es recordata propterea plantabis plantationem fidelem et germen alienum seminabis
ISA|17|11|in die plantationis tuae labrusca et mane semen tuum florebit ablata est messis in die hereditatis et dolebit graviter
ISA|17|12|vae multitudo populorum multorum ut multitudo maris sonantis et tumultus turbarum sicut sonitus aquarum multarum
ISA|17|13|sonabunt populi sicut sonitus aquarum inundantium et increpabit eum et fugiet procul et rapietur sicut pulvis montium a facie venti et sicut turbo coram tempestate
ISA|17|14|in tempore vespere et ecce turbatio in matutino et non subsistet haec est pars eorum qui vastaverunt nos et sors diripientium nos
ISA|18|1|vae terrae cymbalo alarum quae est trans flumina Aethiopiae
ISA|18|2|qui mittit in mari legatos et in vasis papyri super aquas ite angeli veloces ad gentem convulsam et dilaceratam ad populum terribilem post quem non est alius gentem expectantem expectantem et conculcatam cuius diripuerunt flumina terram eius
ISA|18|3|omnes habitatores orbis qui moramini in terra cum elevatum fuerit signum in montibus videbitis et clangorem tubae audietis
ISA|18|4|quia haec dicit Dominus ad me quiescam et considerabo in loco meo sicut meridiana lux clara est et sicut nubes roris in die messis
ISA|18|5|ante messem enim totus effloruit et inmatura perfectio germinabit et praecidentur ramusculi eius falcibus et quae derelicta fuerint abscidentur excutientur
ISA|18|6|et relinquentur simul avibus montium et bestiis terrae et aestate perpetua erunt super eum volucres et omnes bestiae terrae super illum hiemabunt
ISA|18|7|in tempore illo deferetur munus Domino exercituum a populo divulso et dilacerato a populo terribili post quem non fuit alius a gente expectante expectante et conculcata cuius diripuerunt flumina terram eius ad locum nominis Domini exercituum montem Sion
ISA|19|1|onus Aegypti ecce Dominus ascendet super nubem levem et ingredietur Aegyptum et movebuntur simulacra Aegypti a facie eius et cor Aegypti tabescet in medio eius
ISA|19|2|et concurrere faciam Aegyptios adversum Aegyptios et pugnabit vir contra fratrem suum et vir contra amicum suum civitas adversus civitatem regnum adversus regnum
ISA|19|3|et disrumpetur spiritus Aegypti in visceribus eius et consilium eius praecipitabo et interrogabunt simulacra sua et divinos suos et pythones et ariolos
ISA|19|4|et tradam Aegyptum in manu dominorum crudelium et rex fortis dominabitur eorum ait Dominus Deus exercituum
ISA|19|5|et arescet aqua de mari et fluvius desolabitur atque siccabitur
ISA|19|6|et deficient flumina adtenuabuntur et siccabuntur rivi aggerum calamus et iuncus marcescet
ISA|19|7|nudabitur alveus rivi a fonte suo et omnis sementis inrigua siccabitur arescet et non erit
ISA|19|8|et maerebunt piscatores et lugebunt omnes mittentes in flumen hamum et expandentes rete super faciem aquae marcescent
ISA|19|9|confundentur qui operabantur linum pectentes et texentes subtilia
ISA|19|10|et erunt inrigua eius flaccentia omnes qui faciebant lacunas ad capiendos pisces
ISA|19|11|stulti principes Taneos sapientes consiliarii Pharao dederunt consilium insipiens quomodo dicetis Pharaoni filius sapientium ego filius regum antiquorum
ISA|19|12|ubi sunt nunc sapientes tui adnuntient tibi et indicent quid cogitaverit Dominus exercituum super Aegyptum
ISA|19|13|stulti facti sunt principes Taneos emarcuerunt principes Mempheos deceperunt Aegyptum angulum populorum eius
ISA|19|14|Dominus miscuit in medio eius spiritum vertiginis et errare fecerunt Aegyptum in omni opere suo sicut errat ebrius et vomens
ISA|19|15|et non erit Aegypto opus quod faciat caput et caudam incurvantem et refrenantem
ISA|19|16|in die illa erit Aegyptus quasi mulieres et stupebunt et timebunt a facie commotionis manus Domini exercituum quam ipse movebit super eam
ISA|19|17|et erit terra Iuda Aegypto in festivitatem omnis qui illius fuerit recordatus pavebit a facie consilii Domini exercituum quod ipse cogitavit super eam
ISA|19|18|in die illa erunt quinque civitates in terra Aegypti loquentes lingua Chanaan et iurantes per Dominum exercituum civitas Solis vocabitur una
ISA|19|19|in die illa erit altare Domini in medio terrae Aegypti et titulus iuxta terminum eius Domini
ISA|19|20|et erit in signum et in testimonium Domino exercituum in terra Aegypti clamabunt enim ad Dominum a facie tribulantis et mittet eis salvatorem et propugnatorem qui liberet eos
ISA|19|21|et cognoscetur Dominus ab Aegypto et cognoscent Aegyptii Dominum in die illa et colent eum in hostiis et muneribus et vota vovebunt Domino et solvent
ISA|19|22|et percutiet Dominus Aegyptum plaga et sanabit eam et revertentur ad Dominum et placabitur eis et sanabit eos
ISA|19|23|in die illa erit via de Aegypto in Assyrios et intrabit Assyrius Aegyptum et Aegyptius in Assyrios et servient Aegyptii Assur
ISA|19|24|in die illa erit Israhel tertius Aegyptio et Assyrio benedictio in medio terrae
ISA|19|25|cui benedixit Dominus exercituum dicens benedictus populus meus Aegypti et opus manuum mearum Assyrio hereditas autem mea Israhel
ISA|20|1|in anno quo ingressus est Tharthan in Azotum cum misisset eum Sargon rex Assyriorum et pugnasset contra Azotum et cepisset eam
ISA|20|2|in tempore illo locutus est Dominus in manu Isaiae filii Amos dicens vade et solve saccum de lumbis tuis et calciamenta tua tolle de pedibus tuis et fecit sic vadens nudus et disculciatus
ISA|20|3|et dixit Dominus sicut ambulavit servus meus Isaias nudus et disculciatus trium annorum signum et portentum erit super Aegyptum et super Aethiopiam
ISA|20|4|sic minabit rex Assyriorum captivitatem Aegypti et transmigrationem Aethiopiae iuvenum et senum nudam et disculciatam discopertis natibus ignominiam Aegypti
ISA|20|5|et timebunt et confundentur ab Aethiopia spe sua et ab Aegypto gloria sua
ISA|20|6|et dicet habitator insulae huius in die illa ecce haec erat spes nostra ad quos confugimus in auxilium ut liberaret nos a facie regis Assyriorum et quomodo effugere poterimus nos
ISA|21|1|onus deserti maris sicut turbines ab africo veniunt de deserto venit de terra horribili
ISA|21|2|visio dura nuntiata est mihi qui incredulus est infideliter agit et qui depopulator est vastat ascende Aelam obside Mede omnem gemitum eius cessare feci
ISA|21|3|propterea repleti sunt lumbi mei dolore angustia possedit me sicut angustia parientis corrui cum audirem conturbatus sum cum viderem
ISA|21|4|emarcuit cor meum tenebrae stupefecerunt me Babylon dilecta mea posita est mihi in miraculum
ISA|21|5|pone mensam contemplare in specula comedentes bibentes surgite principes arripite clypeum
ISA|21|6|haec enim dixit mihi Dominus vade et pone speculatorem et quodcumque viderit adnuntiet
ISA|21|7|et vidit currum duorum equitum ascensorem asini et ascensorem cameli et contemplatus est diligenter multo intuitu
ISA|21|8|et clamavit leo super specula Domini ego sum stans iugiter per diem et super custodiam meam ego sum stans totis noctibus
ISA|21|9|ecce iste venit ascensor vir bigae equitum et respondit et dixit cecidit cecidit Babylon et omnia sculptilia deorum eius contrita sunt in terram
ISA|21|10|tritura mea et fili areae meae quae audivi a Domino exercituum Deo Israhel adnuntiavi vobis
ISA|21|11|onus Duma ad me clamat ex Seir custos quid de nocte custos quid de nocte
ISA|21|12|dixit custos venit mane et nox si quaeritis quaerite convertimini venite
ISA|21|13|onus in Arabia in saltu ad vesperam dormietis in semitis Dodanim
ISA|21|14|occurrentes sitienti ferte aquam qui habitatis terram austri cum panibus occurrite fugienti
ISA|21|15|a facie enim gladiorum fugerunt a facie gladii inminentis a facie arcus extenti a facie gravis proelii
ISA|21|16|quoniam haec dicit Dominus ad me adhuc in uno anno quasi in anno mercennarii et auferetur omnis gloria Cedar
ISA|21|17|et reliquiae numeri sagittariorum fortium de filiis Cedar inminuentur Dominus enim Deus Israhel locutus est
ISA|22|1|onus vallis Visionis quidnam tibi quoque est quia ascendisti et tu omnis in tecta
ISA|22|2|clamoris plena urbs frequens civitas exultans interfecti tui non interfecti gladio nec mortui in bello
ISA|22|3|cuncti principes tui fugerunt simul dureque ligati sunt omnes qui inventi sunt vincti sunt pariter procul fugerunt
ISA|22|4|propterea dixi recedite a me amare flebo nolite incumbere ut consolemini me super vastitate filiae populi mei
ISA|22|5|dies enim interfectionis et conculcationis et fletuum Domino Deo exercituum in valle Visionis scrutans murum et magnificus super montem
ISA|22|6|et Aelam sumpsit faretram currum hominis equitis et parietem nudavit clypeus
ISA|22|7|et erunt electae valles tuae plenae quadrigarum et equites ponent sedes suas in porta
ISA|22|8|et revelabitur operimentum Iudae et videbis in die illa armamentarium domus saltus
ISA|22|9|et scissuras civitatis David videbitis quia multiplicatae sunt et congregastis aquas piscinae inferioris
ISA|22|10|et domos Hierusalem numerastis et destruxistis domos ad muniendum murum
ISA|22|11|et lacum fecistis inter duos muros et aquam piscinae veteris et non suspexistis ad eum qui fecerat eam et operatorem eius de longe non vidistis
ISA|22|12|et vocavit Dominus Deus exercituum in die illa ad fletum et ad planctum ad calvitium et ad cingulum sacci
ISA|22|13|et ecce gaudium et laetitia occidere vitulos et iugulare arietes comedere carnes et bibere vinum comedamus et bibamus cras enim moriemur
ISA|22|14|et revelata est in auribus meis Domini exercituum si dimittetur iniquitas haec vobis donec moriamini dicit Dominus Deus exercituum
ISA|22|15|haec dicit Dominus Deus exercituum vade ingredere ad eum qui habitat in tabernaculo ad Sobnam praepositum templi
ISA|22|16|quid tu hic aut quasi quis hic quia excidisti tibi hic sepulchrum excidisti in excelso memoriam diligenter in petra tabernaculum tibi
ISA|22|17|ecce Dominus asportari te faciet sicut asportatur gallus gallinacius et quasi amictum sic sublevabit te
ISA|22|18|coronans coronabit te tribulatione quasi pilam mittet te in terram latam et spatiosam ibi morieris et ibi erit currus gloriae tuae ignominia domus Domini tui
ISA|22|19|et expellam te de statione tua et de ministerio tuo deponam te
ISA|22|20|et erit in die illa vocabo servum meum Eliachim filium Helciae
ISA|22|21|et induam illum tunicam tuam et cingulo tuo confortabo eum et potestatem tuam dabo in manu eius et erit quasi pater habitantibus Hierusalem et domui Iuda
ISA|22|22|et dabo clavem domus David super umerum eius et aperiet et non erit qui claudat et claudet et non erit qui aperiat
ISA|22|23|et figam illum paxillum in loco fideli et erit in solium gloriae domui patris sui
ISA|22|24|et suspendent super eum omnem gloriam domus patris eius vasorum diversa genera omne vas parvulum a vasis craterarum usque ad omne vas musicorum
ISA|22|25|in die illo dicit Dominus exercituum auferetur paxillus qui fixus fuerat in loco fideli et frangetur et cadet et peribit quod pependerat in eo quia Dominus locutus est
ISA|23|1|onus Tyri ululate naves maris quia vastata est domus unde venire consueverant de terra Cetthim revelatum est eis
ISA|23|2|tacete qui habitatis in insula negotiatio Sidonis transfretantes mare repleverunt te
ISA|23|3|in aquis multis semen Nili messis fluminis fruges eius et facta est negotiatio gentium
ISA|23|4|erubesce Sidon ait enim mare fortitudo maris dicens non parturivi et non peperi et non enutrivi iuvenes nec ad incrementum perduxi virgines
ISA|23|5|cum auditum fuerit in Aegypto dolebunt cum audierint de Tyro
ISA|23|6|transite maria ululate qui habitatis in insula
ISA|23|7|numquid non haec vestra est quae gloriabatur a diebus pristinis in antiquitate sua ducent eam pedes sui longe ad peregrinandum
ISA|23|8|quis cogitavit hoc super Tyrum quondam coronatam cuius negotiatores principes institores eius incliti terrae
ISA|23|9|Dominus exercituum cogitavit hoc ut detraheret superbiam omnis gloriae et ad ignominiam deduceret universos inclitos terrae
ISA|23|10|transi terram tuam quasi flumen filia maris non est cingulum ultra tibi
ISA|23|11|manum suam extendit super mare conturbavit regna Dominus mandavit adversum Chanaan ut contereret fortes eius
ISA|23|12|et dixit non adicies ultra ut glorieris calumniam sustinens virgo filia Sidonis in Cetthim consurgens transfreta ibi quoque non erit requies tibi
ISA|23|13|ecce terra Chaldeorum talis populus non fuit Assur fundavit eam in captivitatem transduxerunt robustos eius suffoderunt domos eius posuerunt eam in ruinam
ISA|23|14|ululate naves maris quia devastata est fortitudo vestra
ISA|23|15|et erit in die illa in oblivione eris o Tyre septuaginta annis sicut dies regis unius post septuaginta autem annos erit Tyro quasi canticum meretricis
ISA|23|16|sume citharam circui civitatem meretrix oblivioni tradita bene cane frequenta canticum ut memoria tui sit
ISA|23|17|et erit post septuaginta annos visitabit Dominus Tyrum et reducet eam ad mercedes suas et rursum fornicabitur cum universis regnis terrae super faciem terrae
ISA|23|18|et erunt negotiatio eius et mercedes eius sanctificatae Domino non condentur neque reponentur quia his qui habitaverint coram Domino erit negotiatio eius ut manducent in saturitatem et vestiantur usque ad vetustatem
ISA|24|1|ecce Dominus dissipabit terram et nudabit eam et adfliget faciem eius et disperget habitatores eius
ISA|24|2|et erit sicut populus sic sacerdos et sicut servus sic dominus eius sicut ancilla sic domina eius sicut emens sic ille qui vendit sicut fenerator sic is qui mutuum accipit sicut qui repetit sic qui debet
ISA|24|3|dissipatione dissipabitur terra et direptione praedabitur Dominus enim locutus est verbum hoc
ISA|24|4|luxit et defluxit terra et infirmata est defluxit orbis infirmata est altitudo populi terrae
ISA|24|5|et terra interfecta est ab habitatoribus suis quia transgressi sunt leges mutaverunt ius dissipaverunt foedus sempiternum
ISA|24|6|propter hoc maledictio vorabit terram et peccabunt habitatores eius ideoque insanient cultores eius et relinquentur homines pauci
ISA|24|7|luxit vindemia infirmata est vitis ingemuerunt omnes qui laetabantur corde
ISA|24|8|cessavit gaudium tympanorum quievit sonitus laetantium conticuit dulcedo citharae
ISA|24|9|cum cantico non bibent vinum amara erit potio bibentibus illam
ISA|24|10|adtrita est civitas vanitatis clausa est omnis domus nullo introeunte
ISA|24|11|clamor erit super vino in plateis deserta est omnis laetitia translatum est gaudium terrae
ISA|24|12|relicta est in urbe solitudo et calamitas opprimet portas
ISA|24|13|quia haec erunt in medio terrae in medio populorum quomodo si paucae olivae quae remanserunt excutiantur ex olea et racemi cum fuerit finita vindemia
ISA|24|14|hii levabunt vocem suam atque laudabunt cum glorificatus fuerit Dominus hinnient de mari
ISA|24|15|propter hoc in doctrinis glorificate Dominum in insulis maris nomen Domini Dei Israhel
ISA|24|16|a finibus terrae laudes audivimus gloriam iusti et dixi secretum meum mihi secretum meum mihi vae mihi praevaricantes praevaricati sunt et praevaricatione transgressorum praevaricati sunt
ISA|24|17|formido et fovea et laqueus super te qui habitator es terrae
ISA|24|18|et erit qui fugerit a voce formidinis cadet in foveam et qui se explicuerit de fovea tenebitur laqueo quia cataractae de excelsis apertae sunt et concutientur fundamenta terrae
ISA|24|19|confractione confringetur terra contritione conteretur terra commotione commovebitur terra
ISA|24|20|agitatione agitabitur terra sicut ebrius et auferetur quasi tabernaculum unius noctis et gravabit eam iniquitas sua et corruet et non adiciet ut resurgat
ISA|24|21|et erit in die illa visitabit Dominus super militiam caeli in excelso et super reges terrae qui sunt super terram
ISA|24|22|et congregabuntur in congregationem unius fascis in lacum et cludentur ibi in carcerem et post multos dies visitabuntur
ISA|24|23|et erubescet luna et confundetur sol cum regnaverit Dominus exercituum in monte Sion et in Hierusalem et in conspectu senum suorum fuerit glorificatus
ISA|25|1|Domine Deus meus es tu exaltabo te confitebor nomini tuo quoniam fecisti mirabilia cogitationes antiquas fideles amen
ISA|25|2|quia posuisti civitatem in tumulum urbem fortem in ruinam domum alienorum ut non sit civitas et in sempiternum non aedificetur
ISA|25|3|super hoc laudabit te populus fortis civitas gentium robustarum timebit te
ISA|25|4|quia factus es fortitudo pauperi fortitudo egeno in tribulatione sua spes a turbine umbraculum ab aestu spiritus enim robustorum quasi turbo inpellens parietem
ISA|25|5|sicut aestum in siti tumultum alienorum humiliabis et quasi calore sub nube torrente propaginem fortium marcescere facies
ISA|25|6|et faciet Dominus exercituum omnibus populis in monte hoc convivium pinguium convivium vindemiae pinguium medullatorum vindemiae defecatae
ISA|25|7|et praecipitabit in monte isto faciem vinculi conligati super omnes populos et telam quam orditus est super universas nationes
ISA|25|8|praecipitabit mortem in sempiternum et auferet Dominus Deus lacrimam ab omni facie et obprobrium populi sui auferet de universa terra quia Dominus locutus est
ISA|25|9|et dicet in die illa ecce Deus noster iste expectavimus eum et salvabit nos iste Dominus sustinuimus eum exultabimus et laetabimur in salutari eius
ISA|25|10|quia requiescet manus Domini in monte isto et triturabitur Moab sub eo sicuti teruntur paleae in plaustro
ISA|25|11|et extendet manus suas sub eo sicut extendit natans ad natandum et humiliabit gloriam eius cum adlisione manuum eius
ISA|25|12|et munimenta sublimium murorum tuorum concident et humiliabuntur et detrahentur in terram usque ad pulverem
ISA|26|1|in die illa cantabitur canticum istud in terra Iuda urbs fortitudinis nostrae salvator ponetur in ea murus et antemurale
ISA|26|2|aperite portas et ingrediatur gens iusta custodiens veritatem
ISA|26|3|vetus error abiit servabis pacem pacem quia in te speravimus
ISA|26|4|sperastis in Domino in saeculis aeternis in Domino Deo forti in perpetuum
ISA|26|5|quia incurvabit habitantes in excelso civitatem sublimem humiliabit humiliabit eam usque ad terram detrahet eam usque ad pulverem
ISA|26|6|conculcabit eam pes pedes pauperis gressus egenorum
ISA|26|7|semita iusti recta est rectus callis iusti ad ambulandum
ISA|26|8|et in semita iudiciorum tuorum Domine sustinuimus te nomen tuum et memoriale tuum in desiderio animae
ISA|26|9|anima mea desideravit te in nocte sed et spiritu meo in praecordiis meis de mane vigilabo ad te cum feceris iudicia tua in terra iustitiam discent habitatores orbis
ISA|26|10|misereamur impio et non discet iustitiam in terra sanctorum inique gessit et non videbit gloriam Domini
ISA|26|11|Domine exaltetur manus tua et non videant videant et confundantur zelantes populi et ignis hostes tuos devoret
ISA|26|12|Domine dabis pacem nobis omnia enim opera nostra operatus es nobis
ISA|26|13|Domine Deus noster possederunt nos domini absque te tantum in te recordemur nominis tui
ISA|26|14|morientes non vivant gigantes non resurgant propterea visitasti et contrivisti eos et perdidisti omnem memoriam eorum
ISA|26|15|indulsisti genti Domine indulsisti genti numquid glorificatus es elongasti omnes terminos terrae
ISA|26|16|Domine in angustia requisierunt te in tribulatione murmuris doctrina tua eis
ISA|26|17|sicut quae concipit cum adpropinquaverit ad partum dolens clamat in doloribus suis sic facti sumus a facie tua Domine
ISA|26|18|concepimus et quasi parturivimus et peperimus spiritum salutes non fecimus in terra ideo non ceciderunt habitatores terrae
ISA|26|19|vivent mortui tui interfecti mei resurgent expergiscimini et laudate qui habitatis in pulvere quia ros lucis ros tuus et terram gigantum detrahes in ruinam
ISA|26|20|vade populus meus intra in cubicula tua claude ostia tua super te abscondere modicum ad momentum donec pertranseat indignatio
ISA|26|21|ecce enim Dominus egreditur de loco suo ut visitet iniquitatem habitatoris terrae contra eum et revelabit terra sanguinem suum et non operiet ultra interfectos suos
ISA|27|1|in die illo visitabit Dominus in gladio suo duro et grandi et forti super Leviathan serpentem vectem et super Leviathan serpentem tortuosum et occidet cetum qui in mari est
ISA|27|2|in die illa vinea meri cantabit ei
ISA|27|3|ego Dominus qui servo eam repente propinabo ei ne forte visitetur contra eam nocte et die servo eam
ISA|27|4|indignatio non est mihi quis dabit me spinam et veprem in proelio gradiar super eam succendam eam pariter
ISA|27|5|an potius tenebit fortitudinem meam faciet pacem mihi pacem faciet mihi
ISA|27|6|qui egrediuntur impetu ad Iacob florebit et germinabit Israhel et implebunt faciem orbis semine
ISA|27|7|numquid iuxta plagam percutientis se percussit eum aut sicut occidit interfectos eius sic occisus est
ISA|27|8|in mensura contra mensuram cum abiecta fuerit iudicabis eam meditata est in spiritu suo duro per diem aestus
ISA|27|9|idcirco super hoc dimittetur iniquitas domui Iacob et iste omnis fructus ut auferatur peccatum eius cum posuerit omnes lapides altaris sicut lapides cineris adlisos non stabunt luci et delubra
ISA|27|10|civitas enim munita desolata erit speciosa relinquetur et dimittetur quasi desertum ibi pascetur vitulus et ibi accubabit et consumet summitates eius
ISA|27|11|in siccitate messis illius conterentur mulieres venientes et docentes eam non est enim populus sapiens propterea non miserebitur eius qui fecit eum et qui formavit eum non parcet ei
ISA|27|12|et erit in die illa percutiet Dominus ab alveo Fluminis usque ad torrentem Aegypti et vos congregabimini unus et unus filii Israhel
ISA|27|13|et erit in die illa clangetur in tuba magna et venient qui perditi fuerant de terra Assyriorum et qui eiecti erant in terra Aegypti et adorabunt Dominum in monte sancto in Hierusalem
ISA|28|1|vae coronae superbiae ebriis Ephraim et flori decidenti gloriae exultationis eius qui erant in vertice vallis pinguissimae errantes a vino
ISA|28|2|ecce validus et fortis Domini sicut impetus grandinis turbo confringens sicut impetus aquarum multarum inundantium et emissarum super terram spatiosam
ISA|28|3|pedibus conculcabitur corona superbiae ebriorum Ephraim
ISA|28|4|et erit flos decidens gloriae exultationis eius qui est super verticem vallis pinguium quasi temporaneum ante maturitatem autumni quod cum aspexerit videns statim ut manu tenuerit devorabit illud
ISA|28|5|in die illa erit Dominus exercituum corona gloriae et sertum exultationis residuo populi sui
ISA|28|6|et spiritus iudicii sedenti super iudicium et fortitudo revertentibus de bello ad portam
ISA|28|7|verum hii quoque prae vino nescierunt et prae ebrietate erraverunt sacerdos et propheta nescierunt prae ebrietate absorti sunt a vino erraverunt in ebrietate nescierunt videntem ignoraverunt iudicium
ISA|28|8|omnes enim mensae repletae sunt vomitu sordiumque ita ut non esset ultra locus
ISA|28|9|quem docebit scientiam et quem intellegere faciet auditum ablactatos a lacte apulsos ab uberibus
ISA|28|10|quia manda remanda manda remanda expecta reexpecta expecta reexpecta modicum ibi modicum ibi
ISA|28|11|in loquella enim labii et lingua altera loquetur ad populum istum
ISA|28|12|cui dixit haec requies reficite lassum et hoc est meum refrigerium et noluerunt audire
ISA|28|13|et erit eis verbum Domini manda remanda manda remanda expecta reexpecta expecta reexpecta modicum ibi modicum ibi ut vadant et cadant retrorsum et conterantur et inlaqueentur et capiantur
ISA|28|14|propter hoc audite verbum Domini viri inlusores qui dominamini super populum meum qui est in Hierusalem
ISA|28|15|dixistis enim percussimus foedus cum morte et cum inferno fecimus pactum flagellum inundans cum transierit non veniet super nos quia posuimus mendacium spem nostram et mendacio protecti sumus
ISA|28|16|idcirco haec dicit Dominus Deus ecce ego mittam in fundamentis Sion lapidem lapidem probatum angularem pretiosum in fundamento fundatum qui crediderit non festinet
ISA|28|17|et ponam iudicium in pondere et iustitiam in mensura et subvertet grando spem mendacii et protectionem aquae inundabunt
ISA|28|18|et delebitur foedus vestrum cum morte et pactum vestrum cum inferno non stabit flagellum inundans cum transierit eritis ei in conculcationem
ISA|28|19|quandocumque pertransierit tollet vos quoniam mane diluculo pertransibit in die et in nocte et tantummodo sola vexatio intellectum dabit auditui
ISA|28|20|coangustatum est enim stratum ita ut alter decidat et pallium breve utrumque operire non potest
ISA|28|21|sicut enim in monte Divisionum stabit Dominus sicut in valle quae est in Gabao irascetur ut faciat opus suum alienum opus eius ut operetur opus suum peregrinum est opus ab eo
ISA|28|22|et nunc nolite inludere ne forte constringantur vincula vestra consummationem enim et adbreviationem audivi a Domino Deo exercituum super universam terram
ISA|28|23|auribus percipite et audite vocem meam adtendite et audite eloquium meum
ISA|28|24|numquid tota die arabit arans ut serat proscindet et sariet humum suam
ISA|28|25|nonne cum adaequaverit faciem eius seret gith et cyminum sparget et ponet triticum per ordinem et hordeum et milium et viciam in finibus suis
ISA|28|26|et erudiet eum illud in iudicio Deus suus docebit eum illud
ISA|28|27|non enim in serris triturabitur gith nec rota plaustri super cyminum circumiet sed in virga excutietur gith et cyminum in baculo
ISA|28|28|panis autem comminuetur verum non in perpetuum triturans triturabit illum neque vexabit eum rota plaustri nec in ungulis suis comminuet eum
ISA|28|29|et hoc a Domino Deo exercituum exivit ut mirabile faceret consilium et magnificaret iustitiam
ISA|29|1|vae Arihel Arihel civitas quam circumdedit David additus est annus ad annum sollemnitates evolutae sunt
ISA|29|2|et circumvallabo Arihel et erit tristis et maerens et erit mihi quasi Arihel
ISA|29|3|et circumdabo quasi spheram in circuitu tuo et iaciam contra te aggerem et munimenta ponam in obsidionem tuam
ISA|29|4|humiliaberis de terra loqueris et de humo audietur eloquium tuum et erit quasi pythonis de terra vox tua et de humo eloquium tuum mussitabit
ISA|29|5|et erit sicut pulvis tenuis multitudo ventilantium te et sicut favilla pertransiens multitudo eorum qui contra te praevaluerunt
ISA|29|6|eritque repente confestim a Domino exercituum visitabitur in tonitru et commotione terrae et voce magna turbinis et tempestatis et flammae ignis devorantis
ISA|29|7|et erit sicut somnium visionis nocturnae multitudo omnium gentium quae dimicaverunt contra Arihel et omnes qui militaverunt et obsederunt et praevaluerunt adversus eam
ISA|29|8|et sicuti somniat esuriens et comedit cum autem fuerit expertus vacua est anima eius et sicut somniat sitiens et bibit et postquam fuerit expergefactus lassus adhuc sitit et anima eius vacua est sic erit multitudo omnium gentium quae dimicaverunt contra montem Sion
ISA|29|9|obstupescite et admiramini fluctuate et vacillate inebriamini et non a vino movemini et non ebrietate
ISA|29|10|quoniam miscuit vobis Dominus spiritum soporis claudet oculos vestros prophetas et principes vestros qui vident visiones operiet
ISA|29|11|et erit vobis visio omnium sicut verba libri signati quem cum dederint scienti litteras dicent lege istum et respondebit non possum signatus est enim
ISA|29|12|et dabitur liber nescienti litteras diceturque ei lege et respondebit nescio litteras
ISA|29|13|et dixit Dominus eo quod adpropinquat populus iste ore suo et labiis suis glorificat me cor autem eius longe est a me et timuerunt me mandato hominum et doctrinis
ISA|29|14|ideo ecce ego addam ut admirationem faciam populo huic miraculo grandi et stupendo peribit enim sapientia a sapientibus eius et intellectus prudentium eius abscondetur
ISA|29|15|vae qui profundi estis corde ut a Domino abscondatis consilium quorum sunt in tenebris opera et dicunt quis videt nos et quis novit nos
ISA|29|16|perversa est haec vestra cogitatio quasi lutum contra figulum cogitet et dicat opus factori suo non fecisti me et figmentum dicat fictori suo non intellegis
ISA|29|17|nonne adhuc in modico et in brevi convertetur Libanus in Chermel et Chermel in saltum reputabitur
ISA|29|18|et audient in die illa surdi verba libri et de tenebris et caligine oculi caecorum videbunt
ISA|29|19|et addent mites in Domino laetitiam et pauperes homines in Sancto Israhel exultabunt
ISA|29|20|quoniam defecit qui praevalebat consummatus est inlusor et succisi sunt omnes qui vigilabant super iniquitatem
ISA|29|21|qui peccare faciebant homines in verbo et arguentem in porta subplantabant et declinaverunt frustra a iusto
ISA|29|22|propter hoc haec dicit Dominus ad domum Iacob qui redemit Abraham non modo confundetur Iacob nec modo vultus eius erubescet
ISA|29|23|sed cum viderit filios suos opera manuum mearum in medio sui sanctificantes nomen meum et sanctificabunt Sanctum Iacob et Deum Israhel praedicabunt
ISA|29|24|et scient errantes spiritu intellectum et mussitatores discent legem
ISA|30|1|vae filii desertores dicit Dominus ut faceretis consilium et non ex me et ordiremini telam et non per spiritum meum ut adderetur peccatum super peccatum
ISA|30|2|qui ambulatis ut descendatis in Aegyptum et os meum non interrogastis sperantes auxilium in fortitudine Pharao et habentes fiduciam in umbra Aegypti
ISA|30|3|et erit vobis fortitudo Pharaonis in confusionem et fiducia umbrae Aegypti in ignominiam
ISA|30|4|erant enim in Tanis principes tui et nuntii tui usque ad Anes pervenerunt
ISA|30|5|omnes confusi sunt super populo qui eis prodesse non potuit non fuerunt in auxilium et in aliquam utilitatem sed in confusionem et obprobrium
ISA|30|6|onus iumentorum austri in terra tribulationis et angustiae leaena et leo ex eis vipera et regulus volans portantes super umeros iumentorum divitias suas et super gibbum camelorum thesauros suos ad populum qui eis prodesse non poterit
ISA|30|7|Aegyptus enim frustra et vane auxiliabitur ideo clamavi super hoc superbia tantum est quiesce
ISA|30|8|nunc ingressus scribe eis super buxum et in libro diligenter exara illud et erit in die novissimo in testimonium usque ad aeternum
ISA|30|9|populus enim ad iracundiam provocans est et filii mendaces filii nolentes audire legem Domini
ISA|30|10|qui dicunt videntibus nolite videre et aspicientibus nolite aspicere nobis ea quae recta sunt loquimini nobis placentia videte nobis errores
ISA|30|11|auferte a me viam declinate a me semitam cesset a facie nostra Sanctus Israhel
ISA|30|12|propterea haec dicit Sanctus Israhel pro eo quod reprobastis verbum hoc et sperastis in calumniam et tumultum et innixi estis super eo
ISA|30|13|propterea erit vobis iniquitas haec sicut interruptio cadens et requisita in muro excelso quoniam subito dum non speratur veniet contritio eius
ISA|30|14|et comminuetur sicut conteritur lagoena figuli contritione pervalida et non invenietur de fragmentis eius testa in qua portetur igniculus de incendio aut hauriatur parum aquae de fovea
ISA|30|15|quia haec dicit Dominus Deus Sanctus Israhel si revertamini et quiescatis salvi eritis in silentio et in spe erit fortitudo vestra et noluistis
ISA|30|16|et dixistis nequaquam sed ad equos fugiemus ideo fugietis et super veloces ascendemus ideo veloces erunt qui persequentur vos
ISA|30|17|mille homines a facie terroris unius et a facie terroris quinque fugietis donec relinquamini quasi malus navis in vertice montis et quasi signum super collem
ISA|30|18|propterea expectat Dominus ut misereatur vestri et ideo exaltabitur parcens vobis quia Deus iudicii Dominus beati omnes qui expectant eum
ISA|30|19|populus enim Sion habitabit in Hierusalem plorans nequaquam plorabis miserans miserebitur tui ad vocem clamoris tui statim ut audierit respondebit tibi
ISA|30|20|et dabit vobis Dominus panem artum et aquam brevem et non faciet avolare a te ultra doctorem tuum et erunt oculi tui videntes praeceptorem tuum
ISA|30|21|et aures tuae audient verbum post tergum monentis haec via ambulate in ea neque ad dexteram neque ad sinistram
ISA|30|22|et contaminabis lamminas sculptilium argenti tui et vestimentum conflatilis auri tui et disperges ea sicut inmunditiam menstruatae egredere dices ei
ISA|30|23|et dabitur pluvia semini tuo ubicumque seminaveris in terra et panis frugum terrae erit uberrimus et pinguis pascetur in possessione tua in die illo agnus spatiose
ISA|30|24|et tauri tui et pulli asinorum qui operantur terram commixtum migma comedent sic in area ut ventilatum est
ISA|30|25|et erunt super omnem montem excelsum et super omnem collem elevatum rivi currentium aquarum in die interfectionis multorum cum ceciderint turres
ISA|30|26|et erit lux lunae sicut lux solis et lux solis erit septempliciter sicut lux septem dierum in die qua alligaverit Dominus vulnus populi sui et percussuram plagae eius sanaverit
ISA|30|27|ecce nomen Domini venit de longinquo ardens furor eius et gravis ad portandum labia eius repleta sunt indignatione et lingua eius quasi ignis devorans
ISA|30|28|spiritus eius velut torrens inundans usque ad medium colli ad perdendas gentes in nihilum et frenum erroris quod erat in maxillis populorum
ISA|30|29|canticum erit vobis sicut nox sanctificatae sollemnitatis et laetitia cordis sicut qui pergit cum tibia ut intret in montem Domini ad Fortem Israhel
ISA|30|30|et auditam faciet Dominus gloriam vocis suae et terrorem brachii sui ostendet in comminatione furoris et flamma ignis devorantis adlidet in turbine et in lapide grandinis
ISA|30|31|a voce enim Domini pavebit Assur virga percussus
ISA|30|32|et erit transitus virgae fundatus quam requiescere faciet Dominus super eum in tympanis et in citharis et in bellis praecipuis expugnabit eos
ISA|30|33|praeparata est enim ab heri Thofeth a rege praeparata profunda et dilatata nutrimenta eius ignis et ligna multa flatus Domini sicut torrens sulphuris succendens eam
ISA|31|1|vae qui descendunt in Aegyptum ad auxilium in equis sperantes et habentes fiduciam super quadrigis quia multae sunt et super equitibus quia praevalidi nimis et non sunt confisi super Sanctum Israhel et Dominum non requisierunt
ISA|31|2|ipse autem sapiens adduxit malum et verba sua non abstulit et consurget contra domum pessimorum et contra auxilium operantium iniquitatem
ISA|31|3|Aegyptus homo et non deus et equi eorum caro et non spiritus et Dominus inclinabit manum suam et corruet auxiliator et cadet cui praestatur auxilium simulque omnes consumentur
ISA|31|4|quia haec dicit Dominus ad me quomodo si rugiat leo et catulus leonis super praedam suam cum occurrerit ei multitudo pastorum a voce eorum non formidabit et a multitudine eorum non pavebit sic descendet Dominus exercituum ut proelietur super montem Sion et super collem eius
ISA|31|5|sicut aves volantes sic proteget Dominus exercituum Hierusalem protegens et liberans transiens et salvans
ISA|31|6|convertimini sicut in profundum recesseratis filii Israhel
ISA|31|7|in die enim illa abiciet vir idola argenti sui et idola auri sui quae fecerunt vobis manus vestrae in peccatum
ISA|31|8|et cadet Assur in gladio non viri et gladius non hominis vorabit eum et fugiet non a facie gladii et iuvenes eius vectigales erunt
ISA|31|9|et fortitudo eius a terrore transibit et pavebunt fugientes principes eius dixit Dominus cuius ignis est in Sion et caminus eius in Hierusalem
ISA|32|1|ecce in iustitia regnabit rex et principes in iudicio praeerunt
ISA|32|2|et erit vir sicut qui absconditur a vento et celat se a tempestate sicut rivi aquarum in siti et umbra petrae prominentis in terra deserta
ISA|32|3|non caligabunt oculi videntium et aures audientium diligenter auscultabunt
ISA|32|4|et cor stultorum intelleget scientiam et lingua balborum velociter loquetur et plane
ISA|32|5|non vocabitur ultra is qui insipiens est princeps neque fraudulentus appellabitur maior
ISA|32|6|stultus enim fatua loquetur et cor eius faciet iniquitatem ut perficiat simulationem et loquatur ad Dominum fraudulenter et vacuefaciat animam esurientis et potum sitienti auferat
ISA|32|7|fraudulenti vasa pessima sunt ipse enim cogitationes concinnavit ad perdendos mites in sermone mendacii cum loqueretur pauper iudicium
ISA|32|8|princeps vero ea quae digna sunt principe cogitavit et ipse super duces stabit
ISA|32|9|mulieres opulentae surgite et audite vocem meam filiae confidentes percipite auribus eloquium meum
ISA|32|10|post dies et annum et vos conturbabimini confidentes consummata est enim vindemia collectio ultra non veniet
ISA|32|11|obstupescite opulentae conturbamini confidentes exuite vos et confundimini accingite lumbos vestros
ISA|32|12|super ubera plangite super regione desiderabili super vinea fertili
ISA|32|13|super humum populi mei spina et vepres ascendent quanto magis super omnes domos gaudii civitatis exultantis
ISA|32|14|domus enim dimissa est multitudo urbis relicta est tenebrae et palpatio factae sunt super speluncas usque in aeternum gaudium onagrorum pascua gregum
ISA|32|15|donec effundatur super nos spiritus de excelso et erit desertum in Chermel et Chermel in saltum reputabitur
ISA|32|16|et habitabit in solitudine iudicium et iustitia in Chermel sedebit
ISA|32|17|et erit opus iustitiae pax et cultus iustitiae silentium et securitas usque in sempiternum
ISA|32|18|et sedebit populus meus in pulchritudine pacis et in tabernaculis fiduciae et in requie opulenta
ISA|32|19|grando autem in descensione saltus et humilitate humiliabitur civitas
ISA|32|20|beati qui seminatis super omnes aquas inmittentes pedem bovis et asini
ISA|33|1|vae qui praedaris nonne et ipse praedaberis et qui spernis nonne et ipse sperneris cum consummaveris depraedationem depraedaberis cum fatigatus desiveris contemnere contemneris
ISA|33|2|Domine miserere nostri te expectavimus esto brachium eorum in mane et salus nostra in tempore tribulationis
ISA|33|3|a voce angeli fugerunt populi ab exaltatione tua dispersae sunt gentes
ISA|33|4|et congregabuntur spolia vestra sicut colligitur brucus velut cum fossae plenae fuerint de eo
ISA|33|5|magnificatus est Dominus quoniam habitavit in excelso implevit Sion iudicio et iustitia
ISA|33|6|et erit fides in temporibus tuis divitiae salutis sapientia et scientia timor Domini ipse thesaurus eius
ISA|33|7|ecce videntes clamabunt foris angeli pacis amare flebunt
ISA|33|8|dissipatae sunt viae cessavit transiens per semitam irritum factum est pactum proiecit civitates non reputavit homines
ISA|33|9|luxit et elanguit terra confusus est Libanus et obsorduit et factus est Saron sicut desertum et concussa est Basan et Carmelus
ISA|33|10|nunc consurgam dicit Dominus nunc exaltabor nunc sublevabor
ISA|33|11|concipietis ardorem parietis stipulam spiritus vester ut ignis vorabit vos
ISA|33|12|et erunt populi quasi de incendio cinis spinae congregatae igni conburentur
ISA|33|13|audite qui longe estis quae fecerim et cognoscite vicini fortitudinem meam
ISA|33|14|conterriti sunt in Sion peccatores possedit tremor hypocritas quis poterit habitare de vobis cum igne devorante quis habitabit ex vobis cum ardoribus sempiternis
ISA|33|15|qui ambulat in iustitiis et loquitur veritates qui proicit avaritiam ex calumnia et excutit manus suas ab omni munere qui obturat aures suas ne audiat sanguinem et claudit oculos suos ne videat malum
ISA|33|16|iste in excelsis habitabit munimenta saxorum sublimitas eius panis ei datus est aquae eius fideles sunt
ISA|33|17|regem in decore suo videbunt oculi eius cernent terram de longe
ISA|33|18|cor tuum meditabitur timorem ubi est litteratus ubi legis verba ponderans ubi doctor parvulorum
ISA|33|19|populum inpudentem non videbis populum alti sermonis ita ut non possis intellegere disertitudinem linguae eius in quo nulla est sapientia
ISA|33|20|respice Sion civitatem sollemnitatis nostrae oculi tui videbunt Hierusalem habitationem opulentam tabernaculum quod nequaquam transferri poterit nec auferentur clavi eius in sempiternum et omnes funiculi eius non rumpentur
ISA|33|21|quia solummodo ibi magnificus Dominus noster locus fluviorum rivi latissimi et patentes non transibit per eum navis remigum neque trieris magna transgredietur eum
ISA|33|22|Dominus enim iudex noster Dominus legifer noster Dominus rex noster ipse salvabit nos
ISA|33|23|laxati sunt funiculi tui sed non praevalebunt sic erit malus tuus ut dilatare signum non queas tunc dividentur spolia praedarum multarum claudi diripient rapinam
ISA|33|24|nec dicet vicinus elangui populus qui habitat in ea auferetur ab eo iniquitas
ISA|34|1|accedite gentes et audite et populi adtendite audiat terra et plenitudo eius orbis et omne germen eius
ISA|34|2|quia indignatio Domini super omnes gentes et furor super universam militiam eorum interfecit eos et dedit eos in occisionem
ISA|34|3|interfecti eorum proicientur et de cadaveribus eorum ascendet fetor tabescent montes sanguine eorum
ISA|34|4|et tabescet omnis militia caelorum et conplicabuntur sicut liber caeli et omnis militia eorum defluet sicut defluit folium de vinea et de ficu
ISA|34|5|quoniam inebriatus est in caelo gladius meus ecce super Idumeam descendet et super populum interfectionis meae ad iudicium
ISA|34|6|gladius Domini repletus est sanguine incrassatus est adipe de sanguine agnorum et hircorum de sanguine medullatorum arietum victima enim Domini in Bosra et interfectio magna in terra Edom
ISA|34|7|et descendent unicornes cum eis et tauri cum potentibus inebriabitur terra eorum sanguine et humus eorum adipe pinguium
ISA|34|8|quia dies ultionis Domini annus retributionum iudicii Sion
ISA|34|9|et convertentur torrentes eius in picem et humus eius in sulphur et erit terra eius in picem ardentem
ISA|34|10|nocte et die non extinguetur in sempiternum ascendet fumus eius a generatione in generationem desolabitur in saeculum saeculorum non erit transiens per eam
ISA|34|11|et possidebunt illam onocrotalus et ericius et ibis et corvus habitabunt in ea et extendetur super eam mensura ut redigatur ad nihilum et perpendiculum in desolationem
ISA|34|12|nobiles eius non erunt ibi regem potius invocabunt et omnes principes eius erunt in nihilum
ISA|34|13|et orientur in domibus eius spinae et urticae et paliurus in munitionibus eius et erit cubile draconum et pascua strutionum
ISA|34|14|et occurrent daemonia onocentauris et pilosus clamabit alter ad alterum ibi cubavit lamia et invenit sibi requiem
ISA|34|15|ibi habuit foveam ericius et enutrivit catulos et circumfodit et fovit in umbra eius illuc congregati sunt milvi alter ad alterum
ISA|34|16|requirite diligenter in libro Domini et legite unum ex eis non defuit alter ad alterum non quaesivit quia quod ex ore meo procedit ille mandavit et spiritus eius ipse congregavit ea
ISA|34|17|et ipse misit eis sortem et manus eius divisit eam illis in mensuram usque in aeternum possidebunt eam in generatione et generatione habitabunt in ea
ISA|35|1|laetabitur deserta et invia et exultabit solitudo et florebit quasi lilium
ISA|35|2|germinans germinabit et exultabit laetabunda et laudans gloria Libani data est ei decor Carmeli et Saron ipsi videbunt gloriam Domini et decorem Dei nostri
ISA|35|3|confortate manus dissolutas et genua debilia roborate
ISA|35|4|dicite pusillanimis confortamini nolite timere ecce Deus vester ultionem adducet retributionis Deus ipse veniet et salvabit vos
ISA|35|5|tunc aperientur oculi caecorum et aures surdorum patebunt
ISA|35|6|tunc saliet sicut cervus claudus et aperta erit lingua mutorum quia scissae sunt in deserto aquae et torrentes in solitudine
ISA|35|7|et quae erat arida in stagnum et sitiens in fontes aquarum in cubilibus in quibus prius dracones habitabant orietur viror calami et iunci
ISA|35|8|et erit ibi semita et via et via sancta vocabitur non transibit per eam pollutus et haec erit nobis directa via ita ut stulti non errent per eam
ISA|35|9|non erit ibi leo et mala bestia non ascendet per eam nec invenietur ibi et ambulabunt qui liberati fuerint
ISA|35|10|et redempti a Domino convertentur et venient in Sion cum laude et laetitia sempiterna super caput eorum gaudium et laetitiam obtinebunt et fugiet dolor et gemitus
ISA|36|1|et factum est in quartodecimo anno regis Ezechiae ascendit Sennacherib rex Assyriorum super omnes civitates Iuda munitas et cepit eas
ISA|36|2|et misit rex Assyriorum Rabsacen de Lachis in Hierusalem ad regem Ezechiam in manu gravi et stetit in aquaeductu piscinae superioris in via agri Fullonis
ISA|36|3|et egressus est ad eum Eliachim filius Helciae qui erat super domum et Sobna scriba et Ioae filius Asaph a commentariis
ISA|36|4|et dixit ad eos Rabsaces dicite Ezechiae haec dicit rex magnus rex Assyriorum quae est ista fiducia qua confidis
ISA|36|5|aut quo consilio vel fortitudine rebellare disponis super quem habes fiduciam quia recessisti a me
ISA|36|6|ecce confidis super baculum harundineum confractum istum super Aegyptum cui si innisus fuerit homo intrabit in manu eius et perforabit eam sic Pharao rex Aegypti omnibus qui confidunt in eo
ISA|36|7|quod si responderis mihi in Domino Deo nostro confidimus nonne ipse est cuius abstulit Ezechias excelsa et altaria et dixit Iudae et Hierusalem coram altari isto adorabitis
ISA|36|8|et nunc trade te domino meo regi Assyriorum et dabo tibi duo milia equorum nec poteris ex te praebere ascensores eorum
ISA|36|9|et quomodo sustinebis faciem iudicis unius loci ex servis domini mei minoribus quod si confidis in Aegypto in quadriga et in equitibus
ISA|36|10|et nunc numquid sine Domino ascendi ad terram istam ut disperderem eam Dominus dixit ad me ascende super terram istam et disperde eam
ISA|36|11|et dixit Eliachim et Sobna et Ioae ad Rabsacen loquere ad servos tuos syra lingua intellegimus enim ne loquaris ad nos iudaice in auribus populi qui est super murum
ISA|36|12|et dixit ad eos Rabsaces numquid ad dominum tuum et ad te misit me dominus meus ut loquerer omnia verba ista et non potius ad viros qui sedent in muro ut comedant stercora sua et bibant urinam pedum suorum vobiscum
ISA|36|13|et stetit Rabsaces et clamavit voce magna iudaice et dixit audite verba regis magni regis Assyriorum
ISA|36|14|haec dicit rex non seducat vos Ezechias quia non poterit eruere vos
ISA|36|15|et non vobis tribuat fiduciam Ezechias super Domino dicens eruens liberabit nos Dominus non dabitur civitas ista in manu regis Assyriorum
ISA|36|16|nolite audire Ezechiam haec enim dicit rex Assyriorum facite mecum benedictionem et egredimini ad me et comedite unusquisque vineam suam et unusquisque ficum suam et bibite unusquisque aquam cisternae suae
ISA|36|17|donec veniam et tollam vos ad terram quae est ut terra vestra terram frumenti et vini terram panum et vinearum
ISA|36|18|ne conturbet vos Ezechias dicens Dominus liberabit nos numquid liberaverunt dii gentium unusquisque terram suam de manu regis Assyriorum
ISA|36|19|ubi est deus Emath et Arfad ubi est deus Seffarvaim numquid liberaverunt Samariam de manu mea
ISA|36|20|quis est ex omnibus diis terrarum istarum qui eruerit terram suam de manu mea ut eruat Dominus Hierusalem de manu mea
ISA|36|21|et siluerunt et non responderunt ei verbum mandaverat enim rex dicens ne respondeatis ei
ISA|36|22|et ingressus est Eliachim filius Helciae qui erat super domum et Sobna scriba et Ioae filius Asaph a commentariis ad Ezechiam scissis vestibus et nuntiaverunt ei verba Rabsacis
ISA|37|1|et factum est cum audisset rex Ezechias scidit vestimenta sua et obvolutus est sacco et intravit in domum Domini
ISA|37|2|et misit Eliachim qui erat super domum et Sobnam scribam et seniores de sacerdotibus opertos saccis ad Isaiam filium Amos prophetam
ISA|37|3|et dixerunt ad eum haec dicit Ezechias dies tribulationis et correptionis et blasphemiae dies haec quia venerunt filii usque ad partum et virtus non est parienti
ISA|37|4|si quo modo audiat Dominus Deus tuus verba Rabsaces quem misit rex Assyriorum dominus suus ad blasphemandum Deum viventem et obprobrandum sermonibus quos audivit Dominus Deus tuus leva ergo orationem pro reliquiis quae reppertae sunt
ISA|37|5|et venerunt servi regis Ezechiae ad Isaiam
ISA|37|6|et dixit ad eos Isaias haec dicetis domino vestro haec dicit Dominus ne timeas a facie verborum quae audisti quibus blasphemaverunt pueri regis Assyriorum me
ISA|37|7|ecce ego dabo ei spiritum et audiet nuntium et revertetur ad terram suam et corruere eum faciam gladio in terra sua
ISA|37|8|reversus est autem Rabsaces et invenit regem Assyriorum proeliantem adversus Lobna audierat enim quia profectus esset de Lachis
ISA|37|9|et audivit de Tharaca rege Aethiopiae dicentes egressus est ut pugnet contra te quod cum audisset misit nuntios ad Ezechiam dicens
ISA|37|10|haec dicetis Ezechiae regi Iudae loquentes non te decipiat Deus tuus in quo tu confidis dicens non dabitur Hierusalem in manu regis Assyriorum
ISA|37|11|ecce tu audisti omnia quae fecerunt reges Assyriorum omnibus terris quas subverterunt et tu poteris liberari
ISA|37|12|numquid eruerunt eos dii gentium quos subverterunt patres mei Gozan et Aran et Reseph et filios Eden qui erant in Thalassar
ISA|37|13|ubi est rex Emath et rex Arfad et rex urbis Seffarvaim Anahe et Ava
ISA|37|14|et tulit Ezechias libros de manu nuntiorum et legit eos et ascendit in domum Domini et expandit eos Ezechias coram Domino
ISA|37|15|et oravit Ezechias ad Dominum dicens
ISA|37|16|Domine exercituum Deus Israhel qui sedes super cherubin tu es Deus solus omnium regnorum terrae tu fecisti caelum et terram
ISA|37|17|inclina Domine aurem tuam et audi aperi Domine oculos tuos et vide et audi omnia verba Sennacherib quae misit ad blasphemandum Deum viventem
ISA|37|18|vere enim Domine desertas fecerunt reges Assyriorum terras et regiones earum
ISA|37|19|et dederunt deos earum igni non enim erant dii sed opera manuum hominum lignum et lapis et comminuerunt eos
ISA|37|20|et nunc Domine Deus noster salva nos de manu eius et cognoscant omnia regna terrae quia tu es Dominus solus
ISA|37|21|et misit Isaias filius Amos ad Ezechiam dicens haec dicit Dominus Deus Israhel pro quibus rogasti me de Sennacherib rege Assyriorum
ISA|37|22|hoc est verbum quod locutus est Dominus super eum despexit te subsannavit te virgo filia Sion post te caput movit filia Hierusalem
ISA|37|23|cui exprobrasti et quem blasphemasti et super quem exaltasti vocem et levasti altitudinem oculorum tuorum ad Sanctum Israhel
ISA|37|24|in manu servorum tuorum exprobrasti Domino et dixisti in multitudine quadrigarum mearum ego ascendi altitudinem montium iuga Libani et succidam excelsa cedrorum eius electas abietes illius et introibo altitudinem summitatis eius saltum Carmeli eius
ISA|37|25|ego fodi et bibi aquam et exsiccavi vestigio pedis mei omnes rivos aggerum
ISA|37|26|numquid non audisti quae olim fecerim ei ex diebus antiquis ego plasmavi illud et nunc adduxi et factum est in eradicationem collium conpugnantium et civitatum munitarum
ISA|37|27|habitatores earum breviata manu contremuerunt et confusi sunt facti sunt sicut faenum agri et gramen pascuae et herba tectorum quae exaruit antequam maturesceret
ISA|37|28|habitationem tuam et egressum tuum et introitum tuum cognovi et insaniam tuam contra me
ISA|37|29|cum fureres adversum me superbia tua ascendit in aures meas ponam ergo circulum in naribus tuis et frenum in labiis tuis et reducam te in viam per quam venisti
ISA|37|30|tibi autem hoc erit signum comede hoc anno quae sponte nascuntur et in anno secundo pomis vescere in anno autem tertio seminate et metite et plantate vineas et comedite fructum earum
ISA|37|31|et mittet id quod salvatum fuerit de domo Iuda et quod reliquum est radicem deorsum et faciet fructum sursum
ISA|37|32|quia de Hierusalem exibunt reliquiae et salvatio de monte Sion zelus Domini exercituum faciet istud
ISA|37|33|propterea haec dicit Dominus de rege Assyriorum non introibit civitatem hanc et non iaciet ibi sagittam et non occupabit eam clypeus et non mittet in circuitu eius aggerem
ISA|37|34|in via qua venit per eam revertetur et civitatem hanc non ingredietur dicit Dominus
ISA|37|35|et protegam civitatem istam ut salvem eam propter me et propter David servum meum
ISA|37|36|egressus est autem angelus Domini et percussit in castris Assyriorum centum octoginta quinque milia et surrexerunt mane et ecce omnes cadavera mortuorum
ISA|37|37|et egressus est et abiit et reversus est Sennacherib rex Assyriorum et habitavit in Nineve
ISA|37|38|et factum est cum adoraret in templo Nesrach deum suum Adramelech et Sarasar filii eius percusserunt eum gladio fugeruntque in terram Ararat et regnavit Asoraddon filius eius pro eo
ISA|38|1|in diebus illis aegrotavit Ezechias usque ad mortem et introivit ad eum Isaias filius Amos propheta et dixit ei haec dicit Dominus dispone domui tuae quia morieris tu et non vives
ISA|38|2|et convertit Ezechias faciem suam ad parietem et oravit ad Dominum
ISA|38|3|et dixit obsecro Domine memento quaeso quomodo ambulaverim coram te in veritate et in corde perfecto et quod bonum est in oculis tuis fecerim et flevit Ezechias fletu magno
ISA|38|4|et factum est verbum Domini ad Isaiam dicens
ISA|38|5|vade et dic Ezechiae haec dicit Dominus Deus David patris tui audivi orationem tuam vidi lacrimam tuam ecce ego adiciam super dies tuos quindecim annos
ISA|38|6|et de manu regis Assyriorum eruam te et civitatem istam et protegam eam
ISA|38|7|hoc autem tibi erit signum a Domino quia faciet Dominus verbum hoc quod locutus est
ISA|38|8|ecce ego reverti faciam umbram linearum per quas descenderat in horologio Ahaz in sole retrorsum decem lineis et reversus est sol decem lineis per gradus quos descenderat
ISA|38|9|scriptura Ezechiae regis Iuda cum aegrotasset et convaluisset de infirmitate sua
ISA|38|10|ego dixi in dimidio dierum meorum vadam ad portas inferi quaesivi residuum annorum meorum
ISA|38|11|dixi non videbo Dominum Dominum in terra viventium non aspiciam hominem ultra et habitatorem quievit
ISA|38|12|generatio mea ablata est et convoluta est a me quasi tabernaculum pastorum praecisa est velut a texente vita mea dum adhuc ordirer succidit me de mane usque ad vesperam finies me
ISA|38|13|sperabam usque ad mane quasi leo sic contrivit omnia ossa mea de mane usque ad vesperam finies me
ISA|38|14|sicut pullus hirundinis sic clamabo meditabor ut columba adtenuati sunt oculi mei suspicientes in excelsum Domine vim patior sponde pro me
ISA|38|15|quid dicam aut quid respondebit mihi cum ipse fecerit recogitabo omnes annos meos in amaritudine animae meae
ISA|38|16|Domine sic vivitur et in talibus vita spiritus mei corripies me et vivificabis me
ISA|38|17|ecce in pace amaritudo mea amarissima tu autem eruisti animam meam ut non periret proiecisti post tergum tuum omnia peccata mea
ISA|38|18|quia non infernus confitebitur tibi neque mors laudabit te non expectabunt qui descendunt in lacum veritatem tuam
ISA|38|19|vivens vivens ipse confitebitur tibi sicut et ego hodie pater filiis notam faciet veritatem tuam
ISA|38|20|Domine salvum me fac et psalmos nostros cantabimus cunctis diebus vitae nostrae in domo Domini
ISA|38|21|et iussit Isaias ut tollerent massam de ficis et cataplasmarent super vulnus et sanaretur
ISA|38|22|et dixit Ezechias quod erit signum quia ascendam in domo Domini
ISA|39|1|in tempore illo misit Marodach Baladan filius Baladan rex Babylonis libros et munera ad Ezechiam audierat enim quod aegrotasset et convaluisset
ISA|39|2|laetatus est autem super eis Ezechias et ostendit eis cellam aromatum et argenti et auri et odoramentorum et unguenti optimi et omnes apothecas supellectilis suae et universa quae inventa sunt in thesauris eius non fuit verbum quod non ostenderet eis Ezechias in domo sua et in omni potestate sua
ISA|39|3|introiit autem Isaias propheta ad regem Ezechiam et dixit ei quid dixerunt viri isti et unde venerunt ad te et dixit Ezechias de terra longinqua venerunt ad me de Babylone
ISA|39|4|et dixit quid viderunt in domo tua et dixit Ezechias omnia quae in domo mea sunt viderunt non fuit res quam non ostenderim eis in thesauris meis
ISA|39|5|et dixit Isaias ad Ezechiam audi verbum Domini exercituum
ISA|39|6|ecce dies venient et auferentur omnia quae in domo tua sunt et quae thesaurizaverunt patres tui usque ad diem hanc in Babylonem non relinquetur quicquam dicit Dominus
ISA|39|7|et de filiis tuis qui exibunt de te quos genueris tollent et erunt eunuchi in palatio regis Babylonis
ISA|39|8|et dixit Ezechias ad Isaiam bonum verbum Domini quod locutus est et dixit fiat tantum pax et veritas in diebus meis
ISA|40|1|consolamini consolamini populus meus dicit Deus vester
ISA|40|2|loquimini ad cor Hierusalem et avocate eam quoniam conpleta est malitia eius dimissa est iniquitas illius suscepit de manu Domini duplicia pro omnibus peccatis suis
ISA|40|3|vox clamantis in deserto parate viam Domini rectas facite in solitudine semitas Dei nostri
ISA|40|4|omnis vallis exaltabitur et omnis mons et collis humiliabitur et erunt prava in directa et aspera in vias planas
ISA|40|5|et revelabitur gloria Domini et videbit omnis caro pariter quod os Domini locutum est
ISA|40|6|vox dicentis clama et dixi quid clamabo omnis caro faenum et omnis gloria eius quasi flos agri
ISA|40|7|exsiccatum est faenum et cecidit flos quia spiritus Domini sufflavit in eo vere faenum est populus
ISA|40|8|exsiccatum est faenum cecidit flos verbum autem Dei nostri stabit in aeternum
ISA|40|9|super montem excelsum ascende tu quae evangelizas Sion exalta in fortitudine vocem tuam quae evangelizas Hierusalem exalta noli timere dic civitatibus Iudae ecce Deus vester
ISA|40|10|ecce Dominus Deus in fortitudine veniet et brachium eius dominabitur ecce merces eius cum eo et opus illius coram eo
ISA|40|11|sicut pastor gregem suum pascet in brachio suo congregabit agnos et in sinu suo levabit fetas ipse portabit
ISA|40|12|quis mensus est pugillo aquas et caelos palmo ponderavit quis adpendit tribus digitis molem terrae et libravit in pondere montes et colles in statera
ISA|40|13|quis adiuvit spiritum Domini aut quis consiliarius eius fuit et ostendit illi
ISA|40|14|cum quo iniit consilium et instruxit eum et docuit eum semitam iustitiae et erudivit eum scientiam et viam prudentiae ostendit illi
ISA|40|15|ecce gentes quasi stilla situlae et quasi momentum staterae reputatae sunt ecce insulae quasi pulvis exiguus
ISA|40|16|et Libanus non sufficiet ad succendendum et animalia eius non sufficient ad holocaustum
ISA|40|17|omnes gentes quasi non sint sic sunt coram eo et quasi nihilum et inane reputatae sunt ei
ISA|40|18|cui ergo similem fecistis Deum aut quam imaginem ponetis ei
ISA|40|19|numquid sculptile conflavit faber aut aurifex auro figuravit illud et lamminis argenteis argentarius
ISA|40|20|forte lignum et inputribile elegit artifex sapiens quaerit quomodo statuat simulacrum quod non moveatur
ISA|40|21|numquid non scietis numquid non audietis numquid non adnuntiatum est ab initio vobis numquid non intellexistis fundamenta terrae
ISA|40|22|qui sedet super gyrum terrae et habitatores eius sunt quasi lucustae qui extendit velut nihilum caelos et expandit eos sicut tabernaculum ad inhabitandum
ISA|40|23|qui dat secretorum scrutatores quasi non sint iudices terrae velut inane fecit
ISA|40|24|et quidem neque plantatos neque satos neque radicato in terra trunco eorum repente flavit in eos et aruerunt et turbo quasi stipulam auferet eos
ISA|40|25|et cui adsimilastis me et adaequastis dicit Sanctus
ISA|40|26|levate in excelsum oculos vestros et videte quis creavit haec qui educit in numero militiam eorum et omnes ex nomine vocat prae multitudine fortitudinis et roboris virtutisque eius neque unum reliquum fuit
ISA|40|27|quare dicis Iacob et loqueris Israhel abscondita est via mea a Domino et a Deo meo iudicium meum transibit
ISA|40|28|numquid nescis aut non audisti Deus sempiternus Dominus qui creavit terminos terrae non deficiet neque laborabit nec est investigatio sapientiae eius
ISA|40|29|qui dat lasso virtutem et his qui non sunt fortitudinem et robur multiplicat
ISA|40|30|deficient pueri et laborabunt et iuvenes in infirmitate cadent
ISA|40|31|qui autem sperant in Domino mutabunt fortitudinem adsument pinnas sicut aquilae current et non laborabunt ambulabunt et non deficient
ISA|41|1|taceant ad me insulae et gentes mutent fortitudinem accedant et tunc loquantur simul ad iudicium propinquemus
ISA|41|2|quis suscitavit ab oriente iustum vocavit eum ut sequeretur se dabit in conspectu eius gentes et reges obtinebit dabit quasi pulverem gladio eius sicut stipulam vento raptam arcui eius
ISA|41|3|persequetur eos transibit in pace semita in pedibus eius non apparebit
ISA|41|4|quis haec operatus est et fecit vocans generationes ab exordio ego Dominus primus et novissimus ego sum
ISA|41|5|viderunt insulae et timuerunt extrema terrae obstipuerunt adpropinquaverunt et accesserunt
ISA|41|6|unusquisque proximo suo auxiliatur et fratri suo dicit confortare
ISA|41|7|confortabit faber aerarius percutiens malleo eum qui cudebat tunc temporis dicens glutino bonum est et confortavit eum in clavis ut non moveatur
ISA|41|8|et tu Israhel serve meus Iacob quem elegi semen Abraham amici mei
ISA|41|9|in quo adprehendi te ab extremis terrae et a longinquis eius vocavi te et dixi tibi servus meus es tu elegi te et non abieci te
ISA|41|10|ne timeas quia tecum sum ego ne declines quia ego Deus tuus confortavi te et auxiliatus sum tui et suscepi te dextera iusti mei
ISA|41|11|ecce confundentur et erubescent omnes qui pugnant adversum te erunt quasi non sint et peribunt viri qui contradicunt tibi
ISA|41|12|quaeres eos et non invenies viros rebelles tuos erunt quasi non sint et veluti consumptio homines bellantes adversum te
ISA|41|13|quia ego Dominus Deus tuus adprehendens manum tuam dicensque tibi ne timeas ego adiuvi te
ISA|41|14|noli timere vermis Iacob qui mortui estis ex Israhel ego auxiliatus sum tui dicit Dominus et redemptor tuus Sanctus Israhel
ISA|41|15|ego posui te quasi plaustrum triturans novum habens rostra serrantia triturabis montes et comminues et colles quasi pulverem pones
ISA|41|16|ventilabis eos et ventus tollet et turbo disperget eos et tu exultabis in Domino in Sancto Israhel laetaberis
ISA|41|17|egeni et pauperes quaerunt aquas et non sunt lingua eorum siti aruit ego Dominus exaudiam eos Deus Israhel non derelinquam eos
ISA|41|18|aperiam in supinis collibus flumina et in medio camporum fontes ponam desertum in stagna aquarum et terram inviam in rivos aquarum
ISA|41|19|dabo in solitudine cedrum et spinam et myrtum et lignum olivae ponam in deserto abietem ulmum et buxum simul
ISA|41|20|ut videant et sciant et recogitent et intellegant pariter quia manus Domini fecit hoc et Sanctus Israhel creavit illud
ISA|41|21|prope facite iudicium vestrum dicit Dominus adferte si quid forte habetis dixit Rex Iacob
ISA|41|22|accedant et nuntient nobis quaecumque ventura sunt priora quae fuerint nuntiate et ponemus cor nostrum et sciemus novissima eorum et quae ventura sunt indicate nobis
ISA|41|23|adnuntiate quae ventura sunt in futurum et sciemus quia dii estis vos bene quoque aut male si potestis facite et loquamur et videamus simul
ISA|41|24|ecce vos estis ex nihilo et opus vestrum ex eo quod non est abominatio est qui elegit vos
ISA|41|25|suscitavi ab aquilone et venit ab ortu solis vocabit nomen meum et adducet magistratus quasi lutum et velut plastes conculcans humum
ISA|41|26|quis adnuntiavit ab exordio ut sciamus et a principio ut dicamus iustus es non est neque adnuntians neque praedicens neque audiens sermones vestros
ISA|41|27|primus ad Sion dicet ecce adsunt et Hierusalem evangelistam dabo
ISA|41|28|et vidi et non erat neque ex istis quisquam qui iniret consilium et interrogatus responderet verbum
ISA|41|29|ecce omnes iniusti et vana opera eorum ventus et inane simulacra eorum
ISA|42|1|ecce servus meus suscipiam eum electus meus conplacuit sibi in illo anima mea dedi spiritum meum super eum iudicium gentibus proferet
ISA|42|2|non clamabit neque accipiet personam nec audietur foris vox eius
ISA|42|3|calamum quassatum non conteret et linum fumigans non extinguet in veritate educet iudicium
ISA|42|4|non erit tristis neque turbulentus donec ponat in terra iudicium et legem eius insulae expectabunt
ISA|42|5|haec dicit Dominus Deus creans caelos et extendens eos firmans terram et quae germinant ex ea dans flatum populo qui est super eam et spiritum calcantibus eam
ISA|42|6|ego Dominus vocavi te in iustitia et adprehendi manum tuam et servavi et dedi te in foedus populi in lucem gentium
ISA|42|7|ut aperires oculos caecorum et educeres de conclusione vinctum de domo carceris sedentes in tenebris
ISA|42|8|ego Dominus hoc est nomen meum gloriam meam alteri non dabo et laudem meam sculptilibus
ISA|42|9|quae prima fuerant ecce venerunt nova quoque ego adnuntio antequam oriantur audita vobis faciam
ISA|42|10|cantate Domino canticum novum laus eius ab extremis terrae qui descenditis in mare et plenitudo eius insulae et habitatores earum
ISA|42|11|sublevetur desertum et civitates eius in domibus habitabit Cedar laudate habitatores Petrae de vertice montium clamabunt
ISA|42|12|ponent Domino gloriam et laudem eius in insulis nuntiabunt
ISA|42|13|Dominus sicut fortis egredietur sicut vir proeliator suscitabit zelum vociferabitur et clamabit super inimicos suos confortabitur
ISA|42|14|tacui semper silui patiens fui sicut pariens loquar dissipabo et absorbebo simul
ISA|42|15|desertos faciam montes et colles et omne gramen eorum exsiccabo et ponam flumina in insulas et stagna arefaciam
ISA|42|16|et ducam caecos in via quam nesciunt in semitis quas ignoraverunt ambulare eos faciam ponam tenebras coram eis in lucem et prava in recta haec verba feci eis et non dereliqui eos
ISA|42|17|conversi sunt retrorsum confundantur confusione qui confidunt in sculptili qui dicunt conflatili vos dii nostri
ISA|42|18|surdi audite et caeci intuemini ad videndum
ISA|42|19|quis caecus nisi servus meus et surdus nisi ad quem nuntios meos misi quis caecus nisi qui venundatus est quis caecus nisi servus Domini
ISA|42|20|qui vides multa nonne custodies qui apertas habes aures nonne audies
ISA|42|21|et Dominus voluit ut sanctificaret eum et magnificaret legem et extolleret
ISA|42|22|ipse autem populus direptus et vastatus laqueus iuvenum omnes et in domibus carcerum absconditi sunt facti sunt in rapinam nec est qui eruat in direptionem et non est qui dicat redde
ISA|42|23|quis est in vobis qui audiat hoc adtendat et auscultet futura
ISA|42|24|quis dedit in direptionem Iacob et Israhel vastantibus nonne Dominus ipse cui peccavimus et noluerunt in viis eius ambulare et non audierunt legem eius
ISA|42|25|et effudit super eum indignationem furoris sui et forte bellum et conbusit eum in circuitu et non cognovit et succendit eum et non intellexit
ISA|43|1|et nunc haec dicit Dominus creans te Iacob et formans te Israhel noli timere quia redemi te et vocavi nomine tuo meus es tu
ISA|43|2|cum transieris per aquas tecum ero et flumina non operient te cum ambulaveris in igne non conbureris et flamma non ardebit in te
ISA|43|3|quia ego Dominus Deus tuus Sanctus Israhel salvator tuus dedi propitiationem tuam Aegyptum Aethiopiam et Saba pro te
ISA|43|4|ex quo honorabilis factus es in oculis meis et gloriosus ego dilexi te et dabo homines pro te et populos pro anima tua
ISA|43|5|noli timere quoniam tecum ego sum ab oriente adducam semen tuum et ab occidente congregabo te
ISA|43|6|dicam aquiloni da et austro noli prohibere adfer filios meos de longinquo et filias meas ab extremis terrae
ISA|43|7|et omnem qui invocat nomen meum in gloriam meam creavi eum et formavi eum et feci eum
ISA|43|8|educ foras populum caecum et oculos habentem surdum et aures ei sunt
ISA|43|9|omnes gentes congregatae sunt simul et collectae sunt tribus quis in vobis adnuntiet istud et quae prima sunt audire nos faciat dent testes eorum et iustificentur et audiant et dicant vere
ISA|43|10|vos testes mei dicit Dominus et servus meus quem elegi ut sciatis et credatis mihi et intellegatis quia ego ipse sum ante me non est formatus deus et post me non erit
ISA|43|11|ego sum ego sum Dominus et non est absque me salvator
ISA|43|12|ego adnuntiavi et salvavi auditum feci et non fuit in vobis alienus vos testes mei dicit Dominus et ego Deus
ISA|43|13|et ab initio ego ipse et non est qui de manu mea eruat operabor et quis avertet illud
ISA|43|14|haec dicit Dominus redemptor vester Sanctus Israhel propter vos emisi Babylonem et detraxi vectes universos et Chaldeos in navibus suis gloriantes
ISA|43|15|ego Dominus Sanctus vester creans Israhel Rex vester
ISA|43|16|haec dicit Dominus qui dedit in mari viam et in aquis torrentibus semitam
ISA|43|17|qui eduxit quadrigam et equum agmen et robustum simul obdormierunt nec resurgent contriti sunt quasi linum et extincti sunt
ISA|43|18|ne memineritis priorum et antiqua ne intueamini
ISA|43|19|ecce ego facio nova et nunc orientur utique cognoscetis ea ponam in deserto viam et in invio flumina
ISA|43|20|glorificabit me bestia agri dracones et strutiones quia dedi in deserto aquas flumina in invio ut darem potum populo meo electo meo
ISA|43|21|populum istum formavi mihi laudem meam narrabit
ISA|43|22|non me invocasti Iacob nec laborasti in me Israhel
ISA|43|23|non obtulisti mihi arietem holocausti tui et victimis tuis non glorificasti me non te servire feci in oblatione nec laborem tibi praebui in ture
ISA|43|24|non emisti mihi argento calamum et adipe victimarum tuarum non inebriasti me verumtamen servire me fecisti in peccatis tuis praebuisti mihi laborem in iniquitatibus tuis
ISA|43|25|ego sum ego sum ipse qui deleo iniquitates tuas propter me et peccatorum tuorum non recordabor
ISA|43|26|reduc me in memoriam et iudicemur simul narra si quid habes ut iustificeris
ISA|43|27|pater tuus primus peccavit et interpretes tui praevaricati sunt in me
ISA|43|28|et contaminavi principes sanctos dedi ad internicionem Iacob et Israhel in blasphemiam
ISA|44|1|et nunc audi Iacob serve meus et Israhel quem elegi
ISA|44|2|haec dicit Dominus faciens et formans te ab utero auxiliator tuus noli timere serve meus Iacob et Rectissime quem elegi
ISA|44|3|effundam enim aquas super sitientem et fluenta super aridam effundam spiritum meum super semen tuum et benedictionem meam super stirpem tuam
ISA|44|4|et germinabunt inter herbas quasi salices iuxta praeterfluentes aquas
ISA|44|5|iste dicet Domini ego sum et ille vocabit in nomine Iacob et hic scribet manu sua Domino et in nomine Israhel adsimilabitur
ISA|44|6|haec dicit Dominus rex Israhel et redemptor eius Dominus exercituum ego primus et ego novissimus et absque me non est deus
ISA|44|7|quis similis mei vocet et adnuntiet et ordinem exponat mihi ex quo constitui populum antiquum ventura et quae futura sunt adnuntient eis
ISA|44|8|nolite timere neque conturbemini ex tunc audire te feci et adnuntiavi vos estis testes mei numquid est deus absque me et formator quem ego non noverim
ISA|44|9|plastae idoli omnes nihil sunt et amantissima eorum non proderunt eis ipsi sunt testes eorum quia non vident neque intellegunt ut confundantur
ISA|44|10|quis formavit deum et sculptile conflavit ad nihil utile
ISA|44|11|ecce omnes participes eius confundentur fabri enim sunt ex hominibus convenient omnes stabunt et pavebunt et confundentur simul
ISA|44|12|faber ferrarius lima operatus est in prunis et in malleis formavit illud et operatus est in brachio fortitudinis suae esuriet et deficiet non bibet aquam et lassescet
ISA|44|13|artifex lignarius extendit normam formavit illud in runcina fecit illud in angularibus et in circino tornavit illud et fecit imaginem viri quasi speciosum hominem habitantem in domo
ISA|44|14|succidit cedros tulit ilicem et quercum quae steterat inter ligna saltus plantavit pinum quam pluvia nutrivit
ISA|44|15|et facta est hominibus in focum sumpsit ex eis et calefactus est et succendit et coxit panes de reliquo autem operatus est deum et adoravit fecit sculptile et curvatus est ante illud
ISA|44|16|medium eius conbusit igni et de medio eius carnes comedit coxit pulmentum et saturatus est et calefactus est et dixit va calefactus sum vidi focum
ISA|44|17|reliquum autem eius deum fecit sculptile sibi curvatur ante illud et adorat illud et obsecrat dicens libera me quia deus meus es tu
ISA|44|18|nescierunt neque intellexerunt lutati enim sunt ne videant oculi eorum et ne intellegant corde suo
ISA|44|19|non recogitant in mente sua neque cognoscunt neque sentiunt ut dicant medietatem eius conbusi igne et coxi super carbones eius panes coxi carnes et comedi et de reliquo eius idolum faciam ante truncum ligni procidam
ISA|44|20|pars eius cinis est cor insipiens adoravit illud et non liberabit animam suam neque dicet forte mendacium est in dextera mea
ISA|44|21|memento horum Iacob et Israhel quoniam servus meus es tu formavi te servus meus es tu Israhel non oblivisceris mei
ISA|44|22|delevi ut nubem iniquitates tuas et quasi nebulam peccata tua revertere ad me quoniam redemi te
ISA|44|23|laudate caeli quoniam fecit Dominus iubilate extrema terrae resonate montes laudationem saltus et omne lignum eius quoniam redemit Dominus Iacob et Israhel gloriabitur
ISA|44|24|haec dicit Dominus redemptor tuus et formator tuus ex utero ego sum Dominus faciens omnia extendens caelos solus stabiliens terram et nullus mecum
ISA|44|25|irrita faciens signa divinorum et ariolos in furorem vertens convertens sapientes retrorsum et scientiam eorum stultam faciens
ISA|44|26|suscitans verbum servi sui et consilium nuntiorum suorum conplens qui dico Hierusalem habitaberis et civitatibus Iuda aedificabimini et deserta eius suscitabo
ISA|44|27|qui dico profundo desolare et flumina tua arefaciam
ISA|44|28|qui dico Cyro pastor meus es et omnem voluntatem meam conplebis qui dico Hierusalem aedificaberis et templo fundaberis
ISA|45|1|haec dicit Dominus christo meo Cyro cuius adprehendi dexteram ut subiciam ante faciem eius gentes et dorsa regum vertam et aperiam coram eo ianuas et portae non cludentur
ISA|45|2|ego ante te ibo et gloriosos terrae humiliabo portas aereas conteram et vectes ferreos confringam
ISA|45|3|et dabo tibi thesauros absconditos et arcana secretorum ut scias quia ego Dominus qui voco nomen tuum Deus Israhel
ISA|45|4|propter servum meum Iacob et Israhel electum meum et vocavi te in nomine tuo adsimilavi te et non cognovisti me
ISA|45|5|ego Dominus et non est amplius extra me non est deus accinxi te et non cognovisti me
ISA|45|6|ut sciant hii qui ab ortu solis et qui ab occidente quoniam absque me non est ego Dominus et non est alter
ISA|45|7|formans lucem et creans tenebras faciens pacem et creans malum ego Dominus faciens omnia haec
ISA|45|8|rorate caeli desuper et nubes pluant iustum aperiatur terra et germinet salvatorem et iustitia oriatur simul ego Dominus creavi eum
ISA|45|9|vae qui contradicit fictori suo testa de samiis terrae numquid dicet lutum figulo suo quid facis et opus tuum absque manibus est
ISA|45|10|vae qui dicit patri quid generas et mulieri quid parturis
ISA|45|11|haec dicit Dominus Sanctus Israhel plastes eius ventura interrogate me super filios meos et super opus manuum mearum mandastis mihi
ISA|45|12|ego feci terram et hominem super eam creavi ego manus meae tetenderunt caelos et omni militiae eorum mandavi
ISA|45|13|ego suscitavi eum ad iustitiam et omnes vias eius dirigam ipse aedificabit civitatem meam et captivitatem meam dimittet non in pretio neque in muneribus dicit Dominus Deus exercituum
ISA|45|14|haec dicit Dominus labor Aegypti et negotiatio Aethiopiae et Sabaim viri sublimes ad te transibunt et tui erunt post te ambulabunt vincti manicis pergent et te adorabunt teque deprecabuntur tantum in te est Deus et non est absque te deus
ISA|45|15|vere tu es Deus absconditus Deus Israhel salvator
ISA|45|16|confusi sunt et erubuerunt omnes simul abierunt in confusione fabricatores errorum
ISA|45|17|Israhel salvatus est in Domino salute aeterna non confundemini et non erubescetis usque in saeculum saeculi
ISA|45|18|quia haec dicit Dominus creans caelos ipse Deus formans terram et faciens eam ipse plastes eius non in vanum creavit eam ut habitetur formavit eam ego Dominus et non est alius
ISA|45|19|non in abscondito locutus sum in loco terrae tenebroso non dixi semini Iacob frustra quaerite me ego Dominus loquens iustitiam adnuntians recta
ISA|45|20|congregamini et venite et accedite simul qui salvati estis ex gentibus nescierunt qui levant lignum sculpturae suae et rogant deum non salvantem
ISA|45|21|adnuntiate et venite et consiliamini simul quis auditum fecit hoc ab initio ex tunc praedixit illud numquid non ego Dominus et non est ultra Deus absque me Deus iustus et salvans non est praeter me
ISA|45|22|convertimini ad me et salvi eritis omnes fines terrae quia ego Deus et non est alius
ISA|45|23|in memet ipso iuravi egredietur de ore meo iustitiae verbum et non revertetur quia mihi curvabunt omnia genu et iurabit omnis lingua
ISA|45|24|ergo in Domino dicet meae sunt iustitiae et imperium ad eum venient et confundentur omnes qui repugnant ei
ISA|45|25|in Domino iustificabitur et laudabitur omne semen Israhel
ISA|46|1|conflatus est Bel contritus est Nabo facta sunt simulacra eorum bestiis et iumentis onera vestra gravi pondere usque ad lassitudinem
ISA|46|2|contabuerunt et contrita sunt simul non potuerunt salvare portantem et anima eorum in captivitatem ibit
ISA|46|3|audite me domus Iacob et omne residuum domus Israhel qui portamini a meo utero qui gestamini a mea vulva
ISA|46|4|usque ad senectam ego ipse et usque ad canos ego portabo ego feci et ego feram et ego portabo et salvabo
ISA|46|5|cui adsimilastis me et adaequastis et conparastis me et fecistis similem
ISA|46|6|qui confertis aurum de sacculo et argentum statera ponderatis conducentes aurificem ut faciat deum et procidunt et adorant
ISA|46|7|portant illud in umeris gestantes et ponentes in loco suo et stabit ac de loco suo non movebitur sed et cum clamaverint ad eum non audiet de tribulatione non salvabit eos
ISA|46|8|mementote istud et fundamini redite praevaricatores ad cor
ISA|46|9|recordamini prioris saeculi quoniam ego sum Deus et non est ultra Deus nec est similis mei
ISA|46|10|adnuntians ab exordio novissimum et ab initio quae necdum facta sunt dicens consilium meum stabit et omnis voluntas mea fiet
ISA|46|11|vocans ab oriente avem et de terra longinqua virum voluntatis meae et locutus sum et adducam illud creavi et faciam illud
ISA|46|12|audite me duro corde qui longe estis a iustitia
ISA|46|13|prope feci iustitiam meam non elongabitur et salus mea non morabitur dabo in Sion salutem et Israheli gloriam meam
ISA|47|1|descende sede in pulverem virgo filia Babylon sede in terra non est solium filiae Chaldeorum quia ultra non vocaberis mollis et tenera
ISA|47|2|tolle molam et mole farinam denuda turpitudinem tuam discoperi umerum revela crus transi flumina
ISA|47|3|revelabitur ignominia tua et videbitur obprobrium tuum ultionem capiam et non resistet mihi homo
ISA|47|4|redemptor noster Dominus exercituum nomen illius Sanctus Israhel
ISA|47|5|sede tace et intra in tenebras filia Chaldeorum quia non vocaberis ultra domina regnorum
ISA|47|6|iratus sum super populum meum contaminavi hereditatem meam et dedi eos in manu tua non posuisti eis misericordias super senem adgravasti iugum tuum valde
ISA|47|7|et dixisti in sempiternum ero domina non posuisti haec super cor tuum neque recordata es novissimi tui
ISA|47|8|et nunc audi haec delicata et habitans confidenter quae dicis in corde tuo ego sum et non est praeter me amplius non sedebo vidua et ignorabo sterilitatem
ISA|47|9|venient tibi duo haec subito in die una sterilitas et viduitas universa venerunt super te propter multitudinem maleficiorum tuorum et propter duritiam incantatorum tuorum vehementem
ISA|47|10|et fiduciam habuisti in malitia tua et dixisti non est qui videat me sapientia tua et scientia tua haec decepit te et dixisti in corde tuo ego sum et praeter me non est altera
ISA|47|11|veniet super te malum et nescies ortum eius et inruet super te calamitas quam non poteris expiare veniet super te repente miseria quam nescies
ISA|47|12|sta cum incantatoribus tuis et cum multitudine maleficiorum tuorum in quibus laborasti ab adulescentia tua si forte quid prosit tibi aut si possis fieri fortior
ISA|47|13|defecisti in multitudine consiliorum tuorum stent et salvent te augures caeli qui contemplabantur sidera et supputabant menses ut ex eis adnuntiarent ventura tibi
ISA|47|14|ecce facti sunt quasi stipula ignis conbusit eos non liberabunt animam suam de manu flammae non sunt prunae quibus calefiant nec focus ut sedeant ad eum
ISA|47|15|sic facta sunt tibi in quibuscumque laboraveras negotiatores tui ab adulescentia tua unusquisque in via sua erraverunt non est qui salvet te
ISA|48|1|audite hoc domus Iacob qui vocamini nomine Israhel et de aquis Iuda existis qui iuratis in nomine Domini et Dei Israhel recordamini non in veritate neque in iustitia
ISA|48|2|de civitate enim sancta vocati sunt et super Deum Israhel constabiliti sunt Dominus exercituum nomen eius
ISA|48|3|priora ex tunc adnuntiavi et ex ore meo exierunt et audita feci ea repente operatus sum et venerunt
ISA|48|4|scivi enim quia durus es tu et nervus ferreus cervix tua et frons tua aerea
ISA|48|5|praedixi tibi ex tunc antequam venirent indicavi tibi ne forte diceres idola mea fecerunt haec et sculptilia mea et conflatilia mandaverunt ista
ISA|48|6|quae audisti vide omnia vos autem non adnuntiastis audita feci tibi nova ex nunc et conservata quae nescis
ISA|48|7|nunc creata sunt et non ex tunc et ante diem et non audisti ea ne forte dicas ecce cognovi ea
ISA|48|8|neque audisti neque cognovisti neque ex tunc aperta est auris tua scio enim quia praevaricans praevaricabis et transgressorem ex ventre vocavi te
ISA|48|9|propter nomen meum longe faciam furorem meum et laude mea infrenabo te ne intereas
ISA|48|10|ecce excoxi te sed non quasi argentum elegi te in camino paupertatis
ISA|48|11|propter me propter me faciam ut non blasphemer et gloriam meam alteri non dabo
ISA|48|12|audi me Iacob et Israhel quem ego voco ego ipse ego primus et ego novissimus
ISA|48|13|manus quoque mea fundavit terram et dextera mea mensa est caelos ego vocabo eos et stabunt simul
ISA|48|14|congregamini omnes vos et audite quis de eis adnuntiavit haec Dominus dilexit eum faciet voluntatem suam in Babylone et brachium suum in Chaldeis
ISA|48|15|ego ego locutus sum et vocavi eum adduxi eum et directa est via eius
ISA|48|16|accedite ad me et audite hoc non a principio in abscondito locutus sum ex tempore antequam fieret ibi eram et nunc Dominus Deus misit me et spiritus eius
ISA|48|17|haec dicit Dominus redemptor tuus Sanctus Israhel ego Dominus Deus tuus docens te utilia gubernans te in via qua ambulas
ISA|48|18|utinam adtendisses mandata mea facta fuisset sicut flumen pax tua et iustitia tua sicut gurgites maris
ISA|48|19|et fuisset quasi harena semen tuum et stirps uteri tui ut lapilli eius non interisset et non fuisset adtritum nomen eius a facie mea
ISA|48|20|egredimini de Babylone fugite a Chaldeis in voce exultationis adnuntiate auditum facite hoc efferte illud usque ad extrema terrae dicite redemit Dominus servum suum Iacob
ISA|48|21|non sitierunt in deserto cum educeret eos aquam de petra produxit eis et scidit petram et fluxerunt aquae
ISA|48|22|non est pax dicit Dominus impiis
ISA|49|1|audite insulae et adtendite populi de longe Dominus ab utero vocavit me de ventre matris meae recordatus est nominis mei
ISA|49|2|et posuit os meum quasi gladium acutum in umbra manus suae protexit me et posuit me sicut sagittam electam in faretra sua abscondit me
ISA|49|3|et dixit mihi servus meus es tu Israhel quia in te gloriabor
ISA|49|4|et ego dixi in vacuum laboravi sine causa et vane fortitudinem meam consumpsi ergo iudicium meum cum Domino et opus meum cum Deo meo
ISA|49|5|et nunc dicit Dominus formans me ex utero servum sibi ut reducam Iacob ad eum et Israhel non congregabitur et glorificatus sum in oculis Domini et Deus meus factus est fortitudo mea
ISA|49|6|et dixit parum est ut sis mihi servus ad suscitandas tribus Iacob et feces Israhel convertendas dedi te in lucem gentium ut sis salus mea usque ad extremum terrae
ISA|49|7|haec dicit Dominus redemptor Israhel Sanctus eius ad contemptibilem animam ad abominatam gentem ad servum dominorum reges videbunt et consurgent principes et adorabunt propter Dominum quia fidelis est et Sanctum Israhel qui elegit te
ISA|49|8|haec dicit Dominus in tempore placito exaudivi te et in die salutis auxiliatus sum tui et servavi te et dedi te in foedus populi ut suscitares terram et possideres hereditates dissipatas
ISA|49|9|ut diceres his qui vincti sunt exite et his qui in tenebris revelamini super vias pascentur et in omnibus planis pascua eorum
ISA|49|10|non esurient neque sitient et non percutiet eos aestus et sol quia miserator eorum reget eos et ad fontes aquarum portabit eos
ISA|49|11|et ponam omnes montes meos in viam et semitae meae exaltabuntur
ISA|49|12|ecce isti de longe venient et ecce illi ab aquilone et mari et isti de terra australi
ISA|49|13|laudate caeli et exulta terra iubilate montes laudem quia consolatus est Dominus populum suum et pauperum suorum miserebitur
ISA|49|14|et dixit Sion dereliquit me Dominus et Dominus oblitus est mei
ISA|49|15|numquid oblivisci potest mulier infantem suum ut non misereatur filio uteri sui et si illa oblita fuerit ego tamen non obliviscar tui
ISA|49|16|ecce in manibus meis descripsi te muri tui coram oculis meis semper
ISA|49|17|venerunt structores tui destruentes te et dissipantes a te exibunt
ISA|49|18|leva in circuitu oculos tuos et vide omnes isti congregati sunt venerunt tibi vivo ego dicit Dominus quia omnibus his velut ornamento vestieris et circumdabis tibi eos quasi sponsa
ISA|49|19|quia deserta tua et solitudines tuae et terra ruinae tuae nunc angusta erunt prae habitatoribus et longe fugabuntur qui absorbebant te
ISA|49|20|adhuc dicent in auribus tuis filii sterilitatis tuae angustus mihi est locus fac spatium mihi ut habitem
ISA|49|21|et dices in corde tuo quis genuit mihi istos ego sterilis et non pariens transmigrata et captiva et istos quis enutrivit ego destituta et sola et isti ubi hic erant
ISA|49|22|haec dicit Dominus Deus ecce levo ad gentes manum meam et ad populos exaltabo signum meum et adferent filios tuos in ulnis et filias tuas super umeros portabunt
ISA|49|23|et erunt reges nutricii tui et reginae nutrices tuae vultu in terra dimisso adorabunt te et pulverem pedum tuorum lingent et scies quia ego Dominus super quo non confundentur qui expectant eum
ISA|49|24|numquid tolletur a forte praeda aut quod captum fuerit a robusto salvum esse poterit
ISA|49|25|quia haec dicit Dominus equidem et captivitas a forte tolletur et quod ablatum fuerit a robusto salvabitur eos vero qui iudicaverunt te ego iudicabo et filios tuos ego salvabo
ISA|49|26|et cibabo hostes tuos carnibus suis et quasi musto sanguine suo inebriabuntur et sciet omnis caro quia ego Dominus salvans te et redemptor tuus Fortis Iacob
ISA|50|1|haec dicit Dominus quis est hic liber repudii matris vestrae quo dimisi eam aut quis est creditor meus cui vendidi vos ecce in iniquitatibus vestris venditi estis et in sceleribus vestris dimisi matrem vestram
ISA|50|2|quia veni et non erat vir vocavi et non erat qui audiret numquid adbreviata et parvula facta est manus mea ut non possim redimere aut non est in me virtus ad liberandum ecce in increpatione mea desertum faciam mare ponam flumina in siccum conputrescent pisces sine aqua et morientur in siti
ISA|50|3|induam caelos tenebris et saccum ponam operimentum eorum
ISA|50|4|Dominus dedit mihi linguam eruditam ut sciam sustentare eum qui lassus est verbo erigit mane mane erigit mihi aurem ut audiam quasi magistrum
ISA|50|5|Dominus Deus aperuit mihi aurem ego autem non contradico retrorsum non abii
ISA|50|6|corpus meum dedi percutientibus et genas meas vellentibus faciem meam non averti ab increpantibus et conspuentibus
ISA|50|7|Dominus Deus auxiliator meus ideo non sum confusus ideo posui faciem meam ut petram durissimam et scio quoniam non confundar
ISA|50|8|iuxta est qui iustificat me quis contradicet mihi stemus simul quis est adversarius meus accedat ad me
ISA|50|9|ecce Dominus Deus auxiliator meus quis est qui condemnet me ecce omnes quasi vestimentum conterentur tinea comedet eos
ISA|50|10|quis ex vobis timens Dominum audiens vocem servi sui qui ambulavit in tenebris et non est lumen ei speret in nomine Domini et innitatur super Deum suum
ISA|50|11|ecce omnes vos accendentes ignem accincti flammis ambulate in lumine ignis vestri et in flammis quas succendistis de manu mea factum est hoc vobis in doloribus dormietis
ISA|51|1|audite me qui sequimini quod iustum est et quaeritis Dominum adtendite ad petram unde excisi estis et ad cavernam laci de qua praecisi estis
ISA|51|2|adtendite ad Abraham patrem vestrum et ad Sarram quae peperit vos quia unum vocavi eum et benedixi ei et multiplicavi eum
ISA|51|3|consolabitur ergo Dominus et Sion consolabitur omnes ruinas eius et ponet desertum eius quasi delicias et solitudinem eius quasi hortum Domini gaudium et laetitia invenietur in ea gratiarum actio et vox laudis
ISA|51|4|adtendite ad me populus meus et tribus mea me audite quia lex a me exiet et iudicium meum in lucem populorum requiescet
ISA|51|5|prope est iustus meus egressus est salvator meus et brachia mea populos iudicabunt me insulae expectabunt et brachium meum sustinebunt
ISA|51|6|levate in caelum oculos vestros et videte sub terra deorsum quia caeli sicut fumus liquescent et terra sicut vestimentum adteretur et habitatores eius sicut haec interibunt salus autem mea in sempiternum erit et iustitia mea non deficiet
ISA|51|7|audite me qui scitis iustum populus lex mea in corde eorum nolite timere obprobrium hominum et blasphemias eorum ne metuatis
ISA|51|8|sicut enim vestimentum sic comedet eos vermis et sicut lanam sic devorabit eos tinea salus autem mea in sempiternum erit et iustitia mea in generationes generationum
ISA|51|9|consurge consurge induere fortitudinem brachium Domini consurge sicut in diebus antiquis in generationibus saeculorum numquid non tu percussisti superbum vulnerasti draconem
ISA|51|10|numquid non tu siccasti mare aquam abyssi vehementis qui posuisti profundum maris viam ut transirent liberati
ISA|51|11|et nunc qui redempti sunt a Domino revertentur et venient in Sion laudantes et laetitia sempiterna super capita eorum gaudium et laetitiam tenebunt fugiet dolor et gemitus
ISA|51|12|ego ego ipse consolabor vos quis tu ut timeres ab homine mortali et a filio hominis qui quasi faenum ita arescet
ISA|51|13|et oblitus es Domini factoris tui qui tetendit caelos et fundavit terram et formidasti iugiter tota die a facie furoris eius qui te tribulabat et paraverat ad perdendum ubi nunc est furor tribulantis
ISA|51|14|cito veniet gradiens ad aperiendum et non interficiet usque ad internicionem nec deficiet panis eius
ISA|51|15|ego autem sum Dominus Deus tuus qui conturbo mare et intumescunt fluctus eius Dominus exercituum nomen meum
ISA|51|16|posui verba mea in ore tuo et in umbra manus meae protexi te ut plantes caelos et fundes terram et dicas ad Sion populus meus es tu
ISA|51|17|elevare elevare consurge Hierusalem quae bibisti de manu Domini calicem irae eius usque ad fundum calicis soporis bibisti et epotasti usque ad feces
ISA|51|18|non est qui sustentet eam ex omnibus filiis quos genuit et non est qui adprehendat manum eius ex omnibus filiis quos enutrivit
ISA|51|19|duo sunt quae occurrerunt tibi quis contristabitur super te vastitas et contritio et fames et gladius quis consolabitur te
ISA|51|20|filii tui proiecti sunt dormierunt in capite omnium viarum sicut bestia inlaqueata pleni indignatione Domini increpatione Dei tui
ISA|51|21|idcirco audi hoc paupercula et ebria non a vino
ISA|51|22|haec dicit Dominator tuus Dominus et Deus tuus qui pugnavit pro populo suo ecce tuli de manu tua calicem soporis fundum calicis indignationis meae non adicies ut bibas illud ultra
ISA|51|23|et ponam illud in manu eorum qui te humiliaverunt et dixerunt animae tuae incurvare ut transeamus et posuisti ut terram corpus tuum et quasi viam transeuntibus
ISA|52|1|consurge consurge induere fortitudine tua Sion induere vestimentis gloriae tuae Hierusalem civitas sancti quia non adiciet ultra ut pertranseat per te incircumcisus et inmundus
ISA|52|2|excutere de pulvere consurge sede Hierusalem solve vincula colli tui captiva filia Sion
ISA|52|3|quia haec dicit Dominus gratis venundati estis et sine argento redimemini
ISA|52|4|quia haec dicit Dominus Deus in Aegyptum descendit populus meus in principio ut colonus esset ibi et Assur absque ulla causa calumniatus est eum
ISA|52|5|et nunc quid mihi est hic dicit Dominus quoniam ablatus est populus meus gratis dominatores eius inique agunt dicit Dominus et iugiter tota die nomen meum blasphematur
ISA|52|6|propter hoc sciet populus meus nomen meum in die illa quia ego ipse qui loquebar ecce adsum
ISA|52|7|quam pulchri super montes pedes adnuntiantis et praedicantis pacem adnuntiantis bonum praedicantis salutem dicentis Sion regnavit Deus tuus
ISA|52|8|vox speculatorum tuorum levaverunt vocem simul laudabunt quia oculum ad oculum videbunt cum converterit Dominus Sion
ISA|52|9|gaudete et laudate simul deserta Hierusalem quia consolatus est Dominus populum suum redemit Hierusalem
ISA|52|10|paravit Dominus brachium sanctum suum in oculis omnium gentium et videbunt omnes fines terrae salutare Dei nostri
ISA|52|11|recedite recedite exite inde pollutum nolite tangere exite de medio eius mundamini qui fertis vasa Domini
ISA|52|12|quoniam non in tumultu exibitis nec in fuga properabitis praecedet enim vos Dominus et congregabit vos Deus Israhel
ISA|52|13|ecce intelleget servus meus exaltabitur et elevabitur et sublimis erit valde
ISA|52|14|sicut obstipuerunt super te multi sic inglorius erit inter viros aspectus eius et forma eius inter filios hominum
ISA|52|15|iste asperget gentes multas super ipsum continebunt reges os suum quia quibus non est narratum de eo viderunt et qui non audierunt contemplati sunt
ISA|53|1|quis credidit auditui nostro et brachium Domini cui revelatum est
ISA|53|2|et ascendet sicut virgultum coram eo et sicut radix de terra sitienti non est species ei neque decor et vidimus eum et non erat aspectus et desideravimus eum
ISA|53|3|despectum et novissimum virorum virum dolorum et scientem infirmitatem et quasi absconditus vultus eius et despectus unde nec reputavimus eum
ISA|53|4|vere languores nostros ipse tulit et dolores nostros ipse portavit et nos putavimus eum quasi leprosum et percussum a Deo et humiliatum
ISA|53|5|ipse autem vulneratus est propter iniquitates nostras adtritus est propter scelera nostra disciplina pacis nostrae super eum et livore eius sanati sumus
ISA|53|6|omnes nos quasi oves erravimus unusquisque in viam suam declinavit et Dominus posuit in eo iniquitatem omnium nostrum
ISA|53|7|oblatus est quia ipse voluit et non aperuit os suum sicut ovis ad occisionem ducetur et quasi agnus coram tondente obmutescet et non aperiet os suum
ISA|53|8|de angustia et de iudicio sublatus est generationem eius quis enarrabit quia abscisus est de terra viventium propter scelus populi mei percussit eum
ISA|53|9|et dabit impios pro sepultura et divitem pro morte sua eo quod iniquitatem non fecerit neque dolus fuerit in ore eius
ISA|53|10|et Dominus voluit conterere eum in infirmitate si posuerit pro peccato animam suam videbit semen longevum et voluntas Domini in manu eius dirigetur
ISA|53|11|pro eo quod laboravit anima eius videbit et saturabitur in scientia sua iustificabit ipse iustus servus meus multos et iniquitates eorum ipse portabit
ISA|53|12|ideo dispertiam ei plurimos et fortium dividet spolia pro eo quod tradidit in morte animam suam et cum sceleratis reputatus est et ipse peccatum multorum tulit et pro transgressoribus rogavit
ISA|54|1|lauda sterilis quae non paris decanta laudem et hinni quae non pariebas quoniam multi filii desertae magis quam eius quae habebat virum dicit Dominus
ISA|54|2|dilata locum tentorii tui et pelles tabernaculorum tuorum extende ne parcas longos fac funiculos tuos et clavos tuos consolida
ISA|54|3|ad dexteram enim et ad levam penetrabis et semen tuum gentes hereditabit et civitates desertas inhabitabit
ISA|54|4|noli timere quia non confunderis neque erubescas non enim te pudebit quia confusionis adulescentiae tuae oblivisceris et obprobrii viduitatis tuae non recordaberis amplius
ISA|54|5|quia dominabitur tui qui fecit te Dominus exercituum nomen eius et redemptor tuus Sanctus Israhel Deus omnis terrae vocabitur
ISA|54|6|quia ut mulierem derelictam et maerentem spiritu vocavit te Dominus et uxorem ab adulescentia abiectam dixit Deus tuus
ISA|54|7|ad punctum in modico dereliqui te et in miserationibus magnis congregabo te
ISA|54|8|in momento indignationis abscondi faciem meam parumper a te et in misericordia sempiterna misertus sum tui dixit redemptor tuus Dominus
ISA|54|9|sicut in diebus Noe istud mihi est cui iuravi ne inducerem aquas Noe ultra super terram sic iuravi ut non irascar tibi et non increpem te
ISA|54|10|montes enim commovebuntur et colles contremescent misericordia autem mea non recedet et foedus pacis meae non movebitur dixit miserator tuus Dominus
ISA|54|11|paupercula tempestate convulsa absque ulla consolatione ecce ego sternam per ordinem lapides tuos et fundabo te in sapphyris
ISA|54|12|et ponam iaspidem propugnacula tua et portas tuas in lapides sculptos et omnes terminos tuos in lapides desiderabiles
ISA|54|13|universos filios tuos doctos a Domino et multitudinem pacis filiis tuis
ISA|54|14|et in iustitia fundaberis recede procul a calumnia quia non timebis et a pavore quia non adpropinquabit tibi
ISA|54|15|ecce accola veniet qui non erat mecum advena quondam tuus adiungetur tibi
ISA|54|16|ecce ego creavi fabrum sufflantem in igne prunas et proferentem vas in opus suum et ego creavi interfectorem ad disperdendum
ISA|54|17|omne vas quod fictum est contra te non dirigetur et omnem linguam resistentem tibi in iudicio iudicabis haec hereditas servorum Domini et iustitia eorum apud me dicit Dominus
ISA|55|1|o omnes sitientes venite ad aquas et qui non habetis argentum properate emite et comedite venite emite absque argento et absque ulla commutatione vinum et lac
ISA|55|2|quare adpenditis argentum non in panibus et laborem vestrum non in saturitate audite audientes me et comedite bonum et delectabitur in crassitudine anima vestra
ISA|55|3|inclinate aurem vestram et venite ad me audite et vivet anima vestra et feriam vobis pactum sempiternum misericordias David fideles
ISA|55|4|ecce testem populis dedi eum ducem ac praeceptorem gentibus
ISA|55|5|ecce gentem quam nesciebas vocabis et gentes quae non cognoverunt te ad te current propter Dominum Deum tuum et Sanctum Israhel quia glorificavit te
ISA|55|6|quaerite Dominum dum inveniri potest invocate eum dum prope est
ISA|55|7|derelinquat impius viam suam et vir iniquus cogitationes suas et revertatur ad Dominum et miserebitur eius et ad Deum nostrum quoniam multus est ad ignoscendum
ISA|55|8|non enim cogitationes meae cogitationes vestrae neque viae vestrae viae meae dicit Dominus
ISA|55|9|quia sicut exaltantur caeli a terra sic exaltatae sunt viae meae a viis vestris et cogitationes meae a cogitationibus vestris
ISA|55|10|et quomodo descendit imber et nix de caelo et illuc ultra non revertitur sed inebriat terram et infundit eam et germinare eam facit et dat semen serenti et panem comedenti
ISA|55|11|sic erit verbum meum quod egredietur de ore meo non revertetur ad me vacuum sed faciet quaecumque volui et prosperabitur in his ad quae misi illud
ISA|55|12|quia in laetitia egrediemini et in pace deducemini montes et colles cantabunt coram vobis laudem et omnia ligna regionis plaudent manu
ISA|55|13|pro saliunca ascendet abies et pro urtica crescet myrtus et erit Dominus nominatus in signum aeternum quod non auferetur
ISA|56|1|haec dicit Dominus custodite iudicium et facite iustitiam quia iuxta est salus mea ut veniat et iustitia mea ut reveletur
ISA|56|2|beatus vir qui facit hoc et filius hominis qui adprehendit istud custodiens sabbatum ne polluat illud custodiens manus suas ne faciat omne malum
ISA|56|3|et non dicat filius advenae qui adheret Domino dicens separatione dividet me Dominus a populo suo et non dicat eunuchus ecce ego lignum aridum
ISA|56|4|quia haec dicit Dominus eunuchis qui custodierint sabbata mea et elegerint quae volui et tenuerint foedus meum
ISA|56|5|dabo eis in domo mea et in muris meis locum et nomen melius a filiis et filiabus nomen sempiternum dabo eis quod non peribit
ISA|56|6|et filios advenae qui adherent Domino ut colant eum et diligant nomen eius ut sint ei in servos omnem custodientem sabbatum ne polluat illud et tenentem foedus meum
ISA|56|7|adducam eos in montem sanctum meum et laetificabo eos in domo orationis meae holocausta eorum et victimae eorum placebunt mihi super altari meo quia domus mea domus orationis vocabitur cunctis populis
ISA|56|8|ait Dominus Deus qui congregat dispersos Israhel adhuc congregabo ad eum congregatos eius
ISA|56|9|omnes bestiae agri venite ad devorandum universae bestiae saltus
ISA|56|10|speculatores eius caeci omnes nescierunt universi canes muti non valentes latrare videntes vana dormientes et amantes somnia
ISA|56|11|et canes inpudentissimi nescierunt saturitatem ipsi pastores ignoraverunt intellegentiam omnes in viam suam declinaverunt unusquisque ad avaritiam suam a summo usque ad novissimum
ISA|56|12|venite sumamus vinum et impleamur ebrietate et erit sicut hodie sic et cras et multo amplius
ISA|57|1|iustus perit et nemo est qui recogitet in corde suo et viri misericordiae colliguntur quia non est qui intellegat a facie enim malitiae collectus est iustus
ISA|57|2|veniat pax requiescat in cubili suo qui ambulavit in directione sua
ISA|57|3|vos autem accedite huc filii auguratricis semen adulteri et fornicariae
ISA|57|4|super quem lusistis super quem dilatastis os et eiecistis linguam numquid non vos filii scelesti semen mendax
ISA|57|5|qui consolamini in diis subter omne lignum frondosum immolantes parvulos in torrentibus subter inminentes petras
ISA|57|6|in partibus torrentis pars tua haec est sors tua et ipsis effudisti libamen obtulisti sacrificium numquid super his non indignabor
ISA|57|7|super montem excelsum et sublimem posuisti cubile tuum et illuc ascendisti ut immolares hostias
ISA|57|8|et post ostium et retro postem posuisti memoriale tuum quia iuxta me discoperuisti et suscepisti adulterum dilatasti cubile tuum et pepigisti cum eis dilexisti stratum eorum manu aperta
ISA|57|9|et ornasti te regi unguento et multiplicasti pigmenta tua misisti legatos tuos procul et humiliata es usque ad inferos
ISA|57|10|in multitudine viae tuae laborasti non dixisti quiescam vitam manus tuae invenisti propterea non rogasti
ISA|57|11|pro quo sollicita timuisti quia mentita es et mei non es recordata neque cogitasti in corde tuo quia ego tacens et quasi non videns et mei oblita es
ISA|57|12|ego adnuntiabo iustitiam tuam et opera tua non proderunt tibi
ISA|57|13|cum clamaveris liberent te congregati tui et omnes eos auferet ventus tollet aura qui autem fiduciam habet mei hereditabit terram et possidebit montem sanctum meum
ISA|57|14|et dicam viam facite praebete iter declinate de semita auferte offendicula de via populi mei
ISA|57|15|quia haec dicit Excelsus et Sublimis habitans aeternitatem et sanctum nomen eius in excelso et in sancto habitans et cum contrito et humili spiritu ut vivificet spiritum humilium et vivificet cor contritorum
ISA|57|16|non enim in sempiternum litigabo neque usque ad finem irascar quia spiritus a facie mea egredietur et flatus ego faciam
ISA|57|17|propter iniquitatem avaritiae eius iratus sum et percussi eum abscondi et indignatus sum et abiit vagus in via cordis sui
ISA|57|18|vias eius vidi et dimisi eum et reduxi eum et reddidi consolationes ipsi et lugentibus eius
ISA|57|19|creavi fructum labiorum pacem pacem ei qui longe est et qui prope dixit Dominus et sanavi eum
ISA|57|20|impii autem quasi mare fervens quod quiescere non potest et redundant fluctus eius in conculcationem et lutum
ISA|57|21|non est pax dixit Deus meus impiis
ISA|58|1|clama ne cesses quasi tuba exalta vocem tuam et adnuntia populo meo scelera eorum et domui Iacob peccata eorum
ISA|58|2|me etenim de die in diem quaerunt et scire vias meas volunt quasi gens quae iustitiam fecerit et quae iudicium Dei sui non reliquerit rogant me iudicia iustitiae adpropinquare Deo volunt
ISA|58|3|quare ieiunavimus et non aspexisti humiliavimus animam nostram et nescisti ecce in die ieiunii vestri invenitur voluntas et omnes debitores vestros repetitis
ISA|58|4|ecce ad lites et contentiones ieiunatis et percutitis pugno impie nolite ieiunare sicut usque ad hanc diem ut audiatur in excelso clamor vester
ISA|58|5|numquid tale est ieiunium quod elegi per diem adfligere hominem animam suam numquid contorquere quasi circulum caput suum et saccum et cinerem sternere numquid istud vocabis ieiunium et diem acceptabilem Domino
ISA|58|6|nonne hoc est magis ieiunium quod elegi dissolve conligationes impietatis solve fasciculos deprimentes dimitte eos qui confracti sunt liberos et omne onus disrumpe
ISA|58|7|frange esurienti panem tuum et egenos vagosque induc in domum tuam cum videris nudum operi eum et carnem tuam ne despexeris
ISA|58|8|tunc erumpet quasi mane lumen tuum et sanitas tua citius orietur et anteibit faciem tuam iustitia tua et gloria Domini colliget te
ISA|58|9|tunc invocabis et Dominus exaudiet clamabis et dicet ecce adsum si abstuleris de medio tui catenam et desieris digitum extendere et loqui quod non prodest
ISA|58|10|cum effuderis esurienti animam tuam et animam adflictam repleveris orietur in tenebris lux tua et tenebrae tuae erunt sicut meridies
ISA|58|11|et requiem tibi dabit Dominus semper et implebit splendoribus animam tuam et ossa tua liberabit et eris quasi hortus inriguus et sicut fons aquarum cuius non deficient aquae
ISA|58|12|et aedificabuntur in te deserta saeculorum fundamenta generationis et generationis suscitabis et vocaberis aedificator sepium avertens semitas in quietem
ISA|58|13|si averteris a sabbato pedem tuum facere voluntatem tuam in die sancto meo et vocaveris sabbatum delicatum et sanctum Domini gloriosum et glorificaveris eum dum non facis vias tuas et non invenitur voluntas tua ut loquaris sermonem
ISA|58|14|tunc delectaberis super Domino et sustollam te super altitudines terrae et cibabo te hereditate Iacob patris tui os enim Domini locutum est
ISA|59|1|ecce non est adbreviata manus Domini ut salvare nequeat neque adgravata est auris eius ut non exaudiat
ISA|59|2|sed iniquitates vestrae diviserunt inter vos et Deum vestrum et peccata vestra absconderunt faciem eius a vobis ne exaudiret
ISA|59|3|manus enim vestrae pollutae sunt sanguine et digiti vestri iniquitate labia vestra locuta sunt mendacium et lingua vestra iniquitatem fatur
ISA|59|4|non est qui invocet iustitiam neque est qui iudicet vere sed confidunt in nihili et loquuntur vanitates conceperunt laborem et pepererunt iniquitatem
ISA|59|5|ova aspidum ruperunt et telas araneae texuerunt qui comederit de ovis eorum morietur et quod confotum est erumpet in regulum
ISA|59|6|telae eorum non erunt in vestimentum neque operientur operibus suis opera eorum opera inutilia et opus iniquitatis in manibus eorum
ISA|59|7|pedes eorum ad malum currunt et festinant ut effundant sanguinem innocentem cogitationes eorum cogitationes inutiles vastitas et contritio in viis eorum
ISA|59|8|viam pacis nescierunt et non est iudicium in gressibus eorum semitae eorum incurvatae sunt eis omnis qui calcat in ea ignorat pacem
ISA|59|9|propter hoc elongatum est iudicium a nobis et non adprehendet nos iustitia expectavimus lucem et ecce tenebrae splendorem et in tenebris ambulavimus
ISA|59|10|palpavimus sicut caeci parietem et quasi absque oculis adtrectavimus inpegimus meridie quasi in tenebris in caligosis quasi mortui
ISA|59|11|rugiemus quasi ursi omnes et quasi columbae meditantes gememus expectavimus iudicium et non est salutem et elongata est a nobis
ISA|59|12|multiplicatae sunt enim iniquitates nostrae coram te et peccata nostra responderunt nobis quia scelera nostra nobiscum et iniquitates nostras cognovimus
ISA|59|13|peccare et mentiri contra Dominum et aversi sumus ne iremus post tergum Dei nostri ut loqueremur calumniam et transgressionem concepimus et locuti sumus de corde verba mendacii
ISA|59|14|et conversum est retrorsum iudicium et iustitia longe stetit quia corruit in platea veritas et aequitas non potuit ingredi
ISA|59|15|et facta est veritas in oblivione et qui recessit a malo praedae patuit et vidit Dominus et malum apparuit in oculis eius quia non est iudicium
ISA|59|16|et vidit quia non est vir et aporiatus est quia non est qui occurrat et salvavit sibi brachium suum et iustitia eius ipsa confirmavit eum
ISA|59|17|indutus est iustitia ut lorica et galea salutis in capite eius indutus est vestimentis ultionis et opertus est quasi pallio zeli
ISA|59|18|sicut ad vindictam quasi ad retributionem indignationis hostibus suis et vicissitudinem inimicis suis insulis vicem reddet
ISA|59|19|et timebunt qui ab occidente nomen Domini et qui ab ortu solis gloriam eius cum venerit quasi fluvius violentus quem spiritus Domini cogit
ISA|59|20|et venerit Sion redemptor et eis qui redeunt ab iniquitate in Iacob dicit Dominus
ISA|59|21|hoc foedus meum cum eis dicit Dominus spiritus meus qui est in te et verba mea quae posui in ore tuo non recedent de ore tuo et de ore seminis tui et de ore seminis seminis tui dixit Dominus amodo et usque in sempiternum
ISA|60|1|surge inluminare quia venit lumen tuum et gloria Domini super te orta est
ISA|60|2|quia ecce tenebrae operient terram et caligo populos super te autem orietur Dominus et gloria eius in te videbitur
ISA|60|3|et ambulabunt gentes in lumine tuo et reges in splendore ortus tui
ISA|60|4|leva in circuitu oculos tuos et vide omnes isti congregati sunt venerunt tibi filii tui de longe venient et filiae tuae in latere sugent
ISA|60|5|tunc videbis et afflues et mirabitur et dilatabitur cor tuum quando conversa fuerit ad te multitudo maris fortitudo gentium venerit tibi
ISA|60|6|inundatio camelorum operiet te dromedariae Madian et Efa omnes de Saba venient aurum et tus deferentes et laudem Domino adnuntiantes
ISA|60|7|omne pecus Cedar congregabitur tibi arietes Nabaioth ministrabunt tibi offerentur super placabili altari meo et domum maiestatis meae glorificabo
ISA|60|8|qui sunt isti qui ut nubes volant et quasi columbae ad fenestras suas
ISA|60|9|me enim insulae expectant et naves maris in principio ut adducam filios tuos de longe argentum eorum et aurum eorum cum eis nomini Domini Dei tui et Sancto Israhel quia glorificavit te
ISA|60|10|et aedificabunt filii peregrinorum muros tuos et reges eorum ministrabunt tibi in indignatione enim mea percussi te et in reconciliatione mea misertus sum tui
ISA|60|11|et aperientur portae tuae iugiter die et nocte non claudentur ut adferatur ad te fortitudo gentium et reges earum adducantur
ISA|60|12|gens enim et regnum quod non servierit tibi peribit et gentes solitudine vastabuntur
ISA|60|13|gloria Libani ad te veniet abies et buxus et pinus simul ad ornandum locum sanctificationis meae et locum pedum meorum glorificabo
ISA|60|14|et venient ad te curvi filii eorum qui humiliaverunt te et adorabunt vestigia pedum tuorum omnes qui detrahebant tibi et vocabunt te civitatem Domini Sion Sancti Israhel
ISA|60|15|pro eo quod fuisti derelicta et odio habita et non erat qui per te transiret ponam te in superbiam saeculorum gaudium in generationem et generationem
ISA|60|16|et suges lac gentium et mamilla regum lactaberis et scies quia ego Dominus salvans te et redemptor tuus Fortis Iacob
ISA|60|17|pro aere adferam aurum et pro ferro adferam argentum et pro lignis aes et pro lapidibus ferrum et ponam visitationem tuam pacem et praepositos tuos iustitiam
ISA|60|18|non audietur ultra iniquitas in terra tua vastitas et contritio in terminis tuis et occupabit salus muros tuos et portas tuas laudatio
ISA|60|19|non erit tibi amplius sol ad lucendum per diem nec splendor lunae inluminabit te sed erit tibi Dominus in lucem sempiternam et Deus tuus in gloriam tuam
ISA|60|20|non occidet ultra sol tuus et luna tua non minuetur quia Dominus erit in lucem sempiternam et conplebuntur dies luctus tui
ISA|60|21|populus autem tuus omnes iusti in perpetuum hereditabunt terram germen plantationis meae opus manus meae ad glorificandum
ISA|60|22|minimus erit in mille et parvulus in gentem fortissimam ego Dominus in tempore eius subito faciam istud
ISA|61|1|spiritus Domini super me eo quod unxerit Dominus me ad adnuntiandum mansuetis misit me ut mederer contritis corde et praedicarem captivis indulgentiam et clausis apertionem
ISA|61|2|ut praedicarem annum placabilem Domini et diem ultionis Deo nostro ut consolarer omnes lugentes
ISA|61|3|ut ponerem lugentibus Sion et darem eis coronam pro cinere oleum gaudii pro luctu pallium laudis pro spiritu maeroris et vocabuntur in ea fortes iustitiae plantatio Domini ad glorificandum
ISA|61|4|et aedificabunt deserta a saeculo et ruinas antiquas erigent et instaurabunt civitates desertas dissipatas in generationem et generationem
ISA|61|5|et stabunt alieni et pascent pecora vestra et filii peregrinorum agricolae et vinitores vestri erunt
ISA|61|6|vos autem sacerdotes Domini vocabimini ministri Dei nostri dicetur vobis fortitudinem gentium comedetis et in gloria earum superbietis
ISA|61|7|pro confusione vestra duplici et rubore laudabunt partem eorum propter hoc in terra sua duplicia possidebunt laetitia sempiterna erit eis
ISA|61|8|quia ego Dominus diligens iudicium odio habens rapinam in holocausto et dabo opus eorum in veritate et foedus perpetuum feriam eis
ISA|61|9|et scietur in gentibus semen eorum et germen eorum in medio populorum omnes qui viderint eos cognoscent eos quia isti sunt semen cui benedixit Dominus
ISA|61|10|gaudens gaudebo in Domino et exultabit anima mea in Deo meo quia induit me vestimentis salutis et indumento iustitiae circumdedit me quasi sponsum decoratum corona et quasi sponsam ornatam monilibus suis
ISA|61|11|sicut enim terra profert germen suum et sicut hortus semen suum germinat sic Dominus Deus germinabit iustitiam et laudem coram universis gentibus
ISA|62|1|propter Sion non tacebo et propter Hierusalem non quiescam donec egrediatur ut splendor iustus eius et salvator eius ut lampas accendatur
ISA|62|2|et videbunt gentes iustum tuum et cuncti reges inclitum tuum et vocabitur tibi nomen novum quod os Domini nominabit
ISA|62|3|et eris corona gloriae in manu Domini et diadema regni in manu Dei tui
ISA|62|4|non vocaberis ultra Derelicta et terra tua non vocabitur amplius Desolata sed vocaberis Voluntas mea in ea et terra tua Inhabitata quia conplacuit Domino in te et terra tua inhabitabitur
ISA|62|5|habitabit enim iuvenis cum virgine et habitabunt in te filii tui et gaudebit sponsus super sponsam gaudebit super te Deus tuus
ISA|62|6|super muros tuos Hierusalem constitui custodes tota die et tota nocte perpetuo non tacebunt qui reminiscimini Domini ne taceatis
ISA|62|7|et ne detis silentium ei donec stabiliat et donec ponat Hierusalem laudem in terra
ISA|62|8|iuravit Dominus in dextera sua et in brachio fortitudinis suae si dedero triticum tuum ultra cibum inimicis tuis et si biberint filii alieni vinum tuum in quo laborasti
ISA|62|9|quia qui congregabunt illud comedent et laudabunt Dominum et qui conportant illud bibent in atriis sanctis meis
ISA|62|10|transite transite per portas praeparate viam populo planum facite iter et eligite lapides elevate signum ad populos
ISA|62|11|ecce Dominus auditum fecit in extremis terrae dicite filiae Sion ecce salvator tuus venit ecce merces eius cum eo et opus eius coram illo
ISA|62|12|et vocabunt eos Populus sanctus Redempti a Domino tu autem vocaberis Quaesita civitas et non Derelicta
ISA|63|1|quis est iste qui venit de Edom tinctis vestibus de Bosra iste formonsus in stola sua gradiens in multitudine fortitudinis suae ego qui loquor iustitiam et propugnator sum ad salvandum
ISA|63|2|quare ergo rubrum est indumentum tuum et vestimenta tua sicut calcantium in torculari
ISA|63|3|torcular calcavi solus et de gentibus non est vir mecum calcavi eos in furore meo et conculcavi eos in ira mea et aspersus est sanguis eorum super vestimenta mea et omnia indumenta mea inquinavi
ISA|63|4|dies enim ultionis in corde meo annus redemptionis meae venit
ISA|63|5|circumspexi et non erat auxiliator quaesivi et non fuit qui adiuvaret et salvavit mihi brachium meum et indignatio mea ipsa auxiliata est mihi
ISA|63|6|et conculcavi populos in furore meo et inebriavi eos in indignatione mea et detraxi in terra virtutem eorum
ISA|63|7|miserationum Domini recordabor laudem Domini super omnibus quae reddidit nobis Dominus et super multitudinem bonorum domui Israhel quae largitus est eis secundum indulgentiam suam et secundum multitudinem misericordiarum suarum
ISA|63|8|et dixit verumtamen populus meus est filii non negantes et factus est eis salvator
ISA|63|9|in omni tribulatione eorum non est tribulatus et angelus faciei eius salvavit eos in dilectione sua et in indulgentia sua ipse redemit eos et portavit eos et levavit eos cunctis diebus saeculi
ISA|63|10|ipsi autem ad iracundiam provocaverunt et adflixerunt spiritum Sancti eius et conversus est eis in inimicum et ipse debellavit eos
ISA|63|11|et recordatus est dierum saeculi Mosi populi sui ubi est qui eduxit eos de mari cum pastoribus gregis sui ubi est qui posuit in medio eius spiritum Sancti sui
ISA|63|12|qui eduxit ad dexteram Mosen brachio maiestatis suae qui scidit aquas ante eos ut faceret sibi nomen sempiternum
ISA|63|13|qui duxit eos per abyssos quasi equum in deserto non inpingentem
ISA|63|14|quasi animal in campo descendens spiritus Domini ductor eius fuit sic adduxisti populum tuum ut faceres tibi nomen gloriae
ISA|63|15|adtende de caelo et vide de habitaculo sancto tuo et gloriae tuae ubi est zelus tuus et fortitudo tua multitudo viscerum tuorum et miserationum tuarum super me continuerunt se
ISA|63|16|tu enim pater noster et Abraham nescivit nos et Israhel ignoravit nos tu Domine pater noster redemptor noster a saeculo nomen tuum
ISA|63|17|quare errare nos fecisti Domine de viis tuis indurasti cor nostrum ne timeremus te convertere propter servos tuos tribus hereditatis tuae
ISA|63|18|quasi nihilum possederunt populum sanctum tuum hostes nostri conculcaverunt sanctificationem tuam
ISA|63|19|facti sumus quasi in principio cum non dominareris nostri neque invocaretur nomen tuum super nos
ISA|64|1|utinam disrumperes caelos et descenderes a facie tua montes defluerent
ISA|64|2|sicut exustio ignis tabescerent aquae arderent igni ut notum fieret nomen tuum inimicis tuis a facie tua gentes turbarentur
ISA|64|3|cum feceris mirabilia non sustinebimus descendisti et a facie tua montes defluxerunt
ISA|64|4|a saeculo non audierunt neque auribus perceperunt oculus non vidit Deus absque te quae praeparasti expectantibus te
ISA|64|5|occurristi laetanti et facienti iustitiam in viis tuis recordabuntur tui ecce tu iratus es et peccavimus in ipsis fuimus semper et salvabimur
ISA|64|6|et facti sumus ut inmundus omnes nos quasi pannus menstruatae universae iustitiae nostrae et cecidimus quasi folium universi et iniquitates nostrae quasi ventus abstulerunt nos
ISA|64|7|non est qui invocet nomen tuum qui consurgat et teneat te abscondisti faciem tuam a nobis et adlisisti nos in manu iniquitatis nostrae
ISA|64|8|et nunc Domine pater noster es tu nos vero lutum et fictor noster et opera manuum tuarum omnes nos
ISA|64|9|ne irascaris Domine satis et ne ultra memineris iniquitatis ecce respice populus tuus omnes nos
ISA|64|10|civitas sancti tui facta est deserta Sion deserta facta est Hierusalem desolata
ISA|64|11|domus sanctificationis nostrae et gloriae nostrae ubi laudaverunt te patres nostri facta est in exustionem ignis et omnia desiderabilia nostra versa sunt in ruinas
ISA|64|12|numquid super his continebis te Domine tacebis et adfliges nos vehementer
ISA|65|1|quaesierunt me qui ante non interrogabant invenerunt qui non quaesierunt me dixi ecce ego ecce ego ad gentem quae non vocabat nomen meum
ISA|65|2|expandi manus meas tota die ad populum incredulum qui graditur in via non bona post cogitationes suas
ISA|65|3|populus qui ad iracundiam provocat me ante faciem meam semper qui immolant in hortis et sacrificant super lateres
ISA|65|4|qui habitant in sepulchris et in delubris idolorum dormiunt qui comedunt carnem suillam et ius profanum in vasis eorum
ISA|65|5|qui dicunt recede a me non adpropinques mihi quia inmundus es isti fumus erunt in furore meo ignis ardens tota die
ISA|65|6|ecce scriptum est coram me non tacebo sed reddam et retribuam in sinu eorum
ISA|65|7|iniquitates vestras et iniquitates patrum vestrorum simul dicit Dominus qui sacrificaverunt super montes et super colles exprobraverunt mihi et remetiar opus eorum primum in sinu eorum
ISA|65|8|haec dicit Dominus quomodo si inveniatur granum in botro et dicatur ne dissipes illud quoniam benedictio est sic faciam propter servos meos ut non disperdam totum
ISA|65|9|et educam de Iacob semen et de Iuda possidentem montes meos et hereditabunt eam electi mei et servi mei habitabunt ibi
ISA|65|10|et erunt campestria in caulas gregum et vallis Achor in cubile armentorum populo meo qui requisierunt me
ISA|65|11|et vos qui dereliquistis Dominum qui obliti estis montem sanctum meum qui ponitis Fortunae mensam et libatis super eam
ISA|65|12|numerabo vos in gladio et omnes in caede corruetis pro eo quod vocavi et non respondistis locutus sum et non audistis et faciebatis malum in oculis meis et quae nolui elegistis
ISA|65|13|propter hoc haec dicit Dominus Deus ecce servi mei comedent et vos esurietis ecce servi mei bibent et vos sitietis
ISA|65|14|ecce servi mei laetabuntur et vos confundemini ecce servi mei laudabunt prae exultatione cordis et vos clamabitis prae dolore cordis et prae contritione spiritus ululabitis
ISA|65|15|et dimittetis nomen vestrum in iuramentum electis meis et interficiet te Dominus Deus et servos suos vocabit nomine alio
ISA|65|16|in quo qui benedictus est super terram benedicetur in Deo amen et qui iurat in terra iurabit in Deo amen quia oblivioni traditae sunt angustiae priores et quia absconditae sunt ab oculis nostris
ISA|65|17|ecce enim ego creo caelos novos et terram novam et non erunt in memoria priora et non ascendent super cor
ISA|65|18|sed gaudebitis et exultabitis usque in sempiternum in his quae ego creo quia ecce ego creo Hierusalem exultationem et populum eius gaudium
ISA|65|19|et exultabo in Hierusalem et gaudebo in populo meo et non audietur in eo ultra vox fletus et vox clamoris
ISA|65|20|non erit ibi amplius infans dierum et senex qui non impleat dies suos quoniam puer centum annorum morietur et peccator centum annorum maledictus erit
ISA|65|21|et aedificabunt domos et habitabunt et plantabunt vineas et comedent fructum earum
ISA|65|22|non aedificabunt et alius habitabit non plantabunt et alius comedet secundum dies enim ligni erunt dies populi mei et opera manuum eorum inveterabunt
ISA|65|23|electis meis non laborabunt frustra neque generabunt in conturbatione quia semen benedictorum Domini est et nepotes eorum cum eis
ISA|65|24|eritque antequam clament ego exaudiam adhuc illis loquentibus ego audiam
ISA|65|25|lupus et agnus pascentur simul et leo et bos comedent paleas et serpenti pulvis panis eius non nocebunt neque occident in omni monte sancto meo dicit Dominus
ISA|66|1|haec dicit Dominus caelum sedis mea et terra scabillum pedum meorum quae ista domus quam aedificabitis mihi et quis iste locus quietis meae
ISA|66|2|omnia haec manus mea fecit et facta sunt universa ista dicit Dominus ad quem autem respiciam nisi ad pauperculum et contritum spiritu et trementem sermones meos
ISA|66|3|qui immolat bovem quasi qui interficiat virum qui mactat pecus quasi qui excerebret canem qui offert oblationem quasi qui sanguinem suillum offerat qui recordatur turis quasi qui benedicat idolo haec omnia elegerunt in viis suis et in abominationibus suis anima eorum delectata est
ISA|66|4|unde et ego eligam inlusiones eorum et quae timebant adducam eis quia vocavi et non erat qui responderet locutus sum et non audierunt feceruntque malum in oculis meis et quae nolui elegerunt
ISA|66|5|audite verbum Domini qui tremetis ad verbum eius dixerunt fratres vestri odientes vos et abicientes propter nomen meum glorificetur Dominus et videbimus in laetitia vestra ipsi autem confundentur
ISA|66|6|vox populi de civitate vox de templo vox Domini reddentis retributionem inimicis suis
ISA|66|7|antequam parturiret peperit antequam veniret partus eius peperit masculum
ISA|66|8|quis audivit umquam tale et quis vidit huic simile numquid parturiet terra in die una aut parietur gens simul quia parturivit et peperit Sion filios suos
ISA|66|9|numquid ego qui alios parere facio ipse non pariam dicit Dominus si ego qui generationem ceteris tribuo sterilis ero ait Dominus Deus tuus
ISA|66|10|laetamini cum Hierusalem et exultate in ea omnes qui diligitis eam gaudete cum ea gaudio universi qui lugetis super eam
ISA|66|11|ut sugatis et repleamini ab ubere consolationis eius ut mulgeatis et deliciis affluatis ab omnimoda gloria eius
ISA|66|12|quia haec dicit Dominus ecce ego declinabo super eam quasi fluvium pacis et quasi torrentem inundantem gloriam gentium quam sugetis ad ubera portabimini et super genua blandientur vobis
ISA|66|13|quomodo si cui mater blandiatur ita ego consolabor vos et in Hierusalem consolabimini
ISA|66|14|videbitis et gaudebit cor vestrum et ossa vestra quasi herba germinabunt et cognoscetur manus Domini servis eius et indignabitur inimicis suis
ISA|66|15|quia ecce Dominus in igne veniet et quasi turbo quadrigae eius reddere in indignatione furorem suum et increpationem suam in flamma ignis
ISA|66|16|quia in igne Dominus diiudicatur et in gladio suo ad omnem carnem et multiplicabuntur interfecti a Domino
ISA|66|17|qui sanctificabantur et mundos se putabant in hortis post unam intrinsecus qui comedebant carnem suillam et abominationem et murem simul consumentur dicit Dominus
ISA|66|18|ego autem opera eorum et cogitationes eorum venio ut congregem cum omnibus gentibus et linguis et venient et videbunt gloriam meam
ISA|66|19|et ponam in eis signum et mittam ex eis qui salvati fuerint ad gentes in mari in Africa in Lydia tenentes sagittam in Italiam et Graeciam ad insulas longe ad eos qui non audierunt de me et non viderunt gloriam meam et adnuntiabunt gloriam meam gentibus
ISA|66|20|et adducent omnes fratres vestros de cunctis gentibus donum Domino in equis et in quadrigis et in lecticis et in mulis et in carrucis ad montem sanctum meum Hierusalem dicit Dominus quomodo si inferant filii Israhel munus in vase mundo in domum Domini
ISA|66|21|et adsumam ex eis in sacerdotes et in Levitas dicit Dominus
ISA|66|22|quia sicut caeli novi et terra nova quae ego facio stare coram me dicit Dominus sic stabit semen vestrum et nomen vestrum
ISA|66|23|et erit mensis ex mense et sabbatum ex sabbato veniet omnis caro ut adoret coram facie mea dicit Dominus
ISA|66|24|et egredientur et videbunt cadavera virorum qui praevaricati sunt in me vermis eorum non morietur et ignis eorum non extinguetur et erunt usque ad satietatem visionis omni carni
