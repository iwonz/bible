MIC|1|1|The word of the LORD that came to Micah the Morasthite in the days of Jotham, Ahaz, and Hezekiah, kings of Judah, which he saw concerning Samaria and Jerusalem.
MIC|1|2|Hear, all ye people; hearken, O earth, and all that therein is: and let the Lord GOD be witness against you, the LORD from his holy temple.
MIC|1|3|For, behold, the LORD cometh forth out of his place, and will come down, and tread upon the high places of the earth.
MIC|1|4|And the mountains shall be molten under him, and the valleys shall be cleft, as wax before the fire, and as the waters that are poured down a steep place.
MIC|1|5|For the transgression of Jacob is all this, and for the sins of the house of Israel. What is the transgression of Jacob? is it not Samaria? and what are the high places of Judah? are they not Jerusalem?
MIC|1|6|Therefore I will make Samaria as an heap of the field, and as plantings of a vineyard: and I will pour down the stones thereof into the valley, and I will discover the foundations thereof.
MIC|1|7|And all the graven images thereof shall be beaten to pieces, and all the hires thereof shall be burned with the fire, and all the idols thereof will I lay desolate: for she gathered it of the hire of an harlot, and they shall return to the hire of an harlot.
MIC|1|8|Therefore I will wail and howl, I will go stripped and naked: I will make a wailing like the dragons, and mourning as the owls.
MIC|1|9|For her wound is incurable; for it is come unto Judah; he is come unto the gate of my people, even to Jerusalem.
MIC|1|10|Declare ye it not at Gath, weep ye not at all: in the house of Aphrah roll thyself in the dust.
MIC|1|11|Pass ye away, thou inhabitant of Saphir, having thy shame naked: the inhabitant of Zaanan came not forth in the mourning of Bethezel; he shall receive of you his standing.
MIC|1|12|For the inhabitant of Maroth waited carefully for good: but evil came down from the LORD unto the gate of Jerusalem.
MIC|1|13|O thou inhabitant of Lachish, bind the chariot to the swift beast: she is the beginning of the sin to the daughter of Zion: for the transgressions of Israel were found in thee.
MIC|1|14|Therefore shalt thou give presents to Moreshethgath: the houses of Achzib shall be a lie to the kings of Israel.
MIC|1|15|Yet will I bring an heir unto thee, O inhabitant of Mareshah: he shall come unto Adullam the glory of Israel.
MIC|1|16|Make thee bald, and poll thee for thy delicate children; enlarge thy baldness as the eagle; for they are gone into captivity from thee.
MIC|2|1|Woe to them that devise iniquity, and work evil upon their beds! when the morning is light, they practise it, because it is in the power of their hand.
MIC|2|2|And they covet fields, and take them by violence; and houses, and take them away: so they oppress a man and his house, even a man and his heritage.
MIC|2|3|Therefore thus saith the LORD; Behold, against this family do I devise an evil, from which ye shall not remove your necks; neither shall ye go haughtily: for this time is evil.
MIC|2|4|In that day shall one take up a parable against you, and lament with a doleful lamentation, and say, We be utterly spoiled: he hath changed the portion of my people: how hath he removed it from me! turning away he hath divided our fields.
MIC|2|5|Therefore thou shalt have none that shall cast a cord by lot in the congregation of the LORD.
MIC|2|6|Prophesy ye not, say they to them that prophesy: they shall not prophesy to them, that they shall not take shame.
MIC|2|7|O thou that art named the house of Jacob, is the spirit of the LORD straitened? are these his doings? do not my words do good to him that walketh uprightly?
MIC|2|8|Even of late my people is risen up as an enemy: ye pull off the robe with the garment from them that pass by securely as men averse from war.
MIC|2|9|The women of my people have ye cast out from their pleasant houses; from their children have ye taken away my glory for ever.
MIC|2|10|Arise ye, and depart; for this is not your rest: because it is polluted, it shall destroy you, even with a sore destruction.
MIC|2|11|If a man walking in the spirit and falsehood do lie, saying, I will prophesy unto thee of wine and of strong drink; he shall even be the prophet of this people.
MIC|2|12|I will surely assemble, O Jacob, all of thee; I will surely gather the remnant of Israel; I will put them together as the sheep of Bozrah, as the flock in the midst of their fold: they shall make great noise by reason of the multitude of men.
MIC|2|13|The breaker is come up before them: they have broken up, and have passed through the gate, and are gone out by it: and their king shall pass before them, and the LORD on the head of them.
MIC|3|1|And I said, Hear, I pray you, O heads of Jacob, and ye princes of the house of Israel; Is it not for you to know judgment?
MIC|3|2|Who hate the good, and love the evil; who pluck off their skin from off them, and their flesh from off their bones;
MIC|3|3|Who also eat the flesh of my people, and flay their skin from off them; and they break their bones, and chop them in pieces, as for the pot, and as flesh within the caldron.
MIC|3|4|Then shall they cry unto the LORD, but he will not hear them: he will even hide his face from them at that time, as they have behaved themselves ill in their doings.
MIC|3|5|Thus saith the LORD concerning the prophets that make my people err, that bite with their teeth, and cry, Peace; and he that putteth not into their mouths, they even prepare war against him.
MIC|3|6|Therefore night shall be unto you, that ye shall not have a vision; and it shall be dark unto you, that ye shall not divine; and the sun shall go down over the prophets, and the day shall be dark over them.
MIC|3|7|Then shall the seers be ashamed, and the diviners confounded: yea, they shall all cover their lips; for there is no answer of God.
MIC|3|8|But truly I am full of power by the spirit of the LORD, and of judgment, and of might, to declare unto Jacob his transgression, and to Israel his sin.
MIC|3|9|Hear this, I pray you, ye heads of the house of Jacob, and princes of the house of Israel, that abhor judgment, and pervert all equity.
MIC|3|10|They build up Zion with blood, and Jerusalem with iniquity.
MIC|3|11|The heads thereof judge for reward, and the priests thereof teach for hire, and the prophets thereof divine for money: yet will they lean upon the LORD, and say, Is not the LORD among us? none evil can come upon us.
MIC|3|12|Therefore shall Zion for your sake be plowed as a field, and Jerusalem shall become heaps, and the mountain of the house as the high places of the forest.
MIC|4|1|But in the last days it shall come to pass, that the mountain of the house of the LORD shall be established in the top of the mountains, and it shall be exalted above the hills; and people shall flow unto it.
MIC|4|2|And many nations shall come, and say, Come, and let us go up to the mountain of the LORD, and to the house of the God of Jacob; and he will teach us of his ways, and we will walk in his paths: for the law shall go forth of Zion, and the word of the LORD from Jerusalem.
MIC|4|3|And he shall judge among many people, and rebuke strong nations afar off; and they shall beat their swords into plowshares, and their spears into pruninghooks: nation shall not lift up a sword against nation, neither shall they learn war any more.
MIC|4|4|But they shall sit every man under his vine and under his fig tree; and none shall make them afraid: for the mouth of the LORD of hosts hath spoken it.
MIC|4|5|For all people will walk every one in the name of his god, and we will walk in the name of the LORD our God for ever and ever.
MIC|4|6|In that day, saith the LORD, will I assemble her that halteth, and I will gather her that is driven out, and her that I have afflicted;
MIC|4|7|And I will make her that halted a remnant, and her that was cast far off a strong nation: and the LORD shall reign over them in mount Zion from henceforth, even for ever.
MIC|4|8|And thou, O tower of the flock, the strong hold of the daughter of Zion, unto thee shall it come, even the first dominion; the kingdom shall come to the daughter of Jerusalem.
MIC|4|9|Now why dost thou cry out aloud? is there no king in thee? is thy counsellor perished? for pangs have taken thee as a woman in travail.
MIC|4|10|Be in pain, and labour to bring forth, O daughter of Zion, like a woman in travail: for now shalt thou go forth out of the city, and thou shalt dwell in the field, and thou shalt go even to Babylon; there shalt thou be delivered; there the LORD shall redeem thee from the hand of thine enemies.
MIC|4|11|Now also many nations are gathered against thee, that say, Let her be defiled, and let our eye look upon Zion.
MIC|4|12|But they know not the thoughts of the LORD, neither understand they his counsel: for he shall gather them as the sheaves into the floor.
MIC|4|13|Arise and thresh, O daughter of Zion: for I will make thine horn iron, and I will make thy hoofs brass: and thou shalt beat in pieces many people: and I will consecrate their gain unto the LORD, and their substance unto the Lord of the whole earth.
MIC|5|1|Now gather thyself in troops, O daughter of troops: he hath laid siege against us: they shall smite the judge of Israel with a rod upon the cheek.
MIC|5|2|But thou, Bethlehem Ephratah, though thou be little among the thousands of Judah, yet out of thee shall he come forth unto me that is to be ruler in Israel; whose goings forth have been from of old, from everlasting.
MIC|5|3|Therefore will he give them up, until the time that she which travaileth hath brought forth: then the remnant of his brethren shall return unto the children of Israel.
MIC|5|4|And he shall stand and feed in the strength of the LORD, in the majesty of the name of the LORD his God; and they shall abide: for now shall he be great unto the ends of the earth.
MIC|5|5|And this man shall be the peace, when the Assyrian shall come into our land: and when he shall tread in our palaces, then shall we raise against him seven shepherds, and eight principal men.
MIC|5|6|And they shall waste the land of Assyria with the sword, and the land of Nimrod in the entrances thereof: thus shall he deliver us from the Assyrian, when he cometh into our land, and when he treadeth within our borders.
MIC|5|7|And the remnant of Jacob shall be in the midst of many people as a dew from the LORD, as the showers upon the grass, that tarrieth not for man, nor waiteth for the sons of men.
MIC|5|8|And the remnant of Jacob shall be among the Gentiles in the midst of many people as a lion among the beasts of the forest, as a young lion among the flocks of sheep: who, if he go through, both treadeth down, and teareth in pieces, and none can deliver.
MIC|5|9|Thine hand shall be lifted up upon thine adversaries, and all thine enemies shall be cut off.
MIC|5|10|And it shall come to pass in that day, saith the LORD, that I will cut off thy horses out of the midst of thee, and I will destroy thy chariots:
MIC|5|11|And I will cut off the cities of thy land, and throw down all thy strong holds:
MIC|5|12|And I will cut off witchcrafts out of thine hand; and thou shalt have no more soothsayers:
MIC|5|13|Thy graven images also will I cut off, and thy standing images out of the midst of thee; and thou shalt no more worship the work of thine hands.
MIC|5|14|And I will pluck up thy groves out of the midst of thee: so will I destroy thy cities.
MIC|5|15|And I will execute vengeance in anger and fury upon the heathen, such as they have not heard.
MIC|6|1|Hear ye now what the LORD saith; Arise, contend thou before the mountains, and let the hills hear thy voice.
MIC|6|2|Hear ye, O mountains, the LORD's controversy, and ye strong foundations of the earth: for the LORD hath a controversy with his people, and he will plead with Israel.
MIC|6|3|O my people, what have I done unto thee? and wherein have I wearied thee? testify against me.
MIC|6|4|For I brought thee up out of the land of Egypt, and redeemed thee out of the house of servants; and I sent before thee Moses, Aaron, and Miriam.
MIC|6|5|O my people, remember now what Balak king of Moab consulted, and what Balaam the son of Beor answered him from Shittim unto Gilgal; that ye may know the righteousness of the LORD.
MIC|6|6|Wherewith shall I come before the LORD, and bow myself before the high God? shall I come before him with burnt offerings, with calves of a year old?
MIC|6|7|Will the LORD be pleased with thousands of rams, or with ten thousands of rivers of oil? shall I give my firstborn for my transgression, the fruit of my body for the sin of my soul?
MIC|6|8|He hath shewed thee, O man, what is good; and what doth the LORD require of thee, but to do justly, and to love mercy, and to walk humbly with thy God?
MIC|6|9|The LORD's voice crieth unto the city, and the man of wisdom shall see thy name: hear ye the rod, and who hath appointed it.
MIC|6|10|Are there yet the treasures of wickedness in the house of the wicked, and the scant measure that is abominable?
MIC|6|11|Shall I count them pure with the wicked balances, and with the bag of deceitful weights?
MIC|6|12|For the rich men thereof are full of violence, and the inhabitants thereof have spoken lies, and their tongue is deceitful in their mouth.
MIC|6|13|Therefore also will I make thee sick in smiting thee, in making thee desolate because of thy sins.
MIC|6|14|Thou shalt eat, but not be satisfied; and thy casting down shall be in the midst of thee; and thou shalt take hold, but shalt not deliver; and that which thou deliverest will I give up to the sword.
MIC|6|15|Thou shalt sow, but thou shalt not reap; thou shalt tread the olives, but thou shalt not anoint thee with oil; and sweet wine, but shalt not drink wine.
MIC|6|16|For the statutes of Omri are kept, and all the works of the house of Ahab, and ye walk in their counsels; that I should make thee a desolation, and the inhabitants thereof an hissing: therefore ye shall bear the reproach of my people.
MIC|7|1|Woe is me! for I am as when they have gathered the summer fruits, as the grapegleanings of the vintage: there is no cluster to eat: my soul desired the firstripe fruit.
MIC|7|2|The good man is perished out of the earth: and there is none upright among men: they all lie in wait for blood; they hunt every man his brother with a net.
MIC|7|3|That they may do evil with both hands earnestly, the prince asketh, and the judge asketh for a reward; and the great man, he uttereth his mischievous desire: so they wrap it up.
MIC|7|4|The best of them is as a brier: the most upright is sharper than a thorn hedge: the day of thy watchmen and thy visitation cometh; now shall be their perplexity.
MIC|7|5|Trust ye not in a friend, put ye not confidence in a guide: keep the doors of thy mouth from her that lieth in thy bosom.
MIC|7|6|For the son dishonoureth the father, the daughter riseth up against her mother, the daughter in law against her mother in law; a man's enemies are the men of his own house.
MIC|7|7|Therefore I will look unto the LORD; I will wait for the God of my salvation: my God will hear me.
MIC|7|8|Rejoice not against me, O mine enemy: when I fall, I shall arise; when I sit in darkness, the LORD shall be a light unto me.
MIC|7|9|I will bear the indignation of the LORD, because I have sinned against him, until he plead my cause, and execute judgment for me: he will bring me forth to the light, and I shall behold his righteousness.
MIC|7|10|Then she that is mine enemy shall see it, and shame shall cover her which said unto me, Where is the LORD thy God? mine eyes shall behold her: now shall she be trodden down as the mire of the streets.
MIC|7|11|In the day that thy walls are to be built, in that day shall the decree be far removed.
MIC|7|12|In that day also he shall come even to thee from Assyria, and from the fortified cities, and from the fortress even to the river, and from sea to sea, and from mountain to mountain.
MIC|7|13|Notwithstanding the land shall be desolate because of them that dwell therein, for the fruit of their doings.
MIC|7|14|Feed thy people with thy rod, the flock of thine heritage, which dwell solitarily in the wood, in the midst of Carmel: let them feed in Bashan and Gilead, as in the days of old.
MIC|7|15|According to the days of thy coming out of the land of Egypt will I shew unto him marvellous things.
MIC|7|16|The nations shall see and be confounded at all their might: they shall lay their hand upon their mouth, their ears shall be deaf.
MIC|7|17|They shall lick the dust like a serpent, they shall move out of their holes like worms of the earth: they shall be afraid of the LORD our God, and shall fear because of thee.
MIC|7|18|Who is a God like unto thee, that pardoneth iniquity, and passeth by the transgression of the remnant of his heritage? he retaineth not his anger for ever, because he delighteth in mercy.
MIC|7|19|He will turn again, he will have compassion upon us; he will subdue our iniquities; and thou wilt cast all their sins into the depths of the sea.
MIC|7|20|Thou wilt perform the truth to Jacob, and the mercy to Abraham, which thou hast sworn unto our fathers from the days of old.
