GAL|1|1|Paul, an apostle- not from men nor through man, but through Jesus Christ and God the Father, who raised him from the dead-
GAL|1|2|and all the brothers who are with me, To the churches of Galatia:
GAL|1|3|Grace to you and peace from God our Father and the Lord Jesus Christ,
GAL|1|4|who gave himself for our sins to deliver us from the present evil age, according to the will of our God and Father,
GAL|1|5|to whom be the glory forever and ever. Amen.
GAL|1|6|I am astonished that you are so quickly deserting him who called you in the grace of Christ and are turning to a different gospel-
GAL|1|7|not that there is another one, but there are some who trouble you and want to distort the gospel of Christ.
GAL|1|8|But even if we or an angel from heaven should preach to you a gospel contrary to the one we preached to you, let him be accursed.
GAL|1|9|As we have said before, so now I say again: If anyone is preaching to you a gospel contrary to the one you received, let him be accursed.
GAL|1|10|For am I now seeking the approval of man, or of God? Or am I trying to please man? If I were still trying to please man, I would not be a servant of Christ.
GAL|1|11|For I would have you know, brothers, that the gospel that was preached by me is not man's gospel.
GAL|1|12|For I did not receive it from any man, nor was I taught it, but I received it through a revelation of Jesus Christ.
GAL|1|13|For you have heard of my former life in Judaism, how I persecuted the church of God violently and tried to destroy it.
GAL|1|14|And I was advancing in Judaism beyond many of my own age among my people, so extremely zealous was I for the traditions of my fathers.
GAL|1|15|But when he who had set me apart before I was born, and who called me by his grace,
GAL|1|16|was pleased to reveal his Son to me, in order that I might preach him among the Gentiles, I did not immediately consult with anyone;
GAL|1|17|nor did I go up to Jerusalem to those who were apostles before me, but I went away into Arabia, and returned again to Damascus.
GAL|1|18|Then after three years I went up to Jerusalem to visit Cephas and remained with him fifteen days.
GAL|1|19|But I saw none of the other apostles except James the Lord's brother.
GAL|1|20|(In what I am writing to you, before God, I do not lie!)
GAL|1|21|Then I went into the regions of Syria and Cilicia.
GAL|1|22|And I was still unknown in person to the churches of Judea that are in Christ.
GAL|1|23|They only were hearing it said, "He who used to persecute us is now preaching the faith he once tried to destroy."
GAL|1|24|And they glorified God because of me.
GAL|2|1|Then after fourteen years I went up again to Jerusalem with Barnabas, taking Titus along with me.
GAL|2|2|I went up because of a revelation and set before them (though privately before those who seemed influential) the gospel that I proclaim among the Gentiles, in order to make sure I was not running or had not run in vain.
GAL|2|3|But even Titus, who was with me, was not forced to be circumcised, though he was a Greek.
GAL|2|4|Yet because of false brothers secretly brought in- who slipped in to spy out our freedom that we have in Christ Jesus, so that they might bring us into slavery-
GAL|2|5|to them we did not yield in submission even for a moment, so that the truth of the gospel might be preserved for you.
GAL|2|6|And from those who seemed to be influential (what they were makes no difference to me; God shows no partiality)- those, I say, who seemed influential added nothing to me.
GAL|2|7|On the contrary, when they saw that I had been entrusted with the gospel to the uncircumcised, just as Peter had been entrusted with the gospel to the circumcised
GAL|2|8|(for he who worked through Peter for his apostolic ministry to the circumcised worked also through me for mine to the Gentiles),
GAL|2|9|and when James and Cephas and John, who seemed to be pillars, perceived the grace that was given to me, they gave the right hand of fellowship to Barnabas and me, that we should go to the Gentiles and they to the circumcised.
GAL|2|10|Only, they asked us to remember the poor, the very thing I was eager to do.
GAL|2|11|But when Cephas came to Antioch, I opposed him to his face, because he stood condemned.
GAL|2|12|For before certain men came from James, he was eating with the Gentiles; but when they came he drew back and separated himself, fearing the circumcision party.
GAL|2|13|And the rest of the Jews acted hypocritically along with him, so that even Barnabas was led astray by their hypocrisy.
GAL|2|14|But when I saw that their conduct was not in step with the truth of the gospel, I said to Cephas before them all, "If you, though a Jew, live like a Gentile and not like a Jew, how can you force the Gentiles to live like Jews?"
GAL|2|15|We ourselves are Jews by birth and not Gentile sinners;
GAL|2|16|yet we know that a person is not justified by works of the law but through faith in Jesus Christ, so we also have believed in Christ Jesus, in order to be justified by faith in Christ and not by works of the law, because by works of the law no one will be justified.
GAL|2|17|But if, in our endeavor to be justified in Christ, we too were found to be sinners, is Christ then a servant of sin? Certainly not!
GAL|2|18|For if I rebuild what I tore down, I prove myself to be a transgressor.
GAL|2|19|For through the law I died to the law, so that I might live to God. I have been crucified with Christ.
GAL|2|20|It is no longer I who live, but Christ who lives in me. And the life I now live in the flesh I live by faith in the Son of God, who loved me and gave himself for me.
GAL|2|21|I do not nullify the grace of God, for if justification were through the law, then Christ died for no purpose.
GAL|3|1|O foolish Galatians! Who has bewitched you? It was before your eyes that Jesus Christ was publicly portrayed as crucified.
GAL|3|2|Let me ask you only this: Did you receive the Spirit by works of the law or by hearing with faith?
GAL|3|3|Are you so foolish? Having begun by the Spirit, are you now being perfected by the flesh?
GAL|3|4|Did you suffer so many things in vain- if indeed it was in vain?
GAL|3|5|Does he who supplies the Spirit to you and works miracles among you do so by works of the law, or by hearing with faith-
GAL|3|6|just as Abraham "believed God, and it was counted to him as righteousness"?
GAL|3|7|Know then that it is those of faith who are the sons of Abraham.
GAL|3|8|And the Scripture, foreseeing that God would justify the Gentiles by faith, preached the gospel beforehand to Abraham, saying, "In you shall all the nations be blessed."
GAL|3|9|So then, those who are of faith are blessed along with Abraham, the man of faith.
GAL|3|10|For all who rely on works of the law are under a curse; for it is written, "Cursed be everyone who does not abide by all things written in the Book of the Law, and do them."
GAL|3|11|Now it is evident that no one is justified before God by the law, for "The righteous shall live by faith."
GAL|3|12|But the law is not of faith, rather "The one who does them shall live by them."
GAL|3|13|Christ redeemed us from the curse of the law by becoming a curse for us- for it is written, "Cursed is everyone who is hanged on a tree"-
GAL|3|14|so that in Christ Jesus the blessing of Abraham might come to the Gentiles, so that we might receive the promised Spirit through faith.
GAL|3|15|To give a human example, brothers: even with a man-made covenant, no one annuls it or adds to it once it has been ratified.
GAL|3|16|Now the promises were made to Abraham and to his offspring. It does not say, "And to offsprings," referring to many, but referring to one, "And to your offspring," who is Christ.
GAL|3|17|This is what I mean: the law, which came 430 years afterward, does not annul a covenant previously ratified by God, so as to make the promise void.
GAL|3|18|For if the inheritance comes by the law, it no longer comes by promise; but God gave it to Abraham by a promise.
GAL|3|19|Why then the law? It was added because of transgressions, until the offspring should come to whom the promise had been made, and it was put in place through angels by an intermediary.
GAL|3|20|Now an intermediary implies more than one, but God is one.
GAL|3|21|Is the law then contrary to the promises of God? Certainly not! For if a law had been given that could give life, then righteousness would indeed be by the law.
GAL|3|22|But the Scripture imprisoned everything under sin, so that the promise by faith in Jesus Christ might be given to those who believe.
GAL|3|23|Now before faith came, we were held captive under the law, imprisoned until the coming faith would be revealed.
GAL|3|24|So then, the law was our guardian until Christ came, in order that we might be justified by faith.
GAL|3|25|But now that faith has come, we are no longer under a guardian,
GAL|3|26|for in Christ Jesus you are all sons of God, through faith.
GAL|3|27|For as many of you as were baptized into Christ have put on Christ.
GAL|3|28|There is neither Jew nor Greek, there is neither slave nor free, there is neither male nor female, for you are all one in Christ Jesus.
GAL|3|29|And if you are Christ's, then you are Abraham's offspring, heirs according to promise.
GAL|4|1|I mean that the heir, as long as he is a child, is no different from a slave, though he is the owner of everything,
GAL|4|2|but he is under guardians and managers until the date set by his father.
GAL|4|3|In the same way we also, when we were children, were enslaved to the elementary principles of the world.
GAL|4|4|But when the fullness of time had come, God sent forth his Son, born of woman, born under the law,
GAL|4|5|to redeem those who were under the law, so that we might receive adoption as sons.
GAL|4|6|And because you are sons, God has sent the Spirit of his Son into our hearts, crying, "Abba! Father!"
GAL|4|7|So you are no longer a slave, but a son, and if a son, then an heir through God.
GAL|4|8|Formerly, when you did not know God, you were enslaved to those that by nature are not gods.
GAL|4|9|But now that you have come to know God, or rather to be known by God, how can you turn back again to the weak and worthless elementary principles of the world, whose slaves you want to be once more?
GAL|4|10|You observe days and months and seasons and years!
GAL|4|11|I am afraid I may have labored over you in vain.
GAL|4|12|Brothers, I entreat you, become as I am, for I also have become as you are. You did me no wrong.
GAL|4|13|You know it was because of a bodily ailment that I preached the gospel to you at first,
GAL|4|14|and though my condition was a trial to you, you did not scorn or despise me, but received me as an angel of God, as Christ Jesus.
GAL|4|15|What then has become of the blessing you felt? For I testify to you that, if possible, you would have gouged out your eyes and given them to me.
GAL|4|16|Have I then become your enemy by telling you the truth?
GAL|4|17|They make much of you, but for no good purpose. They want to shut you out, that you may make much of them.
GAL|4|18|It is always good to be made much of for a good purpose, and not only when I am present with you,
GAL|4|19|my little children, for whom I am again in the anguish of childbirth until Christ is formed in you!
GAL|4|20|I wish I could be present with you now and change my tone, for I am perplexed about you.
GAL|4|21|Tell me, you who desire to be under the law, do you not listen to the law?
GAL|4|22|For it is written that Abraham had two sons, one by a slave woman and one by a free woman.
GAL|4|23|But the son of the slave was born according to the flesh, while the son of the free woman was born through promise.
GAL|4|24|Now this may be interpreted allegorically: these women are two covenants. One is from Mount Sinai, bearing children for slavery; she is Hagar.
GAL|4|25|Now Hagar is Mount Sinai in Arabia; she corresponds to the present Jerusalem, for she is in slavery with her children.
GAL|4|26|But the Jerusalem above is free, and she is our mother.
GAL|4|27|For it is written, "Rejoice, O barren one who does not bear; break forth and cry aloud, you who are not in labor! For the children of the desolate one will be more than those of the one who has a husband."
GAL|4|28|Now you, brothers, like Isaac, are children of promise.
GAL|4|29|But just as at that time he who was born according to the flesh persecuted him who was born according to the Spirit, so also it is now.
GAL|4|30|But what does the Scripture say? "Cast out the slave woman and her son, for the son of the slave woman shall not inherit with the son of the free woman."
GAL|4|31|So, brothers, we are not children of the slave but of the free woman.
GAL|5|1|For freedom Christ has set us free; stand firm therefore, and do not submit again to a yoke of slavery.
GAL|5|2|Look: I, Paul, say to you that if you accept circumcision, Christ will be of no advantage to you.
GAL|5|3|I testify again to every man who accepts circumcision that he is obligated to keep the whole law.
GAL|5|4|You are severed from Christ, you who would be justified by the law; you have fallen away from grace.
GAL|5|5|For through the Spirit, by faith, we ourselves eagerly wait for the hope of righteousness.
GAL|5|6|For in Christ Jesus neither circumcision nor uncircumcision counts for anything, but only faith working through love.
GAL|5|7|You were running well. Who hindered you from obeying the truth?
GAL|5|8|This persuasion is not from him who calls you.
GAL|5|9|A little leaven leavens the whole lump.
GAL|5|10|I have confidence in the Lord that you will take no other view than mine, and the one who is troubling you will bear the penalty, whoever he is.
GAL|5|11|But if I, brothers, still preach circumcision, why am I still being persecuted? In that case the offense of the cross has been removed.
GAL|5|12|I wish those who unsettle you would emasculate themselves!
GAL|5|13|For you were called to freedom, brothers. Only do not use your freedom as an opportunity for the flesh, but through love serve one another.
GAL|5|14|For the whole law is fulfilled in one word: "You shall love your neighbor as yourself."
GAL|5|15|But if you bite and devour one another, watch out that you are not consumed by one another.
GAL|5|16|But I say, walk by the Spirit, and you will not gratify the desires of the flesh.
GAL|5|17|For the desires of the flesh are against the Spirit, and the desires of the Spirit are against the flesh, for these are opposed to each other, to keep you from doing the things you want to do.
GAL|5|18|But if you are led by the Spirit, you are not under the law.
GAL|5|19|Now the works of the flesh are evident: sexual immorality, impurity, sensuality,
GAL|5|20|idolatry, sorcery, enmity, strife, jealousy, fits of anger, rivalries, dissensions, divisions,
GAL|5|21|envy, drunkenness, orgies, and things like these. I warn you, as I warned you before, that those who do such things will not inherit the kingdom of God.
GAL|5|22|But the fruit of the Spirit is love, joy, peace, patience, kindness, goodness, faithfulness,
GAL|5|23|gentleness, self-control; against such things there is no law.
GAL|5|24|And those who belong to Christ Jesus have crucified the flesh with its passions and desires.
GAL|5|25|If we live by the Spirit, let us also walk by the Spirit.
GAL|5|26|Let us not become conceited, provoking one another, envying one another.
GAL|6|1|Brothers, if anyone is caught in any transgression, you who are spiritual should restore him in a spirit of gentleness. Keep watch on yourself, lest you too be tempted.
GAL|6|2|Bear one another's burdens, and so fulfill the law of Christ.
GAL|6|3|For if anyone thinks he is something, when he is nothing, he deceives himself.
GAL|6|4|But let each one test his own work, and then his reason to boast will be in himself alone and not in his neighbor.
GAL|6|5|For each will have to bear his own load.
GAL|6|6|One who is taught the word must share all good things with the one who teaches.
GAL|6|7|Do not be deceived: God is not mocked, for whatever one sows, that will he also reap.
GAL|6|8|For the one who sows to his own flesh will from the flesh reap corruption, but the one who sows to the Spirit will from the Spirit reap eternal life.
GAL|6|9|And let us not grow weary of doing good, for in due season we will reap, if we do not give up.
GAL|6|10|So then, as we have opportunity, let us do good to everyone, and especially to those who are of the household of faith.
GAL|6|11|See with what large letters I am writing to you with my own hand.
GAL|6|12|It is those who want to make a good showing in the flesh who would force you to be circumcised, and only in order that they may not be persecuted for the cross of Christ.
GAL|6|13|For even those who are circumcised do not themselves keep the law, but they desire to have you circumcised that they may boast in your flesh.
GAL|6|14|But far be it from me to boast except in the cross of our Lord Jesus Christ, by which the world has been crucified to me, and I to the world.
GAL|6|15|For neither circumcision counts for anything, nor uncircumcision, but a new creation.
GAL|6|16|And as for all who walk by this rule, peace and mercy be upon them, and upon the Israel of God.
GAL|6|17|From now on let no one cause me trouble, for I bear on my body the marks of Jesus.
GAL|6|18|The grace of our Lord Jesus Christ be with your spirit, brothers. Amen.
