JOB|1|1|烏斯 地有一個人名叫 約伯 。這人完全、正直、敬畏上帝、遠離惡事。
JOB|1|2|他生了七個兒子，三個女兒。
JOB|1|3|他的家產有七千隻羊，三千匹駱駝，五百對牛，五百匹母驢，並有許多僕婢。這人在東方人中為至大。
JOB|1|4|他的兒子按著日子各在自己家裏擺設宴席，派人去請他們的三個姊妹來，與他們一同吃喝。
JOB|1|5|宴席的日子過了， 約伯 派人去叫他們自潔。他清早起來，按著他們眾人的數目獻燔祭，因為他說：「恐怕我的兒子犯了罪，心中背棄 上帝。」 約伯 常常這樣行。
JOB|1|6|有一天，上帝的眾使者 來侍立在耶和華面前，撒但也來在其中。
JOB|1|7|耶和華對撒但說：「你從哪裏來？」撒但回答耶和華說：「我從地上走來走去，在那裏往返。」
JOB|1|8|耶和華對撒但說：「你曾用心察看我的僕人 約伯 沒有？地上再沒有人像他那樣完全、正直、敬畏上帝、遠離惡事。」
JOB|1|9|撒但回答耶和華說：「 約伯 敬畏上帝，豈是無故呢？
JOB|1|10|你豈不是四面圈上籬笆圍護他和他的家，以及他一切所有的嗎？他手所做的都蒙你賜福，他的家產也在地上增多。
JOB|1|11|但你若伸手毀他一切所有的，他必當面背棄你。」
JOB|1|12|耶和華對撒但說：「看哪，凡他所有的都在你手中；只是不可伸手加害於他。」於是撒但從耶和華面前退出去。
JOB|1|13|有一天， 約伯 的兒女正在他們長兄的家裏吃飯喝酒，
JOB|1|14|有報信的來見 約伯 ，說：「牛正耕地，母驢在旁邊吃草，
JOB|1|15|示巴 人忽然闖來，把牲畜擄去，並用刀殺了僕人；惟有我一人逃脫，來報信給你。」
JOB|1|16|他還說話的時候，又有人來說：「上帝從天上降下火來，把羊群和僕人都吞滅了；惟有我一人逃脫，來報信給你。」
JOB|1|17|他還說話的時候，又有人來說：「 迦勒底 人分成三隊忽然闖來，把駱駝擄去，並用刀殺了僕人；惟有我一人逃脫，來報信給你。」
JOB|1|18|他還說話的時候，又有人來說：「你的兒女正在他們長兄的家裏吃飯喝酒，
JOB|1|19|看哪，有狂風從曠野颳來，襲擊房屋的四角，房屋倒塌在年輕人身上，他們就都死了；惟有我一人逃脫，來報信給你。」
JOB|1|20|約伯 就起來，撕裂外袍，剃了頭，俯伏在地敬拜，
JOB|1|21|說：「我赤身出於母胎，也必赤身歸回；賞賜的是耶和華，收取的也是耶和華。耶和華的名是應當稱頌的。」
JOB|1|22|在這一切的事上， 約伯 並沒有犯罪，也不以上帝為狂妄。
JOB|2|1|又有一天，上帝的眾使者 來侍立在耶和華面前，撒但也來在其中。
JOB|2|2|耶和華問撒但說：「你從哪裏來？」撒但回答說：「我從地上走來走去，在那裏往返。」
JOB|2|3|耶和華對撒但說：「你曾用心察看我的僕人 約伯 沒有？地上再沒有人像他那樣完全、正直、敬畏上帝、遠離惡事。你雖激起我攻擊他，無故吞滅他，他仍然持守他的純正。」
JOB|2|4|撒但回答耶和華說：「人以皮代皮，情願捨去一切所有的，來保全性命。
JOB|2|5|但你若伸手傷他的骨頭和他的肉，他必當面背棄 你。」
JOB|2|6|耶和華對撒但說：「看哪，他在你手中，只要留下他的性命。」
JOB|2|7|於是撒但從耶和華面前退出去，擊打 約伯 ，使他從腳掌到頭頂長毒瘡。
JOB|2|8|約伯 就坐在灰燼中，拿瓦片刮身體。
JOB|2|9|他的妻子對他說：「你仍然持守你的純正嗎？你背棄上帝，死了吧！」
JOB|2|10|約伯 卻對她說：「你說話，正如愚頑的婦人。唉！難道我們從上帝手裏得福，不也受禍嗎？」在這一切的事上， 約伯 並沒有以口犯罪。
JOB|2|11|約伯 的三個朋友， 提幔 人 以利法 、 書亞 人 比勒達 、 拿瑪 人 瑣法 ，聽說這一切的災禍臨到他身上，各人就從自己的地方相約同來，為他悲傷，安慰他。
JOB|2|12|他們遠遠地舉目觀看，認不出他來，就放聲大哭。各人撕裂外袍，向空中撒塵土，落在自己的頭上。
JOB|2|13|他們同他七天七夜坐在地上，一句話也不對他說，因為他們見到了極大的痛苦。
JOB|3|1|此後， 約伯 開口詛咒自己的生日 。
JOB|3|2|約伯 說：
JOB|3|3|「願我生的那日滅沒， 說『懷了男胎』的那夜也滅沒。
JOB|3|4|願那日變為黑暗， 願上帝不從上面尋找它， 願亮光不照於其上。
JOB|3|5|願黑暗和死蔭索取那日， 願密雲停在其上， 願白天的昏暗 恐嚇它。
JOB|3|6|願那夜被幽暗奪取， 不在一年的日子中喜樂， 也不列入月中的數目。
JOB|3|7|看哪，願那夜沒有生育， 其間也沒有歡樂的聲音。
JOB|3|8|願那些詛咒日子且能惹動 力威亞探 的， 詛咒那夜。
JOB|3|9|願那夜黎明的星宿變為黑暗， 盼亮卻不亮， 也不見晨曦破曉 ；
JOB|3|10|因它沒有把懷我胎的門關閉， 也沒有從我的眼中隱藏患難。
JOB|3|11|「我為何不出母胎而死？ 為何不出母腹就氣絕呢？
JOB|3|12|為何有膝蓋接收我？ 為何有奶哺養我呢？
JOB|3|13|不然，我現在已躺臥安睡， 而且，早已長眠安息；
JOB|3|14|與那些為自己重建荒涼之處， 地上的君王和謀士在一起；
JOB|3|15|或與把銀子裝滿房屋， 擁有金子的王子在一起；
JOB|3|16|我為何不像流產的胎兒被埋藏， 如同未見光的嬰孩？
JOB|3|17|在那裏惡人止息攪擾， 在那裏困乏人得享安息，
JOB|3|18|被囚的人同得安逸， 不再聽見監工的聲音。
JOB|3|19|大的小的都在那裏， 奴僕脫離主人得自由。
JOB|3|20|「遭受患難的人為何有光賜給他呢？ 心中愁苦的人為何有生命賜給他呢？
JOB|3|21|他們等死，卻不得死； 求死，勝於求隱藏的珍寶。
JOB|3|22|他們尋見墳墓， 就歡喜快樂，極其高興。
JOB|3|23|這人的道路遮隱， 上帝又四面圍困他。
JOB|3|24|我吃飯前就發出嘆息， 我的唉哼湧出如水。
JOB|3|25|因我所恐懼的臨到我， 我所懼怕的迎向我；
JOB|3|26|我不得安逸，不得平靜， 也不得安息，卻有患難來到。」
JOB|4|1|提幔 人 以利法 回答說：
JOB|4|2|「人想與你說話，你就厭煩嗎？ 但誰能忍住不發言呢？
JOB|4|3|看哪，你素來教導許多人， 又堅固軟弱的手。
JOB|4|4|你的言語曾扶助跌倒的人； 你使軟弱的膝蓋穩固。
JOB|4|5|但現在禍患臨到 你，你就煩躁了； 它挨近你，你就驚惶。
JOB|4|6|你的倚靠不是在於你敬畏上帝嗎？ 你的盼望不是在於你行事純正嗎？
JOB|4|7|「請你追想：無辜的人有誰滅亡？ 正直的人何處被剪除？
JOB|4|8|按我所見，耕罪孽的， 種毒害的，照樣收割。
JOB|4|9|上帝一噓氣，他們就滅亡； 上帝一發怒，他們就消失。
JOB|4|10|獅子吼叫，猛獅咆哮， 少壯獅子的牙齒被敲斷。
JOB|4|11|公獅因缺獵物而死， 母獅的幼獅都離散。
JOB|4|12|「有話暗中傳遞給我， 耳朵聽其微小的聲音。
JOB|4|13|世人沉睡的時候， 從夜間異象的雜念中，
JOB|4|14|恐懼戰兢臨到我身， 使我百骨戰抖。
JOB|4|15|有靈從我面前經過， 我身上的毫毛豎立。
JOB|4|16|那靈停住， 我卻不能辨其形狀； 有形像在我眼前。 我在靜默中聽見有聲音：
JOB|4|17|『必死的人能比上帝公義嗎？ 壯士能比造他的主純潔嗎？
JOB|4|18|看哪，主不信靠他的僕人， 尚且指他的使者為愚昧，
JOB|4|19|何況那些住在泥屋、 根基在塵土裏、 被蛀蟲所毀壞的人呢？
JOB|4|20|早晚之間，他們就被毀滅， 永歸無有，無人理會。
JOB|4|21|他們帳棚的繩索豈不從中拔出來呢？ 他們死，且是無智慧而死。』」
JOB|5|1|「你呼求吧，有誰回答你呢？ 聖者之中，你轉向哪一位呢？
JOB|5|2|憤怒害死愚妄人， 嫉妒殺死愚蠢的人。
JOB|5|3|我曾見愚妄人扎下根， 但我忽然詛咒他的住處。
JOB|5|4|他的兒女遠離穩妥之地， 在城門口被欺壓，無人搭救。
JOB|5|5|他的莊稼被飢餓的人吃盡了， 就是在荊棘裏的也搶去了； 他的財寶被陷阱 張口吞沒了。
JOB|5|6|因為禍患不是從塵土中出來， 患難也不是從土地裏長出。
JOB|5|7|人生出來必遭遇患難， 如同火花 飛騰。
JOB|5|8|「至於我，我必尋求上帝， 把我的事情交託給他。
JOB|5|9|他行大事不可測度， 行奇事不可勝數。
JOB|5|10|他降雨在地面， 賜水於田野。
JOB|5|11|他將卑微的人安置在高處， 將哀痛的人舉到穩妥之地。
JOB|5|12|他破壞通達人的計謀， 使他們手所做的不得成就。
JOB|5|13|他使有智慧的人中了自己的詭計， 叫狡詐人的計謀速速落空。
JOB|5|14|他們白晝遇見黑暗， 午間摸索如在夜間。
JOB|5|15|上帝拯救貧窮人脫離殘暴人的手， 脫離他們口中的刀。
JOB|5|16|這樣，貧寒人有指望， 不義的人閉口無言。
JOB|5|17|「看哪，上帝所懲治的人是有福的！ 所以你不可輕看全能者的管教。
JOB|5|18|因為他打傷，又包紮； 他擊傷，又親手醫治。
JOB|5|19|你六次遭難，他必救你； 就是七次，災禍也無法害你。
JOB|5|20|在饑荒中，他必救你脫離死亡； 在戰爭中，他必救你脫離刀劍的權勢。
JOB|5|21|你必被隱藏，不受口舌之害； 災害臨到，你也不懼怕。
JOB|5|22|對於災害饑饉，你必譏笑； 至於地上的野獸，你也不懼怕。
JOB|5|23|因為你必與田間的石頭立約， 田裏的野獸也必與你和好。
JOB|5|24|你必知道你的帳棚平安， 你查看你的羊圈，一無所失。
JOB|5|25|你也必知道你的後裔眾多， 你的子孫像地上的青草。
JOB|5|26|你必壽高年邁才歸墳墓， 好像禾捆按時收藏。
JOB|5|27|看哪，這道理我們已經考察，本是如此。 你須要聽，要親自明白。」
JOB|6|1|約伯 回答說：
JOB|6|2|「惟願我的煩惱被秤一秤， 我一切的災害放在天平裏，
JOB|6|3|現今都比海沙更重， 所以我說話急躁。
JOB|6|4|因全能者的箭射中了我， 我的靈喝盡其毒； 上帝的驚嚇擺陣攻擊我。
JOB|6|5|野驢有草豈會叫喚？ 牛有飼料豈會吼叫？
JOB|6|6|食物淡而無鹽豈可吃呢？ 蛋白有甚麼滋味呢？
JOB|6|7|那些可厭的食物， 我心不肯挨近。
JOB|6|8|「惟願我得著所求的， 上帝賞賜我所切望的，
JOB|6|9|願上帝把我壓碎， 伸手將我剪除。
JOB|6|10|我因沒有違棄那聖者的言語， 就仍以此為安慰， 在不止息的痛苦中還可歡躍。
JOB|6|11|我有甚麼氣力使我等候？ 我有甚麼結局使我忍耐？
JOB|6|12|我的氣力豈是石頭的氣力？ 我的肉身豈是銅呢？
JOB|6|13|在我裏面豈不是無助嗎？ 智慧豈不是從我心中被趕逐嗎？
JOB|6|14|「灰心的人，他的朋友當以慈愛待他， 因為他將離棄敬畏全能者的心。
JOB|6|15|我的弟兄詭詐，好像河道， 像溪水流過的河床，
JOB|6|16|因結冰而混濁， 有雪藏在其中，
JOB|6|17|暖和的時候就溶化， 炎熱時便從原處乾涸。
JOB|6|18|商隊偏離道路， 上到荒涼之地而死亡。
JOB|6|19|提瑪 的商隊瞻望， 示巴 的旅客等候。
JOB|6|20|他們因希望落空就抱愧， 來到那裏便蒙羞。
JOB|6|21|現在你們正是這樣 ， 看見驚嚇的事就懼怕。
JOB|6|22|我豈說：『請你們供給我， 從你們的財物中送禮給我』？
JOB|6|23|或說：『請你們拯救我脫離敵人的手， 救贖我脫離殘暴人的手』嗎？
JOB|6|24|「請你們指教我，我就不作聲； 我在何事上有錯，請使我明白。
JOB|6|25|正直言語的力量何其大！ 但你們責備是責備甚麼呢？
JOB|6|26|絕望人的講論既然如風， 你們還計劃批駁言語嗎？
JOB|6|27|你們甚至為孤兒抽籤， 把朋友當貨物。
JOB|6|28|「現在，請你們看著我， 我絕不當面說謊。
JOB|6|29|請你們轉意，不要不公義； 請再轉意，正義在我這裏。
JOB|6|30|我的舌頭豈有不公義嗎？ 我的上膛豈不辨奸惡嗎？」
JOB|7|1|「人在世上豈無勞役呢？ 他的日子不像雇工的日子嗎？
JOB|7|2|像奴僕切慕陰涼， 像雇工等待工錢，
JOB|7|3|我也照樣度過虛空的歲月， 愁煩的夜晚指定給我。
JOB|7|4|我躺臥的時候就說： 『我何時可以起來呢？』漫漫長夜， 我總是翻來覆去，直到天亮。
JOB|7|5|我的肉體以蟲子和塵土為衣， 我的皮膚才收了口又流膿。
JOB|7|6|我的日子比織布的梭更快， 都消耗在沒有指望之中。
JOB|7|7|「你要記得，我的生命不過是一口氣， 我的眼睛必不再看見福樂。
JOB|7|8|觀看我的人，他的眼必不看見我； 你的眼目投向我，我卻不在了。
JOB|7|9|雲彩消散而去； 照樣，人下陰間也不再上來。
JOB|7|10|他不再回自己的家， 他自己的地方也不再認得他。
JOB|7|11|「我甚至不封我的口； 我靈愁苦，要發出言語； 我心苦惱，要吐露哀情。
JOB|7|12|我豈是海洋，豈是大魚， 你竟防守著我呢？
JOB|7|13|我若說：『我的床必安慰我， 我的榻必分擔我的苦情』，
JOB|7|14|你就用夢驚擾我， 用異象恐嚇我。
JOB|7|15|甚至我寧可窒息死亡， 勝似留我這副骨頭。
JOB|7|16|我厭棄生命，不願永遠活著。 你任憑我吧，因我的日子都是虛空。
JOB|7|17|人算甚麼，你竟看他為大， 將他放在心上，
JOB|7|18|每早晨鑒察他， 每時刻考驗他？
JOB|7|19|你到何時才轉眼不看我， 任憑我咽下唾沫呢？
JOB|7|20|鑒察人的主啊，我若有罪，於你何妨？ 為何以我當你的箭靶， 使我成為你的重擔呢？
JOB|7|21|為何不赦免我的過犯， 除掉我的罪孽呢？ 我現今要躺臥在塵土中； 你要切切尋找我，我卻不在了。」
JOB|8|1|書亞 人 比勒達 回答說：
JOB|8|2|「這些話你要說到幾時？ 你口中的言語如狂風要到幾時呢？
JOB|8|3|上帝豈能偏離公平？ 全能者豈能偏離公義？
JOB|8|4|或者你的兒女得罪了他， 他就把他們交在過犯的掌控中。
JOB|8|5|你若切切尋求上帝， 向全能者懇求；
JOB|8|6|你若純潔正直， 他必定為你興起， 使你公義的居所興旺。
JOB|8|7|你起初雖然微小， 日後必非常強盛。
JOB|8|8|「請你詢問上代， 思念他們祖先所查究的。
JOB|8|9|我們不過從昨日才有，一無所知， 因我們在世的日子好像影子。
JOB|8|10|他們豈不指教你，告訴你， 說出發自內心的言語呢？
JOB|8|11|「蒲草沒有泥豈能生長？ 蘆荻沒有水豈能長大？
JOB|8|12|它還青翠，沒有割下的時候， 比百樣的草先枯槁。
JOB|8|13|凡忘記上帝的人，路途也是這樣； 不虔敬人的指望要滅沒。
JOB|8|14|他所仰賴的必折斷， 他所倚靠的是蜘蛛網。
JOB|8|15|他要倚靠房屋，房屋卻站立不住； 他要抓住房屋，房屋卻不能存留。
JOB|8|16|他在日光之下茂盛， 嫩枝在園中蔓延；
JOB|8|17|他的根盤繞石堆， 鑽入石縫 。
JOB|8|18|他若從本地被拔出， 那地就不認識他，說：『我沒有見過你。』
JOB|8|19|看哪，這就是他道路中的喜樂， 以後必另有人從塵土而生。
JOB|8|20|看哪，上帝必不丟棄完全人， 也不扶助邪惡人的手。
JOB|8|21|他還要以喜笑充滿你的口， 以歡呼充滿你的嘴唇。
JOB|8|22|恨惡你的要披戴羞愧， 惡人的帳棚必歸於無有。」
JOB|9|1|約伯 回答說：
JOB|9|2|「我真的知道是這樣， 但人在上帝前怎能成為義呢？
JOB|9|3|人若想要與他爭辯， 千次中也不能回答一次。
JOB|9|4|他心裏有智慧，且大有能力。 誰向上帝剛硬而得平安呢？
JOB|9|5|他把山挪移，山卻不知， 他在怒氣中，把山翻倒。
JOB|9|6|他使地震動，離其本位， 地的柱子就搖撼。
JOB|9|7|他吩咐太陽，太陽就不出來， 又封住眾星。
JOB|9|8|他獨自鋪張諸天， 步行在海浪之上。
JOB|9|9|他造北斗、參星、昴星， 以及南方的星宿 ；
JOB|9|10|他行大事不可測度， 行奇事不可勝數。
JOB|9|11|看哪，他從我旁邊經過，我看不見； 他走過，我沒有察覺他。
JOB|9|12|看哪，他奪去，誰能阻擋他？ 誰敢對他說：『你做甚麼呢？』
JOB|9|13|「上帝必不收回他的怒氣， 扶助 拉哈伯 的，屈身在上帝以下。
JOB|9|14|既是這樣，我怎敢回答他， 怎敢在他之前選擇辯詞呢？
JOB|9|15|我雖有義，也不能回答， 我要向那審判我的懇求。
JOB|9|16|我若呼求，縱然他應允我， 我仍不信他會側耳聽我的聲音。
JOB|9|17|他用暴風 摧折我， 無故加增我的損傷。
JOB|9|18|他不容我喘一口氣， 倒使我飽受苦惱。
JOB|9|19|若論力量，看哪，他真有能力！ 若論審判，『誰能傳我呢？』
JOB|9|20|我雖有義，我的口要定我有罪； 我雖完全，他必證明我為彎曲。
JOB|9|21|我雖完全，不顧自己； 我厭棄我的性命。
JOB|9|22|所以我說，都是一樣； 完全人和惡人，他都滅絕。
JOB|9|23|若災禍忽然帶來死亡， 他必戲笑無辜人的苦難。
JOB|9|24|世界交在惡人手中； 他蒙蔽世界審判官的臉， 若不是他，那麼是誰呢？
JOB|9|25|「我的日子比奔跑者更快， 急速過去，不見福樂。
JOB|9|26|我的日子如蒲草船掠過， 如鷹俯衝抓食。
JOB|9|27|我若說：『我要忘記我的苦情， 強顏歡笑』，
JOB|9|28|我就因一切的愁苦而懼怕； 我知道你必不以我為無辜。
JOB|9|29|我必被定罪， 我何必徒然勞苦呢？
JOB|9|30|我若用雪水洗身， 用鹼潔淨我的手掌，
JOB|9|31|你還要把我扔在坑裏， 我的衣服都憎惡我。
JOB|9|32|他不像我是個人，使我可以回答他， 使我們可以一同受審判。
JOB|9|33|我們中間沒有仲裁者， 可以按手在我們兩造之間。
JOB|9|34|願他使他的杖離開我， 不使他的威嚴恐嚇我，
JOB|9|35|我就說話，不懼怕他； 但對我來說，我卻不是這樣。」
JOB|10|1|「我厭惡自己的性命， 任由我述說自己的苦情； 因心裏苦惱，我要說話。
JOB|10|2|我對上帝說，不要定我有罪， 要指示我，你為何與我爭辯？
JOB|10|3|你手所造的，你又欺壓，又藐視， 卻光照惡人的計謀。 這事你以為美嗎？
JOB|10|4|你的眼豈是肉眼？ 你察看豈像人察看嗎？
JOB|10|5|你的日子豈像人的日子， 你的年歲豈像壯士的年歲，
JOB|10|6|你就追問我的罪孽， 尋察我的罪過嗎？
JOB|10|7|其實，你知道我沒有行惡， 也無人能施行拯救，脫離你的手。
JOB|10|8|你的手塑造我，造了我， 但我整個人卻要一起被你吞滅。
JOB|10|9|求你記得，你製造我如泥土， 你還要使我歸回塵土嗎？
JOB|10|10|你不是倒出我來好像奶， 使我凝結如同奶酪嗎？
JOB|10|11|你以皮和肉給我穿上， 用骨與筋把我聯結起來。
JOB|10|12|你將生命和慈愛賜給我， 你也眷顧保全我的靈。
JOB|10|13|然而，你把這些事藏在你心裏， 我知道這是你的旨意。
JOB|10|14|我若犯罪，你就察看我， 並不赦免我的罪。
JOB|10|15|我若行惡，我就有禍了； 我若行義，也不敢抬頭， 而是飽受羞辱， 看見我的痛苦。
JOB|10|16|你如獅子昂首追捕我 ， 又在我身上顯出奇事。
JOB|10|17|你更新你的見證對付我， 向我加增惱怒， 調遣軍隊攻擊我。
JOB|10|18|「你為何使我出母胎呢？ 甚願我當時氣絕，沒有眼睛看見我。
JOB|10|19|這樣，就如從未有過我， 我一出母胎就被送入墳墓。
JOB|10|20|我的日子不是短少嗎？求你停止， 求你放過我 ，使我可以稍得喜樂，
JOB|10|21|就是在我去而不返， 往黑暗和死蔭之地以先。
JOB|10|22|那是烏黑之地， 猶如幽暗的死蔭， 毫無秩序； 發出的光輝也像幽暗。」
JOB|11|1|拿瑪 人 瑣法 回答說：
JOB|11|2|「這許多的話豈不該回答嗎？ 多嘴多舌的人豈可成為義呢？
JOB|11|3|你誇大的話豈能使人不作聲嗎？ 你戲笑的時候豈沒有人使你受辱嗎？
JOB|11|4|你說：『我的教導純全， 我在你眼前是清潔的。』
JOB|11|5|但是，惟願上帝說話， 願他張開嘴唇攻擊你。
JOB|11|6|願他將智慧的奧祕指示你， 因為健全的知識是兩面的。 你當知道，上帝使你忘記你的一些罪孽。
JOB|11|7|你能尋見上帝的奧祕嗎？ 你能尋見全能者的極限嗎？
JOB|11|8|高如諸天，你能做甚麼？ 比陰間深，你能知道甚麼？
JOB|11|9|其量度比地長， 比海更寬。
JOB|11|10|他若經過，把人拘禁， 召集會眾，誰能阻擋他呢？
JOB|11|11|因為他知道虛妄的人； 當他看見罪惡，豈不留意嗎？
JOB|11|12|空虛的人若獲得知識， 野驢生下的駒子也成了人。
JOB|11|13|「至於你，若堅固己心， 又向主舉手；
JOB|11|14|你若遠遠脫離你手中的罪孽， 不容許不義住在你帳棚之中；
JOB|11|15|這樣，你必仰起臉來，毫無瑕疵； 你也必安穩，無所懼怕。
JOB|11|16|你必忘記你的苦楚， 就是想起來，也如流過的水。
JOB|11|17|你在世要升高，比正午更明， 雖有黑暗，仍像早晨。
JOB|11|18|你因有指望就必穩固， 也必四圍察看 ，安然躺下。
JOB|11|19|你躺臥，無人驚嚇， 並有許多人向你求恩。
JOB|11|20|但惡人的眼睛要失明； 他們無路可逃， 他們的指望就是氣絕身亡。」
JOB|12|1|約伯 回答說：
JOB|12|2|「你們果真是人物啊！ 智慧要與你們一同去死。
JOB|12|3|但我也有聰明，跟你們一樣， 並非不及你們。 這些事，誰不知道呢？
JOB|12|4|我這求告上帝、蒙他應允的人 竟成了朋友所譏笑的； 又公義又完全的人竟遭受譏笑。
JOB|12|5|安逸的人心裏藐視災禍， 這災禍在等待失足滑跌的人。
JOB|12|6|強盜的帳棚安寧， 惹上帝發怒的人穩固， 他們把上帝 握在自己手中 。
JOB|12|7|「你問走獸，走獸必指教你； 你問空中的飛鳥，飛鳥必告訴你；
JOB|12|8|或者你與地說話，地必指教你 ； 海中的魚也必向你說明。
JOB|12|9|在這一切當中， 有誰不知道這是耶和華的手做成的呢？
JOB|12|10|凡動物的生命 和人類的氣息都在他手中。
JOB|12|11|耳朵豈不辨別言語， 正如上膛品嘗食物嗎？
JOB|12|12|年老的有智慧， 壽高的有知識。
JOB|12|13|「在上帝有智慧和能力， 他有謀略和知識。
JOB|12|14|看哪，他拆毀，就不能重建； 他拘禁人，人就不得釋放。
JOB|12|15|看哪，他使水止住，水就乾了； 他把水放出，水就淹沒大地。
JOB|12|16|在他有能力和智慧， 走迷的和使人迷路的都屬他。
JOB|12|17|他把謀士剝衣擄去， 使審判官變為愚妄。
JOB|12|18|他解除君王的權勢 ， 用帶子捆住他們的腰。
JOB|12|19|他把祭司剝衣擄去， 使有權能的人傾覆。
JOB|12|20|他廢去忠信者的言論， 奪去長者的見識。
JOB|12|21|他使貴族蒙羞受辱， 放鬆勇士的腰帶。
JOB|12|22|他從黑暗中彰顯深奧的事， 使死蔭顯出光明。
JOB|12|23|他使邦國興旺而又毀滅， 使邦國擴展又被掠奪。
JOB|12|24|他將地上百姓中領袖的聰明奪去， 使他們迷失在荒涼無路之地。
JOB|12|25|他們在無光的黑暗中摸索； 他使他們搖晃像醉酒的人一樣。」
JOB|13|1|「看哪，這一切，我眼都見過； 我耳都聽過，而且明白。
JOB|13|2|你們所知道的，我也知道， 並非不及你們。
JOB|13|3|然而我要對全能者說話， 我願與上帝理論。
JOB|13|4|但你們是編造謊言的， 全都是無用的醫生。
JOB|13|5|惟願你們全然不作聲， 這就是你們的智慧！
JOB|13|6|請你們聽我的答辯， 留心聽我嘴唇的訴求。
JOB|13|7|你們要為上帝說不義的話嗎？ 要為他說詭詐的言語嗎？
JOB|13|8|你們要看上帝的情面嗎？ 要為他爭辯嗎？
JOB|13|9|他查究你們，這豈是好事嗎？ 人欺騙人，你們也要照樣欺騙他嗎？
JOB|13|10|你們若暗中看人的情面， 他必定要責備你們。
JOB|13|11|他的尊榮豈不叫你們懼怕嗎？ 他豈不使驚嚇臨到你們嗎？
JOB|13|12|你們可記念的諺語是灰燼的箴言； 你們的後盾是泥土的後盾。
JOB|13|13|「你們不要向我作聲， 讓我說話，無論如何我都承當。
JOB|13|14|我為何把我的肉掛在我的牙上， 將我的命放在我的手掌中呢？
JOB|13|15|看哪，他要殺我，我毫無指望 ， 然而我還要在他面前辯明我所行的。
JOB|13|16|這要成為我的拯救， 因為不虔誠的人不可到他面前。
JOB|13|17|你們要細聽我的言語， 讓我的申辯入你們耳中。
JOB|13|18|看哪，我已陳明我的案， 知道自己有義。
JOB|13|19|還有誰要和我爭辯， 我現在就緘默不言，氣絕而死。
JOB|13|20|惟有兩件事不要向我施行， 我就不躲開你的面：
JOB|13|21|就是把你的手縮回，遠離我身； 又不使你的威嚴恐嚇我。
JOB|13|22|這樣，你呼叫，我就回答； 或是讓我說話，你回答我。
JOB|13|23|我的罪孽和我的罪有多少呢？ 求你叫我知道我的過犯與我的罪。
JOB|13|24|你為何轉臉， 拿我當仇敵呢？
JOB|13|25|你要驚動被風吹的葉子嗎？ 要追趕枯乾的碎秸嗎？
JOB|13|26|你寫下苦楚對付我， 又使我擔當幼年的罪孽。
JOB|13|27|你把我的腳鎖上木枷， 察看我一切的道路， 為我的腳掌劃定界限。
JOB|13|28|人像滅絕的爛物， 像蟲蛀的衣裳。」
JOB|14|1|「人為婦人所生， 日子短少，多有患難。
JOB|14|2|他出來如花，凋謝而去； 他飛逝如影，不能存留。
JOB|14|3|這樣的人你豈會睜眼看他， 又叫我 來，在你那裏受審嗎？
JOB|14|4|誰能使潔淨出於污穢呢？ 誰也不能！
JOB|14|5|既然人的日子限定， 他的月數在於你， 你劃定他的界限，他不能越過；
JOB|14|6|求你轉眼不看他，使他得歇息， 直到他像雇工享受他的一天。
JOB|14|7|「因樹有指望， 若被砍下，還可發芽， 嫩枝生長不息。
JOB|14|8|樹根若衰老在地裏， 樹幹也死在土中，
JOB|14|9|及至得了水氣，還會發芽， 長出枝條，像新栽的樹一樣。
JOB|14|10|但壯士一死就消逝了； 人一氣絕，他在何處呢？
JOB|14|11|海中的水枯竭， 江河消散乾涸。
JOB|14|12|人一躺下就不再起來， 等到諸天沒有了 ，仍不復醒， 也不能從睡中喚醒。
JOB|14|13|惟願你把我藏在陰間， 把我隱藏，直到你的憤怒過去； 願你為我定下期限，並記得我。
JOB|14|14|壯士若死了能再活嗎？ 我在一切服役的日子中等待， 直到我退伍的時候來到。
JOB|14|15|你呼叫，我就回答你； 你手所做的，你必期待。
JOB|14|16|但如今你數點我的腳步， 不察看我的罪。
JOB|14|17|我的過犯被你密封在囊中， 你遮掩了我的罪孽。
JOB|14|18|「然而，山崩變為無有， 磐石從原處挪移。
JOB|14|19|流水沖蝕石頭， 急流洗去地上的塵土； 你也照樣滅絕人的指望。
JOB|14|20|你終必勝過人，使他消逝； 你改變他的容貌，把他送走。
JOB|14|21|他的兒子得尊榮，他不知道； 他們降為卑，他也不曉得。
JOB|14|22|他只覺得身上疼痛， 心中為自己悲哀。」
JOB|15|1|提幔 人 以利法 回答說：
JOB|15|2|「智慧人豈可用虛空的知識回答， 用東風充滿自己的肚腹呢？
JOB|15|3|他豈可用無益的話， 用無濟於事的言語理論呢？
JOB|15|4|你誠然廢棄敬畏， 不在上帝面前默想。
JOB|15|5|你的罪孽指教你的口； 你選用詭詐人的舌頭。
JOB|15|6|你自己的口定你有罪，並非是我； 你自己的嘴唇見證你的不是。
JOB|15|7|「你是頭一個生下來的人嗎？ 你受造在諸山之先嗎？
JOB|15|8|你曾聽見上帝的密旨嗎？ 你要獨自得盡智慧嗎？
JOB|15|9|甚麼是你知道，我們不知道的呢？ 甚麼是你明白，我們不明白的呢？
JOB|15|10|我們這裏有白髮的和年老的， 比你父親還年長。
JOB|15|11|上帝的安慰和對你溫和的話， 你以為太小嗎？
JOB|15|12|你的心為何失控， 你的眼為何冒火，
JOB|15|13|以致你的靈反對上帝， 你的口說出這樣的言語呢？
JOB|15|14|人是甚麼，竟算為潔淨呢？ 婦人所生的是甚麼，竟算為義呢？
JOB|15|15|看哪，上帝不信任他的眾聖者； 在他眼前，天也不潔淨，
JOB|15|16|何況那污穢可憎， 喝罪孽如水的世人呢！
JOB|15|17|「我指示你，你要聽我； 我要陳述我所看見的，
JOB|15|18|就是智慧人從列祖所受， 傳講而不隱瞞的事。
JOB|15|19|這地惟獨賜給他們， 並沒有外人從他們中間經過。
JOB|15|20|惡人一生的日子絞痛難熬， 殘暴人存留的年數也是如此。
JOB|15|21|驚嚇的聲音常在他耳中； 在平安時，毀滅者必臨到他。
JOB|15|22|他不信自己能從黑暗中轉回； 他被刀劍看守。
JOB|15|23|他飄流在外求食：『哪裏有食物呢？』 他知道黑暗的日子在他手邊預備好了。
JOB|15|24|急難困苦叫他害怕， 而且勝過他，好像君王預備上陣。
JOB|15|25|因他伸手攻擊上帝， 逞強對抗全能者，
JOB|15|26|挺著頸項， 用盾牌堅厚的凸面向全能者直闖；
JOB|15|27|又因他的臉蒙上油脂， 腰上積滿肥肉。
JOB|15|28|他住在荒涼的城鎮， 房屋無人居住， 將成為廢墟。
JOB|15|29|他不得富足， 財物不得常存， 產業在地上也不加增。
JOB|15|30|他不得脫離黑暗， 火焰要把他的嫩枝燒乾； 因上帝口中的氣，他要離去。
JOB|15|31|不要讓他倚靠虛假，欺騙自己， 因虛假必成為他的報應。
JOB|15|32|他的日期未到之先，這事必實現； 他的枝子不得青綠。
JOB|15|33|他必像葡萄樹，葡萄未熟就掉落； 又像橄欖樹，一開花就凋謝。
JOB|15|34|因不敬虔之輩必不能生育， 受賄賂之人的帳棚必被火吞滅。
JOB|15|35|他們所懷的是毒害，所生的是罪孽， 肚腹裏所預備的是詭詐。」
JOB|16|1|約伯 回答說：
JOB|16|2|「這樣的話我聽了許多； 你們全都是使人愁煩的安慰者。
JOB|16|3|如風的言語有窮盡嗎？ 或者甚麼惹動你回答呢？
JOB|16|4|我也能說你們那樣的話， 你們若處在我的景況， 我也可以堆砌言詞攻擊你們， 又可以向你們搖頭。
JOB|16|5|但我必用口堅固你們， 顫動的嘴唇帶來舒解。
JOB|16|6|「我若說話，痛苦仍不得緩解； 我若停止，痛苦就離開我嗎？
JOB|16|7|但現在上帝使我困倦， 你使所有的親友遠離我，
JOB|16|8|你抓住我 ，成為見證起來攻擊我； 我的枯瘦也當著我的面作證。
JOB|16|9|上帝發怒撕裂我，逼迫我， 向我咬牙切齒； 我的敵人怒目瞪我。
JOB|16|10|他們向我大大張口， 打我的耳光羞辱我， 聚在一起攻擊我。
JOB|16|11|上帝把我交給不敬虔的人， 把我扔到惡人的手中。
JOB|16|12|我本是安逸，他折斷我， 掐住我的頸項，把我摔碎， 又立我作他的箭靶。
JOB|16|13|他的弓箭手圍繞我。 他刺破我的腎臟，並不留情， 把我的膽汁傾倒在地上。
JOB|16|14|他使我破裂，破裂又破裂， 如同勇士向我直闖。
JOB|16|15|「我把麻布縫在我的皮膚上， 把我的角放在塵土中。
JOB|16|16|我的臉因哭泣變紅， 我的眼皮上有死蔭。
JOB|16|17|我的手中卻沒有暴力， 我的祈禱也是純潔的。
JOB|16|18|「地啊，不要遮蓋我的血！ 不要讓我的哀求有藏匿之處！
JOB|16|19|現今，看哪，在天有我的見證， 在上有我的保人。
JOB|16|20|我的朋友譏誚我， 我卻向上帝眼淚汪汪。
JOB|16|21|願人可與上帝理論， 如同人與朋友一樣；
JOB|16|22|因為再過幾年， 我必走那往而不返之路。」
JOB|17|1|「我的靈耗盡，我的日子消逝； 墳墓為我預備好了。
JOB|17|2|戲笑的人果真陪伴著我， 我的眼睛盯住他們的悖逆。
JOB|17|3|「願你親自為我付押擔保。 誰還會與我擊掌呢？
JOB|17|4|因你蒙蔽他們的心，使不明理， 所以你必不高舉他們。
JOB|17|5|控告 朋友為了分享產業的， 他兒女的眼睛要失明。
JOB|17|6|「上帝使我成為人群中的笑談， 他們吐唾沫在我臉上。
JOB|17|7|我的眼睛因憂愁昏花， 我的肢體全像影兒。
JOB|17|8|正直人因此必驚奇； 無辜的人要興起攻擊不敬虔之輩。
JOB|17|9|然而，義人要持守所行的道， 手潔的人要力上加力。
JOB|17|10|至於你們眾人，再回來吧！ 你們中間，我找不到一個智慧人。
JOB|17|11|我的日子已經過去了， 我的謀算、我心的願望已經斷絕了。
JOB|17|12|他們以黑夜為白晝， 即使面臨黑暗，以為亮光已近。
JOB|17|13|我若盼望陰間為我的家， 若下榻在黑暗中，
JOB|17|14|若對地府呼叫：『你是我的父親』， 若對蟲呼叫：『你是我的母親、姊妹』，
JOB|17|15|這樣，我的盼望在哪裏呢？ 我所盼望的，誰能看見呢？
JOB|17|16|這盼望要下到陰間的門閂嗎 ？ 要一起在塵土中安息嗎 ？」
JOB|18|1|書亞 人 比勒達 回答說：
JOB|18|2|「你們尋索言語要到幾時呢 ？ 你們要明白，然後我們才說話。
JOB|18|3|我們為何被視為畜生， 在你們眼中看為愚笨 呢？
JOB|18|4|在怒氣中將自己撕裂的人哪， 難道大地要因你見棄、 磐石要挪開原處嗎？
JOB|18|5|「惡人的亮光必要熄滅， 他的火焰必不照耀。
JOB|18|6|他帳棚中的亮光要變黑暗， 他上面的燈也必熄滅。
JOB|18|7|他強橫的腳步必遭阻礙， 他的計謀必將自己絆倒。
JOB|18|8|他因自己的腳陷入網中， 走在纏人的網子上。
JOB|18|9|羅網必抓住他的腳跟， 陷阱必擒獲他。
JOB|18|10|繩索為他藏在土裏， 羈絆為他藏在路上。
JOB|18|11|四面的驚嚇使他害怕， 在他腳跟後面追趕他。
JOB|18|12|他的力量必因飢餓衰敗， 禍患要在他的旁邊等候，
JOB|18|13|侵蝕他肢體的皮膚； 死亡的長子吞吃他的肢體。
JOB|18|14|他要從所倚靠的帳棚被拔出來， 帶到使人驚恐的王那裏。
JOB|18|15|不屬他的必住在他的帳棚裏， 硫磺必撒在他所住之處。
JOB|18|16|下邊，他的根要枯乾； 上邊，他的枝子要剪除。
JOB|18|17|他的稱號 從地上消失， 他的名字不在街上存留。
JOB|18|18|他必從光明中被驅逐到黑暗裏， 他必被趕出世界。
JOB|18|19|他在自己百姓中必無子無孫， 在寄居之地也沒有倖存者。
JOB|18|20|以後的人 要因他的日子驚訝， 以前的人 也被驚駭抓住。
JOB|18|21|不義之人的住處總是這樣， 這就是不認識上帝之人的下場。」
JOB|19|1|約伯 回答說：
JOB|19|2|「你們攪擾我的心， 用言語壓碎我要到幾時呢？
JOB|19|3|你們這十次羞辱我， 苦待我也不以為恥。
JOB|19|4|果真我有錯， 這錯是在於我。
JOB|19|5|若你們真要向我誇大， 以我的羞辱來責備我，
JOB|19|6|就該知道是上帝傾覆我， 用羅網圍繞我。
JOB|19|7|看哪，我喊冤叫屈，卻不蒙應允； 我呼求，卻沒有公正。
JOB|19|8|上帝攔住我的道路，使我不得經過； 他使黑暗籠罩我的路徑。
JOB|19|9|他剝去我的榮光， 摘去我頭上的冠冕。
JOB|19|10|他在四圍攻擊我，我就走了； 他將我的指望如樹拔出。
JOB|19|11|他向我發烈怒， 以我為他的敵人。
JOB|19|12|他的軍隊一齊上來， 修築道路攻擊我， 在我帳棚的四圍安營。
JOB|19|13|「他把我的兄弟隔在遠處， 使我認識的人全然與我生疏。
JOB|19|14|我的親戚都離開了我； 我的密友都忘記了我。
JOB|19|15|在我家寄居的和我的使女， 都當我是陌生人； 我在他們眼中被視為外邦人。
JOB|19|16|我呼喚僕人，他卻不回答； 我必須親口求他。
JOB|19|17|我口的氣味令我妻子厭惡， 我的同胞都憎惡我。
JOB|19|18|連小男孩也藐視我； 我起來，他們都嘲笑我。
JOB|19|19|我的知心朋友都憎惡我； 我平日所愛的人向我翻臉。
JOB|19|20|我的皮和肉緊貼骨頭， 我得以逃脫，僅剩牙齒 。
JOB|19|21|我的朋友啊，可憐我！可憐我！ 因為上帝的手攻擊我。
JOB|19|22|你們為甚麼彷彿上帝逼迫我， 吃我的肉還不滿足呢？
JOB|19|23|「惟願我的言語現在就寫上， 都記錄在書上；
JOB|19|24|用鐵筆和鉛， 刻在磐石上，存到永遠。
JOB|19|25|我知道我的救贖主 活著， 末後他必站在塵土上。
JOB|19|26|我這皮肉滅絕之後 ， 我必在肉體之外 得見上帝。
JOB|19|27|我自己要見他， 親眼要看他，並不像陌生人。 我的心腸在我裏面耗盡了！
JOB|19|28|你們若說：『我們怎麼逼迫他呢？ 事情的根源是在於他 』，
JOB|19|29|你們就當懼怕刀劍， 因為憤怒帶來刀劍的刑罰。 這樣，你們就知道有審判。」
JOB|20|1|拿瑪 人 瑣法 回答說：
JOB|20|2|「這樣，我的思念叫我回答， 因為我心中急躁。
JOB|20|3|我聽見那羞辱我的責備； 我悟性的靈回答我。
JOB|20|4|你豈不知道嗎？亙古以來， 自從人被安置在地，
JOB|20|5|惡人歡樂的聲音是暫時的， 不敬虔人的喜樂不過是轉眼之間。
JOB|20|6|他的尊榮雖達到天上， 頭雖頂到雲中，
JOB|20|7|他必永遠滅亡，像自己的糞一樣。 看見他的人要說：『他在哪裏呢？』
JOB|20|8|他必如夢飛去，不再尋見； 他被趕走，如夜間的異象。
JOB|20|9|親眼見過他的，必不再見他； 他自己的地方也不再見到他。
JOB|20|10|他的兒女要向窮人求恩； 他的手要賠還錢財。
JOB|20|11|他的骨頭雖然滿有年輕的活力， 卻要和他一同躺臥在塵土之中。
JOB|20|12|「他口中以惡為甘甜， 把惡藏在舌頭底下，
JOB|20|13|愛戀不捨， 含在口中。
JOB|20|14|他的食物在肚裏卻要翻轉， 在他裏面成為虺蛇的毒液。
JOB|20|15|他吞了財寶，還要吐出； 上帝要從他腹中掏出來。
JOB|20|16|他必吸飲虺蛇的毒汁， 毒蛇的舌頭必殺他。
JOB|20|17|他不再看見溪流， 流奶與蜜之河。
JOB|20|18|他勞碌得來的要賠還，不得吞下； 賺取了財貨，也不得歡樂。
JOB|20|19|他欺壓窮人，棄之不顧， 強取非自己所蓋的房屋 。
JOB|20|20|「他的肚腹不知安逸， 所貪戀的連一樣也不放過，
JOB|20|21|剩餘的沒有一樣他不吞吃， 所以他的福樂不能長久。
JOB|20|22|他在滿足有餘的時候，必有困苦臨到； 凡受苦楚之人的手必加在他身上。
JOB|20|23|他的肚腹正要滿足的時候， 上帝必將猛烈的憤怒降在他身上； 他正在吃飯的時候， 上帝要將這憤怒如雨降在他身上。
JOB|20|24|他要躲避鐵的武器， 銅弓要將他射透。
JOB|20|25|箭一抽，就從他背上出來， 發亮的箭頭從他膽中出來； 有驚惶臨到他身上。
JOB|20|26|他的財寶隱藏在深沉的黑暗裏； 有非人吹起的火要把他吞滅， 把他帳棚中所剩下的燒燬。
JOB|20|27|天要顯明他的罪孽， 地要興起去攻擊他。
JOB|20|28|他家裏出產的必消失， 在上帝憤怒的日子被沖走。
JOB|20|29|這是惡人從上帝所得的份， 是上帝為他所定的產業。」
JOB|21|1|約伯 回答說：
JOB|21|2|「你們要細心聽我的言語， 這就算是你們的安慰。
JOB|21|3|請寬容我，我又要說話； 說了以後，任憑你嗤笑吧！
JOB|21|4|我豈是向人訴苦？ 我為何不是沒有耐心呢？
JOB|21|5|你們要轉向我而驚奇， 要用手摀口。
JOB|21|6|我每逢思想，心就驚惶， 戰兢抓住我身。
JOB|21|7|惡人為何存活， 得享高壽，勢力強盛呢？
JOB|21|8|他們的後裔與他們一起 ，堅立在他們面前， 他們得以眼見自己的子孫。
JOB|21|9|他們的家宅平安無懼， 上帝的杖不加在他們身上。
JOB|21|10|他們的公牛傳種而不斷絕， 母牛生牛犢而不掉胎。
JOB|21|11|他們打發小男孩出去，多如羊群， 他們的孩子踴躍跳舞。
JOB|21|12|他們隨著琴鼓歌唱， 因簫聲歡喜。
JOB|21|13|他們度日諸事亨通， 在平安中下到陰間。
JOB|21|14|他們對上帝說：『離開我們吧！ 我們不想知道你的道路。
JOB|21|15|全能者是誰，我們何必事奉他呢？ 求告他有甚麼益處呢？』
JOB|21|16|看哪，他們亨通不是靠自己的手； 惡人的計謀離我好遠。
JOB|21|17|「惡人的燈何嘗熄滅？ 患難何嘗臨到他們呢？ 上帝何嘗發怒，把災禍分給他們呢？
JOB|21|18|他們何嘗像風前的碎秸， 如暴風颳去的糠秕呢？
JOB|21|19|上帝為惡人的兒女積蓄罪孽， 不如本人遭報，好使他親自知道。
JOB|21|20|願他親眼看見自己敗亡， 親自飲全能者的憤怒。
JOB|21|21|他的歲月既盡， 他身後還顧他的家嗎？
JOB|21|22|誰能將知識教導上帝呢？ 是他審判那些居高位的。
JOB|21|23|有人至死身體強壯， 盡得平順安逸；
JOB|21|24|他的肚腹充滿奶汁 ， 他的骨髓滋潤。
JOB|21|25|有人至死心中痛苦， 從未嘗過福樂的滋味；
JOB|21|26|他們同樣躺臥於塵土， 蟲子覆蓋他們。
JOB|21|27|「看哪，我知道你們的意念， 並殘害我的計謀。
JOB|21|28|你們說：『權貴的房屋在哪裏？ 惡人住過的帳棚在哪裏？』
JOB|21|29|你們沒有詢問那些過路的人嗎？ 你們不承認他們的證據嗎？
JOB|21|30|就是惡人在患難的日子得存留， 在憤怒的日子得逃脫。
JOB|21|31|他所行的，有誰當面給他說明？ 他所做的，有誰報應他呢？
JOB|21|32|然而他要被抬到墳地， 並有人看守墓穴。
JOB|21|33|他要以谷中的土塊為甘甜； 人人要跟在他後面， 在他前面去的無數。
JOB|21|34|你們怎能以空話安慰我呢？ 你們的對答全都錯謬！」
JOB|22|1|提幔 人 以利法 回答說：
JOB|22|2|「人能使上帝有益嗎？ 智慧人能使他有益嗎？
JOB|22|3|你為人公義，豈能叫全能者喜悅呢？ 你行為完全，豈能使他得利呢？
JOB|22|4|他豈是因你敬畏的心就責備你， 審判你嗎？
JOB|22|5|你的罪惡豈不是大嗎？ 你的罪孽不是沒有窮盡嗎？
JOB|22|6|因你無故強取弟兄的抵押， 剝去赤身者的衣服。
JOB|22|7|疲乏的人，你沒有給他水喝； 飢餓的人，你沒有給他食物。
JOB|22|8|有能力的人得土地； 尊貴的人住在其中。
JOB|22|9|你打發寡婦空手回去， 你折斷孤兒的膀臂。
JOB|22|10|因此，有羅網環繞你， 有恐懼忽然使你驚惶；
JOB|22|11|或有黑暗使你看不見 ， 有洪水淹沒你。
JOB|22|12|「上帝豈不是在高天嗎？ 你看星宿的頂點何其高呢！
JOB|22|13|你說：『上帝知道甚麼？ 他豈能透過幽暗施行審判呢？
JOB|22|14|密雲將他遮蓋，使他不能看見； 他周遊穹蒼。』
JOB|22|15|你要依從上古的道嗎？ 這道是惡人行過的。
JOB|22|16|他們未到時候就被抓去 ； 他們的根基被江河沖去。
JOB|22|17|他們向上帝說：『離開我們吧！』 全能者能把他們怎麼樣呢？
JOB|22|18|然而，是上帝以美物充滿他們的房屋； 惡人的計謀離我好遠！
JOB|22|19|義人看見他們的結局 就歡喜； 無辜的人嗤笑他們：
JOB|22|20|『攻擊我們的果然被剪除， 剩餘的都被火吞滅。』
JOB|22|21|「你要與上帝和好，要和平， 這樣，福氣必臨到你。
JOB|22|22|你當領受他口中的教導， 將他的言語存在心裏。
JOB|22|23|你若歸向全能者，就必得建立。 你要從你帳棚中遠離不義，
JOB|22|24|你要將黃金丟到塵土裏， 將 俄斐 的金子丟在溪河石頭之間；
JOB|22|25|全能者就必作你的黃金， 作你成堆的銀子。
JOB|22|26|那時，你要以全能者為喜樂， 向上帝仰臉。
JOB|22|27|你要向他禱告，他就聽你； 你也要還你的願。
JOB|22|28|你定意要做何事，必然為你成就； 亮光也必照耀你的路。
JOB|22|29|當人降卑，你說：是因驕傲； 眼目謙卑的人，上帝必然拯救。
JOB|22|30|不是無辜的人，上帝尚且要搭救他 ； 他必因你手中的清潔得蒙拯救。」
JOB|23|1|約伯 回答說：
JOB|23|2|「如今我的哀告還算為悖逆； 我雖唉哼，他的手仍然重重責罰我 。
JOB|23|3|惟願我知道哪裏可以尋見上帝， 能到他的臺前，
JOB|23|4|我就在他面前陳明我的案件， 滿口辯訴。
JOB|23|5|我必知道他回答我的言語， 明白他向我所要說的。
JOB|23|6|他豈用大能與我爭辯呢？ 不！他必理會我。
JOB|23|7|在那裏正直人可以與他辯論， 我就必永遠脫離那審判我的。
JOB|23|8|「看哪，我往前走，他不在那裏； 往後退，也沒有察覺他。
JOB|23|9|他在左邊行事，我卻看不見他； 他轉向右邊 ，我也見不到他。
JOB|23|10|然而他知道我所走的路； 他試煉我，我就如純金。
JOB|23|11|我的腳緊跟他的步伐； 我謹守他的道，並不偏離。
JOB|23|12|他嘴唇的命令，我未曾背棄； 我看重他口中的言語，過於我需用的飲食 。
JOB|23|13|只是他心志已定，誰能使他轉意呢？ 他心裏所願的，就行出來。
JOB|23|14|因此，為我所定的，他必做成， 這類的事他還有許多。
JOB|23|15|所以我在他面前驚惶； 我思想就懼怕他。
JOB|23|16|上帝使我喪膽， 全能者使我驚惶。
JOB|23|17|但我並非被黑暗剪除， 只是幽暗遮蓋了我的臉。
JOB|24|1|「為何全能者不定下期限？ 為何認識他的人看不到那些日子呢？
JOB|24|2|有人挪移地界， 搶奪群畜去放牧。
JOB|24|3|他們拉走孤兒的驢， 強取寡婦的牛作抵押。
JOB|24|4|他們使貧窮人離開正道； 世上的困苦人盡都隱藏。
JOB|24|5|看哪，他們如同野驢出到曠野，殷勤尋找食物， 在野地給孩童餬口。
JOB|24|6|他們收割別人田間的莊稼， 摘取惡人剩餘的葡萄。
JOB|24|7|他們終夜赤身無衣， 在寒冷中毫無遮蓋。
JOB|24|8|他們在山上被大雨淋濕， 因沒有避身之處就擁抱磐石。
JOB|24|9|又有人從母懷中搶走孤兒， 在困苦人身上強取抵押品 。
JOB|24|10|困苦人赤身無衣，到處流浪， 餓著肚子扛抬禾捆，
JOB|24|11|他們在圍牆內榨油， 踹壓酒池，自己卻口渴。
JOB|24|12|在城內垂死的人呻吟， 受傷的人哀號； 上帝卻不理會狂妄的事。
JOB|24|13|「又有人背棄光明， 不認識光明的道， 不留在光明的路上。
JOB|24|14|殺人者黎明起來， 殺害困苦人和貧窮人， 夜間又作盜賊。
JOB|24|15|姦夫的眼等候黃昏， 說：『沒有眼睛能見我』， 就把臉蒙住。
JOB|24|16|盜賊黑夜挖洞； 他們白日躲藏， 並不認識光明。
JOB|24|17|他們全都看早晨如死蔭， 因為他們熟悉死蔭的驚駭。
JOB|24|18|「惡人在水面上快速飄盪， 他們在地上所得的產業被詛咒； 無人再回到他們的葡萄園。
JOB|24|19|乾旱炎熱融化雪水； 陰間也如此吞沒犯罪的人。
JOB|24|20|懷他的母胎忘記他； 蟲子要吃他，覺得甘甜； 他不再被人記念； 不義的人必如樹折斷。
JOB|24|21|「他與不懷孕不生育的婦人交往 ， 卻不善待寡婦。
JOB|24|22|然而上帝用能力保全有勢力的人； 那性命難保的人仍然興起。
JOB|24|23|上帝使他安穩，他就有所倚靠； 上帝的眼目看顧他們的道路。
JOB|24|24|他們高升，不過片刻就沒有了； 他們降為卑，被除滅，與眾人一樣 ， 又如穀的穗子被割下。
JOB|24|25|若不是這樣，誰能指證我是說謊的， 以我的言語為毫無根據呢？」
JOB|25|1|書亞 人 比勒達 回答說：
JOB|25|2|「上帝有統治之權，威嚴可畏； 他在高處施行和平。
JOB|25|3|他的軍隊豈能數算？ 他的光向誰不會升起呢 ？
JOB|25|4|這樣，在上帝面前人怎能稱義？ 婦人所生的怎能潔淨？
JOB|25|5|看哪，在上帝眼前，月亮無光， 星宿也不皎潔，
JOB|25|6|更何況是如蟲的人， 如蛆的世人呢！
JOB|26|1|約伯 回答說：
JOB|26|2|「無能的人蒙你何等的幫助！ 膀臂無力的人蒙你何等的拯救！
JOB|26|3|無智慧的人蒙你何等的指教！ 你向他顯出豐富的知識。
JOB|26|4|你向誰發出言語？ 誰的靈從你而出？
JOB|26|5|在大水和水族以下， 陰魂戰兢。
JOB|26|6|在上帝面前，陰間顯露； 冥府 也不得遮掩。
JOB|26|7|上帝將北極鋪在空中， 將大地懸在虛空。
JOB|26|8|他將水包在密雲中， 盛水的雲卻不破裂。
JOB|26|9|他遮蔽寶座的正面， 把他的雲彩鋪在其上。
JOB|26|10|他在水面上劃一圓圈， 直到光明與黑暗的交界。
JOB|26|11|天的柱子震動， 因他的斥責驚奇。
JOB|26|12|他以能力攪動 大海 ， 藉知識打傷 拉哈伯 。
JOB|26|13|他藉自己的靈使天空晴朗； 他的手刺殺爬得快的蛇。
JOB|26|14|看哪，這不過是上帝工作的些微； 我們聽見他的話，是何等細微的聲音！ 他大能的雷聲誰能明白呢？」
JOB|27|1|約伯 繼續發表他的言論說：
JOB|27|2|「我指著奪去我公道的永生上帝， 並使我心中愁苦的全能者起誓：
JOB|27|3|只要我的生命尚在我裏面， 上帝所賜的氣息仍在我鼻孔內，
JOB|27|4|我的唇絕不說不義， 我的舌也不說詭詐。
JOB|27|5|我斷不以你們為義； 我至死不放棄自己的純正！
JOB|27|6|我持定我的義，並不放鬆； 在世的日子，我的心不責備我。
JOB|27|7|「願我的仇敵如惡人一樣； 願那起來攻擊我的，如不義之人一般。
JOB|27|8|不敬虔的人有甚麼指望呢？ 上帝要剪除他，取他的性命。
JOB|27|9|患難臨到他， 上帝豈聽他的呼求？
JOB|27|10|他豈以全能者為樂， 隨時求告上帝呢？
JOB|27|11|上帝手所做的，我要指教你們； 全能者所行的，我也不會隱瞞。
JOB|27|12|看哪，你們自己也都見過， 為何全變為這樣虛妄呢？
JOB|27|13|「這是上帝為惡人所定的份， 殘暴人從全能者所得的產業：
JOB|27|14|倘若他的兒女增多，仍被刀所殺； 他的子孫必不得飽食。
JOB|27|15|他遺留的人必死而埋葬， 他的寡婦也不哀哭。
JOB|27|16|他雖積蓄銀子如塵沙， 堆積衣服如泥土，
JOB|27|17|他儘管堆積，義人卻要穿上， 無辜的人卻要分取銀子。
JOB|27|18|他建造房屋如蟲做窩， 又如守望者所搭的棚。
JOB|27|19|他雖富足躺臥，卻不得收殮 ， 他張開眼睛，就不在了。
JOB|27|20|驚恐如洪水將他追上， 暴風在夜間將他颳去。
JOB|27|21|東風把他吹去，他就走了； 風將他颳離原地。
JOB|27|22|風 無情地擊打他， 他試圖逃脫風的手。
JOB|27|23|風要因他拍掌， 並要發叱聲，使他離開原地。」
JOB|28|1|「銀子有礦； 煉金有場。
JOB|28|2|鐵從土裏開採， 銅從礦石鎔出。
JOB|28|3|人探索黑暗的盡頭， 查究礦石直到極處， 那是幽暗和死蔭；
JOB|28|4|他在無人居住之處開鑿礦穴， 在無足跡之地被遺忘 ， 與人遠離，懸空搖擺。
JOB|28|5|地出產糧食， 地底翻騰如火。
JOB|28|6|地的石頭是藍寶石之處， 那裏還有金沙。
JOB|28|7|鷙鳥不知那條路， 鷹眼也未曾見過。
JOB|28|8|狂傲的野獸未曾踩踏， 猛烈的獅子也未曾經過。
JOB|28|9|「人動手鑿開堅石， 翻倒山的根基，
JOB|28|10|在磐石中鑿出水道， 親眼看見各樣寶物。
JOB|28|11|他封閉河川不得涓滴 ， 使隱藏之物顯露出來。
JOB|28|12|「然而，智慧何處可尋？ 聰明之地在哪裏？
JOB|28|13|智慧的價值 無人能知， 活人之地也無處可尋。
JOB|28|14|深淵說：『不在我裏面。』 滄海說：『不在我這裏。』
JOB|28|15|智慧不可用黃金換取， 也不能用白銀秤她的價值。
JOB|28|16|俄斐 的金子和貴重的紅瑪瑙， 以及藍寶石，不足與她比擬；
JOB|28|17|黃金和玻璃不足與她比較； 純金的器皿不足兌換她。
JOB|28|18|珊瑚、水晶都不值得提； 智慧的價值勝過寶石 。
JOB|28|19|古實 的紅璧璽不足與她比較； 純金也不足與她比擬。
JOB|28|20|「智慧從何處來呢？ 聰明之地在哪裏？
JOB|28|21|她隱藏，遠離眾生的眼目， 她掩蔽，遠離空中的飛鳥。
JOB|28|22|毀滅和死亡說： 『我們風聞其名。』
JOB|28|23|「上帝明白智慧的道路， 知道智慧的所在。
JOB|28|24|因為他鑒察直到地極， 遍觀普天之下，
JOB|28|25|要為風定輕重， 又度量諸水，
JOB|28|26|為雨定律例， 為雷電定道路。
JOB|28|27|那時他看見智慧，就談論她， 堅定她，並且查究她。
JOB|28|28|他對人說：『看哪，敬畏主就是智慧； 遠離惡事就是聰明。』」
JOB|29|1|約伯 繼續發表他的言論說：
JOB|29|2|「惟願我如從前的歲月， 如上帝保護我的日子。
JOB|29|3|那時他的燈照在我頭上， 我藉他的光行過黑暗。
JOB|29|4|在我壯年的時候， 上帝親密的情誼臨到我的帳棚中。
JOB|29|5|全能者仍與我同在， 我的兒女都環繞我。
JOB|29|6|我的腳洗在乳酪當中； 磐石為我流出油河。
JOB|29|7|我出到城門， 在廣場安排座位，
JOB|29|8|年輕人見我而迴避， 老年人起身站立。
JOB|29|9|王子都停止說話， 用手摀口；
JOB|29|10|領袖靜默無聲， 舌頭貼住上膛。
JOB|29|11|耳朵聽見了，稱我有福； 眼睛看見了，就稱讚我。
JOB|29|12|因我拯救了哀求的困苦人 和無人幫助的孤兒。
JOB|29|13|將要滅亡的為我祝福， 我使寡婦心中歡呼。
JOB|29|14|我穿上公義，它遮蔽我； 我的公平如外袍和冠冕。
JOB|29|15|我作瞎子的眼， 瘸子的腳。
JOB|29|16|我作貧窮人的父； 我不認識之人的案件，我也去查明。
JOB|29|17|我打破不義之人的大牙， 從他牙齒中奪走他所搶的。
JOB|29|18|我說：『我要增添我的日子如塵沙， 我必死在自己家中 。
JOB|29|19|我的根伸展到水邊， 露水夜宿我的枝上。
JOB|29|20|我的榮耀在我身上更新， 我的弓在我手中日新。』
JOB|29|21|「人聽我說話而等候， 為我的教導而靜默。
JOB|29|22|我說話之後，他們就不再說； 我的言語滴在他們身上。
JOB|29|23|他們等候我如等雨水， 又張口如切慕春雨。
JOB|29|24|我向他們微笑，他們不敢相信； 他們不使我臉上的光失色。
JOB|29|25|我為他們選擇道路，又坐首位； 我如君王在軍隊中居住， 又如人安慰哀傷的人。」
JOB|30|1|「但如今，比我年輕的人譏笑我； 我曾藐視他們的父親， 不放在我的牧羊犬中。
JOB|30|2|他們的精力既已衰敗， 手中的氣力於我何益？
JOB|30|3|他們因窮乏飢餓，沒有生氣， 在荒廢淒涼的幽暗中啃乾燥之地。
JOB|30|4|他們在草叢之中採鹹草， 羅騰 樹的根成為他們的食物。
JOB|30|5|他們從人群中被趕出， 人追喊他們如賊一般，
JOB|30|6|以致他們住在荒谷， 住在地洞和巖穴中。
JOB|30|7|他們在草叢中叫喚， 在荊棘下擠成一團。
JOB|30|8|這都是愚頑卑微人的兒女； 他們被鞭打，趕出境外。
JOB|30|9|「現在這些人以我為歌曲， 以我為笑談。
JOB|30|10|他們厭惡我，躲避我， 不住地吐唾沫在我臉上。
JOB|30|11|上帝鬆開我的弓弦 使我受苦， 他們就在我面前脫去轡頭。
JOB|30|12|這夥人在我右邊起來， 他們推開我的腳， 築災難之路攻擊我。
JOB|30|13|他們毀壞我的道， 加增我的災害； 他們毋須人幫助。
JOB|30|14|他們來，如同闖進大缺口， 在暴風間滾動。
JOB|30|15|驚恐傾倒在我身上， 我的尊榮被逐如風； 我的福祿如雲飄去。
JOB|30|16|「現在我的心極其悲傷， 困苦的日子將我抓住。
JOB|30|17|夜間，我裏面的骨頭刺痛， 啃著我的沒有止息。
JOB|30|18|我的外衣因大力扭皺 ， 內衣的領子把我勒住。
JOB|30|19|上帝把我扔在淤泥之中， 我就像塵土和灰燼一樣。
JOB|30|20|我呼求你，你不應允我； 我站起來，你只是望著我。
JOB|30|21|你對我變得殘忍， 大能的手追逼我。
JOB|30|22|你把我提到風中，使我乘風而去， 使我消失在烈風之中。
JOB|30|23|我知道你要使我歸於死亡， 到那為眾生所定的陰宅。
JOB|30|24|「然而，人在廢墟豈不伸手？ 遇災難時一定呼救。
JOB|30|25|人遭難的日子，我豈不為他哭泣呢？ 人貧窮的時候，我豈不為他憂愁呢？
JOB|30|26|我仰望福氣，災禍就來到； 我等待光明，黑暗便來臨。
JOB|30|27|我內心煩擾不安， 困苦的日子臨到我身。
JOB|30|28|我在陰暗中行走，沒有日光 ， 我在會眾中站立求救。
JOB|30|29|我與野狗為弟兄， 我跟鴕鳥為同伴。
JOB|30|30|我的皮膚變黑脫落， 我的骨頭因熱燒焦。
JOB|30|31|我的琴音變為哀泣； 我的簫聲變為哭聲。」
JOB|31|1|「我與眼睛立約， 怎能凝望少女呢？
JOB|31|2|從至上的上帝所得之分， 從至高全能者所得之業是甚麼呢？
JOB|31|3|豈不是禍患臨到不義的， 災害臨到作惡的嗎？
JOB|31|4|上帝豈不察看我的道路， 數點我所有的腳步嗎？
JOB|31|5|「我若與虛謊同行， 我腳若緊跟詭詐，
JOB|31|6|願上帝用公道的天平秤我， 願他知道我的純正。
JOB|31|7|我的腳步若偏離正路， 我的心若隨從我眼目， 我的手掌若黏有污穢；
JOB|31|8|願我栽種，別人來吃， 我的農作物連根拔出。
JOB|31|9|「我心若因婦人受迷惑， 在鄰舍的門外等候，
JOB|31|10|就願我妻子給別人推磨， 別人與她同寢。
JOB|31|11|因為這是邪惡的事， 審判官裁定的罪孽。
JOB|31|12|這是一場火，直燒到毀滅 ， 必拔除我一切的家產。
JOB|31|13|「我的僕婢與我爭辯， 我若藐視不聽他們的冤情，
JOB|31|14|上帝興起的時候，我怎樣行呢？ 他察問的時候，我怎樣回答他呢？
JOB|31|15|造我在母腹中的，不也是造了他嗎？ 在母胎中使我們成形的，豈不是同一位嗎？
JOB|31|16|「我若不讓貧寒人遂其所願， 或是叫寡婦眼中失望，
JOB|31|17|或獨自吃自己的食物， 孤兒沒有吃其中些許；
JOB|31|18|從我年輕時，孤兒就與我一同長大，我好像他的父親， 我從出母腹就扶助寡婦 ；
JOB|31|19|我若見人因無衣死亡， 或見貧窮人毫無遮蓋；
JOB|31|20|我若不使他真心為我祝福， 不使他因我羊的毛得暖；
JOB|31|21|我若舉手攻擊孤兒， 因為在城門口見有幫助我的；
JOB|31|22|情願我的肩膀從肩胛骨脫落， 我的膀臂從肱骨折斷。
JOB|31|23|因上帝降的災禍使我恐懼 ， 因他的威嚴，我甚麼都不能。
JOB|31|24|「我若以黃金為我的指望， 對純金說：你是我的倚靠；
JOB|31|25|我若因財物豐裕， 因手多得資財而歡喜；
JOB|31|26|我若見太陽發光， 明月運行，
JOB|31|27|心就暗暗被引誘， 口親吻自己的手；
JOB|31|28|這也是審判官裁定的罪孽， 因為我背棄了至上的上帝。
JOB|31|29|「我若見恨我的遇難就歡喜， 見他遭災就高興；
JOB|31|30|其實我沒有容許口犯罪， 以詛咒要他的性命；
JOB|31|31|若我帳棚中的人未曾說： 『誰不以他的肉食吃飽呢？』
JOB|31|32|我未曾讓旅客在街上過夜， 卻開門迎接行路的人；
JOB|31|33|我若像 亞當 遮掩自己的過犯， 將罪孽藏在懷中；
JOB|31|34|我若因大大懼怕眾人， 又因宗族的藐視而恐懼， 以致我緘默不言，閉門不出；
JOB|31|35|惟願有一位肯聽我！ 看哪，我的記號，願全能者回答我！ 願那與我爭訟的寫下狀詞！
JOB|31|36|我必把它帶在肩上， 綁在頭上為冠冕。
JOB|31|37|我必向上帝述說我腳步的數目， 如同王子進到他面前。
JOB|31|38|「若我的田地喊冤告我， 犁溝也一同哭泣；
JOB|31|39|我若吃地的出產不給銀錢， 或叫地的原主喪命；
JOB|31|40|願蒺藜生長代替麥子， 惡臭的草代替大麥。」 約伯 的話說完了。
JOB|32|1|於是這三個人因 約伯 看自己為義就停止，不再回答他。
JOB|32|2|那時 布西 人， 蘭 族 巴拉迦 的兒子 以利戶 發怒了。他向 約伯 發怒，因 約伯 自以為義，不以上帝為義。
JOB|32|3|他又向 約伯 的三個朋友發怒，因為他們想不出回答的話來，仍以 約伯 為有罪。
JOB|32|4|以利戶 因為他們比自己年老，就等候要與 約伯 說話。
JOB|32|5|以利戶 見這三個人口中無話回答，就發怒。
JOB|32|6|布西 人 巴拉迦 的兒子 以利戶 回答說： 「我年輕，你們年長， 因此我退讓，不敢向你們陳述我的意見。
JOB|32|7|我說：『年長的當先說話； 壽高的當以智慧教導人。』
JOB|32|8|其實，是人裏面的靈， 全能者的氣使人有聰明。
JOB|32|9|壽高的不都有智慧， 年老的不都明白公平。
JOB|32|10|因此我說：『你們要聽我， 我也要陳述我的意見。』
JOB|32|11|「看哪，我等候你們的話， 側耳聽你們的高見； 直到你們找到要說的言語。
JOB|32|12|我留心聽你們， 看哪，你們中間無一人能折服 約伯 ， 回答他的話。
JOB|32|13|你們切不可說：『我們尋得智慧； 上帝能勝他 ，人卻不能。』
JOB|32|14|約伯 沒有用言語與我爭辯； 我也不用你們的話回答他。
JOB|32|15|「他們驚惶不再回答， 一言不發。
JOB|32|16|我豈因他們不說話， 因他們站住不再回答，仍舊等候呢？
JOB|32|17|我也要以我的一番話回答， 我也要陳述我的意見。
JOB|32|18|因為我滿懷言語， 我裏面的靈激動我。
JOB|32|19|看哪，我的肚腹如酒囊沒有氣孔， 又如新皮袋 快要破裂。
JOB|32|20|我要說話，使我舒暢； 我要張開嘴唇回答。
JOB|32|21|我必不看人的情面， 也不奉承人。
JOB|32|22|我不懂得奉承； 不然，造我的主必快快除滅我。」
JOB|33|1|「但是， 約伯 啊，請聽我的言語， 側耳聽我一切的話。
JOB|33|2|看哪，我開口， 我的舌在上膛發言。
JOB|33|3|我的言語要表明心中的正直， 我嘴唇所知道的就誠實地說。
JOB|33|4|上帝的靈造了我， 全能者的氣使我得生。
JOB|33|5|你若能夠，就請回答我； 請你站起來，在我面前陳明。
JOB|33|6|看哪，我在上帝面前與你一樣， 也是用泥土造成的。
JOB|33|7|看哪，我不用威嚴恐嚇你， 也不用勢力重壓你。
JOB|33|8|「其實，你向我耳朵說話， 我聽見你言語的聲音：
JOB|33|9|『我是純潔無過的， 我是無辜的，在我裏面沒有罪孽。
JOB|33|10|看哪，上帝找機會攻擊我， 以我為他的仇敵，
JOB|33|11|把我的腳鎖上木枷， 察看我一切的道路。』
JOB|33|12|「看哪，你這話無理，我要回答你， 因上帝比世人更大。
JOB|33|13|你為何與他爭論： 『他任何事都不向人解答』？
JOB|33|14|上帝說一次、兩次， 人卻不理會。
JOB|33|15|世人在床上沉睡安眠時， 在夢中和夜間的異象裏，
JOB|33|16|上帝就開通世人的耳朵， 把警告印在他們心上 ，
JOB|33|17|好叫人轉離自己的行為， 叫壯士遠離驕傲，
JOB|33|18|攔阻人不陷入地府， 不讓他命喪刀下 。
JOB|33|19|「人在床上被疼痛懲治， 骨頭不住地掙扎，
JOB|33|20|以致生命厭棄食物， 心中厭惡美味。
JOB|33|21|他的肉消瘦，難以看見； 先前看不見的骨頭都凸出來。
JOB|33|22|他的性命臨近地府， 他的生命挨近滅命者。
JOB|33|23|一千天使中， 若有一個作傳話的臨到他， 指示人所當行的事，
JOB|33|24|上帝就施恩給他，說： 『要救贖他 免得下入地府， 我已經得了贖價。
JOB|33|25|他的肉要比孩童的肉更嫩； 他就返老還童。』
JOB|33|26|他向上帝禱告，上帝就悅納他； 他必歡呼朝見上帝的面， 因上帝恢復他的義。
JOB|33|27|他在人前歌唱說： 『我犯了罪，顛倒是非， 卻沒有受該得的報應。
JOB|33|28|上帝救贖我的性命免入地府， 我的生命也必見光。』
JOB|33|29|「看哪，上帝兩次、三次 向人行這一切的事，
JOB|33|30|為要從地府救回人的性命， 使他被生命之光照耀。
JOB|33|31|約伯 啊，你當留心聽我； 不要作聲，我要說話。
JOB|33|32|你若有話說，可以回答我； 你只管說，因我願以你為義。
JOB|33|33|若不然，你當聽我； 不要作聲，我要把智慧教導你。」
JOB|34|1|以利戶 繼續說：
JOB|34|2|「你們智慧人要聽我的言語， 有知識的人要側耳聽我。
JOB|34|3|因為耳朵辨別言語， 好像上膛品嘗食物。
JOB|34|4|我們當選擇公理， 彼此知道何為善。
JOB|34|5|約伯 曾說：『我是公義的， 上帝奪去我的公理。
JOB|34|6|我有理，豈能說謊呢？ 我無過，受的箭傷卻不能醫治。』
JOB|34|7|哪一個人像 約伯 ， 喝譏誚如同喝水呢？
JOB|34|8|他與作惡的結伴， 和惡人同行。
JOB|34|9|他說：『人以上帝為樂， 總是無益。』
JOB|34|10|「所以，你們明理的人要聽我， 上帝斷不致行惡， 全能者斷不致不義。
JOB|34|11|他必按人所做的報應人， 使各人照所行的得報。
JOB|34|12|確實地，上帝必不作惡， 全能者必不偏離公平。
JOB|34|13|誰派他治理大地？ 誰安定全世界呢？
JOB|34|14|他若專心為己， 將靈和氣收歸自己，
JOB|34|15|凡血肉之軀必一同死亡； 世人必歸於塵土。
JOB|34|16|「你若明理，當聽這話， 側耳聽我言語的聲音。
JOB|34|17|難道恨惡公平的可以掌權嗎？ 那有公義、有大能的，你豈可定他有罪呢？
JOB|34|18|你會對君王說：『你是卑鄙的』； 對貴族說：『你們是邪惡的』嗎？
JOB|34|19|他待王子不徇情面， 也不看重富足的過於貧寒的， 因為他們都是他手所造的。
JOB|34|20|一瞬間他們就死亡。 百姓在半夜中被震動而去世； 有權力的被奪去，非藉人手。
JOB|34|21|「上帝的眼目觀看人的道路， 察看他每一腳步。
JOB|34|22|沒有黑暗，沒有死蔭， 能給作惡者在那裏藏身。
JOB|34|23|上帝不必再三傳人 到他面前受審判。
JOB|34|24|他毋須調查就粉碎有大能的人， 指定別人代替他們。
JOB|34|25|所以他知道他們的行為， 使他們在夜間傾倒壓碎。
JOB|34|26|他在眾目睽睽下擊打他們， 如同擊打惡人。
JOB|34|27|因為他們轉離不跟從他， 不留心他一切的道，
JOB|34|28|甚至使貧寒人的哀聲達到他那裏； 他也聽了困苦人的哀聲。
JOB|34|29|他安靜，誰能定罪呢？ 他轉臉，誰能見他呢？ 無論一國或一人都是如此。
JOB|34|30|不虔敬的人不得作王， 免得百姓陷入圈套。
JOB|34|31|「有誰對上帝說： 『我受了責罰，必不再犯罪；
JOB|34|32|我所看不明的，求你指教我； 我若行了不義，必不再行』？
JOB|34|33|他因你拒絕不接受， 就隨你的心願施行報應嗎？ 選擇的是你，不是我。 你所知道的，只管說吧！
JOB|34|34|明理的人必對我說， 聽我的智慧人也說：
JOB|34|35|『 約伯 說話沒有知識， 他的言語毫無智慧。』
JOB|34|36|願 約伯 被考驗到底， 因他回答像惡人一樣。
JOB|34|37|他在罪上又加悖逆； 在我們中間引起疑惑 ， 用許多言語輕慢上帝。」
JOB|35|1|以利戶 繼續說：
JOB|35|2|「你以為這話有理， 說：『我在上帝面前是公義的。』
JOB|35|3|你說：『這對你有甚麼益處？ 我不犯罪有甚麼好處呢？』
JOB|35|4|至於我，我要用言語回答你 和跟你一起的朋友。
JOB|35|5|你要向天觀看， 瞻望那高於你的穹蒼。
JOB|35|6|你若犯罪，能使上帝受何害呢？ 你的過犯加增，能使上帝受何損呢？
JOB|35|7|你若是公義，能加增他甚麼呢？ 他從你手裏還接受甚麼呢？
JOB|35|8|你的罪惡只影響像你這類的人； 你的公義也只影響世人。
JOB|35|9|「人因多受欺壓就哀求， 因強權者的膀臂而求救。
JOB|35|10|但無人說：『造我的上帝在哪裏？ 他使人夜間歌唱，
JOB|35|11|教導我們多過地上的走獸， 使我們比空中的飛鳥更聰明。』
JOB|35|12|因為惡人驕傲， 他們在那裏呼求，他卻不回答。
JOB|35|13|虛妄的呼求，上帝必不垂聽； 全能者必不留意。
JOB|35|14|何況你說，你不得見他。 案件就在他面前，你等候他吧。
JOB|35|15|但如今因他未曾發怒降罰， 也一點都不理會狂傲，
JOB|35|16|所以 約伯 開口說虛妄的話， 多多發表無知識的言語。」
JOB|36|1|以利戶 繼續說：
JOB|36|2|「你再給我片時，我就指示你， 因我還有話要為上帝說。
JOB|36|3|我要把我的知識從遠處引來， 我要將公義歸給造我的主。
JOB|36|4|我的言語絕不虛假， 有全備知識的與你同在。
JOB|36|5|「看哪，上帝有大能，並不藐視人； 他的心智能力廣大。
JOB|36|6|他不讓惡人活著， 卻為困苦人伸冤。
JOB|36|7|他的眼目不遠離義人， 卻使他們和君王同坐寶座， 永遠被高舉 。
JOB|36|8|他們若被鎖鏈捆住， 被苦難的繩索纏住，
JOB|36|9|他就向他們指示他們的作為和過犯， 以及他們的狂妄自大。
JOB|36|10|他也開通他們的耳朵來領受教導， 吩咐他們回轉離開罪孽。
JOB|36|11|他們若聽從事奉他， 就必度日亨通， 歷年享福。
JOB|36|12|他們若不聽從，就要被刀殺滅， 無知無識而死。
JOB|36|13|「那心中不敬虔的人積蓄怒氣； 上帝捆綁他們，他們竟不求救。
JOB|36|14|他們必在青年時死亡， 與神廟娼妓一樣喪命。
JOB|36|15|上帝藉著困苦救拔困苦人， 藉所受的欺壓開通他們的耳朵。
JOB|36|16|上帝也必引你脫離患難， 進入寬闊不狹窄之地； 擺在你席上的必滿有肥甘。
JOB|36|17|「但你充滿著惡人的辯辭， 辯辭和審判抓住你。
JOB|36|18|不可讓憤怒觸動你，使你破口謾罵 ； 也不可因贖價大而偏行。
JOB|36|19|你的呼求 和一切的勢力， 果真有用，使你不遭患難嗎？
JOB|36|20|不要切慕黑夜， 就是眾民在本處被除滅的時候。
JOB|36|21|你要謹慎，不可偏向罪孽， 因你選擇罪孽過於苦難。
JOB|36|22|看哪，上帝因他的能力而崇高； 有誰像他那樣作教師呢？
JOB|36|23|誰派定他的道路呢？ 誰能說：『你行了不義』？
JOB|36|24|「你要記得頌讚他的作為， 就是人所歌頌的。
JOB|36|25|他的作為，萬人都看見； 世人也從遠處觀看。
JOB|36|26|看哪，上帝崇高，我們不能知道； 他的年數，不能測度。
JOB|36|27|因他吸取水點， 水點就從雲霧中變成雨；
JOB|36|28|雲彩將雨落下， 沛然降於世人。
JOB|36|29|又有誰能明白密雲如何鋪張， 和上帝行宮的雷聲呢？
JOB|36|30|看哪，他的亮光普照自己的四圍； 他覆蓋海的深處。
JOB|36|31|因他用這些審判 眾民， 又賜豐富的糧食。
JOB|36|32|他以閃電遮手掌， 命令它擊中靶子。
JOB|36|33|所發的雷聲將他顯明， 牲畜也指明要起暴風 。」
JOB|37|1|「因此我心戰兢， 從原處移動。
JOB|37|2|聽啊，聽他轟轟的聲音， 是上帝口中所發的響聲。
JOB|37|3|他發響聲震遍天下， 他的閃電直到地極。
JOB|37|4|隨後，人聽見他的聲音， 是那轟轟的聲音； 他發出威嚴的雷聲， 而不加以遏止。
JOB|37|5|上帝發出奇妙的雷聲； 他行大事，我們不能測透。
JOB|37|6|他對雪說：『要降在地上』； 對大雨和暴雨也是這樣說。
JOB|37|7|他封住各人的手， 叫所造的萬人都知道他的作為。
JOB|37|8|野獸進入穴中， 臥在自己洞內。
JOB|37|9|暴風來自內宮， 寒冷出於狂風。
JOB|37|10|上帝噓氣成冰， 凝結寬闊之水，
JOB|37|11|使密雲盛滿水氣， 烏雲散佈閃電。
JOB|37|12|雲藉著他的指引遊行旋轉， 在世界的地面上行他一切所吩咐的，
JOB|37|13|或為責罰，或為他的地， 或為慈愛，都是他所行的。
JOB|37|14|「 約伯 啊，側耳聽這話， 要站立，思想上帝奇妙的作為。
JOB|37|15|你知道上帝如何安排這些， 如何使雲中的閃電照耀嗎？
JOB|37|16|你知道雲彩如何浮於空中， 知識全備者奇妙的作為嗎？
JOB|37|17|你知道南風使地寂靜， 你的衣服就變為熱嗎？
JOB|37|18|你豈能與上帝同鋪穹蒼， 堅固如同鑄成的鏡子嗎？
JOB|37|19|我們因在黑暗中，不會陳說， 請你指教我們該對他說甚麼。
JOB|37|20|有人告訴他我要說話嗎？ 豈有人說他願被吞滅嗎？
JOB|37|21|「現在，人不得見穹蒼的亮光； 風一吹過，天色晴朗。
JOB|37|22|金色的光輝來自北方， 在上帝那裏有可畏的威嚴。
JOB|37|23|全能者，我們不能測度； 他大有能力，又有公平， 滿有公義，必不苦待人。
JOB|37|24|所以，世人敬畏他； 凡自以為 有智慧的，他都不看顧。」
JOB|38|1|那時，耶和華從旋風中回答 約伯 說：
JOB|38|2|「誰用無知的言語使我的旨意暗昧不明？
JOB|38|3|你要如勇士束腰； 我問你，你可以讓我知道。
JOB|38|4|「我立大地根基的時候，你在哪裏？ 你若明白事理，只管說吧！
JOB|38|5|你知道是誰定地的尺度， 是誰把準繩拉在其上嗎？
JOB|38|6|地的根基安置在何處？ 地的角石是誰安放的？
JOB|38|7|那時，晨星一同歌唱； 上帝的眾使者也都歡呼。
JOB|38|8|「當海水衝出，如出母胎， 誰用門將它關閉呢？
JOB|38|9|是我用雲彩當海的衣服， 用幽暗當包裹它的布，
JOB|38|10|為它定界限， 又安門和閂，
JOB|38|11|說：『你只可到這裏，不可越過； 你狂傲的浪要到此止住。』
JOB|38|12|「你有生以來，曾命定晨光， 曾使黎明知道自己的地位，
JOB|38|13|抓住地的四極， 把惡人從其中驅逐出來嗎？
JOB|38|14|地改變如泥上蓋印， 萬物出現如衣服一樣。
JOB|38|15|亮光不照惡人， 高舉的膀臂也必折斷。
JOB|38|16|「你曾進到海之源， 或在深淵的隱密處行走嗎？
JOB|38|17|死亡的門曾向你顯露嗎？ 死蔭的門你曾見過嗎？
JOB|38|18|地的廣大，你能測透嗎？ 你若全知道，只管說吧！
JOB|38|19|「往光明居所的路在哪裏？ 黑暗的地方在何處？
JOB|38|20|你能將它帶到其領域， 能辨明其居所之路嗎？
JOB|38|21|你知道的，因為那時你已出生， 你活的日子數目也多。
JOB|38|22|「你曾進入雪之庫， 或見過雹的倉嗎？
JOB|38|23|雪雹是我為災難的時候， 為打仗和戰爭的日子所預備。
JOB|38|24|光亮從何路分開？ 東風從何路分散遍地？
JOB|38|25|「誰為大雨分道， 誰為雷電開路，
JOB|38|26|使雨降在無人之地， 在無人居住的曠野，
JOB|38|27|使荒廢淒涼之地得以豐足， 青草得以生長？
JOB|38|28|「雨有父親嗎？ 露珠是誰生的呢？
JOB|38|29|冰出於誰的胎？ 天上的霜是誰生的呢？
JOB|38|30|諸水堅硬如石頭， 深淵之面凝結成冰。
JOB|38|31|「你能為昴星繫結嗎？ 你能為參星解帶嗎？
JOB|38|32|你能按時領出星宿嗎？ 能引導北斗與其眾星嗎？
JOB|38|33|你知道天的定律嗎？ 你能使地歸其權下嗎？
JOB|38|34|「你能向密雲揚起聲來， 使傾盆的雨遮蓋你嗎？
JOB|38|35|你能發出閃電，使它們 行走， 並對你說：『我們在這裏』嗎？
JOB|38|36|誰將智慧放在朱鷺 中？ 誰將聰明賜給雄雞 ？
JOB|38|37|誰能用智慧數算雲彩？ 誰能傾倒天上的瓶呢？
JOB|38|38|那時，塵土聚集成團， 土塊緊緊結連。
JOB|38|39|「你能為母獅抓取獵物， 使少壯的獅子飽足嗎？
JOB|38|40|那時，牠們在洞中蹲伏， 在隱密處埋伏。
JOB|38|41|誰能為烏鴉預備食物呢？ 那時，烏鴉之雛哀求上帝， 因無食物飛來飛去。」
JOB|39|1|「你知道巖石間的野山羊幾時生產嗎？ 你能觀察母鹿下小鹿嗎？
JOB|39|2|你能數算牠們懷胎的月數嗎？ 你知道牠們幾時生產嗎？
JOB|39|3|牠們屈身，生下幼兒， 就解除了陣痛。
JOB|39|4|其子漸漸肥壯，在荒野長大； 牠們出去，不再歸回。
JOB|39|5|「誰放野驢自由？ 誰解開快驢的繩索？
JOB|39|6|我使曠野作牠的住處， 使鹽地當牠的居所。
JOB|39|7|牠嘲笑城內的喧嚷， 不聽趕牲口的喝聲。
JOB|39|8|諸山是牠漫遊的草場， 牠尋找各樣青綠之物。
JOB|39|9|「野牛豈肯服事你？ 豈肯在你的槽旁過夜？
JOB|39|10|你豈能用套繩將野牛繫於犁溝？ 牠豈肯隨你耙鬆山谷之地？
JOB|39|11|你豈可因牠力大就倚靠牠？ 豈可把你的工交給牠做呢？
JOB|39|12|你豈能靠牠把你的穀物運回， 又收聚在你的禾場上嗎？
JOB|39|13|「鴕鳥的翅膀歡然拍動， 但豈是鸛的翎毛和羽毛嗎 ？
JOB|39|14|因牠把蛋留在地上， 使蛋在塵土中得溫暖，
JOB|39|15|卻忘記腳會把蛋踹碎， 野獸會踐踏它。
JOB|39|16|牠粗暴待雛，似乎不是自己生的； 雖徒然勞苦 ，也不懼怕。
JOB|39|17|因為上帝使牠忘記智慧， 也未將悟性分給牠。
JOB|39|18|牠幾時挺身展開翅膀， 就嘲笑馬和騎馬的人。
JOB|39|19|「馬的力量是你所賜的嗎？ 牠頸項上的鬃是你披上的嗎？
JOB|39|20|是你叫牠跳躍像蝗蟲嗎？ 牠噴氣之威嚴使人驚惶。
JOB|39|21|牠用蹄在谷中挖地 ，以能力歡躍； 牠出去迎擊仇敵 。
JOB|39|22|牠嘲笑懼怕，並不驚惶， 也不因刀劍退卻。
JOB|39|23|箭袋在牠身上錚錚有聲， 槍和短槍閃閃發亮。
JOB|39|24|牠震顫激動，將地吞下 ； 一聽角聲就站不住。
JOB|39|25|每逢角聲一響，牠說：『啊哈！』 牠從遠處聞到戰爭的氣息， 聽見軍官如雷的吼聲和吶喊。
JOB|39|26|「鷹展開翅膀向南飛翔， 豈是藉著你的智慧嗎？
JOB|39|27|大鷹上騰在高處搭窩， 豈是聽你的指示嗎？
JOB|39|28|牠住在山巖， 以山峰和堅固之所為家，
JOB|39|29|從那裏窺察食物， 眼睛自遠方瞭望。
JOB|39|30|牠的雛吸血； 被殺的人在哪裏，牠也在哪裏。」
JOB|40|1|耶和華繼續對 約伯 說：
JOB|40|2|「強辯的豈可與全能者爭論？ 與上帝辯駁的可以回答吧！」
JOB|40|3|於是， 約伯 回答耶和華說：
JOB|40|4|「看哪，我是卑賤的！我用甚麼回答你呢？ 我只好用手摀住我的口。
JOB|40|5|我說了一次，就不回答； 說了兩次，不再說了。」
JOB|40|6|於是，耶和華從旋風中回答 約伯 說：
JOB|40|7|「你要如勇士束腰； 我問你，你可以讓我知道。
JOB|40|8|你豈可廢棄我的判斷？ 豈可定我有罪，好顯自己為義嗎？
JOB|40|9|你有上帝那樣的膀臂嗎？ 你能像他那樣發雷聲嗎？
JOB|40|10|「你要以榮耀莊嚴為妝飾， 以尊榮威嚴為衣服。
JOB|40|11|你要發出你滿溢的怒氣， 見一切驕傲的人，使他降卑；
JOB|40|12|你見一切驕傲的人，將他制伏， 把惡人踐踏在原來地方。
JOB|40|13|你將他們一同埋藏在塵土中， 把他們的臉遮蔽在隱密處 。
JOB|40|14|這樣，我也向你承認， 你的右手能救你自己。
JOB|40|15|「看哪，我造河馬， 也造了你； 牠吃草像牛一樣。
JOB|40|16|看哪，牠的力氣在腰間， 能力在肚腹的肌肉上。
JOB|40|17|牠挺直 尾巴如香柏樹， 牠大腿的筋緊密結合。
JOB|40|18|牠的骨頭好像銅管； 牠的肢體彷彿鐵棍。
JOB|40|19|「牠在上帝所造之物中為首， 只有創造牠的能攜刀臨近牠。
JOB|40|20|諸山為牠產出食物， 百獸也在那裏遊玩。
JOB|40|21|牠伏在蓮葉之下， 在蘆葦和沼澤的隱密處。
JOB|40|22|蓮葉的陰影遮蔽牠， 溪旁的柳樹環繞牠。
JOB|40|23|看哪，河水氾濫，牠不慌張； 連 約旦河 漲到牠口邊，牠也安然自若。
JOB|40|24|誰能在牠眼前捉拿牠呢？ 誰能以圈套穿牠鼻子呢？」
JOB|41|1|「你能用魚鉤釣上 力威亞探 嗎？ 能用繩子壓下牠的舌頭嗎？
JOB|41|2|你能用繩索穿牠的鼻子嗎？ 能用鉤子穿牠的腮骨嗎？
JOB|41|3|牠豈向你連連懇求， 向你說溫柔的話嗎？
JOB|41|4|牠豈肯與你立約， 讓你拿牠永遠作奴僕嗎？
JOB|41|5|你豈可拿牠當雀鳥玩耍？ 豈可將牠繫來給你幼女？
JOB|41|6|合夥的魚販豈可拿牠當貨物？ 他們豈可把牠分給商人呢？
JOB|41|7|你能用倒鉤扎滿牠的皮， 能用魚叉叉滿牠的頭嗎？
JOB|41|8|把你的手掌按在牠身上吧！ 想一想與牠搏鬥，你就不再這樣做了！
JOB|41|9|看哪，對牠有指望是徒然的； 一見牠，豈不也喪膽嗎？
JOB|41|10|沒有那麼兇猛的人敢惹牠。 這樣，誰能在我面前站立得住呢？
JOB|41|11|誰能與我對質，使我償還呢？ 天下萬物都是我的。
JOB|41|12|「我不能緘默不提 牠的肢體和力量，以及健美的骨骼。
JOB|41|13|誰能剝牠的外皮？ 誰能進牠的鎧甲之間 呢？
JOB|41|14|誰能開牠的腮頰？ 牠牙齒的四圍是可畏的。
JOB|41|15|牠的背上有一排排的鱗甲 ， 緊緊閉合，封得嚴密。
JOB|41|16|這鱗甲一一相連， 氣不得透入其間，
JOB|41|17|互相連接， 膠結一起，不能分開。
JOB|41|18|牠打噴嚏就發出光來， 牠的眼睛好像晨曦 。
JOB|41|19|從牠口中發出燒著的火把， 有火星飛迸出來；
JOB|41|20|從牠鼻孔冒出煙來， 如燒開的鍋在沸騰 。
JOB|41|21|牠的氣點著煤炭， 有火焰從牠口中發出。
JOB|41|22|牠頸項中存著勁力， 恐懼在牠面前蹦跳。
JOB|41|23|牠的肉塊緊緊結連， 緊貼其身，不能搖動。
JOB|41|24|牠的心結實如石頭， 如下面的磨石那樣結實。
JOB|41|25|牠一起來，神明都恐懼， 因崩潰而驚慌失措。
JOB|41|26|人用刀劍扎牠，是無用的， 槍、標槍、尖槍也一樣。
JOB|41|27|牠以鐵為乾草， 以銅為爛木。
JOB|41|28|箭不能使牠逃走， 牠看彈石如碎秸。
JOB|41|29|牠當棍棒作碎秸， 牠嘲笑短槍的颼颼聲。
JOB|41|30|牠肚腹下面是尖瓦片； 牠如釘耙刮過淤泥。
JOB|41|31|牠使深淵滾沸如鍋， 使海洋如鍋中膏油。
JOB|41|32|牠使走過以後的路發光， 令人覺得深淵如同白髮。
JOB|41|33|塵世上沒有像牠那樣的受造物， 一無所懼。
JOB|41|34|凡高大的，牠盯著看； 牠在一切狂傲的野獸中作王。」
JOB|42|1|約伯 回答耶和華說：
JOB|42|2|「我知道，你萬事都能做； 你的計劃不能攔阻。
JOB|42|3|誰無知使你的旨意隱藏呢？ 因此我說的，我不明白； 這些事太奇妙，是我不知道的。
JOB|42|4|求你聽我，我要說話； 我問你，求你讓我知道。
JOB|42|5|我從前風聞有你， 現在親眼看見你。
JOB|42|6|因此我撤回 ， 在塵土和爐灰中懊悔。」
JOB|42|7|耶和華對 約伯 說話以後，耶和華就對 提幔 人 以利法 說：「我的怒氣向你和你兩個朋友發作，因為你們議論我，不如我的僕人 約伯 說的正確。
JOB|42|8|現在你們要為自己取七頭公牛，七隻公羊，到我的僕人 約伯 那裏去，為自己獻上燔祭，我的僕人 約伯 就為你們祈禱。我必悅納他，不按你們的愚妄處置你們。你們議論我，不如我的僕人 約伯 說的正確。」
JOB|42|9|於是 提幔 人 以利法 、 書亞 人 比勒達 、 拿瑪 人 瑣法 遵照耶和華所吩咐的去做，耶和華就悅納 約伯 。
JOB|42|10|約伯 為他的朋友祈禱。耶和華就使 約伯 從苦境 中轉回，並且耶和華賜給他的比他從前所有的加倍。
JOB|42|11|約伯 的兄弟、姊妹，和以前所認識的人都來到他那裏，在他家裏跟他一同吃飯。他們因耶和華所降於他的一切災禍，都為他悲傷，安慰他。每人送他一塊可錫塔 和一個金環。
JOB|42|12|這樣，耶和華後來賜福給 約伯 比先前更多。他有一萬四千隻羊，六千匹駱駝，一千對牛，一千匹母驢。
JOB|42|13|他也有七個兒子，三個女兒。
JOB|42|14|他給長女起名叫 耶米瑪 ，次女叫 基洗亞 ，三女叫 基連哈樸 。
JOB|42|15|在全地的婦女中找不著像 約伯 的女兒那樣美貌的。她們的父親使她們在兄弟中得產業。
JOB|42|16|此後， 約伯 又活了一百四十年，得見他的四代兒孫。
JOB|42|17|這樣， 約伯 年紀老邁，日子滿足而死。
