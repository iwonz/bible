JUDE|1|1|耶稣基督的仆人、 雅各 的兄弟 犹大 ，写信给那些被召、在父上帝里蒙爱、为耶稣基督保守的人。
JUDE|1|2|愿怜悯、平安 、慈爱多多加给你们！
JUDE|1|3|亲爱的，我一直很迫切地想要写信给你们，论到我们同享的救恩，但我觉得有必要现在就写信劝你们，要为从前一次交付给圣徒的真道竭力奋斗。
JUDE|1|4|因为有些人偷偷地进来，就是早就被判定受惩罚的不虔诚的人，他们把我们上帝的恩典变为放纵情欲的机会，并且不认独一的主宰—我们的主耶稣基督。
JUDE|1|5|这一切的事，你们虽然知道，我却仍要提醒你们：从前主 只一次就 救了他的百姓出 埃及 地，后来却把那些不信的灭绝了。
JUDE|1|6|至于那些不守本位、离开自己住处的天使，主用锁链把他们永远拘留在黑暗里，等候大日子的审判。
JUDE|1|7|同样， 所多玛 、 蛾摩拉 和周围城镇的人也跟着他们一样犯淫乱，随从逆性的情欲，以致遭受永不熄灭之火的惩罚，作为众人的鉴戒。
JUDE|1|8|照样，这些做梦的人也污秽身体，轻慢掌权者，毁谤众尊荣者。
JUDE|1|9|天使长 米迦勒 为 摩西 的尸首与魔鬼争辩的时候，尚且不敢用毁谤的话谴责他，只说：“主责备你吧！”
JUDE|1|10|但这些人毁谤他们所不知道的。他们与那些没有理性的牲畜一样，只做本性所知道的事，败坏了自己。
JUDE|1|11|他们有祸了！因为他们走 该隐 的道路，又为财利往 巴兰 的错谬里直奔，并在 可拉 的背叛中灭亡了。
JUDE|1|12|这样的人是你们爱筵上的污点 ；他们无所惧怕地同你们宴乐，仿佛牧人只顾喂饱自己。他们是无雨的浮云，被风飘荡；是秋天没有果子的树，死而又死，连根被拔出来；
JUDE|1|13|是海里的狂浪，涌出自己可耻的沫子来；是流荡的星，有漆黑的幽暗永远为他们保留着。
JUDE|1|14|亚当 的七世孙 以诺 曾预言这些人说：“看哪，主带着他的千万圣者来临，
JUDE|1|15|要审判众人，证实一切不敬虔的人所妄行一切不敬虔的事，又证实不敬虔的罪人所说顶撞他的刚愎的话。”
JUDE|1|16|这些人喜出怨言，责怪他人，随从自己的情欲而行，口说夸大的话，为自己的利益谄媚人。
JUDE|1|17|亲爱的，至于你们，要记得我们主耶稣基督的使徒从前所说的话。
JUDE|1|18|他们曾对你们说过，末世必有好嘲弄的人随从自己不敬虔的私欲而行。
JUDE|1|19|这就是那些好结党分派、属乎血气、没有圣灵的人。
JUDE|1|20|亲爱的，至于你们，要在至圣的真道上造就自己，藉着圣灵祷告，
JUDE|1|21|保守自己常在上帝的爱中，仰望我们主耶稣基督的怜悯，进入永生。
JUDE|1|22|有些人心中犹疑 ，你们要怜悯 他们；
JUDE|1|23|有些人你们要从火中抢出来，搭救他们 ；有些人你们要存惧怕的心怜悯他们，连那被情欲污染的衣服也要厌恶。
JUDE|1|24|愿那能保守你们不失脚，使你们无瑕无疵、欢欢喜喜站在他荣耀之前的、
JUDE|1|25|我们的救主独一的上帝，藉着我们的主耶稣基督，得享荣耀、威严、能力、权柄，从万古以前，到现今，直到永永远远。阿们！
