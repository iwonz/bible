1KGS|1|1|大衛 王年紀老邁，雖然蓋著外袍，仍不夠暖和。
1KGS|1|2|臣僕對他說：「不如為我主我王找一個年輕的少女，侍立在王面前，照顧王，睡在王的懷中，好使我主我王得暖。」
1KGS|1|3|於是他們在 以色列 全境尋找美貌的少女，找到了一個 書念 女子 亞比煞 ，帶到王那裏。
1KGS|1|4|這少女極其美貌，她照顧王，伺候王，王卻沒有與她親近。
1KGS|1|5|那時， 哈及 的兒子 亞多尼雅 妄自尊大，說：「我要作王」，就為自己預備座車、騎兵，又派五十人在他前頭奔跑。
1KGS|1|6|他父親從來沒有責怪他，說：「你為何這麼做？」他非常俊美，生在 押沙龍 之後。
1KGS|1|7|亞多尼雅 與 洗魯雅 的兒子 約押 和 亞比亞他 祭司商議；他們就順從 亞多尼雅 ，幫助他。
1KGS|1|8|但 撒督 祭司、 耶何耶大 的兒子 比拿雅 、 拿單 先知、 示每 、 利以 ，以及 大衛 自己的勇士 都不順從 亞多尼雅 。
1KGS|1|9|亞多尼雅 在 隱‧羅結 旁 瑣希列 磐石那裏獻牛羊、肥犢為祭，請了他的眾兄弟，就是王的眾兒子，以及所有作王臣僕的 猶大 人。
1KGS|1|10|但他沒有邀請 拿單 先知、 比拿雅 和勇士們，以及他的弟弟 所羅門 。
1KGS|1|11|拿單 對 所羅門 的母親 拔示巴 說：「 哈及 的兒子 亞多尼雅 作王了，你沒有聽見嗎？我們的主 大衛 卻不知道。
1KGS|1|12|現在，來，我給你出個主意，好保全你和你兒子 所羅門 的性命。
1KGS|1|13|你去，進到 大衛 王那裏，對他說：『我主我王啊，你不是曾向使女起誓說：你兒子 所羅門 必接續我作王，他必坐在我的王位上嗎？ 亞多尼雅 怎麼作了王呢？』
1KGS|1|14|看哪，你還在那裏與王說話的時候，我會隨後進去，證實你的話。」
1KGS|1|15|拔示巴 進入內室，到王那裏。那時，王很老了， 書念 女子 亞比煞 正伺候著王。
1KGS|1|16|拔示巴 向王屈身下拜，王說：「你要甚麼？」
1KGS|1|17|她對王說：「我主啊，你曾向使女指著耶和華－你的上帝起誓：『你兒子 所羅門 必接續我作王，他必坐在我的王位上。』
1KGS|1|18|現在，看哪， 亞多尼雅 作王了，你 ，我主我王卻不知道。
1KGS|1|19|他獻許多牛羊、肥犢為祭，請了王的眾兒子和 亞比亞他 祭司，以及 約押 元帥，他卻沒有請王的僕人 所羅門 。
1KGS|1|20|但你 ，我主我王啊， 以色列 眾人的眼目都仰望你，等你告訴他們，在我主我王之後誰坐你的王位。
1KGS|1|21|若不然，我主我王與祖先同睡的時候，我和我兒子 所羅門 必列為罪犯了。」
1KGS|1|22|看哪， 拔示巴 還與王說話的時候， 拿單 先知也進來了。
1KGS|1|23|有人奏告王說：「看哪， 拿單 先知來了。」 拿單 進到王面前，臉伏於地，向王叩拜。
1KGS|1|24|拿單 說：「我主我王，你果真說過『 亞多尼雅 必接續我作王，他要坐在我的王位上』嗎？
1KGS|1|25|他今日下去，獻了許多牛羊、肥犢為祭，請了王的眾兒子和軍官們，以及 亞比亞他 祭司；看哪，他們正在 亞多尼雅 面前吃喝，說：『 亞多尼雅 王萬歲！』
1KGS|1|26|至於我，就是你的僕人，和 撒督 祭司、 耶何耶大 的兒子 比拿雅 、王的僕人 所羅門 ，他都沒有請。
1KGS|1|27|這事果真出於我主我王嗎？王卻沒有告訴僕人們，在我主我王之後誰坐你的王位。」
1KGS|1|28|大衛 王回答說：「召 拔示巴 到我這裏來。」 拔示巴 就來，站在王面前。
1KGS|1|29|王起誓說：「我指著救我性命脫離一切苦難的永生的耶和華起誓。
1KGS|1|30|我既然指著耶和華－ 以色列 的上帝向你起誓說：你兒子 所羅門 必接續我作王，他必繼承我坐在我的王位上，我今日必這樣做。」
1KGS|1|31|於是， 拔示巴 屈身，臉伏於地，向王叩拜，說：「我主 大衛 王萬歲！」
1KGS|1|32|大衛 王又說：「召 撒督 祭司、 拿單 先知、 耶何耶大 的兒子 比拿雅 到我這裏來！」他們就都來到王面前。
1KGS|1|33|王對他們說：「要帶領你們主的僕人，讓我兒子 所羅門 騎我自己的騾子，送他下到 基訓 。
1KGS|1|34|在那裏， 撒督 祭司和 拿單 先知要膏他作 以色列 的王；你們也要吹角，說：『 所羅門 王萬歲！』
1KGS|1|35|你們要跟隨他上來，使他坐在我的王位上，他要接續我作王。我已立他作 以色列 和 猶大 的君王。」
1KGS|1|36|耶何耶大 的兒子 比拿雅 回應王說：「阿們！願耶和華－我主我王的上帝這樣說。
1KGS|1|37|耶和華怎樣與我主我王同在，願他照樣與 所羅門 同在，使他的王位比我主 大衛 王的王位更大。」
1KGS|1|38|於是， 撒督 祭司、 拿單 先知、 耶何耶大 的兒子 比拿雅 ，以及 基利提 人和 比利提 人都下去，讓 所羅門 騎上 大衛 王的騾子，送他到 基訓 。
1KGS|1|39|撒督 祭司從帳幕中取了盛膏油的角來，膏 所羅門 。他們就吹角，眾百姓都說：「 所羅門 王萬歲！」
1KGS|1|40|眾百姓跟隨他上來，吹著笛，大大歡呼，地被他們的聲音震裂。
1KGS|1|41|亞多尼雅 和所有的賓客剛吃完，聽見這聲音； 約押 聽見角聲就說：「城中為何有這響聲呢？」
1KGS|1|42|他正說話的時候，看哪， 亞比亞他 祭司的兒子 約拿單 來了。 亞多尼雅 說：「進來吧！你是個賢明的人，必是來報好消息的。」
1KGS|1|43|約拿單 回答 亞多尼雅 說：「我們的主 大衛 王已經立 所羅門 為王了！
1KGS|1|44|王派 撒督 祭司、 拿單 先知、 耶何耶大 的兒子 比拿雅 ，以及 基利提 人和 比利提 人和 所羅門 一起去，叫他騎上王的騾子。
1KGS|1|45|撒督 祭司和 拿單 先知已經在 基訓 膏他作王了。他們從那裏歡呼著上來，城都震動，這就是你們所聽見的聲音。
1KGS|1|46|所羅門 也已經登上國度的王位了。
1KGS|1|47|王的臣僕也來為我們的主 大衛 王祝福，說：『願上帝使 所羅門 的名比你的名更尊榮，使他的王位比你的王位更大。』王在床上屈身敬拜，
1KGS|1|48|王也這樣說：『耶和華－ 以色列 的上帝是應當稱頌的，因他今日賞賜一個人坐在我的王位上，我也親眼看見了。』」
1KGS|1|49|亞多尼雅 所有的賓客都戰兢，起來，各走各路去了。
1KGS|1|50|亞多尼雅 懼怕 所羅門 ，就起來，去抓住祭壇的翹角。
1KGS|1|51|有人告訴 所羅門 說：「看哪， 亞多尼雅 懼怕 所羅門 王。看哪，他抓住祭壇的翹角，說：『願 所羅門 王先向我起誓，必不用刀殺死僕人。』」
1KGS|1|52|所羅門 說：「他若作賢明的人，連一根頭髮也不致落在地上；他若作惡，必要死亡。」
1KGS|1|53|於是 所羅門 王派人叫 亞多尼雅 從壇上下來，他就來向 所羅門 王下拜。 所羅門 對他說：「你回家去吧！」
1KGS|2|1|大衛 的死期臨近了，就吩咐他兒子 所羅門 說：
1KGS|2|2|「我要走世人必走的路了。你當剛強，作大丈夫，
1KGS|2|3|遵守耶和華－你上帝所吩咐的，照著 摩西 律法上所寫的行耶和華的道，謹守他的律例、誡命、典章、法度，好讓你無論做甚麼，不拘往何處去，盡都亨通。
1KGS|2|4|耶和華必成就他所說關於我的話，說：『你的子孫若謹慎自己的行為，盡心盡意憑信實行在我面前，就不斷有人坐 以色列 的王位。』
1KGS|2|5|你也知道 洗魯雅 的兒子 約押 向我所做的事，他對付 以色列 的兩個元帥， 尼珥 的兒子 押尼珥 和 益帖 的兒子 亞瑪撒 ，殺了他們。他在太平之時，如同戰爭一般，流這二人的血，把這戰爭的血染了他腰間束的帶和腳上穿的鞋。
1KGS|2|6|所以你要照你的智慧去做，不讓他白髮安然下陰間。
1KGS|2|7|你當恩待 基列 人 巴西萊 的眾兒子，請他們常與你同席吃飯，因為我躲避你哥哥 押沙龍 的時候，他們親近我。
1KGS|2|8|看哪，在你這裏有來自 巴戶琳 的 便雅憫 人， 基拉 的兒子 示每 。我到 瑪哈念 去的那日，他用狠毒的言語咒罵我。後來他卻下 約旦河 迎接我，我就指著耶和華向他起誓說：『我必不用刀殺死你。』
1KGS|2|9|但現在你不要以他為無罪。你是有智慧的人，必知道怎樣待他，使他白髮流血下陰間。」
1KGS|2|10|大衛 與他祖先同睡，葬在 大衛城 。
1KGS|2|11|大衛 作 以色列 王四十年：在 希伯崙 作王七年，在 耶路撒冷 作王三十三年。
1KGS|2|12|所羅門 坐他父親 大衛 的王位，他的國度非常穩固。
1KGS|2|13|哈及 的兒子 亞多尼雅 到 所羅門 的母親 拔示巴 那裏， 拔示巴 問他說：「你是為平安來的嗎？」他說：「為平安來的。」
1KGS|2|14|他又說：「我有話對你說。」 拔示巴 說：「你說吧。」
1KGS|2|15|亞多尼雅 說：「你知道這國原是歸我的，全 以色列 也都期望我作王。然而，這國反歸了我兄弟，因這國歸了他是出乎耶和華。
1KGS|2|16|現在我有一件事求你，請你不要推辭。」 拔示巴 對他說：「你說吧。」
1KGS|2|17|他說：「求你請 所羅門 王把 書念 女子 亞比煞 賜我為妻，因他必不拒絕你。」
1KGS|2|18|拔示巴 說：「好，我必為你對王提說。」
1KGS|2|19|於是， 拔示巴 來到 所羅門 王那裏，要為 亞多尼雅 說話。王起來迎接，向她下拜，然後坐在自己的位上，又為王的母親設一座位，她就坐在王的右邊。
1KGS|2|20|拔示巴 說：「我要向你提出一個小小的請求，請你不要回絕我。」王對她說：「母親，請提出來，我必不回絕你。」
1KGS|2|21|拔示巴 說：「請你把 書念 女子 亞比煞 賜給你哥哥 亞多尼雅 為妻。」
1KGS|2|22|所羅門 王回答母親說：「為何替 亞多尼雅 求 書念 女子 亞比煞 呢？可以為他求王國吧！他是我的兄長，不但為他，也為 亞比亞他 祭司和 洗魯雅 的兒子 約押 求吧！ 」
1KGS|2|23|所羅門 王指著耶和華起誓說：「 亞多尼雅 講這話是自己送命，不然，願上帝重重懲罰我。
1KGS|2|24|耶和華堅立我，使我坐在父親 大衛 的王位上，照著他所應許的為我建立家室；現在我指著永生的耶和華起誓， 亞多尼雅 今日必被處死。」
1KGS|2|25|於是 所羅門 王派 耶何耶大 的兒子 比拿雅 去擊殺 亞多尼雅 ，他就死了。
1KGS|2|26|王對 亞比亞他 祭司說：「你回 亞拿突 歸自己的田地去吧！你本是該死的，但因你在我父親 大衛 面前抬過主耶和華的約櫃，又與我父親同受一切苦難，所以我今日不殺死你。」
1KGS|2|27|所羅門 就革除 亞比亞他 ，不讓他作耶和華的祭司。這就應驗了耶和華在 示羅 論 以利 家所說的話。
1KGS|2|28|雖然 約押 沒有擁護 押沙龍 ，卻擁護了 亞多尼雅 ；這消息傳到 約押 那裏，他就逃到耶和華的帳幕，抓住祭壇的翹角。
1KGS|2|29|有人告訴 所羅門 王：「 約押 逃到耶和華的帳幕，看哪，他在祭壇的旁邊。」 所羅門 就派 耶何耶大 的兒子 比拿雅 ，說：「去，殺了他。」
1KGS|2|30|比拿雅 來到耶和華的帳幕，對 約押 說：「王這樣吩咐：『你出來吧！』」他說：「不，我要死在這裏。」 比拿雅 就去回覆王，說：「 約押 這樣說，他這樣回答我。」
1KGS|2|31|王對他說：「你可以照著他的話去做，殺了他，把他葬了，好叫 約押 流無辜人血的罪不歸在我和我的父家。
1KGS|2|32|耶和華必使 約押 的血歸到他自己頭上，因為他擊殺兩個比他又公義又良善的人，就是 尼珥 的兒子 以色列 的元帥 押尼珥 和 益帖 的兒子 猶大 的元帥 亞瑪撒 ，用刀殺了他們，我父親 大衛 卻不知道。
1KGS|2|33|這二人的血必歸到 約押 和他後裔頭上，直到永遠；惟有 大衛 和他的後裔，以及他的家與王位，必從耶和華那裏得平安，直到永遠。」
1KGS|2|34|於是 耶何耶大 的兒子 比拿雅 上去，擊殺 約押 ，殺死他，把他葬在曠野 約押 自己的家裏。
1KGS|2|35|王就立 耶何耶大 的兒子 比拿雅 作元帥，代替 約押 ，又使 撒督 祭司代替 亞比亞他 。
1KGS|2|36|王派人召 示每 來，對他說：「你要在 耶路撒冷 為自己建造房屋，住在那裏，不可從那裏出來到任何地方去。
1KGS|2|37|你當確實知道，你何日出來過 汲淪溪 ，就必定死！你的血必歸到自己頭上。」
1KGS|2|38|示每 對王說：「這話很好！我主我王怎樣說，僕人必照樣做。」於是 示每 住在 耶路撒冷 許多日子。
1KGS|2|39|過了三年， 示每 的兩個奴僕逃到 瑪迦 的兒子 迦特 王 亞吉 那裏去。有人告訴 示每 說：「看哪，你的奴僕在 迦特 。」
1KGS|2|40|示每 起來，備上驢，往 迦特 到 亞吉 那裏去找他的奴僕，從 迦特 帶他的奴僕回來。
1KGS|2|41|有人告訴 所羅門 ：「 示每 出 耶路撒冷 到 迦特 去，又回來了。」
1KGS|2|42|王就派人召 示每 來，對他說：「我豈不是叫你指著耶和華起誓，並且警告你說『你當確實知道，你何日出來到任何地方去，就必定死』嗎？你也對我說：『這話很好，我必聽從。』
1KGS|2|43|你為何不遵守你對耶和華的誓言和我吩咐你的命令呢？」
1KGS|2|44|王又對 示每 說：「你向我父親 大衛 所做的一切惡事，你自己心裏都知道，耶和華必使你的罪惡歸到你自己的頭上。
1KGS|2|45|但 所羅門 王必蒙福， 大衛 的王位必在耶和華面前堅立，直到永遠。」
1KGS|2|46|於是王吩咐 耶何耶大 的兒子 比拿雅 ，他就出去，擊殺 示每 ， 示每 就死了。這樣，國度在 所羅門 的手中鞏固了。
1KGS|3|1|所羅門 與 埃及 王法老結親，娶了法老的女兒，接她進入 大衛城 ，直等到建完了自己的宮和耶和華的殿，以及 耶路撒冷 周圍的城牆。
1KGS|3|2|當那些日子，百姓仍在丘壇獻祭，因為還沒有為耶和華的名建殿。
1KGS|3|3|所羅門 愛耶和華，遵行他父親 大衛 的律例，只是還在丘壇獻祭燒香。
1KGS|3|4|所羅門 王到 基遍 ，在那裏獻祭，因為 基遍 有極大的丘壇。 所羅門 在那壇上獻了一千祭牲為燔祭。
1KGS|3|5|在 基遍 ，耶和華夜間在夢中向 所羅門 顯現；上帝說：「你願我賜你甚麼，你可以求。」
1KGS|3|6|所羅門 說：「你曾向你僕人我父親 大衛 大施慈愛，因為他用忠信、公義、正直的心行在你面前。你又為他存留大慈愛，賜他一個兒子坐在他的王位上，正如今日一樣。
1KGS|3|7|現在，耶和華－我的上帝啊，你使僕人接續我父親 大衛 作王；但我是幼小的孩子，不知道應當怎樣出入。
1KGS|3|8|僕人住在你揀選的百姓中，這百姓之多，多得不可點，不可算。
1KGS|3|9|所以求你賜僕人善於了解的心，可以判斷你的百姓，辨別是非。不然，誰能判斷你這麼多的百姓呢？」
1KGS|3|10|所羅門 因為求這事，就蒙主喜悅。
1KGS|3|11|上帝對他說：「你既然求這事，不為自己求壽、求富，也不求滅絕你仇敵的性命，只求能明辨，可以聽訟，
1KGS|3|12|看哪，我會照你的話去做，看哪，我會賜你智慧和明辨的心，在你以前沒有像你的，在你以後也沒有興起像你的。
1KGS|3|13|你沒有求的，我也賜給你，就是富足、尊榮，使你在世一切的日子，列王中沒有一個能比你的。
1KGS|3|14|你若遵行我的道，謹守我的律例、誡命，正如你父親 大衛 所行的，我必使你長壽。」
1KGS|3|15|所羅門 醒了，看哪，是個夢。他就來到 耶路撒冷 ，站在耶和華的約櫃前，獻燔祭和平安祭，又為眾臣僕擺設宴席。
1KGS|3|16|那時，有兩個妓女來，站在王面前。
1KGS|3|17|一個婦人說：「我主啊，我和這婦人同住一屋。她在屋子裏的時候，我生了一個孩子。
1KGS|3|18|我生了以後第三天，這婦人也生了。我們是一起的，屋子裏除了我們二人之外，再沒有別人在屋子裏。
1KGS|3|19|夜間，這婦人的兒子死了，因為她壓在她的兒子身上。
1KGS|3|20|她半夜起來，趁你使女睡著的時候，從我旁邊把我兒子抱走，放在她懷裏，又把她死的兒子放在我懷裏。
1KGS|3|21|清早，我起來要給我的兒子吃奶，看哪，他死了；早晨我仔細察看他，看哪，他不是我所生的兒子。」
1KGS|3|22|另一個婦人說：「不！我的兒子是活的，你的兒子是死的。」但這一個說：「不！你的兒子是死的，我的兒子是活的。」她們就在王面前爭吵。
1KGS|3|23|王說：「這婦人說：『這是我的兒子，他是活的，你的兒子是死的。』那婦人說：『不！你的兒子是死的，我的兒子是活的。』」
1KGS|3|24|王就說：「給我拿刀來！」人就把刀拿到王面前來。
1KGS|3|25|王說：「把活孩子劈成兩半，一半給這婦人，一半給那婦人。」
1KGS|3|26|活孩子的母親為自己的兒子心急如焚，對王說：「求我主把活孩子給那婦人吧，萬不可殺死他！」那婦人說：「這孩子也不歸我，也不歸你，你們就劈了吧！」
1KGS|3|27|王回應說：「把活孩子給這婦人，萬不可殺死他，因為這婦人是他的母親。」
1KGS|3|28|全 以色列 聽見王這樣判斷，就都敬畏王，因為他們看見他心中有上帝的智慧，能夠斷案。
1KGS|4|1|所羅門 作全 以色列 的王。
1KGS|4|2|這些是他的官員： 撒督 的兒子 亞撒利雅 作祭司，
1KGS|4|3|示沙 的兩個兒子 以利何烈 、 亞希亞 作書記， 亞希律 的兒子 約沙法 作史官，
1KGS|4|4|耶何耶大 的兒子 比拿雅 作元帥， 撒督 和 亞比亞他 作祭司，
1KGS|4|5|拿單 的兒子 亞撒利雅 作宰相， 拿單 的兒子 撒布得 作祭司和王的顧問，
1KGS|4|6|亞希煞 作管家， 亞比大 的兒子 亞多尼蘭 掌管服勞役的工人。
1KGS|4|7|所羅門 在全 以色列 有十二個官員，供給王和王室的食物，每年各人供給一個月。
1KGS|4|8|這些是他們的名字：在 以法蓮 山區有 便‧戶珥 ；
1KGS|4|9|在 瑪迦斯 、 沙賓 、 伯‧示麥 、 以倫‧伯‧哈南 有 便‧底甲 ；
1KGS|4|10|在 亞魯泊 有 便‧希悉 ，他管理 梭哥 和 希弗 全地；
1KGS|4|11|在 多珥 山岡 有 便‧亞比拿達 ，他娶了 所羅門 的女兒 她法 為妻；
1KGS|4|12|在 他納 和 米吉多 ，以及靠近 撒拉他拿 、 耶斯列 下邊的 伯‧善 全地，從 伯‧善 到 亞伯‧米何拉 直到 約緬 的另一邊有 亞希律 的兒子 巴拿 ；
1KGS|4|13|在 基列 的 拉末 有 便‧基別 ，他管理在 基列 的 瑪拿西 子孫 睚珥 的城鎮， 巴珊 的 亞珥歌伯 地的六十座大城，各有城牆和銅閂；
1KGS|4|14|在 瑪哈念 有 易多 的兒子 亞希拿達 ；
1KGS|4|15|在 拿弗他利 有 亞希瑪斯 ，他也娶了 所羅門 的一個女兒 巴實抹 為妻；
1KGS|4|16|在 亞設 和 亞祿 有 戶篩 的兒子 巴拿 ；
1KGS|4|17|在 以薩迦 有 帕路亞 的兒子 約沙法 ；
1KGS|4|18|在 便雅憫 有 以拉 的兒子 示每 ；
1KGS|4|19|在 基列 地，就是 亞摩利 王 西宏 和 巴珊 王 噩 之地，有 烏利 的兒子 基別 ，他一個官員管理這地 。
1KGS|4|20|猶大 人和 以色列 人如同海邊的沙那樣多，都吃喝快樂。
1KGS|4|21|所羅門 統治諸國，從 大河 到 非利士 地，直到 埃及 的邊界。 所羅門 在世的日子，這些國都向他進貢，服事他。
1KGS|4|22|所羅門 每日所用的食物：三十歌珥細麵，六十歌珥粗麵，
1KGS|4|23|十頭肥牛，二十頭草場的牛，一百隻羊，還有鹿、羚羊、麃子，以及肥禽。
1KGS|4|24|所羅門 管理整個 大河 西邊，從 提弗薩 直到 迦薩 ，以及 大河 西邊的諸王，屬他的四境盡都平安。
1KGS|4|25|所羅門 在世的日子，從 但 到 別是巴 ， 猶大 和 以色列 各人都在自己的葡萄樹下和無花果樹下安然居住。
1KGS|4|26|所羅門 擁有給戰車用的四萬個 馬棚，還有一萬二千名騎兵。
1KGS|4|27|這些官員各按自己的月份供給 所羅門 王，以及一切與他同席之人的食物，一無所缺。
1KGS|4|28|他們各按其分，把給馬與快馬吃的大麥和乾草送到指定的地方去。
1KGS|4|29|上帝賜給 所羅門 極大的智慧和聰明，以及寬闊的心，如同海邊的沙。
1KGS|4|30|所羅門 的智慧超過所有東方人的智慧，和 埃及 人一切的智慧。
1KGS|4|31|他的智慧勝過萬人，勝過 以斯拉 人 以探 ，以及 瑪曷 的兒子 希幔 、 甲各 、 達大 。他的名聲傳遍四圍的列國。
1KGS|4|32|他作箴言三千句，詩歌一千零五首。
1KGS|4|33|他講論草木，從 黎巴嫩 的香柏樹直到牆上長的牛膝草，又講論飛禽、走獸、爬行動物和魚類。
1KGS|4|34|地上凡曾聽過他智慧的君王，都派人來；萬民都有人來聽 所羅門 的智慧。
1KGS|5|1|推羅 王 希蘭 是 大衛 平生的好友。 希蘭 聽見 以色列 人膏 所羅門 接續他父親作王，就派臣僕到他那裏。
1KGS|5|2|所羅門 也派人到 希蘭 那裏，說：
1KGS|5|3|「你知道我父親 大衛 因四圍的戰爭，不能為耶和華－他上帝的名建殿，直等到耶和華使仇敵都服在他腳下。
1KGS|5|4|現在耶和華－我的上帝使我四圍太平，沒有仇敵，沒有災禍。
1KGS|5|5|看哪，我吩咐要為耶和華－我上帝的名建殿，是照耶和華向我父親 大衛 說的：『我必使你兒子接續你，坐你的王位，他必為我的名建殿。』
1KGS|5|6|現在，請吩咐人在 黎巴嫩 為我砍伐香柏木，我的僕人必幫助你的僕人。至於你僕人的工錢，我必照你所定的給你。你知道，在我們中間沒有人像 西頓 人那樣擅長砍伐樹木。」
1KGS|5|7|希蘭 聽見 所羅門 的話，就很高興，說：「今日耶和華是應當稱頌的，因為他賜給 大衛 一個有智慧的兒子，治理這眾多的百姓。」
1KGS|5|8|希蘭 送信給 所羅門 ，說：「你派人向我所提的那事，我已聽見了；論到香柏木和松木，我必照你一切的心願去做。
1KGS|5|9|我的僕人必把這木料從 黎巴嫩 運到海裏，我會把它們紮成筏子浮在海上，運到你告訴我的地方，在那裏拆開，你就可以收取；你也要照我的心願做，把食物給我的家。」
1KGS|5|10|於是 希蘭 照 所羅門 的心願，給他香柏木和松木；
1KGS|5|11|所羅門 給 希蘭 二萬歌珥麥子，二十歌珥 搗成的油，作他家的食物。 所羅門 每年都是這樣給 希蘭 。
1KGS|5|12|耶和華照著所應許的賜智慧給 所羅門 。 希蘭 與 所羅門 和平相處，二人彼此立約。
1KGS|5|13|所羅門 王從全 以色列 挑取服勞役的人，徵來的人有三萬，
1KGS|5|14|派他們輪流每月一萬人上 黎巴嫩 去；一個月在 黎巴嫩 ，兩個月在家裏。 亞多尼蘭 管理他們。
1KGS|5|15|所羅門 有七萬扛抬的，八萬在山上鑿石頭的。
1KGS|5|16|此外， 所羅門 有三千三百個監督工作的官長，監管百姓做工。
1KGS|5|17|王下令，他們就鑿出又大又貴重的石頭來，用以立殿的根基。
1KGS|5|18|所羅門 的工匠和 希蘭 的工匠，以及 迦巴勒 人，把石頭鑿好，預備了木料和石頭來建殿。
1KGS|6|1|以色列 人出 埃及 地後四百八十年， 所羅門 作 以色列 王第四年西弗月，就是二月，他開工建造耶和華的殿。
1KGS|6|2|所羅門 王為耶和華所建的殿，長六十肘，寬二十肘，高三十肘。
1KGS|6|3|殿的正堂前走廊長二十肘，與殿的寬度一樣，殿前寬十肘；
1KGS|6|4|他為殿做了有框嵌壁式的窗戶。
1KGS|6|5|靠著殿牆，圍著外殿和內殿的牆，周圍建造了廂房；
1KGS|6|6|下層寬五肘，中層寬六肘，第三層寬七肘。他在殿牆的周圍造坎，免得梁木插入殿牆裏。
1KGS|6|7|殿是用山中鑿成的石頭建的，所以建殿的時候，鎚子、斧子和別樣鐵器的響聲都沒有聽見。
1KGS|6|8|在殿右邊當中的廂房有門，可以從螺旋梯上到中層，再從中層上到第三層。
1KGS|6|9|所羅門 完成殿的建造。他用香柏木作梁木和橫板，遮蓋殿頂。
1KGS|6|10|靠著整個殿所造的廂房，每層高五肘，香柏木的梁板擱在殿的牆坎上。
1KGS|6|11|耶和華的話臨到 所羅門 ，說：
1KGS|6|12|「論到你所建的這殿，你若遵行我的律例，謹守我的典章，遵從我的一切誡命，行在其中，我必向你應驗我所應許你父親 大衛 的話。
1KGS|6|13|我必住在 以色列 人中間，並不丟棄我的百姓 以色列 。」
1KGS|6|14|所羅門 完成殿的建造。
1KGS|6|15|他用香柏木板建造殿的內牆，從殿的地到牆頂 都貼上木板，又用松木板鋪地。
1KGS|6|16|他在殿的後部建了一間內殿，長二十肘，從地到牆 用香柏木板，作為至聖所。
1KGS|6|17|殿，就在內殿的前面 ，長四十肘。
1KGS|6|18|殿裏一點石頭都不顯露，一概用香柏木遮蔽；香柏木上刻著野瓜和綻開的花。
1KGS|6|19|他在殿的中間預備內殿，在那裏安放耶和華的約櫃。
1KGS|6|20|內殿 長二十肘，寬二十肘，高二十肘，都貼上純金。他又用香柏木做壇。
1KGS|6|21|所羅門 用純金貼殿內，又用金鏈子掛在內殿前，內殿也貼上金子。
1KGS|6|22|整個殿都貼上金子，直到貼滿；內殿前的整個壇，也都包上金子。
1KGS|6|23|他在內殿裏用橄欖木做兩個基路伯，各高十肘。
1KGS|6|24|這基路伯的一個翅膀長五肘，另一個翅膀長五肘，從一個翅膀尖到另一個翅膀尖共有十肘；
1KGS|6|25|第二個基路伯也是十肘；兩個基路伯的尺寸、形狀都一樣。
1KGS|6|26|這一個基路伯高十肘，第二個基路伯也是如此。
1KGS|6|27|他把兩個基路伯安在內殿中間。基路伯的翅膀是張開的，這基路伯的一個翅膀挨著這邊的牆，第二個基路伯的一個翅膀挨著那邊的牆，向內的兩個翅膀在殿中間彼此相接。
1KGS|6|28|二基路伯都包上金子。
1KGS|6|29|殿周圍的牆上全都刻著基路伯、棕樹和綻開的花，內外都是如此。
1KGS|6|30|殿的地板都貼上金子，內外都是如此。
1KGS|6|31|他用橄欖木製造內殿的入口、門楣和五邊形的門柱。
1KGS|6|32|在橄欖木做的兩門扇上刻著基路伯、棕樹和綻開的花，都貼上金子。基路伯和棕樹上也灑上金子。
1KGS|6|33|他又為外殿的入口，用橄欖木製造門柱，是四邊形的。
1KGS|6|34|他用松木做兩扇門。這一扇有兩葉摺疊，第二扇也有兩葉 摺疊。
1KGS|6|35|上面刻著基路伯、棕樹和綻開的花，雕刻物都均勻地貼上金子。
1KGS|6|36|他又用三層鑿成的石頭、香柏木一層建造內院。
1KGS|6|37|所羅門 在位第四年西弗月，立了耶和華殿的根基。
1KGS|6|38|到十一年布勒月，就是八月，殿和一切屬殿的都按著樣式造成。他建殿共用了七年。
1KGS|7|1|所羅門 為自己建造宮殿，十三年方才建成整座宮殿。
1KGS|7|2|他建造 黎巴嫩林宮 ，長一百肘，寬五十肘，高三十肘，有四行香柏木柱，柱上有香柏木橫梁；
1KGS|7|3|廂房以上覆蓋著香柏木，在四十五根柱子之上，每行十五根。
1KGS|7|4|窗戶有三排，三排的窗與窗相對。
1KGS|7|5|所有的門和門柱都有四方形的框，共有三行，彼此相對。
1KGS|7|6|他建造有柱子的廳，長五十肘，寬三十肘。在這前面有走廊，前面有柱子和頂蓋 。
1KGS|7|7|他又建造一個有座位的廳，就是審判廳，他在那裏審判；這廳的地板從這邊到那邊都鋪上香柏木。
1KGS|7|8|廳後面的院內有 所羅門 自己住的宮殿，都用同樣的建造方式。 所羅門 又為所娶法老的女兒建造一座宮，建造方式與這廳一樣。
1KGS|7|9|建造這一切所用的石頭都是貴重的，按著尺寸鑿成，用鋸子裏外鋸齊；從根基直到房檐，從外頭直到大院，都是如此。
1KGS|7|10|根基是貴重的大石頭，有長十肘的，有長八肘的；
1KGS|7|11|上面有香柏木和按著尺寸鑿成的貴重石頭。
1KGS|7|12|大院周圍有鑿成的石頭三層、香柏木板一層，都照耶和華殿的內院和殿的走廊的樣式。
1KGS|7|13|所羅門 王派人從 推羅 把 戶蘭 接來。
1KGS|7|14|他是 拿弗他利 支派中一個寡婦的兒子，父親是 推羅 人，是作銅匠的。 戶蘭 滿有智慧、聰明、技能，善作各樣的銅器。他來到 所羅門 王那裏，為王做一切的工。
1KGS|7|15|戶蘭 製造兩根銅柱，一根高十八肘，第二根柱子用繩子量，周圍是十二肘 ；
1KGS|7|16|他做了兩個柱頂安在柱上，是用銅鑄造的，一個柱頂高五肘，第二個柱頂也高五肘。
1KGS|7|17|柱子頂上有裝飾的網子和編成的鏈子，一個柱頂有七個，第二個柱頂也有七個。
1KGS|7|18|他做了柱子 ，第一根柱子的柱頂上，周圍有兩行網子在柱子 上面遮蓋柱頂，第二根柱頂也是這樣做。
1KGS|7|19|走廊柱子頂上的柱頂高四肘，刻著百合花。
1KGS|7|20|兩根柱子上面有柱頂，柱頂靠近網子的圓凸面上，有石榴的行列環繞著，共二百個，第二個柱頂也是如此。
1KGS|7|21|他把兩根柱子立在殿的走廊前：右邊立一根，起名叫 雅斤 ；左邊立一根，起名叫 波阿斯 。
1KGS|7|22|柱頂上刻著百合花。這樣，柱子的工程就完畢了。
1KGS|7|23|他又鑄一個銅海，周圍是圓的，直徑十肘，高五肘，用繩子量周圍是三十肘。
1KGS|7|24|銅海邊緣下面的周圍有野瓜的形狀，每肘十個，共兩行，繞著銅海，是造銅海的時候鑄上去的。
1KGS|7|25|銅海安在十二頭銅牛上：三頭向北，三頭向西，三頭向南，三頭向東。銅海安在牛上，牛尾都向內。
1KGS|7|26|銅海厚一掌，邊如杯邊，像百合花，容量是二千罷特。
1KGS|7|27|他用銅製造十個盆座，每座長四肘，寬四肘，高三肘。
1KGS|7|28|銅座的造法是這樣：周圍各有嵌邊，嵌邊裝在框架中。
1KGS|7|29|裝在框架中的嵌邊上有獅子和牛，以及基路伯。框架上有小座，獅子和牛的上面和下面有錘成的花紋浮雕。
1KGS|7|30|每座有四個銅輪和銅軸，它有四個支架在盆以下，這些支架是鑄成的，各邊都有花紋。
1KGS|7|31|它的口在柱頂裏，向上高一肘，口是圓的，做法如座一樣，直徑是一肘半，口上也有雕工。嵌邊是方形的，不是圓的。
1KGS|7|32|四個輪子在嵌邊以下，輪軸與座相連，每輪高一肘半。
1KGS|7|33|輪的樣式如同車的輪子；軸、輞、輻、轂都是鑄成的。
1KGS|7|34|每個座四邊有四個盆形的支架，這些支架是與座從一整塊鑄成的。
1KGS|7|35|座頂有圓架，高半肘；座頂有支柱和嵌邊，是與座從一整塊鑄成的。
1KGS|7|36|他在支柱和嵌邊上，每個空處刻上基路伯、獅子和棕樹，周圍有花紋。
1KGS|7|37|他按照這樣的做法造了十個盆座，它們的鑄法、尺寸、樣式全都相同。
1KGS|7|38|他又造十個銅盆，每盆的容量四十罷特，直徑四肘。在十個座上，每座安設一盆。
1KGS|7|39|他把五個安置在殿的右邊，五個安置在殿的左邊，又把銅海安置在殿的右旁，在東南邊。
1KGS|7|40|戶蘭 又造了盆、鏟子和盤子。這樣， 戶蘭 為 所羅門 王做完了耶和華殿一切的工：
1KGS|7|41|兩根柱子和柱子頂上兩個如碗的柱頂，以及蓋著如碗柱頂的兩個網子；
1KGS|7|42|四百個石榴，安在兩個網子上，每網兩行石榴，蓋著柱子上面兩個如碗的柱頂；
1KGS|7|43|十個盆座和其上的十個盆；
1KGS|7|44|銅海和其下的十二頭牛；
1KGS|7|45|盆、鏟子、盤子。 戶蘭 給 所羅門 王為耶和華殿造的這一切器皿都是用光亮的銅，
1KGS|7|46|是王在 約旦 平原、 疏割 和 撒拉但 中間的泥巴地鑄成的。
1KGS|7|47|所羅門 允許這一切器皿不過秤，因為所用的銅太多，重量無法計算。
1KGS|7|48|所羅門 又為耶和華的殿造了各樣的器皿：金壇和獻供餅的金供桌；
1KGS|7|49|內殿前的純金燈臺，右邊五個，左邊五個，以及其上的花、燈盞、燈剪，都是金的；
1KGS|7|50|純金的杯、鉗子、盤子、勺子 、火盆，以及聖殿的最裏面，就是至聖所的門樞和外殿的門樞，都是金的。
1KGS|7|51|所羅門 王做完了耶和華殿一切的工，就把他父親 大衛 分別為聖的金銀和器皿都帶來，放在耶和華殿的庫房裏。
1KGS|8|1|那時， 所羅門 召集 以色列 的長老、各支派的領袖和 以色列 人的族長到 耶路撒冷 ， 所羅門 王那裏，要把耶和華的約櫃從 大衛城 ，就是 錫安 ，接上來。
1KGS|8|2|以他念月，就是七月，在節期時，所有的 以色列 人都聚集到 所羅門 王那裏。
1KGS|8|3|以色列 眾長老一來到，祭司就抬起約櫃。
1KGS|8|4|祭司和 利未 人將耶和華的約櫃請上來，又把會幕和會幕一切的聖器皿都帶上來。
1KGS|8|5|所羅門 王和聚集到他那裏的 以色列 全會眾一同在約櫃前獻牛羊為祭，多得不可勝數，無法計算。
1KGS|8|6|祭司將耶和華的約櫃請進內殿，就是至聖所，安置在兩個基路伯的翅膀底下約櫃的地方。
1KGS|8|7|基路伯張開翅膀在約櫃上面的地方，從上面遮住約櫃和抬櫃的槓。
1KGS|8|8|這槓很長，從內殿前的聖所可以看見槓頭，從外面卻看不見。這槓直到今日還在那裏。
1KGS|8|9|約櫃裏沒有別的，只有兩塊石版，就是 以色列 人出 埃及 地，耶和華與他們立約的時候， 摩西 在 何烈山 放在那裏的。
1KGS|8|10|祭司從聖所出來的時候，有雲充滿耶和華的殿，
1KGS|8|11|祭司因雲彩的緣故不能站立供職，因為耶和華的榮光充滿了耶和華的殿。
1KGS|8|12|那時， 所羅門 說： 「耶和華曾說要住在幽暗之處 。
1KGS|8|13|我的確為你建了一座雄偉的殿宇， 作為你永遠居住的地方。」
1KGS|8|14|王轉過臉來為 以色列 全會眾祝福， 以色列 全會眾都站立。
1KGS|8|15|所羅門 說：「耶和華－ 以色列 的上帝是應當稱頌的！因他親口向我父 大衛 應許的，也親手成就了；他曾說：
1KGS|8|16|『自從那日我領我百姓 以色列 出 埃及 以來，我未曾在 以色列 各支派中選擇一城，在那裏為我的名建造殿宇，但我揀選 大衛 治理我的百姓 以色列 。』
1KGS|8|17|我父 大衛 的心意是要為耶和華－ 以色列 上帝的名建殿。
1KGS|8|18|耶和華卻對我父 大衛 說：『你有心為我的名建殿，這心意是好的；
1KGS|8|19|但你不可建殿，惟有你親生的兒子才可為我的名建殿。』
1KGS|8|20|現在耶和華實現了他所應許的話，使我接續我父 大衛 坐 以色列 的王位，正如耶和華所說的，我也為耶和華－ 以色列 上帝的名建造了這殿。
1KGS|8|21|我也在那裏為約櫃預備一處。約櫃那裏有耶和華的約，就是他領我們列祖出 埃及 地的時候，與他們所立的約。」
1KGS|8|22|所羅門 當著 以色列 全會眾，站在耶和華的壇前，向天舉手，
1KGS|8|23|說：「耶和華－ 以色列 的上帝啊，天上地下沒有神明可與你相比！你向那些盡心行在你面前的僕人守約施慈愛，
1KGS|8|24|這約是你向你僕人 大衛 守的，是你應許他的。你親口應許，親手成就，正如今日一樣。
1KGS|8|25|耶和華－ 以色列 的上帝啊，你向你僕人我父 大衛 應許說：『你的子孫若謹慎自己的行為，在我面前行事像你所行的一樣，就不斷有人在我面前坐 以色列 的王位。』現在求你信守這話。
1KGS|8|26|以色列 的上帝啊，現在求你成就向你僕人我父 大衛 所應許的話。
1KGS|8|27|「上帝果真住在地上嗎？看哪，天和天上的天尚且不足容納你，何況我所建的這殿呢？
1KGS|8|28|惟求耶和華－我的上帝垂顧僕人的禱告祈求，俯聽僕人今日在你面前的祈禱呼求。
1KGS|8|29|願你的眼目晝夜看顧這殿，就是你說要作為你名的居所；求你垂聽禱告，你僕人向此處的禱告。
1KGS|8|30|你僕人和你百姓 以色列 向此處祈禱的時候，求你在你天上的居所垂聽，垂聽而赦免。
1KGS|8|31|「人若得罪鄰舍，有人強迫他，要他起誓，他來到這殿，在你的壇前起誓，
1KGS|8|32|求你在天上垂聽、處理，向你的僕人施行審判，定惡人有罪，照他所行的報應在他頭上；定義人為義，照他的義賞賜他。
1KGS|8|33|「你的百姓 以色列 若得罪你，敗在仇敵面前，卻又歸向你，宣認你的名，在這殿裏向你祈求禱告，
1KGS|8|34|求你在天上垂聽，赦免你百姓 以色列 的罪，使他們歸回你賜給他們列祖的地。
1KGS|8|35|「你的百姓若得罪了你，你使天閉塞不下雨；他們若向此處禱告，宣認你的名，因你的懲罰而離開他們的罪，
1KGS|8|36|求你在天上垂聽，赦免你僕人你百姓 以色列 的罪，將當行的善道教導他們，並降雨在你的地，就是你賜給你百姓為業之地。
1KGS|8|37|「這地若有饑荒、瘟疫、焚風 、霉爛、蝗蟲、螞蚱，或有仇敵圍困這地的 城門，無論遭遇甚麼災禍疾病，
1KGS|8|38|你的百姓 以色列 ，或眾人或一人，內心知道有禍，向這殿舉手，無論祈求甚麼，禱告甚麼，
1KGS|8|39|求你在天上你的居所垂聽、赦免、處理。因為你知道人心，惟有你知道世人的心，求你照各人所行的一切待他們，
1KGS|8|40|使他們在你賜給我們列祖的土地上一生一世敬畏你。
1KGS|8|41|「論到不屬你百姓 以色列 的外邦人，若為你的名從遠方而來，
1KGS|8|42|他們因聽見你的大名和大能的手，以及伸出來的膀臂，來向這殿禱告，
1KGS|8|43|求你在天上你的居所垂聽，照著外邦人向你所求的一切而行，使地上萬民都認識你的名，敬畏你，像你的百姓 以色列 一樣，又使他們知道我所建造的是稱為你名下的殿。
1KGS|8|44|「你的百姓若奉你的派遣出去，無論往何處與仇敵爭戰，他們若向耶和華所選擇的城，以及我為你名所建造的這殿禱告，
1KGS|8|45|求你在天上垂聽他們的禱告祈求，為他們伸張正義。
1KGS|8|46|「你的百姓若得罪你，因為沒有人不犯罪，你向他們發怒，把他們交在仇敵面前，擄他們的人把他們帶到仇敵之地，或遠或近，
1KGS|8|47|他們若在被擄之地那裏回心轉意，在擄掠者之地悔改，向你懇求說：『我們有罪了，我們悖逆了，我們作惡了』；
1KGS|8|48|他們若在擄他們的仇敵之地盡心盡性歸向你，又向自己的地，就是你賜給他們列祖的地和你所選擇的城，以及我為你名所建造的這殿禱告，
1KGS|8|49|求你在天上你的居所垂聽他們的禱告祈求，為他們伸張正義，
1KGS|8|50|饒恕得罪你的子民，赦免他們向你所犯一切的過犯，使他們在擄他們的人面前蒙憐憫。
1KGS|8|51|因為他們是你的子民，你的產業，是你從 埃及 ，從鐵爐中領出來的。
1KGS|8|52|願你的眼目看顧僕人和你百姓 以色列 的祈求；他們無論何時向你呼求，願你垂聽。
1KGS|8|53|主耶和華啊，你將他們從地上萬民中分別出來作你的產業，是照著你領我們列祖出 埃及 的時候，藉你僕人 摩西 所應許的。」
1KGS|8|54|所羅門 在耶和華的壇前屈膝跪著，向天舉手；他在耶和華面前禱告祈求完畢的時候，就起來，
1KGS|8|55|站著，大聲為 以色列 全會眾祝福，說：
1KGS|8|56|「耶和華是應當稱頌的！因為他照著一切所應許的賜平安給他的百姓 以色列 ，凡藉他僕人 摩西 應許賜福的話，一句都沒有落空。
1KGS|8|57|願耶和華－我們的上帝與我們同在，像與我們列祖同在一樣，不撇下我們，不丟棄我們，
1KGS|8|58|使我們的心歸向他，遵行他一切的道，謹守他吩咐我們列祖的誡命、律例、典章。
1KGS|8|59|願我在耶和華面前祈求的這些話，晝夜靠近耶和華－我們的上帝，好讓他每日為他僕人和他百姓 以色列 伸張正義，
1KGS|8|60|使地上的萬民都知道惟獨耶和華是上帝，沒有別的了。
1KGS|8|61|所以你們當向耶和華－我們的上帝存純正的心，遵行他的律例，謹守他的誡命，如同今日一樣。」
1KGS|8|62|王和全 以色列 一同在耶和華面前獻祭。
1KGS|8|63|所羅門 向耶和華獻平安祭，二萬二千頭牛，十二萬隻羊。這樣，王和全 以色列 為耶和華的殿行了奉獻之禮。
1KGS|8|64|當日，王因耶和華殿前的銅壇太小，容不下燔祭、素祭和平安祭牲的脂肪，就將耶和華殿前院子的中間分別為聖，在那裏獻燔祭、素祭和平安祭牲的脂肪。
1KGS|8|65|那時 所羅門 守節，從 哈馬口 直到 埃及 溪谷的 以色列 眾人都與他同在一起，成了一個盛大的會，在耶和華－我們的上帝面前七日又七日，共十四日。
1KGS|8|66|第八日，王遣散百姓；他們都為王祝福。他們為耶和華向他僕人 大衛 和他百姓 以色列 所施的一切恩惠都心中喜樂，愉快地各回自己的帳棚去了。
1KGS|9|1|所羅門 建造耶和華的殿和王宮，以及一切所想要建造的都完畢了，
1KGS|9|2|耶和華第二次向 所羅門 顯現，如先前在 基遍 向他顯現一樣。
1KGS|9|3|耶和華對他說：「我已聽了你在我面前的禱告和祈求，將你所建的這殿分別為聖，使我的名永遠立在那裏；我的眼、我的心也必時常在那裏。
1KGS|9|4|你若以純正的心和正直行在我面前，效法你父 大衛 所行的，遵行我一切所吩咐你的，謹守我的律例典章，
1KGS|9|5|我就必堅固你在 以色列 國度的王位，直到永遠，正如我應許你父 大衛 說：『你的子孫必不斷有人坐 以色列 的王位。』
1KGS|9|6|倘若你們和你們的子孫轉去不跟從我，不守我擺在你們面前的誡命律例，去事奉別神，敬拜它們，
1KGS|9|7|我就必把 以色列 從我賜給他們的地上剪除，也必從我面前捨棄那為我名所分別為聖的殿，使 以色列 在萬民中成為笑柄，被人譏誚。
1KGS|9|8|這殿雖然崇高 ，將來凡經過的人必驚訝，嗤笑，說：『耶和華為何向這地和這殿如此行呢？』
1KGS|9|9|人必說：『因為此地的人離棄領他們祖先出 埃及 地的耶和華－他們的上帝，去親近別神，敬拜事奉它們，所以耶和華使這一切災禍臨到他們。』」
1KGS|9|10|所羅門 建造耶和華殿和王宮這兩座殿宇，用了二十年才完成。
1KGS|9|11|推羅 王 希蘭 曾照 所羅門 所要的資助他香柏木、松木和金子， 所羅門 王就把 加利利 地的二十座城給了 希蘭 。
1KGS|9|12|希蘭 從 推羅 出來，察看 所羅門 給他的城鎮，看不順眼，
1KGS|9|13|就說：「我兄啊，你給我的是甚麼城鎮呢？」他就給這些城鎮起名叫 迦步勒 地，直到今日。
1KGS|9|14|希蘭 曾給 所羅門 一百二十他連得金子。
1KGS|9|15|所羅門 王挑取服勞役的工人，為要建造耶和華的殿、自己的宮、 米羅 、 耶路撒冷 的城牆、 夏瑣 、 米吉多 和 基色 。
1KGS|9|16|先前 埃及 王法老上來攻取 基色 ，用火焚燒，殺了城內居住的 迦南 人，把城賜給他的女兒，就是 所羅門 的妻子，作為嫁妝。
1KGS|9|17|所羅門 建造 基色 、 下伯‧和崙 、
1KGS|9|18|巴拉 ，和位於境內曠野的 達莫 。
1KGS|9|19|所羅門 建造一切的儲貨城、戰車城、戰馬城，以及他所想要建造的，在 耶路撒冷 、 黎巴嫩 和自己治理全國中的一切建設。
1KGS|9|20|至於所有剩下的百姓，不屬 以色列 人的 亞摩利 人、 赫 人、 比利洗 人、 希未 人、 耶布斯 人，
1KGS|9|21|那些 以色列 人在當地不能滅盡的人， 所羅門 徵召他們剩下的後代作服勞役的奴僕，直到今日。
1KGS|9|22|惟有 以色列 人， 所羅門 不使他們作奴僕，而是作他的戰士、臣僕、官長、軍官、戰車長、騎兵長。
1KGS|9|23|這些是 所羅門 工程的五百五十個監工，他們在百姓中監管作工的人。
1KGS|9|24|法老的女兒從 大衛城 上到 所羅門 為她建造的宮裏。那時， 所羅門 才建造 米羅 。
1KGS|9|25|所羅門 每年三次在他為耶和華所築的壇上獻燔祭和平安祭，又在耶和華面前的壇上燒香。這樣，他完成了建殿。
1KGS|9|26|所羅門 王在 以東 地 紅海 邊，靠近 以祿 的 以旬‧迦別 製造船隻。
1KGS|9|27|希蘭 派他的僕人，就是熟悉航海的船員，與 所羅門 的僕人一同坐船航海。
1KGS|9|28|他們到了 俄斐 ，從那裏得了四百二十他連得金子，運到 所羅門 王那裏。
1KGS|10|1|示巴 女王聽見 所羅門 因耶和華的名所得的名聲，就來要用難題考問 所羅門 。
1KGS|10|2|她帶著很多的隨從來到 耶路撒冷 ，有駱駝馱著香料、極多金子和寶石。她來到 所羅門 那裏，向他提出心中所有的問題。
1KGS|10|3|所羅門 回答了她所有的問題，沒有一個問題太難，王不能向她解答的。
1KGS|10|4|示巴 女王看見 所羅門 一切的智慧，和他所建造的宮殿，
1KGS|10|5|席上的食物，坐著的群臣，侍立的僕人，他們的服裝，和他的司酒長，以及他在耶和華殿裏所獻的燔祭 ，就詫異得神不守舍。
1KGS|10|6|她對王說：「我在本國所聽到的話，論到你的事和你的智慧是真的！
1KGS|10|7|我本來不信那些話，及至我來親眼看見了，看哪，人所告訴我的還不到一半，你的智慧和你的福分超過我所聽見的傳聞。
1KGS|10|8|你的人 是有福的！你這些僕人常侍立在你面前、聽你智慧的話是有福的！
1KGS|10|9|耶和華－你的上帝是應當稱頌的！他喜愛你，使你坐 以色列 的王位，因為他永遠愛 以色列 ，所以立你作王，使你秉公行義。」
1KGS|10|10|於是， 示巴 女王把一百二十他連得金子、極多的香料和寶石送給 所羅門 王；送來的香料，從來沒有像 示巴 女王送給他的那麼多。
1KGS|10|11|希蘭 的船隻也從 俄斐 運了金子來，又從 俄斐 運了許多檀香木和寶石來。
1KGS|10|12|王用檀香木為耶和華的殿和王宮做欄杆，又為歌唱的人做琴瑟。以後再沒有這樣的檀香木運進來，也再沒有人見過，直到如今。
1KGS|10|13|所羅門 王除了照自己的厚意餽贈 示巴 女王之外，凡她所提出的一切要求， 所羅門 王都送給她。於是女王和她臣僕轉回，到本國去了。
1KGS|10|14|所羅門 每年所得的金子，重六百六十六他連得；
1KGS|10|15|另外還有來自商人 和做生意的商品，以及 阿拉伯 諸王和各地省長的。
1KGS|10|16|所羅門 王用錘出來的金子打成二百面盾牌，每面盾牌用六百舍客勒金子；
1KGS|10|17|又用錘出來的金子打成三百面小盾牌，每面小盾牌用三彌那金子。王把它們放在 黎巴嫩林宮 裏。
1KGS|10|18|王又製造一個大的象牙寶座，包上純金。
1KGS|10|19|寶座有六層臺階，座的後背是圓的，座位之處兩旁有扶手，靠近扶手有兩隻獅子站立。
1KGS|10|20|六層臺階上有十二隻獅子站立，分站左邊和右邊；任何國度都沒有這樣做的。
1KGS|10|21|所羅門 王一切的飲器都是金的， 黎巴嫩林宮 裏所有的器皿都是純金的。在 所羅門 的日子，銀子算不了甚麼。
1KGS|10|22|王有 他施 船隻與 希蘭 的船隻一同航海， 他施 船隻每三年一次把金、銀、象牙、猿猴、孔雀 運回來。
1KGS|10|23|所羅門 王的財寶與智慧勝過地上的眾王。
1KGS|10|24|全地都求見 所羅門 的面，要聽上帝放在他心裏的智慧。
1KGS|10|25|他們各帶貢物，就是銀器、金器、衣服、兵器、香料、馬、騾子，每年都有一定的數量。
1KGS|10|26|所羅門 聚集戰車騎兵；他有一千四百輛戰車，一萬二千名騎兵，安置在屯車城，在 耶路撒冷 的王那裏。
1KGS|10|27|王在 耶路撒冷 使銀子多如石頭，香柏木多如 謝非拉 的桑樹。
1KGS|10|28|所羅門 的馬是從 埃及 和 科威 運來的，是王的商人按著定價從 科威 買來的。
1KGS|10|29|從 埃及 進口的戰車，每輛六百舍客勒銀子，馬每匹一百五十舍客勒； 赫 人眾王和 亞蘭 諸王的戰車和馬，也是經由他們的手出口的。
1KGS|11|1|所羅門 王在法老的女兒之外，又寵愛許多外邦女子，就是 摩押 女子、 亞捫 女子、 以東 女子、 西頓 女子、 赫 人女子。
1KGS|11|2|論到這些國的人，耶和華曾吩咐 以色列 人說：「你們不可跟他們通婚，他們也不可跟你們在一起，因為他們一定會誘惑你們的心去隨從他們的神明。」 所羅門 卻為了愛，緊緊跟從他們。
1KGS|11|3|所羅門 娶七百個公主，三百個妃嬪。這些妻妾誘惑他的心。
1KGS|11|4|所羅門 年老的時候，他的妻妾誘惑他的心去隨從別神，不像他父親 大衛 以純正的心順服耶和華－他的上帝。
1KGS|11|5|所羅門 隨從 西頓 人的女神 亞斯她錄 和 亞捫 人可憎的 米勒公 。
1KGS|11|6|所羅門 行耶和華眼中看為惡的事，不像他父親 大衛 專心順從耶和華。
1KGS|11|7|那時， 所羅門 為 摩押 可憎的 基抹 和 亞捫 人可憎的 摩洛 ，在 耶路撒冷 對面的山上建造丘壇。
1KGS|11|8|他為所有的妻妾，就是那些向自己神明燒香獻祭的外邦女子，也是這樣做。
1KGS|11|9|耶和華向 所羅門 發怒，因為他的心偏離了向他顯現兩次的耶和華－ 以色列 的上帝。
1KGS|11|10|耶和華曾吩咐他這件事，不可隨從別神，他卻沒有遵守耶和華所吩咐的。
1KGS|11|11|所以耶和華對他說：「你既然是這樣，不遵守我所吩咐你守的約和律例，我必定把國度撕裂離開你，將它賜給你的大臣。
1KGS|11|12|然而，因你父親 大衛 的緣故，我不在你的日子行這事，而要從你兒子的手中撕裂這國。
1KGS|11|13|只是我不撕裂全國，卻要因我僕人 大衛 和我所選擇的 耶路撒冷 ，保留一個支派給你的兒子。」
1KGS|11|14|耶和華使 以東 人 哈達 興起，作 所羅門 的敵人；他是 以東 王的後裔。
1KGS|11|15|大衛 在 以東 的時候， 約押 元帥上去埋葬陣亡的人，殺了 以東 所有的男丁。
1KGS|11|16|約押 和 以色列 眾人在 以東 住了六個月，直到把 以東 的男丁盡都剪除。
1KGS|11|17|那時 哈達 還是幼童；他和他父親的臣僕，以及幾個 以東 人逃往 埃及 。
1KGS|11|18|他們從 米甸 起行，到了 巴蘭 ，再從 巴蘭 帶著幾個人來到 埃及 ，到 埃及 王法老那裏。法老給他房屋，吩咐給他糧食，又把地賜給他。
1KGS|11|19|哈達 在法老眼前大蒙恩寵，法老就把王后 答比匿 的妹妹嫁給他。
1KGS|11|20|答比匿 的妹妹給 哈達 生了一個兒子，叫 基努拔 。 答比匿 使 基努拔 在法老的宮裏斷奶， 基努拔 就與法老的眾子一同住在法老的宮裏。
1KGS|11|21|哈達 在 埃及 聽見 大衛 與他祖先同睡， 約押 元帥也死了，就對法老說：「請你讓我走，我要回本國去。」
1KGS|11|22|法老對他說：「你在我這裏有甚麼缺乏？看哪，你竟想要回你本國去！」他說：「我沒有缺乏甚麼，只是懇求王准我回去。」
1KGS|11|23|上帝又使 以利亞大 的兒子 利遜 興起，作 所羅門 的敵人。他曾逃避主人 瑣巴 王 哈大底謝 。
1KGS|11|24|大衛 擊殺 瑣巴 人的時候， 利遜 召集了一群人，自己作他們的領袖。他們往 大馬士革 ，住在那裏，在 大馬士革 建立王國。
1KGS|11|25|所羅門 活著的時候，除了 哈達 為患之外， 利遜 也作 以色列 的敵人。他憎恨 以色列 ，作了 亞蘭 人的王。
1KGS|11|26|尼八 的兒子 耶羅波安 也舉起手來攻擊王。他是 所羅門 的臣僕， 以法蓮 支派的 洗利達 人；他母親是個寡婦，名叫 洗魯阿 。
1KGS|11|27|他舉手攻擊王是因先前 所羅門 建造 米羅 ，修補他父親 大衛城 缺口的這件事。
1KGS|11|28|耶羅波安 是個大有才能的人。 所羅門 見這青年殷勤，就派他監管 約瑟 家所有服勞役的工人。
1KGS|11|29|那時， 耶羅波安 出了 耶路撒冷 ， 示羅 人 亞希雅 先知在路上遇見他； 亞希雅 身上穿著一件新衣。田野中只有他們二人，沒有其他的人。
1KGS|11|30|亞希雅 拿起穿在自己身上的新衣，把它撕成十二片，
1KGS|11|31|對 耶羅波安 說：「你可以拿十片。耶和華－ 以色列 的上帝如此說：『看哪，我必從 所羅門 手裏撕裂這國，把十個支派賜給你。
1KGS|11|32|我因我僕人 大衛 和我在 以色列 眾支派中所選擇的 耶路撒冷城 的緣故，仍為 所羅門 留一個支派。
1KGS|11|33|因為他們 離棄我，敬拜 西頓 人的女神 亞斯她錄 、 摩押 的神明 基抹 和 亞捫 人的神明 米勒公 ，沒有像他父親 大衛 一樣遵從我的道，行我眼中看為正的事，守我的律例典章。
1KGS|11|34|但我不從他手裏奪走整個國家，卻使他在活著的日子作君王，是因我所揀選的僕人 大衛 遵守我的誡命律例。
1KGS|11|35|我必從他兒子手裏將王國奪走，賜給你十個支派，
1KGS|11|36|只留一個支派給他的兒子，使我僕人 大衛 在我所選擇立我名的 耶路撒冷城 那裏，在我面前常有燈光。
1KGS|11|37|我選你，使你照你心裏一切所願的作王，成為 以色列 的王。
1KGS|11|38|你若聽從我一切所吩咐你的，遵行我的道，行我眼中看為正的事，謹守我的律例誡命，像我僕人 大衛 所行的，我就與你同在，為你立堅固的家，像我為 大衛 所立的一樣，將 以色列 賜給你。
1KGS|11|39|我必因這事使 大衛 的後裔遭受患難，但不是永遠的。』」
1KGS|11|40|所羅門 想要殺 耶羅波安 ， 耶羅波安 起身逃往 埃及 。他到了 埃及 王 示撒 那裏，就住在 埃及 ，直到 所羅門 死了。
1KGS|11|41|所羅門 其餘的事，凡他所做的和他的智慧，不都寫在《所羅門記》上嗎？
1KGS|11|42|所羅門 在 耶路撒冷 作全 以色列 的王四十年。
1KGS|11|43|所羅門 與他祖先同睡，葬在他父親 大衛 的城裏，他兒子 羅波安 接續他作王。
1KGS|12|1|羅波安 往 示劍 去，因 以色列 眾人都到了 示劍 ，要立他作王。
1KGS|12|2|尼八 的兒子 耶羅波安 先前躲避 所羅門 王，逃往 埃及 ，住在那裏。他還在 埃及 ，聽見了這事 ，
1KGS|12|3|以色列 人派人去請他來。 耶羅波安 就和 以色列 全會眾來，與 羅波安 談話，說：
1KGS|12|4|「你父親使我們負重軛，現在求你減輕你父親所加給我們的苦工和重軛，我們就服事你。」
1KGS|12|5|羅波安 對他們說：「你們走吧，過三天再來見我。」百姓就走了。
1KGS|12|6|羅波安 的父親 所羅門 在世的日子，有侍立在他面前的長者， 羅波安 王和他們商議，說：「你們出個主意，好把話帶回給這百姓。」
1KGS|12|7|他們對他說：「現在王若像僕人一樣服事這百姓，用好話回覆他們，他們就永遠作王的僕人了。」
1KGS|12|8|王不採納長者給他出的主意，卻和那些與他一同長大、在他面前侍立的年輕人商議。
1KGS|12|9|他對他們說：「這百姓對我說：『你父親使我們負重軛，求你減輕一些。』你們出個甚麼主意，我們好把話帶回給他們。」
1KGS|12|10|那些與他一同長大的年輕人對他說：「這百姓對王說：『你父親使我們負重軛，求你給我們減輕一些。』王要對他們如此說：『我的小指頭比我父親的腰還粗呢！
1KGS|12|11|我父親使你們負重軛，現在我必使你們負更重的軛！我父親用鞭子懲罰你們，我要用蠍子懲罰你們！』」
1KGS|12|12|耶羅波安 和眾百姓遵照王所說「你們第三天再來見我」的話，第三天來到 羅波安 那裏。
1KGS|12|13|王嚴厲地回答百姓，不採納長者給他出的主意。
1KGS|12|14|他照著年輕人所出的主意對他們說：「我父親使你們負重軛，我必使你們負更重的軛！我父親用鞭子懲罰你們，我卻要用蠍子懲罰你們！」
1KGS|12|15|王不依從百姓，因這事件是出於耶和華，為要應驗耶和華藉 示羅 人 亞希雅 對 尼八 的兒子 耶羅波安 所說的話。
1KGS|12|16|以色列 眾人見王不依從他們，百姓就回話給王，說： 「我們在 大衛 中有甚麼份呢？ 我們在 耶西 的兒子中沒有產業！ 以色列 啊，回你的帳棚去吧！ 大衛 啊，現在你顧自己的家吧！」 於是， 以色列 人都回自己的帳棚去了；
1KGS|12|17|至於住 猶大 城鎮的 以色列 人， 羅波安 仍作他們的王。
1KGS|12|18|羅波安 王派監管勞役的 亞多蘭 去， 以色列 眾人用石頭打他，他就死了。 羅波安 王急忙上車，逃回 耶路撒冷 去了。
1KGS|12|19|這樣， 以色列 背叛 大衛 家，直到今日。
1KGS|12|20|以色列 眾人聽見 耶羅波安 回來了，就派人去請他到會眾那裏，立他作全 以色列 的王。除了 猶大 支派，沒有跟從 大衛 家的。
1KGS|12|21|羅波安 來到 耶路撒冷 ，召集了 猶大 全家和 便雅憫 支派的人共十八萬，都是精選的戰士，要與 以色列 家打仗，好將王國奪回，歸 所羅門 的兒子 羅波安 。
1KGS|12|22|但上帝的話臨到神人 示瑪雅 ，說：
1KGS|12|23|「你去告訴 所羅門 的兒子 猶大 王 羅波安 ， 猶大 和 便雅憫 全家，以及其餘的百姓，說：
1KGS|12|24|『耶和華如此說：你們不可上去與你們的弟兄 以色列 人打仗。你們各自回家去吧！因為這事是出於我。』」眾人就聽從耶和華的話，遵照耶和華的話回去了。
1KGS|12|25|耶羅波安 在 以法蓮 山區建了 示劍 ，住在其中，又從 示劍 出去，建了 毗努伊勒 。
1KGS|12|26|耶羅波安 心裏說：「現在，這國恐怕仍會歸 大衛 家；
1KGS|12|27|這百姓若上 耶路撒冷 去，在耶和華的殿裏獻祭，他們的心必歸向他們的主 猶大 王 羅波安 。他們會殺了我，仍歸 猶大 王 羅波安 。」
1KGS|12|28|耶羅波安 王就籌劃，鑄造了兩個金牛犢，對眾百姓說：「你們上 耶路撒冷 去實在夠久了。 以色列 啊，看哪，這是領你出 埃及 地的神明。」
1KGS|12|29|他把一個安置在 伯特利 ，另一個安置在 但 。
1KGS|12|30|這事使百姓陷入罪裏，因為他們甚至到 但 去拜那牛犢。
1KGS|12|31|耶羅波安 在一些丘壇建神殿，立不屬 利未 人的平民百姓為祭司。
1KGS|12|32|耶羅波安 定八月十五日為節期，像在 猶大 的節期一樣，自己上壇獻祭。他在 伯特利 這樣做，向他所鑄的牛犢獻祭，又把他所立丘壇的祭司安置在 伯特利 。
1KGS|12|33|他在八月十五日，就是他自己心中所定的月份，在 伯特利 上到自己所造的祭壇；他為 以色列 人定了一個節期，親自上壇燒香。
1KGS|13|1|看哪，有一個神人遵照耶和華的話從 猶大 來到 伯特利 。 耶羅波安 正站在壇旁燒香；
1KGS|13|2|神人遵照耶和華的話向壇呼叫，說：「壇哪，壇哪！耶和華如此說：『看哪， 大衛 家必生一個兒子，名叫 約西亞 ，他必將在你上面燒香的丘壇祭司，宰殺在你上面，人的骨頭也必燒在你上面。』」
1KGS|13|3|當日，神人設個預兆，說：「這是耶和華說的預兆：『看哪，這壇必破裂，壇上的灰必傾倒出來。』」
1KGS|13|4|耶羅波安 王聽見神人向 伯特利 的壇呼叫的話，就從壇上伸手，說：「拿住他！」王向神人所伸的手卻萎縮了，不能彎回。
1KGS|13|5|壇也破裂了，壇上的灰傾倒出來，正如神人遵照耶和華的話所設的預兆。
1KGS|13|6|王對神人說：「請你為我禱告，向耶和華－你的上帝懇求恩惠，使我的手復原。」於是神人向耶和華懇求，王的手就復原了，如平常一樣。
1KGS|13|7|王對神人說：「請你跟我回宮，讓你恢復心力，我必給你賞賜。」
1KGS|13|8|神人對王說：「你就是把你一半的王宮給我，我也不跟你進去，也不在這地方吃飯喝水，
1KGS|13|9|因為耶和華的話這樣吩咐我說：『不可吃飯喝水，也不可從你去的原路回來。』」
1KGS|13|10|於是神人從別的路回去，不從他到 伯特利 來的原路回去。
1KGS|13|11|有一個老先知住在 伯特利 ，他的兒子來，把神人當日在 伯特利 所做的一切事和他向王所說的話，都告訴了父親。
1KGS|13|12|父親對他們說：「神人從哪條路去了呢？」他的兒子都看到 從 猶大 來的神人所去的路。
1KGS|13|13|老先知吩咐兒子說：「你們為我備驢。」他們備好了驢，他就騎上，
1KGS|13|14|去追神人，遇見神人坐在橡樹底下，就對他說：「你是不是從 猶大 來的神人？」他說：「是我。」
1KGS|13|15|老先知對他說：「請你跟我一起回家吃飯。」
1KGS|13|16|神人說：「我不能跟你回去，與你同行，也不能在這地方跟你一起吃飯喝水，
1KGS|13|17|因為有耶和華的話吩咐我說：『你在那裏不可吃飯喝水，也不可從你去的原路回來。』」
1KGS|13|18|老先知對他說：「我也是先知，和你一樣。有天使遵照耶和華的話對我說：『你去帶他一同回你的家，給他吃飯喝水。』」老先知在欺騙他。
1KGS|13|19|於是神人跟老先知回去，在他家裏吃飯喝水。
1KGS|13|20|他們坐席的時候，耶和華的話臨到那帶神人回來的先知，
1KGS|13|21|他就對從 猶大 來的神人宣告說：「耶和華如此說：『你既違背耶和華的指示，不遵守耶和華－你上帝的命令，
1KGS|13|22|反倒回來，在耶和華禁止你吃飯喝水的地方吃了飯喝了水，因此你的屍體必不得葬在你祖先的墳墓裏。』」
1KGS|13|23|神人吃喝完了，老先知為他帶回來的先知備驢。
1KGS|13|24|神人就去了，在路上有隻獅子遇見他，把他咬死。他的屍體倒在路上，驢站在屍體旁邊，獅子也站在屍體旁邊。
1KGS|13|25|看哪，有人經過，看見屍體倒在路上，獅子站在屍體旁邊，就來到老先知所住的城裏述說這事。
1KGS|13|26|那帶神人回來的先知聽見了，就說：「這是那違背了耶和華指示的神人，所以耶和華把他交給獅子；獅子撕裂他，咬死他，正如耶和華對他說的話。」
1KGS|13|27|老先知吩咐他兒子說：「你們為我備驢。」他們就備了驢。
1KGS|13|28|他去了，發現神人的屍體倒在路上，驢和獅子站在屍體旁邊，獅子卻沒有吃屍體，也沒有撕裂驢。
1KGS|13|29|老先知把神人的屍體抬起，馱在驢上，帶回自己的城裏，要為他哀哭，為他安葬。
1KGS|13|30|老先知把屍體葬在自己的墳裏，為他哀哭，說：「哀哉！我的弟兄啊！」
1KGS|13|31|安葬之後，老先知對他兒子說：「我死了，你們要把我葬在神人所葬的墳裏，使我的屍骨在他的屍骨旁邊，
1KGS|13|32|因為他遵照耶和華的話，指著 伯特利 的壇和 撒瑪利亞 各城丘壇神殿所宣告的話必定應驗。」
1KGS|13|33|這事以後， 耶羅波安 仍不離開他的惡道，立平民百姓為丘壇的祭司；凡願意的，他都分別為聖，立為丘壇的祭司。
1KGS|13|34|這事使 耶羅波安 的家陷入罪裏，甚至他的家被剪除，從地面上消滅了。
1KGS|14|1|那時， 耶羅波安 的兒子 亞比雅 病了。
1KGS|14|2|耶羅波安 對他的妻子說：「你起來改裝，使人認不出你是 耶羅波安 的妻子。你往 示羅 去，看哪，那裏有先知 亞希雅 ，他曾告訴我說，你必作這百姓的王。
1KGS|14|3|現在你手裏要帶十個餅、幾個薄餅和一瓶蜜到他那裏去，他必告訴你，孩子會怎樣。」
1KGS|14|4|耶羅波安 的妻子就照樣做，起身往 示羅 去，到了 亞希雅 的家。 亞希雅 因年紀老邁，兩眼發直，不能看見。
1KGS|14|5|耶和華對 亞希雅 說：「看哪， 耶羅波安 的妻子來問你她兒子的事，因她兒子病了，你當如此如此告訴她。她進來的時候會扮成別的婦人。」
1KGS|14|6|她剛進門， 亞希雅 聽見她的腳步聲，就說：「 耶羅波安 的妻子，進來吧！你為何扮成別的婦人呢？我奉差遣將凶信告訴你。
1KGS|14|7|你回去告訴 耶羅波安 說：『耶和華－ 以色列 的上帝如此說：我從百姓中提拔了你，立你作我百姓 以色列 的君王，
1KGS|14|8|將 大衛 家的國撕裂，賜給你，你卻不效法我僕人 大衛 ，遵守我的誡命，全心順從我，行我眼中看為正的事。
1KGS|14|9|你反倒行惡，比在你之前所有的人更嚴重；你離開了我，為自己立了別神，鑄了偶像，惹我發怒，將我丟在背後。
1KGS|14|10|因此，看哪，我必使災禍臨到 耶羅波安 的家，把屬 耶羅波安 的男丁，無論是奴役的、自由的，都從 以色列 中剪除。我必除滅 耶羅波安 的家，如同人掃除糞土，直到消滅。
1KGS|14|11|凡屬 耶羅波安 的人，死在城中的必被狗吃，死在田野的必被空中的鳥吃。這是耶和華說的。』
1KGS|14|12|你起身回家去吧！你的腳一進城，孩子就死了。
1KGS|14|13|以色列 眾人必為他哀哭，為他安葬。凡屬 耶羅波安 的人，只有他可以葬入墳墓，因為在 耶羅波安 的家中，只有他向耶和華－ 以色列 的上帝表現出好的行為。
1KGS|14|14|耶和華必另立一王治理 以色列 ，這一天，他必剪除 耶羅波安 的家；甚麼時候呢？現在就是了。
1KGS|14|15|耶和華必擊打 以色列 ，使他們搖動，像水中的蘆葦一樣，又將他們從耶和華賜給他們列祖的美地上拔出來，分散在 大河 那邊，因為他們造了 亞舍拉 ，惹耶和華發怒。
1KGS|14|16|因 耶羅波安 所犯的罪，又因他使 以色列 陷入罪裏，耶和華必將 以色列 交出來。」
1KGS|14|17|耶羅波安 的妻子起身回去，到了 得撒 ，剛到門檻，孩子就死了。
1KGS|14|18|以色列 眾人為他安葬，為他哀哭，正如耶和華藉他僕人 亞希雅 先知所說的話。
1KGS|14|19|耶羅波安 其餘的事，他怎樣打仗，怎樣作王，看哪，都寫在《以色列諸王記》上。
1KGS|14|20|耶羅波安 作王二十二年，就與他祖先同睡，他兒子 拿答 接續他作王。
1KGS|14|21|所羅門 的兒子 羅波安 作 猶大 王。他登基的時候年四十一歲，在 耶路撒冷 ，就是耶和華從 以色列 眾支派中所選擇立他名的城，作王十七年。 羅波安 的母親名叫 拿瑪 ，是 亞捫 人。
1KGS|14|22|猶大 人行耶和華眼中看為惡的事，以所犯的罪惹動他的妒忌，比他們的祖先所犯的一切更嚴重。
1KGS|14|23|因為他們在各高岡上，各青翠樹下築丘壇，立柱像和 亞舍拉 。
1KGS|14|24|國中也有男的廟妓。他們效法耶和華在 以色列 人面前所趕出的外邦人，行一切可憎惡的事。
1KGS|14|25|羅波安 王第五年， 埃及 王 示撒 上來攻打 耶路撒冷 ，
1KGS|14|26|奪了耶和華殿和王宮裏的寶物，盡都帶走，又奪走 所羅門 製造的一切金盾牌。
1KGS|14|27|羅波安 王製造銅盾牌代替那些金盾牌，交給看守王宮宮門的護衛長看管。
1KGS|14|28|每逢王進耶和華的殿，護衛兵就舉起這些盾牌；隨後仍將盾牌送回護衛室。
1KGS|14|29|羅波安 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？
1KGS|14|30|羅波安 與 耶羅波安 時常交戰。
1KGS|14|31|羅波安 與他祖先同睡，與他祖先同葬在 大衛城 。他母親名叫 拿瑪 ，是 亞捫 人，他兒子 亞比央 接續他作王。
1KGS|15|1|尼八 的兒子 耶羅波安 王十八年， 亞比央 登基作 猶大 王，
1KGS|15|2|在 耶路撒冷 作王三年。他母親名叫 瑪迦 ，是 押沙龍 的女兒。
1KGS|15|3|亞比央 行他父親從前所犯一切的罪，他的心不像他曾祖父 大衛 以純正的心順服耶和華－他的上帝。
1KGS|15|4|然而耶和華－他的上帝因 大衛 的緣故，仍使大衛在 耶路撒冷 有燈光，立他兒子接續他作王，又堅立 耶路撒冷 。
1KGS|15|5|因為 大衛 除了 赫 人 烏利亞 那件事，都行耶和華眼中看為正的事，一生沒有違背耶和華一切所吩咐的。
1KGS|15|6|羅波安 在世的日子常與 耶羅波安 交戰。
1KGS|15|7|亞比央 其餘的事，凡他所做的，不都寫在《猶大列王記》上嗎？ 亞比央 常與 耶羅波安 交戰。
1KGS|15|8|亞比央 與他祖先同睡，葬在 大衛城 ，他兒子 亞撒 接續他作王。
1KGS|15|9|以色列 王 耶羅波安 第二十年， 亞撒 登基作 猶大 王，
1KGS|15|10|在 耶路撒冷 作王四十一年。他祖母名叫 瑪迦 ，是 押沙龍 的女兒。
1KGS|15|11|亞撒 效法他的高祖父 大衛 行耶和華眼中看為正的事，
1KGS|15|12|從國中除去男的廟妓，又除掉他祖先所造的一切偶像。
1KGS|15|13|他甚至廢了他祖母 瑪迦 太后的位，因 瑪迦 造了可憎的 亞舍拉 。 亞撒 砍下她的偶像，在 汲淪溪 邊燒了，
1KGS|15|14|只是丘壇還沒有廢去。 亞撒 一生向耶和華存純正的心。
1KGS|15|15|亞撒 將他父親所分別為聖與自己所分別為聖的金銀和器皿都奉到耶和華的殿裏。
1KGS|15|16|亞撒 和 以色列 王 巴沙 在世的日子常常交戰。
1KGS|15|17|以色列 王 巴沙 上來攻擊 猶大 ，修築 拉瑪 ，不許人從 猶大 王 亞撒 那裏出入。
1KGS|15|18|於是 亞撒 把耶和華殿和王宮府庫裏所剩下的金銀都交在他臣僕手中，派他們到住在 大馬士革 的 亞蘭 王，就是 希旬 的孫子， 他伯利門 的兒子 便‧哈達 那裏去，說：
1KGS|15|19|「你父曾與我父立約，我與你也要這樣立約。看哪，我把金銀送給你作禮物，請你廢掉你與 以色列 王 巴沙 所立的約，使他從我這裏撤退。」
1KGS|15|20|便‧哈達 聽從了 亞撒 王，就派遣他的軍官去攻打 以色列 的城鎮，攻下了 以雲 、 但 、 亞伯‧伯‧瑪迦 、全 基尼烈 、 拿弗他利 全地。
1KGS|15|21|巴沙 聽見了，就停工不修築 拉瑪 ，仍住在 得撒 。
1KGS|15|22|於是 亞撒 王向 猶大 眾人宣佈，不准任何人推辭，吩咐他們運走 巴沙 修築 拉瑪 所用的石頭和木料。 亞撒 王用它們來修築 便雅憫 的 迦巴 和 米斯巴 。
1KGS|15|23|亞撒 其餘的事，他英勇的事蹟，凡他所做的，以及他所建築的城鎮，不都寫在《猶大列王記》上嗎？只是 亞撒 年老的時候患有腳疾。
1KGS|15|24|亞撒 與他祖先同睡，與他祖先同葬在 大衛城 ，他兒子 約沙法 接續他作王。
1KGS|15|25|猶大 王 亞撒 第二年， 耶羅波安 的兒子 拿答 登基作 以色列 王二年，
1KGS|15|26|拿答 行耶和華眼中看為惡的事，行他父親所行的道，犯他父親使 以色列 陷入罪裏的那罪。
1KGS|15|27|以薩迦 人 亞希雅 的兒子 巴沙 背叛 拿答 ，在 非利士 人的 基比頓 殺了他，那時 拿答 和 以色列 眾人正圍困 基比頓 。
1KGS|15|28|猶大 王 亞撒 第三年， 巴沙 殺了 拿答 ，篡了他的位。
1KGS|15|29|巴沙 一作王就殺了 耶羅波安 全家， 耶羅波安 家凡有氣息的，一個也沒有留下，都殺滅了，正如耶和華藉他僕人 示羅 人 亞希雅 所說的話。
1KGS|15|30|這是因為 耶羅波安 所犯的罪，他使 以色列 陷入罪裏，激怒了耶和華－ 以色列 的上帝。
1KGS|15|31|拿答 其餘的事，凡他所做的，不都寫在《以色列諸王記》上嗎？
1KGS|15|32|亞撒 和 以色列 王 巴沙 在世的日子常常交戰。
1KGS|15|33|猶大 王 亞撒 第三年， 亞希雅 的兒子 巴沙 在 得撒 登基，作全 以色列 的王二十四年。
1KGS|15|34|他行耶和華眼中看為惡的事，行 耶羅波安 所行的道，犯他使 以色列 陷入罪裏的那罪。
1KGS|16|1|耶和華的話臨到 哈拿尼 的兒子 耶戶 ，責備 巴沙 說：
1KGS|16|2|「我既從塵埃中提拔你，立你作我百姓 以色列 的君王，你竟行 耶羅波安 所行的道，使我的百姓 以色列 陷入罪裏，以他們的罪惹我發怒，
1KGS|16|3|看哪，我必除盡 巴沙 和他的家，使你的家像 尼八 的兒子 耶羅波安 的家一樣。
1KGS|16|4|凡屬 巴沙 的人，死在城中的必被狗吃，死在田野的必被空中的鳥吃。」
1KGS|16|5|巴沙 其餘的事，凡他所做的和他英勇的事蹟，不都寫在《以色列諸王記》上嗎？
1KGS|16|6|巴沙 與他祖先同睡，葬在 得撒 ，他兒子 以拉 接續他作王。
1KGS|16|7|耶和華的話臨到 哈拿尼 的兒子 耶戶 先知，責備 巴沙 和他的家，因他行耶和華眼中看為惡的一切事，以他手所做的惹耶和華發怒，像 耶羅波安 的家一樣，又因他殺了 耶羅波安 全家。
1KGS|16|8|猶大 王 亞撒 第二十六年， 巴沙 的兒子 以拉 在 得撒 登基，作 以色列 王二年。
1KGS|16|9|他的大臣 心利 ，就是管理他一半戰車的軍官背叛他。當他在 得撒 ，在王宮的管家 亞雜 家裏喝醉的時候，
1KGS|16|10|心利 進去擊殺他，把他殺死，篡了他的位。這是 猶大 王 亞撒 第二十七年的事。
1KGS|16|11|心利 一坐上王位就殺了 巴沙 全家，連他的親屬和朋友，一個男丁也沒有留下。
1KGS|16|12|心利 滅絕 巴沙 全家，正如耶和華藉 耶戶 先知責備 巴沙 的話。
1KGS|16|13|這是因為 巴沙 和他兒子 以拉 的一切罪，就是他們使 以色列 陷入罪裏的那罪，以虛無的神明 惹耶和華－ 以色列 的上帝發怒。
1KGS|16|14|以拉 其餘的事，凡他所做的，不都寫在《以色列諸王記》上嗎？
1KGS|16|15|猶大 王 亞撒 第二十七年， 心利 在 得撒 作王七日。那時軍兵正安營圍攻 非利士 人的 基比頓 。
1KGS|16|16|軍兵在營中聽說 心利 已經背叛，殺了王， 以色列 眾人當日就在營中立 暗利 元帥作 以色列 王。
1KGS|16|17|暗利 率領 以色列 眾人，從 基比頓 上去，圍困 得撒 。
1KGS|16|18|心利 見城被攻陷，就進了王宮的堡壘，放火焚燒宮殿，自焚而死。
1KGS|16|19|這是因為他犯罪，行耶和華眼中看為惡的事，行 耶羅波安 所行的道，犯他使 以色列 陷入罪裏的那罪。
1KGS|16|20|心利 其餘的事和他背叛的事，不都寫在《以色列諸王記》上嗎？
1KGS|16|21|那時， 以色列 百姓分為兩半：一半隨從 基納 的兒子 提比尼 ，要擁立他作王；另一半隨從 暗利 。
1KGS|16|22|但隨從 暗利 的百姓勝過隨從 基納 兒子 提比尼 的百姓。 提比尼 死了， 暗利 就作了王。
1KGS|16|23|猶大 王 亞撒 第三十一年， 暗利 登基作 以色列 王十二年；他在 得撒 作王六年。
1KGS|16|24|暗利 用二他連得銀子向 撒瑪 買了 撒瑪利亞山 ，在山上建城，按著山的原主 撒瑪 的名，給所建的城起名叫 撒瑪利亞 。
1KGS|16|25|暗利 行耶和華眼中看為惡的事，比他以前所有的王作惡更嚴重。
1KGS|16|26|因為他行了 尼八 的兒子 耶羅波安 所行的道，犯他使 以色列 陷入罪裏的那罪，以虛無的神明惹耶和華－ 以色列 的上帝發怒。
1KGS|16|27|暗利 其餘的事，他所做的和所顯出的英勇事蹟，不都寫在《以色列諸王記》上嗎？
1KGS|16|28|暗利 與他祖先同睡，葬在 撒瑪利亞 ，他兒子 亞哈 接續他作王。
1KGS|16|29|猶大 王 亞撒 第三十八年， 暗利 的兒子 亞哈 登基作 以色列 王。 暗利 的兒子 亞哈 在 撒瑪利亞 作 以色列 王二十二年。
1KGS|16|30|暗利 的兒子 亞哈 行耶和華眼中看為惡的事，比他以前所有的王更嚴重。
1KGS|16|31|他犯了 尼八 的兒子 耶羅波安 所犯的罪，還當作是小事，又娶了 西頓 王 謁巴力 的女兒 耶洗別 為妻，去事奉 巴力 ，敬拜它，
1KGS|16|32|又在 撒瑪利亞 建 巴力廟 ，在廟裏為 巴力 築壇。
1KGS|16|33|亞哈 又造 亞舍拉 ，他所做的惹耶和華－ 以色列 的上帝發怒，比他以前所有的 以色列 王更嚴重。
1KGS|16|34|亞哈 的日子， 伯特利 人 希伊勒 重修 耶利哥 。立根基的時候，他喪了長子 亞比蘭 ；安門的時候，他喪了幼子 西割 ，正如耶和華藉 嫩 的兒子 約書亞 所說的話。
1KGS|17|1|住在 基列 的 提斯比 人 以利亞 對 亞哈 說：「我指著所事奉永生的耶和華－ 以色列 的上帝起誓，這幾年我若不禱告，必不降露水，也不下雨。」
1KGS|17|2|耶和華的話臨到 以利亞 ，說：
1KGS|17|3|「你離開這裏往東去，躲在 約旦河 東邊的 基立溪 旁。
1KGS|17|4|你要喝那溪裏的水，我已吩咐烏鴉在那裏供養你。」
1KGS|17|5|於是 以利亞 去了，他遵照耶和華的話做，去住在 約旦河 東的 基立溪 旁。
1KGS|17|6|烏鴉早上給他叼餅和肉來，晚上也有餅和肉，他又喝溪裏的水。
1KGS|17|7|過了些日子溪水乾了，因為雨沒有下在地上。
1KGS|17|8|耶和華的話臨到他，說：
1KGS|17|9|「你起身到 西頓 的 撒勒法 去，住在那裏，看哪，我已吩咐那裏的一個寡婦供養你。」
1KGS|17|10|以利亞 就起身往 撒勒法 去。他到了城門，看哪，有一個寡婦在那裏撿柴。 以利亞 呼喚她說：「請你用器皿取點水來給我喝。」
1KGS|17|11|她去取水的時候， 以利亞 又呼喚她說：「請你手裏也拿點餅來給我。」
1KGS|17|12|她說：「我指著永生的耶和華－你的上帝起誓，我沒有餅，罈內只有一把麵，瓶裏只有一點油。看哪，我去找兩根柴，帶回家為我和我兒子做餅。我們吃了，就等死吧！」
1KGS|17|13|以利亞 對她說：「不要怕！你去照你所說的做吧！只要先為我做一個小餅，拿來給我，然後為你和你的兒子做餅；
1KGS|17|14|因為耶和華－ 以色列 的上帝如此說：『罈內的麵必不用盡，瓶裏的油必不短缺，直到耶和華使雨降在地上的日子。』」
1KGS|17|15|婦人就照 以利亞 的話去做。她和 以利亞 ，以及她家中的人，吃了許多日子。
1KGS|17|16|罈內的麵果然沒有用盡，瓶裏的油也不短缺，正如耶和華藉 以利亞 所說的話。
1KGS|17|17|這事以後，那婦人，就是那家的女主人，她的兒子病了，病得很重，甚至沒有氣息。
1KGS|17|18|婦人對 以利亞 說：「神人哪，我跟你有甚麼關係，你竟到我這裏來，使上帝記起我的罪，以致我的兒子死了呢？」
1KGS|17|19|以利亞 對她說：「把你兒子交給我。」 以利亞 就從婦人懷中接過孩子來，抱到他所住的頂樓，放在自己的床上。
1KGS|17|20|他求告耶和華說：「耶和華－我的上帝啊，我寄居在這寡婦的家裏，你卻降禍於她，使她的兒子死了嗎？」
1KGS|17|21|以利亞 三次伏在孩子的身上，求告耶和華說：「耶和華－我的上帝啊，求你使這孩子的生命歸回給他吧！」
1KGS|17|22|耶和華聽了 以利亞 的呼求，孩子的生命歸回給他，他就活了。
1KGS|17|23|以利亞 把孩子從樓上抱下來，進了房間交給他母親，說：「看，你的兒子活了！」
1KGS|17|24|婦人對 以利亞 說：「現在我知道你是神人，耶和華藉你口所說的話是真的。」
1KGS|18|1|過了許多日子，到了第三年，耶和華的話臨到 以利亞 ，說：「你去，讓 亞哈 看見你，我要降雨在地面上。」
1KGS|18|2|以利亞 就去，要讓 亞哈 見到他。那時， 撒瑪利亞 的饑荒非常嚴重。
1KGS|18|3|亞哈 召來他的管家 俄巴底 。 俄巴底 非常敬畏耶和華。
1KGS|18|4|耶洗別 殺耶和華先知的時候， 俄巴底 把一百個先知藏了，每五十人藏在一個洞裏，拿餅和水供養他們。
1KGS|18|5|亞哈 對 俄巴底 說：「我們要走遍這地，到一切水泉旁和一切溪邊，或者能找到青草，可以救活馬和騾子，免得喪失一些牲畜。」
1KGS|18|6|於是二人分地巡查， 亞哈 獨自走一路， 俄巴底 獨自走另一路。
1KGS|18|7|俄巴底 在路上時，看哪， 以利亞 遇見他。 俄巴底 認出他來，就臉伏於地，說：「你是我主 以利亞 嗎？」
1KGS|18|8|以利亞 對他說：「我是。你去，告訴你主人說：『看哪， 以利亞 在這裏。』」
1KGS|18|9|俄巴底 說：「僕人犯了甚麼罪，你竟要把我交在 亞哈 手裏，使他殺我呢？
1KGS|18|10|我指著永生的耶和華－你的上帝起誓，無論哪一邦哪一國，我主都派人去找你。若他們說：『不在這裏』，他就叫那邦那國的人起誓說，他們實在找不到你。
1KGS|18|11|現在你說：『你去告訴你主人說，看哪， 以利亞 在這裏』；
1KGS|18|12|恐怕我一離開你，耶和華的靈就把你提到我所不知道的地方去。這樣，我去告訴 亞哈 ，他若找不到你，就必殺我。僕人是自幼敬畏耶和華的。
1KGS|18|13|耶洗別 殺耶和華先知的時候，我把耶和華的一百個先知藏了，每五十人藏在一個洞裏，拿餅和水供養他們，難道沒有人把我做的這事告訴我主嗎？
1KGS|18|14|現在你說：『你去告訴你主人說，看哪， 以利亞 在這裏』，他一定會殺我。」
1KGS|18|15|以利亞 說：「我指著所事奉永生的萬軍之耶和華起誓，我今日要讓 亞哈 見到我。」
1KGS|18|16|於是 俄巴底 去迎見 亞哈 ，告訴他這事。 亞哈 就去見 以利亞 。
1KGS|18|17|亞哈 見了 以利亞 ，就說：「真的是你嗎？你這使 以色列 遭殃的人！」
1KGS|18|18|以利亞 說：「使 以色列 遭殃的不是我，而是你和你的父家，因為你們離棄耶和華的誡命 ，去隨從 巴力 。
1KGS|18|19|現在你要派人去召集 以色列 眾人，以及 耶洗別 所供養的四百五十個 巴力 的先知和四百個 亞舍拉 的先知，叫他們都上 迦密山 到我這裏來。」
1KGS|18|20|亞哈 就派人到 以色列 眾人那裏，召集先知上 迦密山 。
1KGS|18|21|以利亞 近前來對眾百姓說：「你們心持二意要到幾時呢？如果耶和華是上帝，就當順從耶和華；如果是 巴力 ，就當順從 巴力 。」百姓一言不答。
1KGS|18|22|以利亞 對百姓說：「作耶和華先知的只剩下我一個； 巴力 的先知卻有四百五十人。
1KGS|18|23|請給我們兩頭牛犢， 巴力 的先知可以為自己挑選一頭牛犢，切成小塊，放在柴上，不要點火；我也預備一頭牛犢放在柴上，也不點火。
1KGS|18|24|你們求告你們神明的名，我也求告耶和華的名。那應允禱告降火的就是上帝。」眾百姓回答說：「好主意。」
1KGS|18|25|以利亞 對 巴力 的先知說：「因為你們人多，先挑選一頭牛犢，預備好了，求告你們神明的名，卻不要點火。」
1KGS|18|26|他們把所給他們的牛犢預備好了，從早晨到中午，求告 巴力 的名說：「 巴力 啊，求你應允我們！」卻沒有聲音，也沒有回應。他們就在所築的壇四圍蹦跳。
1KGS|18|27|到了正午， 以利亞 嘲笑他們，說：「大聲求告吧！因為它是神明，它或許在默想，或許正忙著 ，或許在路上，或許在睡覺，它該醒過來了。」
1KGS|18|28|他們大聲求告，按著他們的儀式，用刀槍刺割自己，直到渾身流血。
1KGS|18|29|中午過去了，他們狂呼亂叫，直到獻晚祭的時候，卻沒有聲音，沒有回應的，也沒有理睬的。
1KGS|18|30|以利亞 對眾百姓說：「你們到我這裏來。」眾百姓就到他那裏，他把那已經毀壞了的耶和華的壇修好。
1KGS|18|31|以利亞 按照 雅各 子孫支派的數目，取了十二塊石頭；耶和華的話曾臨到 雅各 ，說：「你的名要叫 以色列 。」
1KGS|18|32|以利亞 用這些石頭為耶和華的名築一座壇，在壇的四圍挖溝，可容納二細亞穀種。
1KGS|18|33|他又在壇上擺好了柴，把牛犢切成小塊放在柴上，說：「你們用四個桶盛滿水，倒在燔祭和柴上。」
1KGS|18|34|他又說：「倒第二次。」他們就倒第二次。他又說：「倒第三次。」他們就倒第三次。
1KGS|18|35|水流到壇的四圍，溝裏也滿了水。
1KGS|18|36|到了獻晚祭的時候，先知 以利亞 近前來，說：「耶和華－ 亞伯拉罕 、 以撒 、 以色列 的上帝啊，求你今日使人知道你是 以色列 的上帝，我是你的僕人，我遵照你的話做這一切事。
1KGS|18|37|求你應允我，耶和華啊，應允我，使這百姓知道你－耶和華是上帝，是你叫他們回心轉意的。」
1KGS|18|38|於是，耶和華降下火來，燒盡燔祭、木柴、石頭、塵土，又燒乾了溝裏的水。
1KGS|18|39|眾百姓看見了，就臉伏於地，說：「耶和華是上帝！耶和華是上帝！」
1KGS|18|40|以利亞 對他們說：「拿住 巴力 的先知，不讓任何人逃走！」眾人就拿住他們。 以利亞 帶他們到 基順河 邊，在那裏殺了他們。
1KGS|18|41|以利亞 對 亞哈 說：「你現在可以上去吃喝，因為有暴雨的響聲了。」
1KGS|18|42|亞哈 就上去吃喝。 以利亞 上了 迦密山 頂，屈身在地，把臉伏在兩膝之中。
1KGS|18|43|他對僕人說：「你上去，向海觀看。」僕人就上去觀看，說：「沒有甚麼。」 以利亞 說：「你再去。」如此七次。
1KGS|18|44|第七次，僕人說：「看哪，有一小片雲從海裏上來，好像人的手掌那麼大。」 以利亞 說：「你上去告訴 亞哈 ，當套車下去，免得被雨阻擋。」
1KGS|18|45|霎時間，天因風雲黑暗，降下大雨。 亞哈 就坐上車，往 耶斯列 去了。
1KGS|18|46|耶和華的手按在 以利亞 身上，他就束上腰，奔在 亞哈 前頭，一路到 耶斯列 。
1KGS|19|1|亞哈 把 以利亞 一切所做的和他用刀殺眾先知的事都告訴 耶洗別 。
1KGS|19|2|耶洗別 就派使者到 以利亞 那裏，說：「明日約這時候，我若不使你的性命像那些人的性命一樣，願神明重重懲罰我。」
1KGS|19|3|以利亞 害怕 ，就起來逃命，到了 猶大 的 別是巴 ，把僕人留在那裏。
1KGS|19|4|他自己在曠野走了一日的路程，來到一棵羅騰 樹下，就坐在那裏求死，說：「耶和華啊，現在夠了！求你取我的性命吧，因為我不比我的祖先好。」
1KGS|19|5|他躺在羅騰樹下睡著了。看哪，有一個天使拍他，對他說：「起來吃吧！」
1KGS|19|6|他觀看，看哪，頭旁有燒熱的石頭烤的餅和一壺水，他就吃了喝了，又再躺下。
1KGS|19|7|耶和華的使者回來，第二次拍他，說：「起來吃吧！因為你要走的路很遠。」
1KGS|19|8|他就起來吃了喝了，仗著這飲食的力走了四十晝夜，到了上帝的山，就是 何烈山 。
1KGS|19|9|他在那裏進了一個洞，在洞中過夜。看哪，耶和華的話臨到他，說：「 以利亞 ，你在這裏做甚麼？」
1KGS|19|10|他說：「我為耶和華－萬軍之上帝大發熱心，因為 以色列 人背棄了你的約，毀壞了你的壇，用刀殺了你的先知，只剩下我一人，他們還要追殺我。」
1KGS|19|11|耶和華說：「你出來站在山上，在耶和華面前。」看哪，耶和華從那裏經過。在耶和華面前有烈風大作，山崩石裂，耶和華卻不在風中；風後有地震，耶和華也不在其中；
1KGS|19|12|地震後有火，耶和華也不在火中；火以後，有輕微細小的聲音。
1KGS|19|13|以利亞 聽見，就用外衣蒙臉，出來站在洞口。聽啊，有聲音向他說：「 以利亞 ，你在這裏做甚麼？」
1KGS|19|14|他說：「我為耶和華－萬軍之上帝大發熱心，因為 以色列 人背棄了你的約，毀壞了你的壇，用刀殺了你的先知，只剩下我一人，他們還要追殺我。」
1KGS|19|15|耶和華對他說：「去吧，從原路回去，往 大馬士革 的曠野去。到了那裏，你要膏 哈薛 作 亞蘭 王，
1KGS|19|16|又膏 寧示 的孫子 耶戶 作 以色列 王，並膏 亞伯‧米何拉 人 沙法 的兒子 以利沙 作先知接續你。
1KGS|19|17|將來逃過 哈薛 之刀的，必被 耶戶 所殺；逃過 耶戶 之刀的，必被 以利沙 所殺。
1KGS|19|18|但我在 以色列 中留下七千人，是未曾向 巴力 屈膝，未曾親吻 巴力 的。」
1KGS|19|19|於是， 以利亞 離開那裏走了，遇見 沙法 的兒子 以利沙 ；他正在耕田，在他前頭有十二對牛，自己趕著第十二對。 以利亞 經過他，把自己的外衣搭在他身上。
1KGS|19|20|以利沙 就離開牛，跑到 以利亞 那裏，說：「請你讓我先與父母吻別，然後我就跟隨你。」 以利亞 對他說：「因我對你所做的事，你去吧，然後回來。 」
1KGS|19|21|以利沙 離開他回去，宰了一對牛，用套牛的器具煮肉給百姓吃，隨後就起身跟隨 以利亞 ，服事他。
1KGS|20|1|亞蘭 王 便‧哈達 召集他的全軍，率領三十二個王，帶著馬和戰車，上來圍困 撒瑪利亞 ，要攻打它。
1KGS|20|2|他派使者進城到 以色列 王 亞哈 那裏，對他說：「 便‧哈達 如此說：
1KGS|20|3|『你的金銀都要歸我，你妻妾兒女中最美的也要歸我。』」
1KGS|20|4|以色列 王回答說：「我主我王啊，就照著你的話，我和我所有的都歸你。」
1KGS|20|5|使者又來說：「 便‧哈達 如此說：『我已派人到你那裏，要你把你的金銀、妻妾、兒女都歸我。』
1KGS|20|6|但明日約在這時候，我還要派臣僕到你那裏，搜查你的家和你僕人的家，你眼中一切所喜愛的都由他們的手拿走。」
1KGS|20|7|以色列 王召了國內所有的長老來，說：「你們要知道，看哪，這人是來找麻煩的！他派人到我這裏來，要我的妻妾、兒女和金銀，我並沒有拒絕他。」
1KGS|20|8|所有的長老和眾百姓對王說：「不要聽從他，也不要答應他。」
1KGS|20|9|以色列 王對 便‧哈達 的使者說：「你們告訴我主我王說：『王頭一次派人向僕人所要的一切，僕人都依從，但這事我不能依從。』」使者就去回覆 便‧哈達 。
1KGS|20|10|便‧哈達 又派人到 亞哈 那裏，說：「 撒瑪利亞 的塵土若足夠跟從我的軍兵每人手拿一把，願神明重重懲罰我！」
1KGS|20|11|以色列 王回答說：「你們告訴他說，『剛束上腰帶的，不要像已卸下的那樣誇口。』」
1KGS|20|12|便‧哈達 和諸王正在帳幕裏喝酒，聽見這話，就對他臣僕說：「擺陣吧！」他們就擺陣攻城。
1KGS|20|13|看哪，一個先知靠近 以色列 王 亞哈 ，說：「耶和華如此說：『這一大群人你看見了嗎？看哪，今日我必把他們交在你手裏，你就知道我是耶和華。』」
1KGS|20|14|亞哈 說：「藉著誰呢？」他說：「耶和華如此說：『藉著跟從省長的年輕人。』」 亞哈 說：「誰要開戰呢？」他說：「你！」
1KGS|20|15|於是 亞哈 數點跟從省長的年輕人，共二百三十二名，然後又數點 以色列 的眾軍兵，共七千名。
1KGS|20|16|中午，他們出了城； 便‧哈達 和幫助他的三十二個王正在帳幕裏暢飲。
1KGS|20|17|跟從省長的年輕人先出城。 便‧哈達 派人去，他們回報說：「有人從 撒瑪利亞 出來了。」
1KGS|20|18|他說：「他們若為求和出來，要活捉他們，若為打仗出來，也要活捉他們。」
1KGS|20|19|跟從省長的年輕人，和跟隨他們的軍兵，都出了城，
1KGS|20|20|各人遇見敵人就擊殺。 亞蘭 人逃跑， 以色列 人追趕他們； 亞蘭 王 便‧哈達 騎著馬和騎兵一同逃跑。
1KGS|20|21|以色列 王出城攻擊 馬和戰車，大大擊殺 亞蘭 人。
1KGS|20|22|那先知靠近 以色列 王，對他說：「去吧，你當自強，看清楚，也要知道你所要做的事，因為再過一年， 亞蘭 王會上來攻擊你。」
1KGS|20|23|亞蘭 王的臣僕對他說：「他們的神是山神，所以他們勝過我們。但在平原與他們打仗，我們一定勝過他們。
1KGS|20|24|王當做這樣的事，把諸王革去，派軍官代替他們，
1KGS|20|25|又照著王喪失軍兵的數目，再招募一支軍隊，馬補馬，車補車。然後在平原與他們打仗，我們一定勝過他們。」王就聽臣僕的話，照樣去做。
1KGS|20|26|過了一年， 便‧哈達 果然召集 亞蘭 人上 亞弗 去，要與 以色列 人打仗。
1KGS|20|27|以色列 人也召集軍兵，預備食物，去迎戰 亞蘭 人。 以色列 人對著他們安營，好像兩小群的山羊； 亞蘭 人卻佈滿了地面。
1KGS|20|28|有神人靠近，對 以色列 王說：「耶和華如此說：『 亞蘭 人既說我－耶和華是山神，不是平原之神，我必將這一大群人全都交在你手中，你們就知道我是耶和華。』」
1KGS|20|29|以色列 人與 亞蘭 人相對安營七日，到第七日兩軍開戰。那一日 以色列 人殺了 亞蘭 的十萬步兵，
1KGS|20|30|其餘的都逃向 亞弗 ，到了城裏，城牆倒塌，壓死了剩下的二萬七千人。 便‧哈達 也逃入城內，藏在嚴密的內室裏。
1KGS|20|31|他的臣僕對他說：「看哪，我們聽說 以色列 家的王都是仁慈的王；讓我們腰束麻布，頭套繩索，出去到 以色列 王那裏，也許他會存留王的性命。」
1KGS|20|32|於是他們腰束麻布，頭套繩索，來到 以色列 王那裏，說：「王的僕人 便‧哈達 說：『求王饒我一命。』」 亞哈 說：「他還活著嗎？他是我的兄弟。」
1KGS|20|33|這些人正在探測吉凶，就立即抓住他的話說：「 便‧哈達 是王的兄弟！」王說：「你們去請他來。」 便‧哈達 出來到王那裏，王就請他上車。
1KGS|20|34|便‧哈達 對王說：「我父從你父那裏所奪的城鎮，我必歸還給你。你可以在 大馬士革 為你自己設立街市，像我父在 撒瑪利亞 所設立的一樣。」 亞哈 說：「我照此立約，放你回去。」王就與他立約，放了他。
1KGS|20|35|有一個人是先知的門徒，遵照耶和華的話對他同伴說：「你打我吧！」那人不肯打他。
1KGS|20|36|他就對那人說：「你既不聽從耶和華的話，看哪，你一離開我，必有獅子咬死你。」那人一離開他，果然遇見獅子，把他咬死了。
1KGS|20|37|先知的門徒又遇見一個人，對他說：「你打我吧！」那人就打他，把他打傷。
1KGS|20|38|那先知就去了，用頭巾蒙眼，改了裝，在路旁等候王。
1KGS|20|39|王從那裏經過，他向王呼叫說：「僕人出戰的時候，看哪，有人轉過來，帶了一個人到我這裏來，說：『你要看守這人，若他真的失蹤了，你的性命必代替他的性命，否則，你就要交出一他連得銀子來。』
1KGS|20|40|僕人正在到處忙碌的時候，那人就不見了。」 以色列 王對他說：「你自己決定了，就必照樣判你。」
1KGS|20|41|他急忙除掉蒙眼的頭巾， 以色列 王就認出他是一個先知。
1KGS|20|42|他對王說：「耶和華如此說：『因你把我決定要消滅的人從你手中放走，所以你的命必代替他的命，你的百姓必代替他的百姓。』」
1KGS|20|43|於是 以色列 王生氣，憂悶地回 撒瑪利亞 ，到自己的宮去了。
1KGS|21|1|這些事以後，又有一事。 耶斯列 人 拿伯 在 耶斯列 有一個葡萄園，靠近 撒瑪利亞 ， 亞哈 王的宮。
1KGS|21|2|亞哈 對 拿伯 說：「把你的葡萄園給我作菜園，因為它靠近我的宮，我就把更好的葡萄園換給你。你若要銀子，我就按著價錢給你。」
1KGS|21|3|拿伯 對 亞哈 說：「耶和華不准我把我祖先留下的產業給你。」
1KGS|21|4|亞哈 因 耶斯列 人 拿伯 說「我不把我祖先留下的產業給你」，就生氣，憂悶地回宮，躺在床上，臉轉向內，也不吃飯。
1KGS|21|5|耶洗別 王后來對他說：「你為甚麼心裏這樣生氣，不吃飯呢？」
1KGS|21|6|他對王后說：「我向 耶斯列 人 拿伯 說：『把你的葡萄園按價錢賣給我，或是你願意，我可以把別的葡萄園換給你。』他卻說：『我不把我的葡萄園給你。』」
1KGS|21|7|耶洗別 王后對王說：「你現在是不是治理 以色列 國呢？只管起來，心裏暢暢快快地吃飯，我會把 耶斯列 人 拿伯 的葡萄園給你。」
1KGS|21|8|於是王后以 亞哈 的名義寫信，蓋上王的印，把信送給那些與 拿伯 同城居住的長老和貴族。
1KGS|21|9|她在信上寫著說：「你們當宣告禁食，叫 拿伯 坐在百姓的高位上，
1KGS|21|10|又叫兩個無賴坐在 拿伯 對面，作證告他說：『你詛咒了上帝和王。』然後把他拉出去用石頭打死。」
1KGS|21|11|那些與 拿伯 同城居住的長老和貴族，照 耶洗別 送給他們的信去做。正如她送的信上所寫，
1KGS|21|12|他們宣告禁食，叫 拿伯 坐在百姓的高位上。
1KGS|21|13|有兩個無賴來，坐在 拿伯 對面。無賴當著百姓作證告他說：「 拿伯 詛咒上帝和王了！」眾人就把他拉到城外，用石頭打他，他就死了。
1KGS|21|14|於是他們派人到 耶洗別 那裏，說：「 拿伯 被石頭打死了。」
1KGS|21|15|耶洗別 聽見 拿伯 被石頭打死，就對 亞哈 說：「你起來，去取得 耶斯列 人 拿伯 不肯出價賣給你的葡萄園吧！因為 拿伯 不在了，他已經死了。」
1KGS|21|16|亞哈 聽見 拿伯 死了，就起來，下去要取得 耶斯列 人 拿伯 的葡萄園。
1KGS|21|17|耶和華的話臨到 提斯比 人 以利亞 ，說：
1KGS|21|18|「你起來，去見在 撒瑪利亞 的 以色列 王 亞哈 。看哪，他下去要取得 拿伯 的葡萄園，他正在那園裏。
1KGS|21|19|你要對他說：『耶和華如此說：你殺了人，還要取得他的產業嗎？』又要對他說：『耶和華如此說：狗在何處舔 拿伯 的血，狗也必在何處舔你的血。』」
1KGS|21|20|亞哈 對 以利亞 說：「我的仇敵啊，你找到我了嗎？」他說：「我找到你了。因為你出賣自己，行了耶和華眼中看為惡的事。
1KGS|21|21|耶和華說：『看哪，我必使災禍臨到你，把你除滅。 以色列 中凡屬 亞哈 的男丁，無論是奴役的、自由的，我都要剪除。
1KGS|21|22|我必使你的家像 尼八 的兒子 耶羅波安 的家，又像 亞希雅 的兒子 巴沙 的家，因為你惹我發怒，又使 以色列 陷入罪裏。』
1KGS|21|23|論到 耶洗別 ，耶和華說：『狗必在 耶斯列 的城郭 吃 耶洗別 。
1KGS|21|24|凡屬 亞哈 的人，死在城中的必被狗吃，死在田野的必被空中的鳥吃。』」
1KGS|21|25|（只是從來沒有像 亞哈 的，因他受 耶洗別 王后的唆使，出賣自己，行了耶和華眼中看為惡的事。
1KGS|21|26|他行了最可憎的事，隨從偶像，正如耶和華在 以色列 人面前趕出的 亞摩利 人所行的一切。）
1KGS|21|27|亞哈 聽見這些話，就撕裂衣服，禁食，貼身穿著麻布，也睡在麻布上，沮喪地走來走去。
1KGS|21|28|耶和華的話臨到 提斯比 人 以利亞 ，說：
1KGS|21|29|「 亞哈 在我面前這樣謙卑，你看見了嗎？因為他在我面前謙卑，所以在他的日子，我不降這禍；到他兒子的時候，我必降這禍於他的家。」
1KGS|22|1|亞蘭 和 以色列 之間連續三年沒有戰爭。
1KGS|22|2|到了第三年， 猶大 王 約沙法 下去見 以色列 王。
1KGS|22|3|以色列 王對臣僕說：「你們不知道 基列 的 拉末 是屬我們的嗎？我們豈可不採取行動，把它從 亞蘭 王手裏奪回來呢？」
1KGS|22|4|亞哈 問 約沙法 說：「你肯同我去攻打 基列 的 拉末 嗎？」 約沙法 對 以色列 王說：「你我不分彼此，我的軍隊就是你的軍隊，我的馬就是你的馬。」
1KGS|22|5|約沙法 對 以色列 王說：「請你先求問耶和華的話。」
1KGS|22|6|於是 以色列 王召集先知，約有四百人，問他們說：「我可以上去攻打 基列 的 拉末 嗎？還是不要上去呢？」他們說：「可以上去，因為主必將那城交在王的手裏。」
1KGS|22|7|約沙法 說：「這裏還有沒有耶和華的先知，我們好求問他呢？」
1KGS|22|8|以色列 王對 約沙法 說：「還有一個人，是 音拉 的兒子 米該雅 ，我們可以託他求問耶和華。只是我真的很恨他，因為他對我說預言，從不說吉言，總是說凶信。」 約沙法 說：「請王不要這麼說。」
1KGS|22|9|以色列 王召了一個官員來，說：「你快去，把 音拉 的兒子 米該雅 召來。」
1KGS|22|10|以色列 王和 猶大 王 約沙法 在 撒瑪利亞 城門前的禾場，各穿朝服，坐在寶座上，所有的先知都在他們面前說預言。
1KGS|22|11|基拿拿 的兒子 西底家 造了鐵角，說：「耶和華如此說：『你要用這些角牴觸 亞蘭 人，直到將他們滅盡。』」
1KGS|22|12|所有的先知也都這樣預言說：「可以上 基列 的 拉末 去，必然得勝，因為耶和華必將那城交在王的手中。」
1KGS|22|13|那去召 米該雅 的使者對他說：「看哪，眾先知都異口同聲向王說吉言，你也跟他們說一樣的話，說吉言吧！」
1KGS|22|14|米該雅 說：「我指著永生的耶和華起誓，耶和華向我說甚麼，我就說甚麼。」
1KGS|22|15|米該雅 來到王那裏，王問他：「 米該雅 ，我們可以上去攻打 基列 的 拉末 嗎？還是不要上去呢？」他對王說：「你可以上去，必然得勝，耶和華必將那城交在王的手中。」
1KGS|22|16|王對他說：「我要你發誓多少次，你才會奉耶和華的名向我說實話呢？」
1KGS|22|17|米該雅 說：「我看見 以色列 眾人散佈在山上，如同沒有牧人的羊群一般。耶和華說：『這些人沒有主人，他們可以平安地各自回家去。』」
1KGS|22|18|以色列 王對 約沙法 說：「我豈沒有告訴你，這人對我說預言，從不說吉言，只說凶信嗎？」
1KGS|22|19|米該雅 說：「因此你要聽耶和華的話！我看見耶和華坐在寶座上，天上的萬軍侍立在他左右。
1KGS|22|20|耶和華說：『誰去引誘 亞哈 上 基列 的 拉末 去陣亡呢？』這個這樣說，那個那樣說。
1KGS|22|21|隨後有一個靈出來，站在耶和華面前，說：『我去引誘他。』
1KGS|22|22|耶和華問他：『用甚麼方法呢？』他說：『我要出去，在他眾先知的口中成為謊言的靈。』耶和華說：『這樣，你去引誘他，必能成功。你出去，照樣做吧！』
1KGS|22|23|現在，看哪，耶和華使謊言的靈入了你所有的這些先知的口，並且耶和華已經宣告要降禍於你。」
1KGS|22|24|基拿拿 的兒子 西底家 前來，打 米該雅 一巴掌，說：「耶和華的靈從哪裏離開我向你說話呢？」
1KGS|22|25|米該雅 說：「看哪，你進入嚴密的內室躲藏的那日，就必看見。」
1KGS|22|26|以色列 王說：「把 米該雅 帶走，交回給 亞們 市長和 約阿施 王子。
1KGS|22|27|你們要說：『王如此說，把這個人關在監獄裏，使他受苦，吃不飽喝不足，直等到我平安回來。』」
1KGS|22|28|米該雅 說：「你若真的能平安回來，那就是耶和華沒有藉我說這話了。」他又說：「眾百姓啊，你們都要聽！」
1KGS|22|29|以色列 王和 猶大 王 約沙法 上 基列 的 拉末 去。
1KGS|22|30|以色列 王對 約沙法 說：「我要改裝上陣，你可以仍穿王袍。」 以色列 王就改裝上陣去了。
1KGS|22|31|亞蘭 王吩咐他的三十二個戰車長說：「你們不要與他們的大將或小兵交戰，只要單單攻擊 以色列 王。」
1KGS|22|32|那些戰車長看見 約沙法 就說：「這一定是 以色列 王！」他們轉過去與他交戰， 約沙法 就呼喊起來。
1KGS|22|33|戰車長見他不是 以色列 王，就轉身不追他了。
1KGS|22|34|有一人開弓，並不知情，箭恰巧射入 以色列 王鎧甲的縫裏。王對駕車的說：「我受重傷了，你掉過車來，載我離開戰場！」
1KGS|22|35|那日，戰況越來越猛，有人扶著王站在戰車上，面對 亞蘭 人。到了傍晚，王就死了，血從傷處流入車底。
1KGS|22|36|約在日落的時候，有喊聲傳遍軍中，說：「大家各歸本城，各歸本地吧！」
1KGS|22|37|王死了，人把他送到 撒瑪利亞 ，葬在 撒瑪利亞 。
1KGS|22|38|他們在 撒瑪利亞 的水池旁洗他的車，有狗來舔他的血，有妓女在那裏洗澡，正如耶和華所說的話。
1KGS|22|39|亞哈 其餘的事，凡他所做的、他所修造的象牙宮和所建築的一切城鎮，不都寫在《以色列諸王記》上嗎？
1KGS|22|40|亞哈 與他祖先同睡，他兒子 亞哈謝 接續他作王。
1KGS|22|41|以色列 王 亞哈 第四年， 亞撒 的兒子 約沙法 登基作 猶大 王。
1KGS|22|42|約沙法 登基的時候年三十五歲，在 耶路撒冷 作王二十五年。他母親名叫 阿蘇巴 ，是 示利希 的女兒。
1KGS|22|43|約沙法 效法他父親 亞撒 所行的道，不偏離左右，行耶和華眼中看為正的事。只是丘壇還沒有廢去，百姓仍在那裏獻祭燒香。
1KGS|22|44|約沙法 與 以色列 王和平相處。
1KGS|22|45|約沙法 其餘的事和他所行的英勇事蹟，以及他的戰役，不都寫在《猶大列王記》上嗎？
1KGS|22|46|約沙法 把他父親 亞撒 的日子所剩下男的廟妓都從國中除去了。
1KGS|22|47|那時 以東 沒有立王，由總督治理。
1KGS|22|48|約沙法 造了 他施 船隻，要往 俄斐 去，把金子運來，卻沒有啟航，因為船在 以旬‧迦別 毀壞了。
1KGS|22|49|亞哈 的兒子 亞哈謝 對 約沙法 說：「讓我的僕人和你的僕人坐船同去吧！」 約沙法 卻不肯。
1KGS|22|50|約沙法 與他祖先同睡，與他祖先同葬在 大衛城 ，他兒子 約蘭 接續他作王。
1KGS|22|51|猶大 王 約沙法 第十七年， 亞哈 的兒子 亞哈謝 在 撒瑪利亞 登基作 以色列 王；他作 以色列 王二年。
1KGS|22|52|他行耶和華眼中看為惡的事，行他父母的道，又行 尼八 的兒子 耶羅波安 的道，使 以色列 陷入罪裏。
1KGS|22|53|他事奉 巴力 ，敬拜它，惹耶和華－ 以色列 的上帝發怒，正如他父親一切所行的。
