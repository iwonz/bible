PS|1|1|Блажен муж, который не ходит на совет нечестивых и не стоит на пути грешных и не сидит в собрании развратителей,
PS|1|2|но в законе Господа воля его, и о законе Его размышляет он день и ночь!
PS|1|3|И будет он как дерево, посаженное при потоках вод, которое приносит плод свой во время свое, и лист которого не вянет; и во всем, что он ни делает, успеет.
PS|1|4|Не так – нечестивые; но они – как прах, возметаемый ветром.
PS|1|5|Потому не устоят нечестивые на суде, и грешники – в собрании праведных.
PS|1|6|Ибо знает Господь путь праведных, а путь нечестивых погибнет.
PS|2|1|Псалом Давида. Зачем мятутся народы, и племена замышляют тщетное?
PS|2|2|Восстают цари земли, и князья совещаются вместе против Господа и против Помазанника Его.
PS|2|3|"Расторгнем узы их, и свергнем с себя оковы их".
PS|2|4|Живущий на небесах посмеется, Господь поругается им.
PS|2|5|Тогда скажет им во гневе Своем и яростью Своею приведет их в смятение:
PS|2|6|"Я помазал Царя Моего над Сионом, святою горою Моею;
PS|2|7|возвещу определение: Господь сказал Мне: Ты Сын Мой; Я ныне родил Тебя;
PS|2|8|проси у Меня, и дам народы в наследие Тебе и пределы земли во владение Тебе;
PS|2|9|Ты поразишь их жезлом железным; сокрушишь их, как сосуд горшечника".
PS|2|10|Итак вразумитесь, цари; научитесь, судьи земли!
PS|2|11|Служите Господу со страхом и радуйтесь с трепетом.
PS|2|12|Почтите Сына, чтобы Он не прогневался, и чтобы вам не погибнуть в пути [вашем], ибо гнев Его возгорится вскоре. Блаженны все, уповающие на Него.
PS|3|1|Псалом Давида, когда он бежал от Авессалома, сына своего.
PS|3|2|Господи! как умножились враги мои! Многие восстают на меня
PS|3|3|многие говорят душе моей: "нет ему спасения в Боге".
PS|3|4|Но Ты, Господи, щит предо мною, слава моя, и Ты возносишь голову мою.
PS|3|5|Гласом моим взываю к Господу, и Он слышит меня со святой горы Своей.
PS|3|6|Ложусь я, сплю и встаю, ибо Господь защищает меня.
PS|3|7|Не убоюсь тем народа, которые со всех сторон ополчились на меня.
PS|3|8|Восстань, Господи! спаси меня, Боже мой! ибо Ты поражаешь в ланиту всех врагов моих; сокрушаешь зубы нечестивых.
PS|3|9|От Господа спасение. Над народом Твоим благословение Твое.
PS|4|1|Начальнику хора. На струнных [орудиях]. Псалом Давида.
PS|4|2|Когда я взываю, услышь меня, Боже правды моей! В тесноте Ты давал мне простор. Помилуй меня и услышь молитву мою.
PS|4|3|Сыны мужей! доколе слава моя будет в поругании? доколе будете любить суету и искать лжи?
PS|4|4|Знайте, что Господь отделил для Себя святаго Своего; Господь слышит, когда я призываю Его.
PS|4|5|Гневаясь, не согрешайте: размыслите в сердцах ваших на ложах ваших, и утишитесь;
PS|4|6|приносите жертвы правды и уповайте на Господа.
PS|4|7|Многие говорят: "кто покажет нам благо?" Яви нам свет лица Твоего, Господи!
PS|4|8|Ты исполнил сердце мое веселием с того времени, как у них хлеб и вино умножились.
PS|4|9|Спокойно ложусь я и сплю, ибо Ты, Господи, един даешь мне жить в безопасности.
PS|5|1|Начальнику хора. На духовых [орудиях]. Псалом Давида.
PS|5|2|Услышь, Господи, слова мои, уразумей помышления мои.
PS|5|3|Внемли гласу вопля моего, Царь мой и Бог мой! ибо я к Тебе молюсь.
PS|5|4|Господи! рано услышь голос мой, – рано предстану пред Тобою, и буду ожидать,
PS|5|5|ибо Ты Бог, не любящий беззакония; у Тебя не водворится злой;
PS|5|6|нечестивые не пребудут пред очами Твоими: Ты ненавидишь всех, делающих беззаконие.
PS|5|7|Ты погубишь говорящих ложь; кровожадного и коварного гнушается Господь.
PS|5|8|А я, по множеству милости Твоей, войду в дом Твой, поклонюсь святому храму Твоему в страхе Твоем.
PS|5|9|Господи! путеводи меня в правде Твоей, ради врагов моих; уровняй предо мною путь Твой.
PS|5|10|Ибо нет в устах их истины: сердце их – пагуба, гортань их – открытый гроб, языком своим льстят.
PS|5|11|Осуди их, Боже, да падут они от замыслов своих; по множеству нечестия их, отвергни их, ибо они возмутились против Тебя.
PS|5|12|И возрадуются все уповающие на Тебя, вечно будут ликовать, и Ты будешь покровительствовать им; и будут хвалиться Тобою любящие имя Твое.
PS|5|13|Ибо Ты благословляешь праведника, Господи; благоволением, как щитом, венчаешь его.
PS|6|1|Начальнику хора. На восьмиструнном. Псалом Давида.
PS|6|2|Господи! не в ярости Твоей обличай меня и не во гневе Твоем наказывай меня.
PS|6|3|Помилуй меня, Господи, ибо я немощен; исцели меня, Господи, ибо кости мои потрясены;
PS|6|4|и душа моя сильно потрясена; Ты же, Господи, доколе?
PS|6|5|Обратись, Господи, избавь душу мою, спаси меня ради милости Твоей,
PS|6|6|ибо в смерти нет памятования о Тебе: во гробе кто будет славить Тебя?
PS|6|7|Утомлен я воздыханиями моими: каждую ночь омываю ложе мое, слезами моими омочаю постель мою.
PS|6|8|Иссохло от печали око мое, обветшало от всех врагов моих.
PS|6|9|Удалитесь от меня все, делающие беззаконие, ибо услышал Господь голос плача моего,
PS|6|10|услышал Господь моление мое; Господь примет молитву мою.
PS|6|11|Да будут постыжены и жестоко поражены все враги мои; да возвратятся и постыдятся мгновенно.
PS|7|1|Плачевная песнь, которую Давид воспел Господу по делу Хуса, из племени Вениаминова.
PS|7|2|Господи, Боже мой! на Тебя я уповаю; спаси меня от всех гонителей моих и избавь меня;
PS|7|3|да не исторгнет он, подобно льву, души моей, терзая, когда нет избавляющего.
PS|7|4|Господи, Боже мой! если я что сделал, если есть неправда в руках моих,
PS|7|5|если я платил злом тому, кто был со мною в мире, – я, который спасал даже того, кто без причины стал моим врагом, –
PS|7|6|то пусть враг преследует душу мою и настигнет, пусть втопчет в землю жизнь мою, и славу мою повергнет в прах.
PS|7|7|Восстань, Господи, во гневе Твоем; подвигнись против неистовства врагов моих, пробудись для меня на суд, который Ты заповедал, –
PS|7|8|сонм людей станет вокруг Тебя; над ним поднимись на высоту.
PS|7|9|Господь судит народы. Суди меня, Господи, по правде моей и по непорочности моей во мне.
PS|7|10|Да прекратится злоба нечестивых, а праведника подкрепи, ибо Ты испытуешь сердца и утробы, праведный Боже!
PS|7|11|Щит мой в Боге, спасающем правых сердцем.
PS|7|12|Бог – судия праведный, и Бог, всякий день строго взыскивающий,
PS|7|13|если [кто] не обращается. Он изощряет Свой меч, напрягает лук Свой и направляет его,
PS|7|14|приготовляет для него сосуды смерти, стрелы Свои делает палящими.
PS|7|15|Вот, [нечестивый] зачал неправду, был чреват злобою и родил себе ложь;
PS|7|16|рыл ров, и выкопал его, и упал в яму, которую приготовил:
PS|7|17|злоба его обратится на его голову, и злодейство его упадет на его темя.
PS|7|18|Славлю Господа по правде Его и пою имени Господа Всевышнего.
PS|8|1|Начальнику хора. На Гефском [орудии]. Псалом Давида.
PS|8|2|Господи, Боже наш! как величественно имя Твое по всей земле! Слава Твоя простирается превыше небес!
PS|8|3|Из уст младенцев и грудных детей Ты устроил хвалу, ради врагов Твоих, дабы сделать безмолвным врага и мстителя.
PS|8|4|Когда взираю я на небеса Твои – дело Твоих перстов, на луну и звезды, которые Ты поставил,
PS|8|5|то что [есть] человек, что Ты помнишь его, и сын человеческий, что Ты посещаешь его?
PS|8|6|Не много Ты умалил его пред Ангелами: славою и честью увенчал его;
PS|8|7|поставил его владыкою над делами рук Твоих; все положил под ноги его:
PS|8|8|овец и волов всех, и также полевых зверей,
PS|8|9|птиц небесных и рыб морских, все, преходящее морскими стезями.
PS|8|10|Господи, Боже наш! Как величественно имя Твое по всей земле!
PS|9|1|Начальнику хора. По смерти Лабена. Псалом Давида.
PS|9|2|Буду славить [Тебя], Господи, всем сердцем моим, возвещать все чудеса Твои.
PS|9|3|Буду радоваться и торжествовать о Тебе, петь имени Твоему, Всевышний.
PS|9|4|Когда враги мои обращены назад, то преткнутся и погибнут пред лицем Твоим,
PS|9|5|ибо Ты производил мой суд и мою тяжбу; Ты воссел на престоле, Судия праведный.
PS|9|6|Ты вознегодовал на народы, погубил нечестивого, имя их изгладил на веки и веки.
PS|9|7|У врага совсем не стало оружия, и города Ты разрушил; погибла память их с ними.
PS|9|8|Но Господь пребывает вовек; Он приготовил для суда престол Свой,
PS|9|9|и Он будет судить вселенную по правде, совершит суд над народами по правоте.
PS|9|10|И будет Господь прибежищем угнетенному, прибежищем во времена скорби;
PS|9|11|и будут уповать на Тебя знающие имя Твое, потому что Ты не оставляешь ищущих Тебя, Господи.
PS|9|12|Пойте Господу, живущему на Сионе, возвещайте между народами дела Его,
PS|9|13|ибо Он взыскивает за кровь; помнит их, не забывает вопля угнетенных.
PS|9|14|Помилуй меня, Господи; воззри на страдание мое от ненавидящих меня, – Ты, Который возносишь меня от врат смерти,
PS|9|15|чтобы я возвещал все хвалы Твои во вратах дщери Сионовой: буду радоваться о спасении Твоем.
PS|9|16|Обрушились народы в яму, которую выкопали; в сети, которую скрыли они, запуталась нога их.
PS|9|17|Познан был Господь по суду, который Он совершил; нечестивый уловлен делами рук своих.
PS|9|18|Да обратятся нечестивые в ад, – все народы, забывающие Бога.
PS|9|19|Ибо не навсегда забыт будет нищий, и надежда бедных не до конца погибнет.
PS|9|20|Восстань, Господи, да не преобладает человек, да судятся народы пред лицем Твоим.
PS|9|21|Наведи, Господи, страх на них; да знают народы, что человеки они.
PS|9|22|Для чего, Господи, стоишь вдали, скрываешь Себя во время скорби?
PS|9|23|По гордости своей нечестивый преследует бедного: да уловятся они ухищрениями, которые сами вымышляют.
PS|9|24|Ибо нечестивый хвалится похотью души своей; корыстолюбец ублажает себя.
PS|9|25|В надмении своем нечестивый пренебрегает Господа: "не взыщет"; во всех помыслах его: "нет Бога!"
PS|9|26|Во всякое время пути его гибельны; суды Твои далеки для него; на всех врагов своих он смотрит с пренебрежением;
PS|9|27|говорит в сердце своем: "не поколеблюсь; в род и род не приключится [мне] зла";
PS|9|28|уста его полны проклятия, коварства и лжи; под языком – его мучение и пагуба;
PS|9|29|сидит в засаде за двором, в потаенных местах убивает невинного; глаза его подсматривают за бедным;
PS|9|30|подстерегает в потаенном месте, как лев в логовище; подстерегает в засаде, чтобы схватить бедного; хватает бедного, увлекая в сети свои;
PS|9|31|сгибается, прилегает, – и бедные падают в сильные когти его;
PS|9|32|говорит в сердце своем: "забыл Бог, закрыл лице Свое, не увидит никогда".
PS|9|33|Восстань, Господи, Боже [мой], вознеси руку Твою, не забудь угнетенных.
PS|9|34|Зачем нечестивый пренебрегает Бога, говоря в сердце своем: "Ты не взыщешь"?
PS|9|35|Ты видишь, ибо Ты взираешь на обиды и притеснения, чтобы воздать Твоею рукою. Тебе предает себя бедный; сироте Ты помощник.
PS|9|36|Сокруши мышцу нечестивому и злому, так чтобы искать и не найти его нечестия.
PS|9|37|Господь – царь на веки, навсегда; исчезнут язычники с земли Его.
PS|9|38|Господи! Ты слышишь желания смиренных; укрепи сердце их; открой ухо Твое,
PS|9|39|чтобы дать суд сироте и угнетенному, да не устрашает более человек на земле.
PS|10|1|Начальнику хора. Псалом Давида. На Господа уповаю; как же вы говорите душе моей: "улетай на гору вашу, [как] птица"?
PS|10|2|Ибо вот, нечестивые натянули лук, стрелу свою приложили к тетиве, чтобы во тьме стрелять в правых сердцем.
PS|10|3|Когда разрушены основания, что сделает праведник?
PS|10|4|Господь во святом храме Своем, Господь, – престол Его на небесах, очи Его зрят; вежды Его испытывают сынов человеческих.
PS|10|5|Господь испытывает праведного, а нечестивого и любящего насилие ненавидит душа Его.
PS|10|6|Дождем прольет Он на нечестивых горящие угли, огонь и серу; и палящий ветер – их доля из чаши;
PS|10|7|ибо Господь праведен, любит правду; лице Его видит праведника.
PS|11|1|Начальнику хора. На восьмиструнном. Псалом Давида.
PS|11|2|Спаси, Господи, ибо не стало праведного, ибо нет верных между сынами человеческими.
PS|11|3|Ложь говорит каждый своему ближнему; уста льстивы, говорят от сердца притворного.
PS|11|4|Истребит Господь все уста льстивые, язык велеречивый,
PS|11|5|[тех], которые говорят: "языком нашим пересилим, уста наши с нами; кто нам господин"?
PS|11|6|Ради страдания нищих и воздыхания бедных ныне восстану, говорит Господь, поставлю в безопасности того, кого уловить хотят.
PS|11|7|Слова Господни – слова чистые, серебро, очищенное от земли в горниле, семь раз переплавленное.
PS|11|8|Ты, Господи, сохранишь их, соблюдешь от рода сего вовек.
PS|11|9|Повсюду ходят нечестивые, когда ничтожные из сынов человеческих возвысились.
PS|12|1|Начальнику хора. Псалом Давида.
PS|12|2|Доколе, Господи, будешь забывать меня вконец, доколе будешь скрывать лице Твое от меня?
PS|12|3|Доколе мне слагать советы в душе моей, скорбь в сердце моем день [и ночь]? Доколе врагу моему возноситься надо мною?
PS|12|4|Призри, услышь меня, Господи Боже мой! Просвети очи мои, да не усну я [сном] смертным;
PS|12|5|да не скажет враг мой: "я одолел его". Да не возрадуются гонители мои, если я поколеблюсь.
PS|12|6|Я же уповаю на милость Твою; сердце мое возрадуется о спасении Твоем; воспою Господу, облагодетельствовавшему меня.
PS|13|1|Начальнику хора. Псалом Давида. Сказал безумец в сердце своем: "нет Бога". Они развратились, совершили гнусные дела; нет делающего добро.
PS|13|2|Господь с небес призрел на сынов человеческих, чтобы видеть, есть ли разумеющий, ищущий Бога.
PS|13|3|Все уклонились, сделались равно непотребными; нет делающего добро, нет ни одного.
PS|13|4|Неужели не вразумятся все, делающие беззаконие, съедающие народ мой, [как] едят хлеб, и не призывающие Господа?
PS|13|5|Там убоятся они страха, ибо Бог в роде праведных.
PS|13|6|Вы посмеялись над мыслью нищего, что Господь упование его.
PS|13|7|"Кто даст с Сиона спасение Израилю!" Когда Господь возвратит пленение народа Своего, тогда возрадуется Иаков и возвеселится Израиль.
PS|14|1|Псалом Давида. Господи! кто может пребывать в жилище Твоем? кто может обитать на святой горе Твоей?
PS|14|2|Тот, кто ходит непорочно и делает правду, и говорит истину в сердце своем;
PS|14|3|кто не клевещет языком своим, не делает искреннему своему зла и не принимает поношения на ближнего своего
PS|14|4|тот, в глазах которого презрен отверженный, но который боящихся Господа славит; кто клянется, [хотя бы] злому, и не изменяет;
PS|14|5|кто серебра своего не отдает в рост и не принимает даров против невинного. Поступающий так не поколеблется вовек.
PS|15|1|Песнь Давида. Храни меня, Боже, ибо я на Тебя уповаю.
PS|15|2|Я сказал Господу: Ты – Господь мой; блага мои Тебе не нужны.
PS|15|3|К святым, которые на земле, и к дивным [Твоим] – к ним все желание мое.
PS|15|4|Пусть умножаются скорби у тех, которые текут к [богу] чужому; я не возлию кровавых возлияний их и не помяну имен их устами моими.
PS|15|5|Господь есть часть наследия моего и чаши моей. Ты держишь жребий мой.
PS|15|6|Межи мои прошли по прекрасным [местам], и наследие мое приятно для меня.
PS|15|7|Благословлю Господа, вразумившего меня; даже и ночью учит меня внутренность моя.
PS|15|8|Всегда видел я пред собою Господа, ибо Он одесную меня; не поколеблюсь.
PS|15|9|От того возрадовалось сердце мое и возвеселился язык мой; даже и плоть моя успокоится в уповании,
PS|15|10|ибо Ты не оставишь души моей в аде и не дашь святому Твоему увидеть тление,
PS|15|11|Ты укажешь мне путь жизни: полнота радостей пред лицем Твоим, блаженство в деснице Твоей вовек.
PS|16|1|Молитва Давида. Услышь, Господи, правду, внемли воплю моему, прими мольбу из уст нелживых.
PS|16|2|От Твоего лица суд мне да изыдет; да воззрят очи Твои на правоту.
PS|16|3|Ты испытал сердце мое, посетил меня ночью, искусил меня и ничего не нашел; от мыслей моих не отступают уста мои.
PS|16|4|В делах человеческих, по слову уст Твоих, я охранял себя от путей притеснителя.
PS|16|5|Утверди шаги мои на путях Твоих, да не колеблются стопы мои.
PS|16|6|К Тебе взываю я, ибо Ты услышишь меня, Боже; приклони ухо Твое ко мне, услышь слова мои.
PS|16|7|Яви дивную милость Твою, Спаситель уповающих [на Тебя] от противящихся деснице Твоей.
PS|16|8|Храни меня, как зеницу ока; в тени крыл Твоих укрой меня
PS|16|9|от лица нечестивых, нападающих на меня, – от врагов души моей, окружающих меня:
PS|16|10|они заключились в туке своем, надменно говорят устами своими.
PS|16|11|На всяком шагу нашем ныне окружают нас; они устремили глаза свои, чтобы низложить [меня] на землю;
PS|16|12|они подобны льву, жаждущему добычи, подобны скимну, сидящему в местах скрытных.
PS|16|13|Восстань, Господи, предупреди их, низложи их. Избавь душу мою от нечестивого мечом Твоим,
PS|16|14|от людей – рукою Твоею, Господи, от людей мира, которых удел в [этой] жизни, которых чрево Ты наполняешь из сокровищниц Твоих; сыновья их сыты и оставят остаток детям своим.
PS|16|15|А я в правде буду взирать на лице Твое; пробудившись, буду насыщаться образом Твоим.
PS|17|1|Начальнику хора. Раба Господня Давида, который произнес слова песни сей к Господу, когда Господь избавил его от рук всех врагов его и от руки Саула. И он сказал:
PS|17|2|Возлюблю тебя, Господи, крепость моя!
PS|17|3|Господь – твердыня моя и прибежище мое, Избавитель мой, Бог мой, – скала моя; на Него я уповаю; щит мой, рог спасения моего и убежище мое.
PS|17|4|Призову достопоклоняемого Господа и от врагов моих спасусь.
PS|17|5|Объяли меня муки смертные, и потоки беззакония устрашили меня;
PS|17|6|цепи ада облегли меня, и сети смерти опутали меня.
PS|17|7|В тесноте моей я призвал Господа и к Богу моему воззвал. И Он услышал от чертога Своего голос мой, и вопль мой дошел до слуха Его.
PS|17|8|Потряслась и всколебалась земля, дрогнули и подвиглись основания гор, ибо разгневался [Бог];
PS|17|9|поднялся дым от гнева Его и из уст Его огонь поядающий; горячие угли [сыпались] от Него.
PS|17|10|Наклонил Он небеса и сошел, – и мрак под ногами Его.
PS|17|11|И воссел на Херувимов и полетел, и понесся на крыльях ветра.
PS|17|12|И мрак сделал покровом Своим, сению вокруг Себя мрак вод, облаков воздушных.
PS|17|13|От блистания пред Ним бежали облака Его, град и угли огненные.
PS|17|14|Возгремел на небесах Господь, и Всевышний дал глас Свой, град и угли огненные.
PS|17|15|Пустил стрелы Свои и рассеял их, множество молний, и рассыпал их.
PS|17|16|И явились источники вод, и открылись основания вселенной от грозного [гласа] Твоего, Господи, от дуновения духа гнева Твоего.
PS|17|17|Он простер [руку] с высоты и взял меня, и извлек меня из вод многих;
PS|17|18|избавил меня от врага моего сильного и от ненавидящих меня, которые были сильнее меня.
PS|17|19|Они восстали на меня в день бедствия моего, но Господь был мне опорою.
PS|17|20|Он вывел меня на пространное место и избавил меня, ибо Он благоволит ко мне.
PS|17|21|Воздал мне Господь по правде моей, по чистоте рук моих вознаградил меня,
PS|17|22|ибо я хранил пути Господни и не был нечестивым пред Богом моим;
PS|17|23|ибо все заповеди Его предо мною, и от уставов Его я не отступал.
PS|17|24|Я был непорочен пред Ним и остерегался, чтобы не согрешить мне;
PS|17|25|и воздал мне Господь по правде моей, по чистоте рук моих пред очами Его.
PS|17|26|С милостивым Ты поступаешь милостиво, с мужем искренним – искренно,
PS|17|27|с чистым – чисто, а с лукавым – по лукавству его,
PS|17|28|ибо Ты людей угнетенных спасаешь, а очи надменные унижаешь.
PS|17|29|Ты возжигаешь светильник мой, Господи; Бог мой просвещает тьму мою.
PS|17|30|С Тобою я поражаю войско, с Богом моим восхожу на стену.
PS|17|31|Бог! – Непорочен путь Его, чисто слово Господа; щит Он для всех, уповающих на Него.
PS|17|32|Ибо кто Бог, кроме Господа, и кто защита, кроме Бога нашего?
PS|17|33|Бог препоясывает меня силою и устрояет мне верный путь;
PS|17|34|делает ноги мои, как оленьи, и на высотах моих поставляет меня;
PS|17|35|научает руки мои брани, и мышцы мои сокрушают медный лук.
PS|17|36|Ты дал мне щит спасения Твоего, и десница Твоя поддерживает меня, и милость Твоя возвеличивает меня.
PS|17|37|Ты расширяешь шаг мой подо мною, и не колеблются ноги мои.
PS|17|38|Я преследую врагов моих и настигаю их, и не возвращаюсь, доколе не истреблю их;
PS|17|39|поражаю их, и они не могут встать, падают под ноги мои,
PS|17|40|ибо Ты препоясал меня силою для войны и низложил под ноги мои восставших на меня;
PS|17|41|Ты обратил ко мне тыл врагов моих, и я истребляю ненавидящих меня:
PS|17|42|они вопиют, но нет спасающего; ко Господу, – но Он не внемлет им;
PS|17|43|я рассеваю их, как прах пред лицем ветра, как уличную грязь попираю их.
PS|17|44|Ты избавил меня от мятежа народа, поставил меня главою иноплеменников; народ, которого я не знал, служит мне;
PS|17|45|по одному слуху о мне повинуются мне; иноплеменники ласкательствуют предо мною;
PS|17|46|иноплеменники бледнеют и трепещут в укреплениях своих.
PS|17|47|Жив Господь и благословен защитник мой! Да будет превознесен Бог спасения моего,
PS|17|48|Бог, мстящий за меня и покоряющий мне народы,
PS|17|49|и избавляющий меня от врагов моих! Ты вознес меня над восстающими против меня и от человека жестокого избавил меня.
PS|17|50|За то буду славить Тебя, Господи, между иноплеменниками и буду петь имени Твоему,
PS|17|51|величественно спасающий царя и творящий милость помазаннику Твоему Давиду и потомству его вовеки.
PS|18|1|Начальнику хора. Псалом Давида.
PS|18|2|Небеса проповедуют славу Божию, и о делах рук Его вещает твердь.
PS|18|3|День дню передает речь, и ночь ночи открывает знание.
PS|18|4|Нет языка, и нет наречия, где не слышался бы голос их.
PS|18|5|По всей земле проходит звук их, и до пределов вселенной слова их. Он поставил в них жилище солнцу,
PS|18|6|и оно выходит, как жених из брачного чертога своего, радуется, как исполин, пробежать поприще:
PS|18|7|от края небес исход его, и шествие его до края их, и ничто не укрыто от теплоты его.
PS|18|8|Закон Господа совершен, укрепляет душу; откровение Господа верно, умудряет простых.
PS|18|9|Повеления Господа праведны, веселят сердце; заповедь Господа светла, просвещает очи.
PS|18|10|Страх Господень чист, пребывает вовек. Суды Господни истина, все праведны;
PS|18|11|они вожделеннее золота и даже множества золота чистого, слаще меда и капель сота;
PS|18|12|и раб Твой охраняется ими, в соблюдении их великая награда.
PS|18|13|Кто усмотрит погрешности свои? От тайных [моих] очисти меня
PS|18|14|и от умышленных удержи раба Твоего, чтобы не возобладали мною. Тогда я буду непорочен и чист от великого развращения.
PS|18|15|Да будут слова уст моих и помышление сердца моего благоугодны пред Тобою, Господи, твердыня моя и Избавитель мой!
PS|19|1|Начальнику хора. Псалом Давида.
PS|19|2|Да услышит тебя Господь в день печали, да защитит тебя имя Бога Иаковлева.
PS|19|3|Да пошлет тебе помощь из Святилища и с Сиона да подкрепит тебя.
PS|19|4|Да воспомянет все жертвоприношения твои и всесожжение твое да соделает тучным.
PS|19|5|Да даст тебе по сердцу твоему и все намерения твои да исполнит.
PS|19|6|Мы возрадуемся о спасении твоем и во имя Бога нашего поднимем знамя. Да исполнит Господь все прошения твои.
PS|19|7|Ныне познал я, что Господь спасает помазанника Своего, отвечает ему со святых небес Своих могуществом спасающей десницы Своей.
PS|19|8|Иные колесницами, иные конями, а мы именем Господа Бога нашего хвалимся:
PS|19|9|они поколебались и пали, а мы встали и стоим прямо.
PS|19|10|Господи! спаси царя и услышь нас, когда будем взывать [к Тебе].
PS|20|1|Начальнику хора. Псалом Давида.
PS|20|2|Господи! силою Твоею веселится царь и о спасении Твоем безмерно радуется.
PS|20|3|Ты дал ему, чего желало сердце его, и прошения уст его не отринул,
PS|20|4|ибо Ты встретил его благословениями благости, возложил на голову его венец из чистого золота.
PS|20|5|Он просил у Тебя жизни; Ты дал ему долгоденствие на век и век.
PS|20|6|Велика слава его в спасении Твоем; Ты возложил на него честь и величие.
PS|20|7|Ты положил на него благословения на веки, возвеселил его радостью лица Твоего,
PS|20|8|ибо царь уповает на Господа, и во благости Всевышнего не поколеблется.
PS|20|9|Рука Твоя найдет всех врагов Твоих, десница Твоя найдет ненавидящих Тебя.
PS|20|10|Во время гнева Твоего Ты сделаешь их, как печь огненную; во гневе Своем Господь погубит их, и пожрет их огонь.
PS|20|11|Ты истребишь плод их с земли и семя их – из среды сынов человеческих,
PS|20|12|ибо они предприняли против Тебя злое, составили замыслы, но не могли [выполнить их].
PS|20|13|Ты поставишь их целью, из луков Твоих пустишь стрелы в лице их.
PS|20|14|Вознесись, Господи, силою Твоею: мы будем воспевать и прославлять Твое могущество.
PS|21|1|Начальнику хора. При появлении зари. Псалом Давида.
PS|21|2|Боже мой! Боже мой! для чего Ты оставил меня? Далеки от спасения моего слова вопля моего.
PS|21|3|Боже мой! я вопию днем, – и Ты не внемлешь мне, ночью, – и нет мне успокоения.
PS|21|4|Но Ты, Святый, живешь среди славословий Израиля.
PS|21|5|На Тебя уповали отцы наши; уповали, и Ты избавлял их;
PS|21|6|к Тебе взывали они, и были спасаемы; на Тебя уповали, и не оставались в стыде.
PS|21|7|Я же червь, а не человек, поношение у людей и презрение в народе.
PS|21|8|Все, видящие меня, ругаются надо мною, говорят устами, кивая головою:
PS|21|9|"он уповал на Господа; пусть избавит его, пусть спасет, если он угоден Ему".
PS|21|10|Но Ты извел меня из чрева, вложил в меня упование у грудей матери моей.
PS|21|11|На Тебя оставлен я от утробы; от чрева матери моей Ты – Бог мой.
PS|21|12|Не удаляйся от меня, ибо скорбь близка, а помощника нет.
PS|21|13|Множество тельцов обступили меня; тучные Васанские окружили меня,
PS|21|14|раскрыли на меня пасть свою, как лев, алчущий добычи и рыкающий.
PS|21|15|Я пролился, как вода; все кости мои рассыпались; сердце мое сделалось, как воск, растаяло посреди внутренности моей.
PS|21|16|Сила моя иссохла, как черепок; язык мой прильпнул к гортани моей, и Ты свел меня к персти смертной.
PS|21|17|Ибо псы окружили меня, скопище злых обступило меня, пронзили руки мои и ноги мои.
PS|21|18|Можно было бы перечесть все кости мои; а они смотрят и делают из меня зрелище;
PS|21|19|делят ризы мои между собою и об одежде моей бросают жребий.
PS|21|20|Но Ты, Господи, не удаляйся от меня; сила моя! поспеши на помощь мне;
PS|21|21|избавь от меча душу мою и от псов одинокую мою;
PS|21|22|спаси меня от пасти льва и от рогов единорогов, услышав, [избавь] меня.
PS|21|23|Буду возвещать имя Твое братьям моим, посреди собрания восхвалять Тебя.
PS|21|24|Боящиеся Господа! восхвалите Его. Все семя Иакова! прославь Его. Да благоговеет пред Ним все семя Израиля,
PS|21|25|ибо Он не презрел и не пренебрег скорби страждущего, не скрыл от него лица Своего, но услышал его, когда сей воззвал к Нему.
PS|21|26|О Тебе хвала моя в собрании великом; воздам обеты мои пред боящимися Его.
PS|21|27|Да едят бедные и насыщаются; да восхвалят Господа ищущие Его; да живут сердца ваши во веки!
PS|21|28|Вспомнят, и обратятся к Господу все концы земли, и поклонятся пред Тобою все племена язычников,
PS|21|29|ибо Господне есть царство, и Он – Владыка над народами.
PS|21|30|Будут есть и поклоняться все тучные земли; преклонятся пред Ним все нисходящие в персть и не могущие сохранить жизни своей.
PS|21|31|Потомство [мое] будет служить Ему, и будет называться Господним вовек:
PS|21|32|придут и будут возвещать правду Его людям, которые родятся, что сотворил Господь.
PS|22|1|Псалом Давида. Господь – Пастырь мой; я ни в чем не буду нуждаться:
PS|22|2|Он покоит меня на злачных пажитях и водит меня к водам тихим,
PS|22|3|подкрепляет душу мою, направляет меня на стези правды ради имени Своего.
PS|22|4|Если я пойду и долиною смертной тени, не убоюсь зла, потому что Ты со мной; Твой жезл и Твой посох – они успокаивают меня.
PS|22|5|Ты приготовил предо мною трапезу в виду врагов моих; умастил елеем голову мою; чаша моя преисполнена.
PS|22|6|Так, благость и милость да сопровождают меня во все дни жизни моей, и я пребуду в доме Господнем многие дни.
PS|23|1|Псалом Давида. Господня – земля и что наполняет ее, вселенная и все живущее в ней,
PS|23|2|ибо Он основал ее на морях и на реках утвердил ее.
PS|23|3|Кто взойдет на гору Господню, или кто станет на святом месте Его?
PS|23|4|Тот, у которого руки неповинны и сердце чисто, кто не клялся душею своею напрасно и не божился ложно, –
PS|23|5|[тот] получит благословение от Господа и милость от Бога, Спасителя своего.
PS|23|6|Таков род ищущих Его, ищущих лица Твоего, Боже Иакова!
PS|23|7|Поднимите, врата, верхи ваши, и поднимитесь, двери вечные, и войдет Царь славы!
PS|23|8|Кто сей Царь славы? – Господь крепкий и сильный, Господь, сильный в брани.
PS|23|9|Поднимите, врата, верхи ваши, и поднимитесь, двери вечные, и войдет Царь славы!
PS|23|10|Кто сей Царь славы? – Господь сил, Он – царь славы.
PS|24|1|Псалом Давида. К Тебе, Господи, возношу душу мою.
PS|24|2|Боже мой! на Тебя уповаю, да не постыжусь, да не восторжествуют надо мною враги мои,
PS|24|3|да не постыдятся и все надеющиеся на Тебя: да постыдятся беззаконнующие втуне.
PS|24|4|Укажи мне, Господи, пути Твои и научи меня стезям Твоим.
PS|24|5|Направь меня на истину Твою и научи меня, ибо Ты Бог спасения моего; на Тебя надеюсь всякий день.
PS|24|6|Вспомни щедроты Твои, Господи, и милости Твои, ибо они от века.
PS|24|7|Грехов юности моей и преступлений моих не вспоминай; по милости Твоей вспомни меня Ты, ради благости Твоей, Господи!
PS|24|8|Благ и праведен Господь, посему наставляет грешников на путь,
PS|24|9|направляет кротких к правде, и научает кротких путям Своим.
PS|24|10|Все пути Господни – милость и истина к хранящим завет Его и откровения Его.
PS|24|11|Ради имени Твоего, Господи, прости согрешение мое, ибо велико оно.
PS|24|12|Кто есть человек, боящийся Господа? Ему укажет Он путь, который избрать.
PS|24|13|Душа его пребудет во благе, и семя его наследует землю.
PS|24|14|Тайна Господня – боящимся Его, и завет Свой Он открывает им.
PS|24|15|Очи мои всегда к Господу, ибо Он извлекает из сети ноги мои.
PS|24|16|Призри на меня и помилуй меня, ибо я одинок и угнетен.
PS|24|17|Скорби сердца моего умножились; выведи меня из бед моих,
PS|24|18|призри на страдание мое и на изнеможение мое и прости все грехи мои.
PS|24|19|Посмотри на врагов моих, как много их, и [какою] лютою ненавистью они ненавидят меня.
PS|24|20|Сохрани душу мою и избавь меня, да не постыжусь, что я на Тебя уповаю.
PS|24|21|Непорочность и правота да охраняют меня, ибо я на Тебя надеюсь.
PS|24|22|Избавь, Боже, Израиля от всех скорбей его.
PS|25|1|Псалом Давида. Рассуди меня, Господи, ибо я ходил в непорочности моей, и, уповая на Господа, не поколеблюсь.
PS|25|2|Искуси меня, Господи, и испытай меня; расплавь внутренности мои и сердце мое,
PS|25|3|ибо милость Твоя пред моими очами, и я ходил в истине Твоей,
PS|25|4|не сидел я с людьми лживыми, и с коварными не пойду;
PS|25|5|возненавидел я сборище злонамеренных, и с нечестивыми не сяду;
PS|25|6|буду омывать в невинности руки мои и обходить жертвенник Твой, Господи,
PS|25|7|чтобы возвещать гласом хвалы и поведать все чудеса Твои.
PS|25|8|Господи! возлюбил я обитель дома Твоего и место жилища славы Твоей.
PS|25|9|Не погуби души моей с грешниками и жизни моей с кровожадными,
PS|25|10|у которых в руках злодейство, и которых правая рука полна мздоимства.
PS|25|11|А я хожу в моей непорочности; избавь меня, и помилуй меня.
PS|25|12|Моя нога стоит на прямом [пути]; в собраниях благословлю Господа.
PS|26|1|Псалом Давида. Господь – свет мой и спасение мое: кого мне бояться? Господь крепость жизни моей: кого мне страшиться?
PS|26|2|Если будут наступать на меня злодеи, противники и враги мои, чтобы пожрать плоть мою, то они сами преткнутся и падут.
PS|26|3|Если ополчится против меня полк, не убоится сердце мое; если восстанет на меня война, и тогда буду надеяться.
PS|26|4|Одного просил я у Господа, того только ищу, чтобы пребывать мне в доме Господнем во все дни жизни моей, созерцать красоту Господню и посещать храм Его,
PS|26|5|ибо Он укрыл бы меня в скинии Своей в день бедствия, скрыл бы меня в потаенном месте селения Своего, вознес бы меня на скалу.
PS|26|6|Тогда вознеслась бы голова моя над врагами, окружающими меня; и я принес бы в Его скинии жертвы славословия, стал бы петь и воспевать пред Господом.
PS|26|7|Услышь, Господи, голос мой, которым я взываю, помилуй меня и внемли мне.
PS|26|8|Сердце мое говорит от Тебя: "ищите лица Моего"; и я буду искать лица Твоего, Господи.
PS|26|9|Не скрой от меня лица Твоего; не отринь во гневе раба Твоего. Ты был помощником моим; не отвергни меня и не оставь меня, Боже, Спаситель мой!
PS|26|10|ибо отец мой и мать моя оставили меня, но Господь примет меня.
PS|26|11|Научи меня, Господи, пути Твоему и наставь меня на стезю правды, ради врагов моих;
PS|26|12|не предавай меня на произвол врагам моим, ибо восстали на меня свидетели лживые и дышат злобою.
PS|26|13|Но я верую, что увижу благость Господа на земле живых.
PS|26|14|Надейся на Господа, мужайся, и да укрепляется сердце твое, и надейся на Господа.
PS|27|1|Псалом Давида. К тебе, Господи, взываю: твердыня моя! не будь безмолвен для меня, чтобы при безмолвии Твоем я не уподобился нисходящим в могилу.
PS|27|2|Услышь голос молений моих, когда я взываю к Тебе, когда поднимаю руки мои к святому храму Твоему.
PS|27|3|Не погуби меня с нечестивыми и с делающими неправду, которые с ближними своими говорят о мире, а в сердце у них зло.
PS|27|4|Воздай им по делам их, по злым поступкам их; по делам рук их воздай им, отдай им заслуженное ими.
PS|27|5|За то, что они невнимательны к действиям Господа и к делу рук Его, Он разрушит их и не созиждет их.
PS|27|6|Благословен Господь, ибо Он услышал голос молений моих.
PS|27|7|Господь – крепость моя и щит мой; на Него уповало сердце мое, и Он помог мне, и возрадовалось сердце мое; и я прославлю Его песнью моею.
PS|27|8|Господь – крепость народа Своего и спасительная защита помазанника Своего.
PS|27|9|Спаси народ Твой и благослови наследие Твое; паси их и возвышай их во веки!
PS|28|1|Псалом Давида. Воздайте Господу, сыны Божии, воздайте Господу славу и честь,
PS|28|2|воздайте Господу славу имени Его; поклонитесь Господу в благолепном святилище [Его].
PS|28|3|Глас Господень над водами; Бог славы возгремел, Господь над водами многими.
PS|28|4|Глас Господа силен, глас Господа величествен.
PS|28|5|Глас Господа сокрушает кедры; Господь сокрушает кедры Ливанские
PS|28|6|и заставляет их скакать подобно тельцу, Ливан и Сирион, подобно молодому единорогу.
PS|28|7|Глас Господа высекает пламень огня.
PS|28|8|Глас Господа потрясает пустыню; потрясает Господь пустыню Кадес.
PS|28|9|Глас Господа разрешает от бремени ланей и обнажает леса; и во храме Его все возвещает о [Его] славе.
PS|28|10|Господь восседал над потопом, и будет восседать Господь царем вовек.
PS|28|11|Господь даст силу народу Своему, Господь благословит народ Свой миром.
PS|29|1|Псалом Давида; песнь при обновлении дома.
PS|29|2|Превознесу Тебя, Господи, что Ты поднял меня и не дал моим врагам восторжествовать надо мною.
PS|29|3|Господи, Боже мой! я воззвал к Тебе, и Ты исцелил меня.
PS|29|4|Господи! Ты вывел из ада душу мою и оживил меня, чтобы я не сошел в могилу.
PS|29|5|Пойте Господу, святые Его, славьте память святыни Его,
PS|29|6|ибо на мгновение гнев Его, на [всю] жизнь благоволение Его: вечером водворяется плач, а на утро радость.
PS|29|7|И я говорил в благоденствии моем: "не поколеблюсь вовек".
PS|29|8|По благоволению Твоему, Господи, Ты укрепил гору мою; но Ты сокрыл лице Твое, [и] я смутился.
PS|29|9|[Тогда] к Тебе, Господи, взывал я, и Господа умолял:
PS|29|10|"что пользы в крови моей, когда я сойду в могилу? будет ли прах славить Тебя? будет ли возвещать истину Твою?
PS|29|11|услышь, Господи, и помилуй меня; Господи! будь мне помощником".
PS|29|12|И Ты обратил сетование мое в ликование, снял с меня вретище и препоясал меня веселием,
PS|29|13|да славит Тебя душа моя и да не умолкает. Господи, Боже мой! буду славить Тебя вечно.
PS|30|1|Начальнику хора. Псалом Давида.
PS|30|2|На Тебя, Господи, уповаю, да не постыжусь вовек; по правде Твоей избавь меня;
PS|30|3|приклони ко мне ухо Твое, поспеши избавить меня. Будь мне каменною твердынею, домом прибежища, чтобы спасти меня,
PS|30|4|ибо Ты каменная гора моя и ограда моя; ради имени Твоего води меня и управляй мною.
PS|30|5|Выведи меня из сети, которую тайно поставили мне, ибо Ты крепость моя.
PS|30|6|В Твою руку предаю дух мой; Ты избавлял меня, Господи, Боже истины.
PS|30|7|Ненавижу почитателей суетных идолов, но на Господа уповаю.
PS|30|8|Буду радоваться и веселиться о милости Твоей, потому что Ты призрел на бедствие мое, узнал горесть души моей
PS|30|9|и не предал меня в руки врага; поставил ноги мои на пространном месте.
PS|30|10|Помилуй меня, Господи, ибо тесно мне; иссохло от горести око мое, душа моя и утроба моя.
PS|30|11|Истощилась в печали жизнь моя и лета мои в стенаниях; изнемогла от грехов моих сила моя, и кости мои иссохли.
PS|30|12|От всех врагов моих я сделался поношением даже у соседей моих и страшилищем для знакомых моих; видящие меня на улице бегут от меня.
PS|30|13|Я забыт в сердцах, как мертвый; я – как сосуд разбитый,
PS|30|14|ибо слышу злоречие многих; отвсюду ужас, когда они сговариваются против меня, умышляют исторгнуть душу мою.
PS|30|15|А я на Тебя, Господи, уповаю; я говорю: Ты – мой Бог.
PS|30|16|В Твоей руке дни мои; избавь меня от руки врагов моих и от гонителей моих.
PS|30|17|Яви светлое лице Твое рабу Твоему; спаси меня милостью Твоею.
PS|30|18|Господи! да не постыжусь, что я к Тебе взываю; нечестивые же да посрамятся, да умолкнут в аде.
PS|30|19|Да онемеют уста лживые, которые против праведника говорят злое с гордостью и презреньем.
PS|30|20|Как много у Тебя благ, которые Ты хранишь для боящихся Тебя и которые приготовил уповающим на Тебя пред сынами человеческими!
PS|30|21|Ты укрываешь их под покровом лица Твоего от мятежей людских, скрываешь их под сенью от пререкания языков.
PS|30|22|Благословен Господь, что явил мне дивную милость Свою в укрепленном городе!
PS|30|23|В смятении моем я думал: "отвержен я от очей Твоих"; но Ты услышал голос молитвы моей, когда я воззвал к Тебе.
PS|30|24|Любите Господа, все праведные Его; Господь хранит верных и поступающим надменно воздает с избытком.
PS|30|25|Мужайтесь, и да укрепляется сердце ваше, все надеющиеся на Господа!
PS|31|1|Псалом Давида. Учение. Блажен, кому отпущены беззакония, и чьи грехи покрыты!
PS|31|2|Блажен человек, которому Господь не вменит греха, и в чьем духе нет лукавства!
PS|31|3|Когда я молчал, обветшали кости мои от вседневного стенания моего,
PS|31|4|ибо день и ночь тяготела надо мною рука Твоя; свежесть моя исчезла, как в летнюю засуху.
PS|31|5|Но я открыл Тебе грех мой и не скрыл беззакония моего; я сказал: "исповедаю Господу преступления мои", и Ты снял с меня вину греха моего.
PS|31|6|За то помолится Тебе каждый праведник во время благопотребное, и тогда разлитие многих вод не достигнет его.
PS|31|7|Ты покров мой: Ты охраняешь меня от скорби, окружаешь меня радостями избавления.
PS|31|8|"Вразумлю тебя, наставлю тебя на путь, по которому тебе идти; буду руководить тебя, око Мое над тобою".
PS|31|9|"Не будьте как конь, как лошак несмысленный, которых челюсти нужно обуздывать уздою и удилами, чтобы они покорялись тебе".
PS|31|10|Много скорбей нечестивому, а уповающего на Господа окружает милость.
PS|31|11|Веселитесь о Господе и радуйтесь, праведные; торжествуйте, все правые сердцем.
PS|32|1|Радуйтесь, праведные, о Господе: правым прилично славословить.
PS|32|2|Славьте Господа на гуслях, пойте Ему на десятиструнной псалтири;
PS|32|3|пойте Ему новую песнь; пойте Ему стройно, с восклицанием,
PS|32|4|ибо слово Господне право и все дела Его верны.
PS|32|5|Он любит правду и суд; милости Господней полна земля.
PS|32|6|Словом Господа сотворены небеса, и духом уст Его – все воинство их:
PS|32|7|Он собрал, будто груды, морские воды, положил бездны в хранилищах.
PS|32|8|Да боится Господа вся земля; да трепещут пред Ним все живущие во вселенной,
PS|32|9|ибо Он сказал, – и сделалось; Он повелел, – и явилось.
PS|32|10|Господь разрушает советы язычников, уничтожает замыслы народов.
PS|32|11|Совет же Господень стоит вовек; помышления сердца Его – в род и род.
PS|32|12|Блажен народ, у которого Господь есть Бог, – племя, которое Он избрал в наследие Себе.
PS|32|13|С небес призирает Господь, видит всех сынов человеческих;
PS|32|14|с престола, на котором восседает, Он призирает на всех, живущих на земле:
PS|32|15|Он создал сердца всех их и вникает во все дела их.
PS|32|16|Не спасется царь множеством воинства; исполина не защитит великая сила.
PS|32|17|Ненадежен конь для спасения, не избавит великою силою своею.
PS|32|18|Вот, око Господне над боящимися Его и уповающими на милость Его,
PS|32|19|что Он душу их спасет от смерти и во время голода пропитает их.
PS|32|20|Душа наша уповает на Господа: Он – помощь наша и защита наша;
PS|32|21|о Нем веселится сердце наше, ибо на святое имя Его мы уповали.
PS|32|22|Да будет милость Твоя, Господи, над нами, как мы уповаем на Тебя.
PS|33|1|Псалом Давида, когда он притворился безумным пред Авимелехом и был изгнан от него и удалился.
PS|33|2|Благословлю Господа во всякое время; хвала Ему непрестанно в устах моих.
PS|33|3|Господом будет хвалиться душа моя; услышат кроткие и возвеселятся.
PS|33|4|Величайте Господа со мною, и превознесем имя Его вместе.
PS|33|5|Я взыскал Господа, и Он услышал меня, и от всех опасностей моих избавил меня.
PS|33|6|Кто обращал взор к Нему, те просвещались, и лица их не постыдятся.
PS|33|7|Сей нищий воззвал, – и Господь услышал и спас его от всех бед его.
PS|33|8|Ангел Господень ополчается вокруг боящихся Его и избавляет их.
PS|33|9|Вкусите, и увидите, как благ Господь! Блажен человек, который уповает на Него!
PS|33|10|Бойтесь Господа, святые Его, ибо нет скудости у боящихся Его.
PS|33|11|Скимны бедствуют и терпят голод, а ищущие Господа не терпят нужды ни в каком благе.
PS|33|12|Придите, дети, послушайте меня: страху Господню научу вас.
PS|33|13|Хочет ли человек жить и любит ли долгоденствие, чтобы видеть благо?
PS|33|14|Удерживай язык свой от зла и уста свои от коварных слов.
PS|33|15|Уклоняйся от зла и делай добро; ищи мира и следуй за ним.
PS|33|16|Очи Господни [обращены] на праведников, и уши Его – к воплю их.
PS|33|17|Но лице Господне против делающих зло, чтобы истребить с земли память о них.
PS|33|18|Взывают [праведные], и Господь слышит, и от всех скорбей их избавляет их.
PS|33|19|Близок Господь к сокрушенным сердцем и смиренных духом спасет.
PS|33|20|Много скорбей у праведного, и от всех их избавит его Господь.
PS|33|21|Он хранит все кости его; ни одна из них не сокрушится.
PS|33|22|Убьет грешника зло, и ненавидящие праведного погибнут.
PS|33|23|Избавит Господь душу рабов Своих, и никто из уповающих на Него не погибнет.
PS|34|1|Псалом Давида. Учение. Вступись, Господи, в тяжбу с тяжущимися со мною, побори борющихся со мною;
PS|34|2|возьми щит и латы и восстань на помощь мне;
PS|34|3|обнажи мечь и прегради [путь] преследующим меня; скажи душе моей: "Я – спасение твое!"
PS|34|4|Да постыдятся и посрамятся ищущие души моей; да обратятся назад и покроются бесчестием умышляющие мне зло;
PS|34|5|да будут они, как прах пред лицем ветра, и Ангел Господень да прогоняет [их];
PS|34|6|да будет путь их темен и скользок, и Ангел Господень да преследует их,
PS|34|7|ибо они без вины скрыли для меня яму – сеть свою, без вины выкопали [ее] для души моей.
PS|34|8|Да придет на него гибель неожиданная, и сеть его, которую он скрыл [для меня], да уловит его самого; да впадет в нее на погибель.
PS|34|9|А моя душа будет радоваться о Господе, будет веселиться о спасении от Него.
PS|34|10|Все кости мои скажут: "Господи! кто подобен Тебе, избавляющему слабого от сильного, бедного и нищего от грабителя его?"
PS|34|11|Восстали на меня свидетели неправедные: чего я не знаю, о том допрашивают меня;
PS|34|12|воздают мне злом за добро, сиротством душе моей.
PS|34|13|Я во время болезни их одевался во вретище, изнурял постом душу мою, и молитва моя возвращалась в недро мое.
PS|34|14|Я поступал, как бы это был друг мой, брат мой; я ходил скорбный, с поникшею головою, как бы оплакивающий мать.
PS|34|15|А когда я претыкался, они радовались и собирались; собирались ругатели против меня, не знаю за что, поносили и не переставали;
PS|34|16|с лицемерными насмешниками скрежетали на меня зубами своими.
PS|34|17|Господи! долго ли будешь смотреть [на это]? Отведи душу мою от злодейств их, от львов – одинокую мою.
PS|34|18|Я прославлю Тебя в собрании великом, среди народа многочисленного восхвалю Тебя,
PS|34|19|чтобы не торжествовали надо мною враждующие против меня неправедно, и не перемигивались глазами ненавидящие меня безвинно;
PS|34|20|ибо не о мире говорят они, но против мирных земли составляют лукавые замыслы;
PS|34|21|расширяют на меня уста свои; говорят: "хорошо! хорошо! видел глаз наш".
PS|34|22|Ты видел, Господи, не умолчи; Господи! не удаляйся от меня.
PS|34|23|Подвигнись, пробудись для суда моего, для тяжбы моей, Боже мой и Господи мой!
PS|34|24|Суди меня по правде Твоей, Господи, Боже мой, и да не торжествуют они надо мною;
PS|34|25|да не говорят в сердце своем: "хорошо! по душе нашей!" Да не говорят: "мы поглотили его".
PS|34|26|Да постыдятся и посрамятся все, радующиеся моему несчастью; да облекутся в стыд и позор величающиеся надо мною.
PS|34|27|Да радуются и веселятся желающие правоты моей и говорят непрестанно: "да возвеличится Господь, желающий мира рабу Своему!"
PS|34|28|И язык мой будет проповедывать правду Твою и хвалу Твою всякий день.
PS|35|1|Начальнику хора. Раба Господня Давида.
PS|35|2|Нечестие беззаконного говорит в сердце моем: нет страха Божия пред глазами его,
PS|35|3|ибо он льстит себе в глазах своих, будто отыскивает беззаконие свое, чтобы возненавидеть его;
PS|35|4|слова уст его – неправда и лукавство; не хочет он вразумиться, чтобы делать добро;
PS|35|5|на ложе своем замышляет беззаконие, становится на путь недобрый, не гнушается злом.
PS|35|6|Господи! милость Твоя до небес, истина Твоя до облаков!
PS|35|7|Правда Твоя, как горы Божии, и судьбы Твои – бездна великая! Человеков и скотов хранишь Ты, Господи!
PS|35|8|Как драгоценна милость Твоя, Боже! Сыны человеческие в тени крыл Твоих покойны:
PS|35|9|насыщаются от тука дома Твоего, и из потока сладостей Твоих Ты напояешь их,
PS|35|10|ибо у Тебя источник жизни; во свете Твоем мы видим свет.
PS|35|11|Продли милость Твою к знающим Тебя и правду Твою к правым сердцем,
PS|35|12|да не наступит на меня нога гордыни, и рука грешника да не изгонит меня:
PS|35|13|там пали делающие беззаконие, низринуты и не могут встать.
PS|36|1|Псалом Давида. Не ревнуй злодеям, не завидуй делающим беззаконие,
PS|36|2|ибо они, как трава, скоро будут подкошены и, как зеленеющий злак, увянут.
PS|36|3|Уповай на Господа и делай добро; живи на земле и храни истину.
PS|36|4|Утешайся Господом, и Он исполнит желания сердца твоего.
PS|36|5|Предай Господу путь твой и уповай на Него, и Он совершит,
PS|36|6|и выведет, как свет, правду твою и справедливость твою, как полдень.
PS|36|7|Покорись Господу и надейся на Него. Не ревнуй успевающему в пути своем, человеку лукавствующему.
PS|36|8|Перестань гневаться и оставь ярость; не ревнуй до того, чтобы делать зло,
PS|36|9|ибо делающие зло истребятся, уповающие же на Господа наследуют землю.
PS|36|10|Еще немного, и не станет нечестивого; посмотришь на его место, и нет его.
PS|36|11|А кроткие наследуют землю и насладятся множеством мира.
PS|36|12|Нечестивый злоумышляет против праведника и скрежещет на него зубами своими:
PS|36|13|Господь же посмевается над ним, ибо видит, что приходит день его.
PS|36|14|Нечестивые обнажают меч и натягивают лук свой, чтобы низложить бедного и нищего, чтобы пронзить [идущих] прямым путем:
PS|36|15|меч их войдет в их же сердце, и луки их сокрушатся.
PS|36|16|Малое у праведника – лучше богатства многих нечестивых,
PS|36|17|ибо мышцы нечестивых сокрушатся, а праведников подкрепляет Господь.
PS|36|18|Господь знает дни непорочных, и достояние их пребудет вовек:
PS|36|19|не будут они постыжены во время лютое и во дни голода будут сыты;
PS|36|20|а нечестивые погибнут, и враги Господни, как тук агнцев, исчезнут, в дыме исчезнут.
PS|36|21|Нечестивый берет взаймы и не отдает, а праведник милует и дает,
PS|36|22|ибо благословенные Им наследуют землю, а проклятые Им истребятся.
PS|36|23|Господом утверждаются стопы [такого] человека, и Он благоволит к пути его:
PS|36|24|когда он будет падать, не упадет, ибо Господь поддерживает его за руку.
PS|36|25|Я был молод и состарился, и не видал праведника оставленным и потомков его просящими хлеба:
PS|36|26|он всякий день милует и взаймы дает, и потомство его в благословение будет.
PS|36|27|Уклоняйся от зла, и делай добро, и будешь жить вовек:
PS|36|28|ибо Господь любит правду и не оставляет святых Своих; вовек сохранятся они; и потомство нечестивых истребится.
PS|36|29|Праведники наследуют землю и будут жить на ней вовек.
PS|36|30|Уста праведника изрекают премудрость, и язык его произносит правду.
PS|36|31|Закон Бога его в сердце у него; не поколеблются стопы его.
PS|36|32|Нечестивый подсматривает за праведником и ищет умертвить его;
PS|36|33|но Господь не отдаст его в руки его и не допустит обвинить его, когда он будет судим.
PS|36|34|Уповай на Господа и держись пути Его: и Он вознесет тебя, чтобы ты наследовал землю; и когда будут истребляемы нечестивые, ты увидишь.
PS|36|35|Видел я нечестивца грозного, расширявшегося, подобно укоренившемуся многоветвистому дереву;
PS|36|36|но он прошел, и вот нет его; ищу его и не нахожу.
PS|36|37|Наблюдай за непорочным и смотри на праведного, ибо будущность [такого] человека есть мир;
PS|36|38|а беззаконники все истребятся; будущность нечестивых погибнет.
PS|36|39|От Господа спасение праведникам, Он – защита их во время скорби;
PS|36|40|и поможет им Господь и избавит их; избавит их от нечестивых и спасет их, ибо они на Него уповают.
PS|37|1|Псалом Давида. В воспоминание.
PS|37|2|Господи! не в ярости Твоей обличай меня и не во гневе Твоем наказывай меня,
PS|37|3|ибо стрелы Твои вонзились в меня, и рука Твоя тяготеет на мне.
PS|37|4|Нет целого места в плоти моей от гнева Твоего; нет мира в костях моих от грехов моих,
PS|37|5|ибо беззакония мои превысили голову мою, как тяжелое бремя отяготели на мне,
PS|37|6|смердят, гноятся раны мои от безумия моего.
PS|37|7|Я согбен и совсем поник, весь день сетуя хожу,
PS|37|8|ибо чресла мои полны воспалениями, и нет целого места в плоти моей.
PS|37|9|Я изнемог и сокрушен чрезмерно; кричу от терзания сердца моего.
PS|37|10|Господи! пред Тобою все желания мои, и воздыхание мое не сокрыто от Тебя.
PS|37|11|Сердце мое трепещет; оставила меня сила моя, и свет очей моих, – и того нет у меня.
PS|37|12|Друзья мои и искренние отступили от язвы моей, и ближние мои стоят вдали.
PS|37|13|Ищущие же души моей ставят сети, и желающие мне зла говорят о погибели [моей] и замышляют всякий день козни;
PS|37|14|а я, как глухой, не слышу, и как немой, который не открывает уст своих;
PS|37|15|и стал я, как человек, который не слышит и не имеет в устах своих ответа,
PS|37|16|ибо на Тебя, Господи, уповаю я; Ты услышишь, Господи, Боже мой.
PS|37|17|И я сказал: да не восторжествуют надо мною [враги мои]; когда колеблется нога моя, они величаются надо мною.
PS|37|18|Я близок к падению, и скорбь моя всегда предо мною.
PS|37|19|Беззаконие мое я сознаю, сокрушаюсь о грехе моем.
PS|37|20|А враги мои живут и укрепляются, и умножаются ненавидящие меня безвинно;
PS|37|21|и воздающие мне злом за добро враждуют против меня за то, что я следую добру.
PS|37|22|Не оставь меня, Господи, Боже мой! Не удаляйся от меня;
PS|37|23|поспеши на помощь мне, Господи, Спаситель мой!
PS|38|1|Начальнику хора, Идифуму. Псалом Давида.
PS|38|2|Я сказал: буду я наблюдать за путями моими, чтобы не согрешать мне языком моим; буду обуздывать уста мои, доколе нечестивый предо мною.
PS|38|3|Я был нем и безгласен, и молчал [даже] о добром; и скорбь моя подвиглась.
PS|38|4|Воспламенилось сердце мое во мне; в мыслях моих возгорелся огонь; я стал говорить языком моим:
PS|38|5|скажи мне, Господи, кончину мою и число дней моих, какое оно, дабы я знал, какой век мой.
PS|38|6|Вот, Ты дал мне дни, [как] пяди, и век мой как ничто пред Тобою. Подлинно, совершенная суета – всякий человек живущий.
PS|38|7|Подлинно, человек ходит подобно призраку; напрасно он суетится, собирает и не знает, кому достанется то.
PS|38|8|И ныне чего ожидать мне, Господи? надежда моя – на Тебя.
PS|38|9|От всех беззаконий моих избавь меня, не предавай меня на поругание безумному.
PS|38|10|Я стал нем, не открываю уст моих; потому что Ты соделал это.
PS|38|11|Отклони от меня удары Твои; я исчезаю от поражающей руки Твоей.
PS|38|12|Если Ты обличениями будешь наказывать человека за преступления, то рассыплется, как от моли, краса его. Так, суетен всякий человек!
PS|38|13|Услышь, Господи, молитву мою и внемли воплю моему; не будь безмолвен к слезам моим, ибо странник я у Тебя [и] пришлец, как и все отцы мои.
PS|38|14|Отступи от меня, чтобы я мог подкрепиться, прежде нежели отойду и не будет меня.
PS|39|1|Начальнику хора. Псалом Давида.
PS|39|2|Твердо уповал я на Господа, и Он приклонился ко мне и услышал вопль мой;
PS|39|3|извлек меня из страшного рва, из тинистого болота, и поставил на камне ноги мои и утвердил стопы мои;
PS|39|4|и вложил в уста мои новую песнь – хвалу Богу нашему. Увидят многие и убоятся и будут уповать на Господа.
PS|39|5|Блажен человек, который на Господа возлагает надежду свою и не обращается к гордым и к уклоняющимся ко лжи.
PS|39|6|Много соделал Ты, Господи, Боже мой: о чудесах и помышлениях Твоих о нас – кто уподобится Тебе! – хотел бы я проповедывать и говорить, но они превышают число.
PS|39|7|Жертвы и приношения Ты не восхотел; Ты открыл мне уши; всесожжения и жертвы за грех Ты не потребовал.
PS|39|8|Тогда я сказал: вот, иду; в свитке книжном написано о мне:
PS|39|9|я желаю исполнить волю Твою, Боже мой, и закон Твой у меня в сердце.
PS|39|10|Я возвещал правду Твою в собрании великом; я не возбранял устам моим: Ты, Господи, знаешь.
PS|39|11|Правды Твоей не скрывал в сердце моем, возвещал верность Твою и спасение Твое, не утаивал милости Твоей и истины Твоей пред собранием великим.
PS|39|12|Не удерживай, Господи, щедрот Твоих от меня; милость Твоя и истина Твоя да охраняют меня непрестанно,
PS|39|13|ибо окружили меня беды неисчислимые; постигли меня беззакония мои, так что видеть не могу: их более, нежели волос на голове моей; сердце мое оставило меня.
PS|39|14|Благоволи, Господи, избавить меня; Господи! поспеши на помощь мне.
PS|39|15|Да постыдятся и посрамятся все, ищущие погибели душе моей! Да будут обращены назад и преданы посмеянию желающие мне зла!
PS|39|16|Да смятутся от посрамления своего говорящие мне: "хорошо! хорошо!"
PS|39|17|Да радуются и веселятся Тобою все ищущие Тебя, и любящие спасение Твое да говорят непрестанно: "велик Господь!"
PS|39|18|Я же беден и нищ, но Господь печется о мне. Ты – помощь моя и избавитель мой, Боже мой! не замедли.
PS|40|1|Начальнику хора. Псалом Давида.
PS|40|2|Блажен, кто помышляет о бедном! В день бедствия избавит его Господь.
PS|40|3|Господь сохранит его и сбережет ему жизнь; блажен будет он на земле. И Ты не отдашь его на волю врагов его.
PS|40|4|Господь укрепит его на одре болезни его. Ты изменишь все ложе его в болезни его.
PS|40|5|Я сказал: Господи! помилуй меня, исцели душу мою, ибо согрешил я пред Тобою.
PS|40|6|Враги мои говорят обо мне злое: "когда он умрет и погибнет имя его?"
PS|40|7|И если приходит кто видеть меня, говорит ложь; сердце его слагает в себе неправду, и он, выйдя вон, толкует.
PS|40|8|Все ненавидящие меня шепчут между собою против меня, замышляют на меня зло:
PS|40|9|"слово велиала пришло на него; он слег; не встать ему более".
PS|40|10|Даже человек мирный со мною, на которого я полагался, который ел хлеб мой, поднял на меня пяту.
PS|40|11|Ты же, Господи, помилуй меня и восставь меня, и я воздам им.
PS|40|12|Из того узнаю, что Ты благоволишь ко мне, если враг мой не восторжествует надо мною,
PS|40|13|а меня сохранишь в целости моей и поставишь пред лицем Твоим на веки.
PS|40|14|Благословен Господь Бог Израилев от века и до века! Аминь, аминь!
PS|41|1|Начальнику хора. Учение. Сынов Кореевых.
PS|41|2|Как лань желает к потокам воды, так желает душа моя к Тебе, Боже!
PS|41|3|Жаждет душа моя к Богу крепкому, живому: когда приду и явлюсь пред лице Божие!
PS|41|4|Слезы мои были для меня хлебом день и ночь, когда говорили мне всякий день: "где Бог твой?"
PS|41|5|Вспоминая об этом, изливаю душу мою, потому что я ходил в многолюдстве, вступал с ними в дом Божий со гласом радости и славословия празднующего сонма.
PS|41|6|Что унываешь ты, душа моя, и что смущаешься? Уповай на Бога, ибо я буду еще славить Его, Спасителя моего и Бога моего.
PS|41|7|Унывает во мне душа моя; посему я воспоминаю о Тебе с земли Иорданской, с Ермона, с горы Цоар.
PS|41|8|Бездна бездну призывает голосом водопадов Твоих; все воды Твои и волны Твои прошли надо мною.
PS|41|9|Днем явит Господь милость Свою, и ночью песнь Ему у меня, молитва к Богу жизни моей.
PS|41|10|Скажу Богу, заступнику моему: для чего Ты забыл меня? Для чего я сетуя хожу от оскорблений врага?
PS|41|11|Как бы поражая кости мои, ругаются надо мною враги мои, когда говорят мне всякий день: "где Бог твой?"
PS|41|12|Что унываешь ты, душа моя, и что смущаешься? Уповай на Бога, ибо я буду еще славить Его, Спасителя моего и Бога моего.
PS|42|1|Суди меня, Боже, и вступись в тяжбу мою с народом недобрым. От человека лукавого и несправедливого избавь меня,
PS|42|2|ибо Ты Бог крепости моей. Для чего Ты отринул меня? для чего я сетуя хожу от оскорблений врага?
PS|42|3|Пошли свет Твой и истину Твою; да ведут они меня и приведут на святую гору Твою и в обители Твои.
PS|42|4|И подойду я к жертвеннику Божию, к Богу радости и веселия моего, и на гуслях буду славить Тебя, Боже, Боже мой!
PS|42|5|Что унываешь ты, душа моя, и что смущаешься? Уповай на Бога; ибо я буду еще славить Его, Спасителя моего и Бога моего.
PS|43|1|Начальнику хора. Учение. Сынов Кореевых.
PS|43|2|Боже, мы слышали ушами своими, отцы наши рассказывали нам о деле, какое Ты соделал во дни их, во дни древние:
PS|43|3|Ты рукою Твоею истребил народы, а их насадил; поразил племена и изгнал их;
PS|43|4|ибо они не мечом своим приобрели землю, и не их мышца спасла их, но Твоя десница и Твоя мышца и свет лица Твоего, ибо Ты благоволил к ним.
PS|43|5|Боже, Царь мой! Ты – тот же; даруй спасение Иакову.
PS|43|6|С Тобою избодаем рогами врагов наших; во имя Твое попрем ногами восстающих на нас:
PS|43|7|ибо не на лук мой уповаю, и не меч мой спасет меня;
PS|43|8|но Ты спасешь нас от врагов наших, и посрамишь ненавидящих нас.
PS|43|9|О Боге похвалимся всякий день, и имя Твое будем прославлять вовек.
PS|43|10|Но ныне Ты отринул и посрамил нас, и не выходишь с войсками нашими;
PS|43|11|обратил нас в бегство от врага, и ненавидящие нас грабят нас;
PS|43|12|Ты отдал нас, как овец, на съедение и рассеял нас между народами;
PS|43|13|без выгоды Ты продал народ Твой и не возвысил цены его;
PS|43|14|отдал нас на поношение соседям нашим, на посмеяние и поругание живущим вокруг нас;
PS|43|15|Ты сделал нас притчею между народами, покиванием головы между иноплеменниками.
PS|43|16|Всякий день посрамление мое предо мною, и стыд покрывает лице мое
PS|43|17|от голоса поносителя и клеветника, от взоров врага и мстителя:
PS|43|18|все это пришло на нас, но мы не забыли Тебя и не нарушили завета Твоего.
PS|43|19|Не отступило назад сердце наше, и стопы наши не уклонились от пути Твоего,
PS|43|20|когда Ты сокрушил нас в земле драконов и покрыл нас тенью смертною.
PS|43|21|Если бы мы забыли имя Бога нашего и простерли руки наши к богу чужому,
PS|43|22|то не взыскал ли бы сего Бог? Ибо Он знает тайны сердца.
PS|43|23|Но за Тебя умерщвляют нас всякий день, считают нас за овец, [обреченных] на заклание.
PS|43|24|Восстань, что спишь, Господи! пробудись, не отринь навсегда.
PS|43|25|Для чего скрываешь лице Твое, забываешь скорбь нашу и угнетение наше?
PS|43|26|ибо душа наша унижена до праха, утроба наша прильнула к земле.
PS|43|27|Восстань на помощь нам и избавь нас ради милости Твоей.
PS|44|1|Начальнику хора. На [музыкальном орудии] Шошан. Учение. Сынов Кореевых. Песнь любви.
PS|44|2|Излилось из сердца моего слово благое; я говорю: песнь моя о Царе; язык мой – трость скорописца.
PS|44|3|Ты прекраснее сынов человеческих; благодать излилась из уст Твоих; посему благословил Тебя Бог на веки.
PS|44|4|Препояшь Себя по бедру мечом Твоим, Сильный, славою Твоею и красотою Твоею,
PS|44|5|и в сем украшении Твоем поспеши, воссядь на колесницу ради истины и кротости и правды, и десница Твоя покажет Тебе дивные дела.
PS|44|6|Остры стрелы Твои; – народы падут пред Тобою, – они – в сердце врагов Царя.
PS|44|7|Престол Твой, Боже, вовек; жезл правоты – жезл царства Твоего.
PS|44|8|Ты возлюбил правду и возненавидел беззаконие, посему помазал Тебя, Боже, Бог Твой елеем радости более соучастников Твоих.
PS|44|9|Все одежды Твои, как смирна и алой и касия; из чертогов слоновой кости увеселяют Тебя.
PS|44|10|Дочери царей между почетными у Тебя; стала царица одесную Тебя в Офирском золоте.
PS|44|11|Слыши, дщерь, и смотри, и приклони ухо твое, и забудь народ твой и дом отца твоего.
PS|44|12|И возжелает Царь красоты твоей; ибо Он Господь твой, и ты поклонись Ему.
PS|44|13|И дочь Тира с дарами, и богатейшие из народа будут умолять лице Твое.
PS|44|14|Вся слава дщери Царя внутри; одежда ее шита золотом;
PS|44|15|в испещренной одежде ведется она к Царю; за нею ведутся к Тебе девы, подруги ее,
PS|44|16|приводятся с весельем и ликованьем, входят в чертог Царя.
PS|44|17|Вместо отцов Твоих, будут сыновья Твои; Ты поставишь их князьями по всей земле.
PS|44|18|Сделаю имя Твое памятным в род и род; посему народы будут славить Тебя во веки и веки.
PS|45|1|Начальнику хора. Сынов Кореевых. На [музыкальном] [орудии] Аламоф. Песнь.
PS|45|2|Бог нам прибежище и сила, скорый помощник в бедах,
PS|45|3|посему не убоимся, хотя бы поколебалась земля, и горы двинулись в сердце морей.
PS|45|4|Пусть шумят, вздымаются воды их, трясутся горы от волнения их.
PS|45|5|Речные потоки веселят град Божий, святое жилище Всевышнего.
PS|45|6|Бог посреди его; он не поколеблется: Бог поможет ему с раннего утра.
PS|45|7|Восшумели народы; двинулись царства: [Всевышний] дал глас Свой, и растаяла земля.
PS|45|8|Господь сил с нами, Бог Иакова заступник наш.
PS|45|9|Придите и видите дела Господа, – какие произвел Он опустошения на земле:
PS|45|10|прекращая брани до края земли, сокрушил лук и переломил копье, колесницы сжег огнем.
PS|45|11|Остановитесь и познайте, что Я – Бог: буду превознесен в народах, превознесен на земле.
PS|45|12|Господь сил с нами, заступник наш Бог Иакова.
PS|46|1|Начальнику хора. Сынов Кореевых. Псалом.
PS|46|2|Восплещите руками все народы, воскликните Богу гласом радости;
PS|46|3|ибо Господь Всевышний страшен, – великий Царь над всею землею;
PS|46|4|покорил нам народы и племена под ноги наши;
PS|46|5|избрал нам наследие наше, красу Иакова, которого возлюбил.
PS|46|6|Восшел Бог при восклицаниях, Господь при звуке трубном.
PS|46|7|Пойте Богу нашему, пойте; пойте Царю нашему, пойте,
PS|46|8|ибо Бог – Царь всей земли; пойте все разумно.
PS|46|9|Бог воцарился над народами, Бог воссел на святом престоле Своем;
PS|46|10|Князья народов собрались к народу Бога Авраамова, ибо щиты земли – Божии; Он превознесен [над ними].
PS|47|1|Песнь. Псалом. Сынов Кореевых.
PS|47|2|Велик Господь и всехвален во граде Бога нашего, на святой горе Его.
PS|47|3|Прекрасная возвышенность, радость всей земли гора Сион; на северной стороне [ее] город великого Царя.
PS|47|4|Бог в жилищах его ведом, как заступник:
PS|47|5|ибо вот, сошлись цари и прошли все мимо;
PS|47|6|увидели и изумились, смутились и обратились в бегство;
PS|47|7|страх объял их там и мука, как у женщин в родах;
PS|47|8|восточным ветром Ты сокрушил Фарсийские корабли.
PS|47|9|Как слышали мы, так и увидели во граде Господа сил, во граде Бога нашего: Бог утвердит его на веки.
PS|47|10|Мы размышляли, Боже, о благости Твоей посреди храма Твоего.
PS|47|11|Как имя Твое, Боже, так и хвала Твоя до концов земли; десница Твоя полна правды.
PS|47|12|Да веселится гора Сион, да радуются дщери Иудейские ради судов Твоих, [Господи].
PS|47|13|Пойдите вокруг Сиона и обойдите его, пересчитайте башни его;
PS|47|14|обратите сердце ваше к укреплениям его, рассмотрите домы его, чтобы пересказать грядущему роду,
PS|47|15|ибо сей Бог есть Бог наш на веки и веки: Он будет вождем нашим до самой смерти.
PS|48|1|Начальнику хора. Сынов Кореевых. Псалом.
PS|48|2|Слушайте сие, все народы; внимайте сему, все живущие во вселенной, –
PS|48|3|и простые и знатные, богатый, равно как бедный.
PS|48|4|Уста мои изрекут премудрость, и размышления сердца моего – знание.
PS|48|5|Приклоню ухо мое к притче, на гуслях открою загадку мою:
PS|48|6|"для чего бояться мне во дни бедствия, [когда] беззаконие путей моих окружит меня?"
PS|48|7|Надеющиеся на силы свои и хвалящиеся множеством богатства своего!
PS|48|8|человек никак не искупит брата своего и не даст Богу выкупа за него:
PS|48|9|дорога цена искупления души их, и не будет того вовек,
PS|48|10|чтобы остался [кто] жить навсегда и не увидел могилы.
PS|48|11|Каждый видит, что и мудрые умирают, равно как и невежды и бессмысленные погибают и оставляют имущество свое другим.
PS|48|12|В мыслях у них, что домы их вечны, и что жилища их в род и род, и земли свои они называют своими именами.
PS|48|13|Но человек в чести не пребудет; он уподобится животным, которые погибают.
PS|48|14|Этот путь их есть безумие их, хотя последующие за ними одобряют мнение их.
PS|48|15|Как овец, заключат их в преисподнюю; смерть будет пасти их, и наутро праведники будут владычествовать над ними; сила их истощится; могила – жилище их.
PS|48|16|Но Бог избавит душу мою от власти преисподней, когда примет меня.
PS|48|17|Не бойся, когда богатеет человек, когда слава дома его умножается:
PS|48|18|ибо умирая не возьмет ничего; не пойдет за ним слава его;
PS|48|19|хотя при жизни он ублажает душу свою, и прославляют тебя, что ты удовлетворяешь себе,
PS|48|20|но он пойдет к роду отцов своих, которые никогда не увидят света.
PS|48|21|Человек, который в чести и неразумен, подобен животным, которые погибают.
PS|49|1|Псалом Асафа. Бог Богов, Господь возглаголал и призывает землю, от восхода солнца до запада.
PS|49|2|С Сиона, который есть верх красоты, является Бог,
PS|49|3|грядет Бог наш, и не в безмолвии: пред Ним огонь поядающий, и вокруг Его сильная буря.
PS|49|4|Он призывает свыше небо и землю, судить народ Свой:
PS|49|5|"соберите ко Мне святых Моих, вступивших в завет со Мною при жертве".
PS|49|6|И небеса провозгласят правду Его, ибо судия сей есть Бог.
PS|49|7|"Слушай, народ Мой, Я буду говорить; Израиль! Я буду свидетельствовать против тебя: Я Бог, твой Бог.
PS|49|8|Не за жертвы твои Я буду укорять тебя; всесожжения твои всегда предо Мною;
PS|49|9|не приму тельца из дома твоего, ни козлов из дворов твоих,
PS|49|10|ибо Мои все звери в лесу, и скот на тысяче гор,
PS|49|11|знаю всех птиц на горах, и животные на полях предо Мною.
PS|49|12|Если бы Я взалкал, то не сказал бы тебе, ибо Моя вселенная и все, что наполняет ее.
PS|49|13|Ем ли Я мясо волов и пью ли кровь козлов?
PS|49|14|Принеси в жертву Богу хвалу и воздай Всевышнему обеты твои,
PS|49|15|и призови Меня в день скорби; Я избавлю тебя, и ты прославишь Меня".
PS|49|16|Грешнику же говорит Бог: "что ты проповедуешь уставы Мои и берешь завет Мой в уста твои,
PS|49|17|а сам ненавидишь наставление Мое и слова Мои бросаешь за себя?
PS|49|18|когда видишь вора, сходишься с ним, и с прелюбодеями сообщаешься;
PS|49|19|уста твои открываешь на злословие, и язык твой сплетает коварство;
PS|49|20|сидишь и говоришь на брата твоего, на сына матери твоей клевещешь;
PS|49|21|ты это делал, и Я молчал; ты подумал, что Я такой же, как ты. Изобличу тебя и представлю пред глаза твои [грехи твои].
PS|49|22|Уразумейте это, забывающие Бога, дабы Я не восхитил, – и не будет избавляющего.
PS|49|23|Кто приносит в жертву хвалу, тот чтит Меня, и кто наблюдает за путем своим, тому явлю Я спасение Божие".
PS|50|1|Начальнику хора. Псалом Давида,
PS|50|2|Когда приходил к нему пророк Нафан, после того, как Давид вошел к Вирсавии.
PS|50|3|Помилуй меня, Боже, по великой милости Твоей, и по множеству щедрот Твоих изгладь беззакония мои.
PS|50|4|Многократно омой меня от беззакония моего, и от греха моего очисти меня,
PS|50|5|ибо беззакония мои я сознаю, и грех мой всегда предо мною.
PS|50|6|Тебе, Тебе единому согрешил я и лукавое пред очами Твоими сделал, так что Ты праведен в приговоре Твоем и чист в суде Твоем.
PS|50|7|Вот, я в беззаконии зачат, и во грехе родила меня мать моя.
PS|50|8|Вот, Ты возлюбил истину в сердце и внутрь меня явил мне мудрость.
PS|50|9|Окропи меня иссопом, и буду чист; омой меня, и буду белее снега.
PS|50|10|Дай мне услышать радость и веселие, и возрадуются кости, Тобою сокрушенные.
PS|50|11|Отврати лице Твое от грехов моих и изгладь все беззакония мои.
PS|50|12|Сердце чистое сотвори во мне, Боже, и дух правый обнови внутри меня.
PS|50|13|Не отвергни меня от лица Твоего и Духа Твоего Святаго не отними от меня.
PS|50|14|Возврати мне радость спасения Твоего и Духом владычественным утверди меня.
PS|50|15|Научу беззаконных путям Твоим, и нечестивые к Тебе обратятся.
PS|50|16|Избавь меня от кровей, Боже, Боже спасения моего, и язык мой восхвалит правду Твою.
PS|50|17|Господи! отверзи уста мои, и уста мои возвестят хвалу Твою:
PS|50|18|ибо жертвы Ты не желаешь, – я дал бы ее; к всесожжению не благоволишь.
PS|50|19|Жертва Богу – дух сокрушенный; сердца сокрушенного и смиренного Ты не презришь, Боже.
PS|50|20|Облагодетельствуй по благоволению Твоему Сион; воздвигни стены Иерусалима:
PS|50|21|тогда благоугодны будут Тебе жертвы правды, возношение и всесожжение; тогда возложат на алтарь Твой тельцов.
PS|51|1|Начальнику хора. Учение Давида,
PS|51|2|после того, как приходил Доик Идумеянин и донес Саулу и сказал ему, что Давид пришел в дом Ахимелеха.
PS|51|3|Что хвалишься злодейством, сильный? милость Божия всегда [со мною;]
PS|51|4|гибель вымышляет язык твой; как изощренная бритва, он [у] [тебя], коварный!
PS|51|5|ты любишь больше зло, нежели добро, больше ложь, нежели говорить правду;
PS|51|6|ты любишь всякие гибельные речи, язык коварный:
PS|51|7|за то Бог сокрушит тебя вконец, изринет тебя и исторгнет тебя из жилища [твоего] и корень твой из земли живых.
PS|51|8|Увидят праведники и убоятся, посмеются над ним [и скажут]:
PS|51|9|"вот человек, который не в Боге полагал крепость свою, а надеялся на множество богатства своего, укреплялся в злодействе своем".
PS|51|10|А я, как зеленеющая маслина, в доме Божием, и уповаю на милость Божию во веки веков,
PS|51|11|вечно буду славить Тебя за то, что Ты соделал, и уповать на имя Твое, ибо оно благо пред святыми Твоими.
PS|52|1|Начальнику хора. На духовом [орудии]. Учение Давида.
PS|52|2|Сказал безумец в сердце своем: "нет Бога". Развратились они и совершили гнусные преступления; нет делающего добро.
PS|52|3|Бог с небес призрел на сынов человеческих, чтобы видеть, есть ли разумеющий, ищущий Бога.
PS|52|4|Все уклонились, сделались равно непотребными; нет делающего добро, нет ни одного.
PS|52|5|Неужели не вразумятся делающие беззаконие, съедающие народ мой, [как] едят хлеб, и не призывающие Бога?
PS|52|6|Там убоятся они страха, где нет страха, ибо рассыплет Бог кости ополчающихся против тебя. Ты постыдишь их, потому что Бог отверг их.
PS|52|7|Кто даст с Сиона спасение Израилю! Когда Бог возвратит пленение народа Своего, тогда возрадуется Иаков и возвеселится Израиль.
PS|53|1|Начальнику хора. На струнных [орудиях]. Учение Давида,
PS|53|2|когда пришли Зифеи и сказали Саулу: "не у нас ли скрывается Давид?"
PS|53|3|Боже! именем Твоим спаси меня, и силою Твоею суди меня.
PS|53|4|Боже! услышь молитву мою, внемли словам уст моих,
PS|53|5|ибо чужие восстали на меня, и сильные ищут души моей; они не имеют Бога пред собою.
PS|53|6|Вот, Бог помощник мой; Господь подкрепляет душу мою.
PS|53|7|Он воздаст за зло врагам моим; истиною Твоею истреби их.
PS|53|8|Я усердно принесу Тебе жертву, прославлю имя Твое, Господи, ибо оно благо,
PS|53|9|ибо Ты избавил меня от всех бед, и на врагов моих смотрело око мое.
PS|54|1|Начальнику хора. На струнных [орудиях]. Учение Давида.
PS|54|2|Услышь, Боже, молитву мою и не скрывайся от моления моего;
PS|54|3|внемли мне и услышь меня; я стенаю в горести моей, и смущаюсь
PS|54|4|от голоса врага, от притеснения нечестивого, ибо они возводят на меня беззаконие и в гневе враждуют против меня.
PS|54|5|Сердце мое трепещет во мне, и смертные ужасы напали на меня;
PS|54|6|страх и трепет нашел на меня, и ужас объял меня.
PS|54|7|И я сказал: "кто дал бы мне крылья, как у голубя? я улетел бы и успокоился бы;
PS|54|8|далеко удалился бы я, и оставался бы в пустыне;
PS|54|9|поспешил бы укрыться от вихря, от бури".
PS|54|10|Расстрой, Господи, и раздели языки их, ибо я вижу насилие и распри в городе;
PS|54|11|днем и ночью ходят они кругом по стенам его; злодеяния и бедствие посреди его;
PS|54|12|посреди его пагуба; обман и коварство не сходят с улиц его:
PS|54|13|ибо не враг поносит меня, – это я перенес бы; не ненавистник мой величается надо мною, – от него я укрылся бы;
PS|54|14|но ты, который был для меня то же, что я, друг мой и близкий мой,
PS|54|15|с которым мы разделяли искренние беседы и ходили вместе в дом Божий.
PS|54|16|Да найдет на них смерть; да сойдут они живыми в ад, ибо злодейство в жилищах их, посреди их.
PS|54|17|Я же воззову к Богу, и Господь спасет меня.
PS|54|18|Вечером и утром и в полдень буду умолять и вопиять, и Он услышит голос мой,
PS|54|19|избавит в мире душу мою от восстающих на меня, ибо их много у меня;
PS|54|20|услышит Бог, и смирит их от века Живущий, потому что нет в них перемены; они не боятся Бога,
PS|54|21|простерли руки свои на тех, которые с ними в мире, нарушили союз свой;
PS|54|22|уста их мягче масла, а в сердце их вражда; слова их нежнее елея, но они суть обнаженные мечи.
PS|54|23|Возложи на Господа заботы твои, и Он поддержит тебя. Никогда не даст Он поколебаться праведнику.
PS|54|24|Ты, Боже, низведешь их в ров погибели; кровожадные и коварные не доживут и до половины дней своих. А я на Тебя, [Господи], уповаю.
PS|55|1|Начальнику хора. О голубице, безмолвствующей в удалении. Писание Давида, когда Филистимляне захватили его в Гефе.
PS|55|2|Помилуй меня, Боже! ибо человек хочет поглотить меня; нападая всякий день, теснит меня.
PS|55|3|Враги мои всякий день ищут поглотить меня, ибо много восстающих на меня, о, Всевышний!
PS|55|4|Когда я в страхе, на Тебя я уповаю.
PS|55|5|В Боге восхвалю я слово Его; на Бога уповаю, не боюсь; что сделает мне плоть?
PS|55|6|Всякий день извращают слова мои; все помышления их обо мне – на зло:
PS|55|7|собираются, притаиваются, наблюдают за моими пятами, чтобы уловить душу мою.
PS|55|8|Неужели они избегнут воздаяния за неправду [свою]? Во гневе низложи, Боже, народы.
PS|55|9|У Тебя исчислены мои скитания; положи слезы мои в сосуд у Тебя, – не в книге ли они Твоей?
PS|55|10|Враги мои обращаются назад, когда я взываю к Тебе, из этого я узнаю, что Бог за меня.
PS|55|11|В Боге восхвалю я слово [Его], в Господе восхвалю слово [Его].
PS|55|12|На Бога уповаю, не боюсь; что сделает мне человек?
PS|55|13|На мне, Боже, обеты Тебе; Тебе воздам хвалы,
PS|55|14|ибо Ты избавил душу мою от смерти, да и ноги мои от преткновения, чтобы я ходил пред лицем Божиим во свете живых.
PS|56|1|Начальнику хора. Не погуби. Писание Давида, когда он убежал от Саула в пещеру.
PS|56|2|Помилуй меня, Боже, помилуй меня, ибо на Тебя уповает душа моя, и в тени крыл Твоих я укроюсь, доколе не пройдут беды.
PS|56|3|Воззову к Богу Всевышнему, Богу, благодетельствующему мне;
PS|56|4|Он пошлет с небес и спасет меня; посрамит ищущего поглотить меня; пошлет Бог милость Свою и истину Свою.
PS|56|5|Душа моя среди львов; я лежу среди дышущих пламенем, среди сынов человеческих, у которых зубы – копья и стрелы, и у которых язык – острый меч.
PS|56|6|Будь превознесен выше небес, Боже, и над всею землею да будет слава Твоя!
PS|56|7|Приготовили сеть ногам моим; душа моя поникла; выкопали предо мною яму, и [сами] упали в нее.
PS|56|8|Готово сердце мое, Боже, готово сердце мое: буду петь и славить.
PS|56|9|Воспрянь, слава моя, воспрянь, псалтирь и гусли! Я встану рано.
PS|56|10|Буду славить Тебя, Господи, между народами; буду воспевать Тебя среди племен,
PS|56|11|ибо до небес велика милость Твоя и до облаков истина Твоя.
PS|56|12|Будь превознесен выше небес, Боже, и над всею землею да будет слава Твоя!
PS|57|1|Начальнику хора. Не погуби. Писание Давида.
PS|57|2|Подлинно ли правду говорите вы, судьи, и справедливо судите, сыны человеческие?
PS|57|3|Беззаконие составляете в сердце, кладете на весы злодеяния рук ваших на земле.
PS|57|4|С самого рождения отступили нечестивые, от утробы [матери] заблуждаются, говоря ложь.
PS|57|5|Яд у них – как яд змеи, как глухого аспида, который затыкает уши свои
PS|57|6|и не слышит голоса заклинателя, самого искусного в заклинаниях.
PS|57|7|Боже! сокруши зубы их в устах их; разбей, Господи, челюсти львов!
PS|57|8|Да исчезнут, как вода протекающая; когда напрягут стрелы, пусть они будут как переломленные.
PS|57|9|Да исчезнут, как распускающаяся улитка; да не видят солнца, как выкидыш женщины.
PS|57|10|Прежде нежели котлы ваши ощутят горящий терн, и свежее и обгоревшее да разнесет вихрь.
PS|57|11|Возрадуется праведник, когда увидит отмщение; омоет стопы свои в крови нечестивого.
PS|57|12|И скажет человек: "подлинно есть плод праведнику! итак есть Бог, судящий на земле!"
PS|58|1|Начальнику хора. Не погуби. Писание Давида, когда Саул послал стеречь дом его, чтобы умертвить его.
PS|58|2|Избавь меня от врагов моих, Боже мой! защити меня от восстающих на меня;
PS|58|3|избавь меня от делающих беззаконие; спаси от кровожадных,
PS|58|4|ибо вот, они подстерегают душу мою; собираются на меня сильные не за преступление мое и не за грех мой, Господи;
PS|58|5|без вины [моей] сбегаются и вооружаются; подвигнись на помощь мне и воззри.
PS|58|6|Ты, Господи, Боже сил, Боже Израилев, восстань посетить все народы, не пощади ни одного из нечестивых беззаконников:
PS|58|7|вечером возвращаются они, воют, как псы, и ходят вокруг города;
PS|58|8|вот они изрыгают хулу языком своим; в устах их мечи: "ибо", [думают они], "кто слышит?"
PS|58|9|Но Ты, Господи, посмеешься над ними; Ты посрамишь все народы.
PS|58|10|Сила – у них, но я к Тебе прибегаю, ибо Бог – заступник мой.
PS|58|11|Бог мой, милующий меня, предварит меня; Бог даст мне смотреть на врагов моих.
PS|58|12|Не умерщвляй их, чтобы не забыл народ мой; расточи их силою Твоею и низложи их, Господи, защитник наш.
PS|58|13|Слово языка их есть грех уст их, да уловятся они в гордости своей за клятву и ложь, которую произносят.
PS|58|14|Расточи их во гневе, расточи, чтобы их не было; и да познают, что Бог владычествует над Иаковом до пределов земли.
PS|58|15|Пусть возвращаются вечером, воют, как псы, и ходят вокруг города;
PS|58|16|пусть бродят, чтобы найти пищу, и несытые проводят ночи.
PS|58|17|А я буду воспевать силу Твою и с раннего утра провозглашать милость Твою, ибо Ты был мне защитою и убежищем в день бедствия моего.
PS|58|18|Сила моя! Тебя буду воспевать я, ибо Бог – заступник мой, Бог мой, милующий меня.
PS|59|1|Начальнику хора. На [музыкальном орудии] Шушан–Эдуф. Писание Давида для изучения,
PS|59|2|когда он воевал с Сириею Месопотамскою и с Сириею Цованскою, и когда Иоав, возвращаясь, поразил двенадцать тысяч Идумеев в долине Соляной.
PS|59|3|Боже! Ты отринул нас, Ты сокрушил нас, Ты прогневался: обратись к нам.
PS|59|4|Ты потряс землю, разбил ее: исцели повреждения ее, ибо она колеблется.
PS|59|5|Ты дал испытать народу твоему жестокое, напоил нас вином изумления.
PS|59|6|Даруй боящимся Тебя знамя, чтобы они подняли его ради истины,
PS|59|7|чтобы избавились возлюбленные Твои; спаси десницею Твоею и услышь меня.
PS|59|8|Бог сказал во святилище Своем: "восторжествую, разделю Сихем и долину Сокхоф размерю:
PS|59|9|Мой Галаад, Мой Манассия, Ефрем крепость главы Моей, Иуда скипетр Мой,
PS|59|10|Моав умывальная чаша Моя; на Едома простру сапог Мой. Восклицай Мне, земля Филистимская!"
PS|59|11|Кто введет меня в укрепленный город? Кто доведет меня до Едома?
PS|59|12|Не Ты ли, Боже, [Который] отринул нас, и не выходишь, Боже, с войсками нашими?
PS|59|13|Подай нам помощь в тесноте, ибо защита человеческая суетна.
PS|59|14|С Богом мы окажем силу, Он низложит врагов наших.
PS|60|1|Начальнику хора. На струнном [орудии]. Псалом Давида.
PS|60|2|Услышь, Боже, вопль мой, внемли молитве моей!
PS|60|3|От конца земли взываю к Тебе в унынии сердца моего; возведи меня на скалу, для меня недосягаемую,
PS|60|4|ибо Ты прибежище мое, Ты крепкая защита от врага.
PS|60|5|Да живу я вечно в жилище Твоем и покоюсь под кровом крыл Твоих,
PS|60|6|ибо Ты, Боже, услышал обеты мои и дал [мне] наследие боящихся имени Твоего.
PS|60|7|Приложи дни ко дням царя, лета его [продли] в род и род,
PS|60|8|да пребудет он вечно пред Богом; заповедуй милости и истине охранять его.
PS|60|9|И я буду петь имени Твоему вовек, исполняя обеты мои всякий день.
PS|61|1|Начальнику хора Идифумова. Псалом Давида.
PS|61|2|Только в Боге успокаивается душа моя: от Него спасение мое.
PS|61|3|Только Он – твердыня моя, спасение мое, убежище мое: не поколеблюсь более.
PS|61|4|Доколе вы будете налегать на человека? Вы будете низринуты, все вы, как наклонившаяся стена, как ограда пошатнувшаяся.
PS|61|5|Они задумали свергнуть его с высоты, прибегли ко лжи; устами благословляют, а в сердце своем клянут.
PS|61|6|Только в Боге успокаивайся, душа моя! ибо на Него надежда моя.
PS|61|7|Только Он – твердыня моя и спасение мое, убежище мое: не поколеблюсь.
PS|61|8|В Боге спасение мое и слава моя; крепость силы моей и упование мое в Боге.
PS|61|9|Народ! надейтесь на Него во всякое время; изливайте пред Ним сердце ваше: Бог нам прибежище.
PS|61|10|Сыны человеческие – только суета; сыны мужей – ложь; если положить их на весы, все они вместе легче пустоты.
PS|61|11|Не надейтесь на грабительство и не тщеславьтесь хищением; когда богатство умножается, не прилагайте [к нему] сердца.
PS|61|12|Однажды сказал Бог, и дважды слышал я это, что сила у Бога,
PS|61|13|и у Тебя, Господи, милость, ибо Ты воздаешь каждому по делам его.
PS|62|1|Псалом Давида, когда он был в пустыне Иудейской.
PS|62|2|Боже! Ты Бог мой, Тебя от ранней зари ищу я; Тебя жаждет душа моя, по Тебе томится плоть моя в земле пустой, иссохшей и безводной,
PS|62|3|чтобы видеть силу Твою и славу Твою, как я видел Тебя во святилище:
PS|62|4|ибо милость Твоя лучше, нежели жизнь. Уста мои восхвалят Тебя.
PS|62|5|Так благословлю Тебя в жизни моей; во имя Твое вознесу руки мои.
PS|62|6|Как туком и елеем насыщается душа моя, и радостным гласом восхваляют Тебя уста мои,
PS|62|7|когда я вспоминаю о Тебе на постели моей, размышляю о Тебе в [ночные] стражи,
PS|62|8|ибо Ты помощь моя, и в тени крыл Твоих я возрадуюсь;
PS|62|9|к Тебе прилепилась душа моя; десница Твоя поддерживает меня.
PS|62|10|А те, которые ищут погибели душе моей, сойдут в преисподнюю земли;
PS|62|11|Сразят их силою меча; достанутся они в добычу лисицам.
PS|62|12|Царь же возвеселится о Боге, восхвален будет всякий, клянущийся Им, ибо заградятся уста говорящих неправду.
PS|63|1|Начальнику хора. Псалом Давида.
PS|63|2|Услышь, Боже, голос мой в молитве моей, сохрани жизнь мою от страха врага;
PS|63|3|укрой меня от замысла коварных, от мятежа злодеев,
PS|63|4|которые изострили язык свой, как меч; напрягли лук свой – язвительное слово,
PS|63|5|чтобы втайне стрелять в непорочного; они внезапно стреляют в него и не боятся.
PS|63|6|Они утвердились в злом намерении, совещались скрыть сеть, говорили: кто их увидит?
PS|63|7|Изыскивают неправду, делают расследование за расследованием даже до внутренней жизни человека и до глубины сердца.
PS|63|8|Но поразит их Бог стрелою: внезапно будут они уязвлены;
PS|63|9|языком своим они поразят самих себя; все, видящие их, удалятся [от них].
PS|63|10|И убоятся все человеки, и возвестят дело Божие, и уразумеют, что это Его дело.
PS|63|11|А праведник возвеселится о Господе и будет уповать на Него; и похвалятся все правые сердцем.
PS|64|1|Начальнику хора. Псалом Давида для пения.
PS|64|2|Тебе, Боже, принадлежит хвала на Сионе, и Тебе воздастся обет [в Иерусалиме].
PS|64|3|Ты слышишь молитву; к Тебе прибегает всякая плоть.
PS|64|4|Дела беззаконий превозмогают меня; Ты очистишь преступления наши.
PS|64|5|Блажен, кого Ты избрал и приблизил, чтобы он жил во дворах Твоих. Насытимся благами дома Твоего, святаго храма Твоего.
PS|64|6|Страшный в правосудии, услышь нас, Боже, Спаситель наш, упование всех концов земли и находящихся в море далеко,
PS|64|7|поставивший горы силою Своею, препоясанный могуществом,
PS|64|8|укрощающий шум морей, шум волн их и мятеж народов!
PS|64|9|И убоятся знамений Твоих живущие на пределах [земли]. Утро и вечер возбудишь к славе [Твоей].
PS|64|10|Ты посещаешь землю и утоляешь жажду ее, обильно обогащаешь ее: поток Божий полон воды; Ты приготовляешь хлеб, ибо так устроил ее;
PS|64|11|напояешь борозды ее, уравниваешь глыбы ее, размягчаешь ее каплями дождя, благословляешь произрастания ее;
PS|64|12|венчаешь лето благости Твоей, и стези Твои источают тук,
PS|64|13|источают на пустынные пажити, и холмы препоясываются радостью;
PS|64|14|луга одеваются стадами, и долины покрываются хлебом, восклицают и поют.
PS|65|1|Начальнику хора. Песнь. Воскликните Богу, вся земля.
PS|65|2|Пойте славу имени Его, воздайте славу, хвалу Ему.
PS|65|3|Скажите Богу: как страшен Ты в делах Твоих! По множеству силы Твоей, покорятся Тебе враги Твои.
PS|65|4|Вся земля да поклонится Тебе и поет Тебе, да поет имени Твоему.
PS|65|5|Придите и воззрите на дела Бога, страшного в делах над сынами человеческими.
PS|65|6|Он превратил море в сушу; через реку перешли стопами, там веселились мы о Нем.
PS|65|7|Могуществом Своим владычествует Он вечно; очи Его зрят на народы, да не возносятся мятежники.
PS|65|8|Благословите, народы, Бога нашего и провозгласите хвалу Ему.
PS|65|9|Он сохранил душе нашей жизнь и ноге нашей не дал поколебаться.
PS|65|10|Ты испытал нас, Боже, переплавил нас, как переплавляют серебро.
PS|65|11|Ты ввел нас в сеть, положил оковы на чресла наши,
PS|65|12|посадил человека на главу нашу. Мы вошли в огонь и в воду, и Ты вывел нас на свободу.
PS|65|13|Войду в дом Твой со всесожжениями, воздам Тебе обеты мои,
PS|65|14|которые произнесли уста мои и изрек язык мой в скорби моей.
PS|65|15|Всесожжения тучные вознесу Тебе с воскурением тука овнов, принесу в жертву волов и козлов.
PS|65|16|Придите, послушайте, все боящиеся Бога, и я возвещу [вам], что сотворил Он для души моей.
PS|65|17|Я воззвал к Нему устами моими и превознес Его языком моим.
PS|65|18|Если бы я видел беззаконие в сердце моем, то не услышал бы меня Господь.
PS|65|19|Но Бог услышал, внял гласу моления моего.
PS|65|20|Благословен Бог, Который не отверг молитвы моей и не отвратил от меня милости Своей.
PS|66|1|Начальнику хора. На струнных [орудиях]. Псалом. Песнь.
PS|66|2|Боже! будь милостив к нам и благослови нас, освети нас лицем Твоим,
PS|66|3|дабы познали на земле путь Твой, во всех народах спасение Твое.
PS|66|4|Да восхвалят Тебя народы, Боже; да восхвалят Тебя народы все.
PS|66|5|Да веселятся и радуются племена, ибо Ты судишь народы праведно и управляешь на земле племенами.
PS|66|6|Да восхвалят Тебя народы, Боже, да восхвалят Тебя народы все.
PS|66|7|Земля дала плод свой; да благословит нас Бог, Бог наш.
PS|66|8|Да благословит нас Бог, и да убоятся Его все пределы земли.
PS|67|1|Начальнику хора. Псалом Давида. Песнь.
PS|67|2|Да восстанет Бог, и расточатся враги Его, и да бегут от лица Его ненавидящие Его.
PS|67|3|Как рассеивается дым, Ты рассей их; как тает воск от огня, так нечестивые да погибнут от лица Божия.
PS|67|4|А праведники да возвеселятся, да возрадуются пред Богом и восторжествуют в радости.
PS|67|5|Пойте Богу нашему, пойте имени Его, превозносите Шествующего на небесах; имя Ему: Господь, и радуйтесь пред лицем Его.
PS|67|6|Отец сирот и судья вдов Бог во святом Своем жилище.
PS|67|7|Бог одиноких вводит в дом, освобождает узников от оков, а непокорные остаются в знойной пустыне.
PS|67|8|Боже! когда Ты выходил пред народом Твоим, когда Ты шествовал пустынею,
PS|67|9|земля тряслась, даже небеса таяли от лица Божия, и этот Синай – от лица Бога, Бога Израилева.
PS|67|10|Обильный дождь проливал Ты, Боже, на наследие Твое, и когда оно изнемогало от труда, Ты подкреплял его.
PS|67|11|Народ Твой обитал там; по благости Твоей, Боже, Ты готовил [необходимое] для бедного.
PS|67|12|Господь даст слово: провозвестниц великое множество.
PS|67|13|Цари воинств бегут, бегут, а сидящая дома делит добычу.
PS|67|14|Расположившись в уделах [своих], вы стали, как голубица, которой крылья покрыты серебром, а перья чистым золотом:
PS|67|15|когда Всемогущий рассеял царей на сей [земле], она забелела, как снег на Селмоне.
PS|67|16|Гора Божия – гора Васанская! гора высокая – гора Васанская!
PS|67|17|что вы завистливо смотрите, горы высокие, на гору, на которой Бог благоволит обитать и будет Господь обитать вечно?
PS|67|18|Колесниц Божиих тьмы, тысячи тысяч; среди их Господь на Синае, во святилище.
PS|67|19|Ты восшел на высоту, пленил плен, принял дары для человеков, так чтоб и из противящихся могли обитать у Господа Бога.
PS|67|20|Благословен Господь всякий день. Бог возлагает на нас бремя, но Он же и спасает нас.
PS|67|21|Бог для нас – Бог во спасение; во власти Господа Вседержителя врата смерти.
PS|67|22|Но Бог сокрушит голову врагов Своих, волосатое темя закоснелого в своих беззакониях.
PS|67|23|Господь сказал: "от Васана возвращу, выведу из глубины морской,
PS|67|24|чтобы ты погрузил ногу твою, как и псы твои язык свой, в крови врагов".
PS|67|25|Видели шествие Твое, Боже, шествие Бога моего, Царя моего во святыне:
PS|67|26|впереди шли поющие, позади играющие на орудиях, в средине девы с тимпанами:
PS|67|27|"в собраниях благословите [Бога Господа], вы – от семени Израилева!"
PS|67|28|Там Вениамин младший – князь их; князья Иудины – владыки их, князья Завулоновы, князья Неффалимовы.
PS|67|29|Бог твой предназначил тебе силу. Утверди, Боже, то, что Ты соделал для нас!
PS|67|30|Ради храма Твоего в Иерусалиме цари принесут Тебе дары.
PS|67|31|Укроти зверя в тростнике, стадо волов среди тельцов народов, хвалящихся слитками серебра; рассыпь народы, желающие браней.
PS|67|32|Придут вельможи из Египта; Ефиопия прострет руки свои к Богу.
PS|67|33|Царства земные! пойте Богу, воспевайте Господа,
PS|67|34|шествующего на небесах небес от века. Вот, Он дает гласу Своему глас силы.
PS|67|35|Воздайте славу Богу! величие Его – над Израилем, и могущество Его – на облаках.
PS|67|36|Страшен Ты, Боже, во святилище Твоем. Бог Израилев – Он дает силу и крепость народу [Своему]. Благословен Бог!
PS|68|1|Начальнику хора. На Шошанниме. Псалом Давида.
PS|68|2|Спаси меня, Боже, ибо воды дошли до души [моей].
PS|68|3|Я погряз в глубоком болоте, и не на чем стать; вошел во глубину вод, и быстрое течение их увлекает меня.
PS|68|4|Я изнемог от вопля, засохла гортань моя, истомились глаза мои от ожидания Бога [моего].
PS|68|5|Ненавидящих меня без вины больше, нежели волос на голове моей; враги мои, преследующие меня несправедливо, усилились; чего я не отнимал, то должен отдать.
PS|68|6|Боже! Ты знаешь безумие мое, и грехи мои не сокрыты от Тебя.
PS|68|7|Да не постыдятся во мне все, надеющиеся на Тебя, Господи, Боже сил. Да не посрамятся во мне ищущие Тебя, Боже Израилев,
PS|68|8|ибо ради Тебя несу я поношение, и бесчестием покрывают лице мое.
PS|68|9|Чужим стал я для братьев моих и посторонним для сынов матери моей,
PS|68|10|ибо ревность по доме Твоем снедает меня, и злословия злословящих Тебя падают на меня;
PS|68|11|и плачу, постясь душею моею, и это ставят в поношение мне;
PS|68|12|и возлагаю на себя вместо одежды вретище, – и делаюсь для них притчею;
PS|68|13|о мне толкуют сидящие у ворот, и поют в песнях пьющие вино.
PS|68|14|А я с молитвою моею к Тебе, Господи; во время благоугодное, Боже, по великой благости Твоей услышь меня в истине спасения Твоего;
PS|68|15|извлеки меня из тины, чтобы не погрязнуть мне; да избавлюсь от ненавидящих меня и от глубоких вод;
PS|68|16|да не увлечет меня стремление вод, да не поглотит меня пучина, да не затворит надо мною пропасть зева своего.
PS|68|17|Услышь меня, Господи, ибо блага милость Твоя; по множеству щедрот Твоих призри на меня;
PS|68|18|не скрывай лица Твоего от раба Твоего, ибо я скорблю; скоро услышь меня;
PS|68|19|приблизься к душе моей, избавь ее; ради врагов моих спаси меня.
PS|68|20|Ты знаешь поношение мое, стыд мой и посрамление мое: враги мои все пред Тобою.
PS|68|21|Поношение сокрушило сердце мое, и я изнемог, ждал сострадания, но нет его, – утешителей, но не нахожу.
PS|68|22|И дали мне в пищу желчь, и в жажде моей напоили меня уксусом.
PS|68|23|Да будет трапеза их сетью им, и мирное пиршество их – западнею;
PS|68|24|да помрачатся глаза их, чтоб им не видеть, и чресла их расслабь навсегда;
PS|68|25|излей на них ярость Твою, и пламень гнева Твоего да обымет их;
PS|68|26|жилище их да будет пусто, и в шатрах их да не будет живущих,
PS|68|27|ибо, кого Ты поразил, они [еще] преследуют, и страдания уязвленных Тобою умножают.
PS|68|28|Приложи беззаконие к беззаконию их, и да не войдут они в правду Твою;
PS|68|29|да изгладятся они из книги живых и с праведниками да не напишутся.
PS|68|30|А я беден и страдаю; помощь Твоя, Боже, да восставит меня.
PS|68|31|Я буду славить имя Бога [моего] в песни, буду превозносить Его в славословии,
PS|68|32|и будет это благоугоднее Господу, нежели вол, нежели телец с рогами и с копытами.
PS|68|33|Увидят [это] страждущие и возрадуются. И оживет сердце ваше, ищущие Бога,
PS|68|34|ибо Господь внемлет нищим и не пренебрегает узников Своих.
PS|68|35|Да восхвалят Его небеса и земля, моря и все движущееся в них;
PS|68|36|ибо спасет Бог Сион, создаст города Иудины, и поселятся там и наследуют его,
PS|68|37|и потомство рабов Его утвердится в нем, и любящие имя Его будут поселяться на нем.
PS|69|1|Начальнику хора. Псалом Давида. В воспоминание.
PS|69|2|Поспеши, Боже, избавить меня, [поспеши], Господи, на помощь мне.
PS|69|3|Да постыдятся и посрамятся ищущие души моей! Да будут обращены назад и преданы посмеянию желающие мне зла!
PS|69|4|Да будут обращены назад за поношение меня говорящие [мне]: "хорошо! хорошо!"
PS|69|5|Да возрадуются и возвеселятся о Тебе все, ищущие Тебя, и любящие спасение Твое да говорят непрестанно: "велик Бог!"
PS|69|6|Я же беден и нищ; Боже, поспеши ко мне! Ты помощь моя и Избавитель мой; Господи! не замедли.
PS|70|1|На Тебя, Господи, уповаю, да не постыжусь вовек.
PS|70|2|По правде Твоей избавь меня и освободи меня; приклони ухо Твое ко мне и спаси меня.
PS|70|3|Будь мне твердым прибежищем, куда я всегда мог бы укрываться; Ты заповедал спасти меня, ибо твердыня моя и крепость моя – Ты.
PS|70|4|Боже мой! избавь меня из руки нечестивого, из руки беззаконника и притеснителя,
PS|70|5|ибо Ты – надежда моя, Господи Боже, упование мое от юности моей.
PS|70|6|На Тебе утверждался я от утробы; Ты извел меня из чрева матери моей; Тебе хвала моя не престанет.
PS|70|7|Для многих я был как бы дивом, но Ты твердая моя надежда.
PS|70|8|Да наполнятся уста мои хвалою, [чтобы воспевать] всякий день великолепие Твое.
PS|70|9|Не отвергни меня во время старости; когда будет оскудевать сила моя, не оставь меня,
PS|70|10|ибо враги мои говорят против меня, и подстерегающие душу мою советуются между собою,
PS|70|11|говоря: "Бог оставил его; преследуйте и схватите его, ибо нет избавляющего".
PS|70|12|Боже! не удаляйся от меня; Боже мой! поспеши на помощь мне.
PS|70|13|Да постыдятся и исчезнут враждующие против души моей, да покроются стыдом и бесчестием ищущие мне зла!
PS|70|14|А я всегда буду уповать [на Тебя] и умножать всякую хвалу Тебе.
PS|70|15|Уста мои будут возвещать правду Твою, всякий день благодеяния Твои; ибо я не знаю им числа.
PS|70|16|Войду в [размышление] о силах Господа Бога; воспомяну правду Твою – единственно Твою.
PS|70|17|Боже! Ты наставлял меня от юности моей, и доныне я возвещаю чудеса Твои.
PS|70|18|И до старости, и до седины не оставь меня, Боже, доколе не возвещу силы Твоей роду сему и всем грядущим могущества Твоего.
PS|70|19|Правда Твоя, Боже, до превыспренних; великие дела соделал Ты; Боже, кто подобен Тебе?
PS|70|20|Ты посылал на меня многие и лютые беды, но и опять оживлял меня и из бездн земли опять выводил меня.
PS|70|21|Ты возвышал меня и утешал меня.
PS|70|22|И я буду славить Тебя на псалтири, Твою истину, Боже мой; буду воспевать Тебя на гуслях, Святый Израилев!
PS|70|23|Радуются уста мои, когда я пою Тебе, и душа моя, которую Ты избавил;
PS|70|24|и язык мой всякий день будет возвещать правду Твою, ибо постыжены и посрамлены ищущие мне зла.
PS|71|1|О Соломоне. Боже! даруй царю Твой суд и сыну царя Твою правду,
PS|71|2|да судит праведно людей Твоих и нищих Твоих на суде;
PS|71|3|да принесут горы мир людям и холмы правду;
PS|71|4|да судит нищих народа, да спасет сынов убогого и смирит притеснителя, –
PS|71|5|и будут бояться Тебя, доколе пребудут солнце и луна, в роды родов.
PS|71|6|Он сойдет, как дождь на скошенный луг, как капли, орошающие землю;
PS|71|7|во дни его процветет праведник, и будет обилие мира, доколе не престанет луна;
PS|71|8|он будет обладать от моря до моря и от реки до концов земли;
PS|71|9|падут пред ним жители пустынь, и враги его будут лизать прах;
PS|71|10|цари Фарсиса и островов поднесут ему дань; цари Аравии и Савы принесут дары;
PS|71|11|и поклонятся ему все цари; все народы будут служить ему;
PS|71|12|ибо он избавит нищего, вопиющего и угнетенного, у которого нет помощника.
PS|71|13|Будет милосерд к нищему и убогому, и души убогих спасет;
PS|71|14|от коварства и насилия избавит души их, и драгоценна будет кровь их пред очами его;
PS|71|15|и будет жить, и будут давать ему от золота Аравии, и будут молиться о нем непрестанно, всякий день благословлять его;
PS|71|16|будет обилие хлеба на земле, наверху гор; плоды его будут волноваться, как [лес] на Ливане, и в городах размножатся люди, как трава на земле;
PS|71|17|будет имя его вовек; доколе пребывает солнце, будет передаваться имя его; и благословятся в нем [племена], все народы ублажат его.
PS|71|18|Благословен Господь Бог, Бог Израилев, един творящий чудеса,
PS|71|19|и благословенно имя славы Его вовек, и наполнится славою Его вся земля. Аминь и аминь.
PS|71|20|Кончились молитвы Давида, сына Иесеева.
PS|72|1|Псалом Асафа. Как благ Бог к Израилю, к чистым сердцем!
PS|72|2|А я – едва не пошатнулись ноги мои, едва не поскользнулись стопы мои, –
PS|72|3|я позавидовал безумным, видя благоденствие нечестивых,
PS|72|4|ибо им нет страданий до смерти их, и крепки силы их;
PS|72|5|на работе человеческой нет их, и с [прочими] людьми не подвергаются ударам.
PS|72|6|От того гордость, как ожерелье, обложила их, и дерзость, [как] наряд, одевает их;
PS|72|7|выкатились от жира глаза их, бродят помыслы в сердце;
PS|72|8|над всем издеваются, злобно разглашают клевету, говорят свысока;
PS|72|9|поднимают к небесам уста свои, и язык их расхаживает по земле.
PS|72|10|Потому туда же обращается народ Его, и пьют воду полною чашею,
PS|72|11|и говорят: "как узнает Бог? и есть ли ведение у Вышнего?"
PS|72|12|И вот, эти нечестивые благоденствуют в веке сем, умножают богатство.
PS|72|13|так не напрасно ли я очищал сердце мое и омывал в невинности руки мои,
PS|72|14|и подвергал себя ранам всякий день и обличениям всякое утро?
PS|72|15|[Но] если бы я сказал: "буду рассуждать так", – то я виновен был бы пред родом сынов Твоих.
PS|72|16|И думал я, как бы уразуметь это, но это трудно было в глазах моих,
PS|72|17|доколе не вошел я во святилище Божие и не уразумел конца их.
PS|72|18|Так! на скользких путях поставил Ты их и низвергаешь их в пропасти.
PS|72|19|Как нечаянно пришли они в разорение, исчезли, погибли от ужасов!
PS|72|20|Как сновидение по пробуждении, так Ты, Господи, пробудив [их], уничтожишь мечты их.
PS|72|21|Когда кипело сердце мое, и терзалась внутренность моя,
PS|72|22|тогда я был невежда и не разумел; как скот был я пред Тобою.
PS|72|23|Но я всегда с Тобою: Ты держишь меня за правую руку;
PS|72|24|Ты руководишь меня советом Твоим и потом примешь меня в славу.
PS|72|25|Кто мне на небе? и с Тобою ничего не хочу на земле.
PS|72|26|Изнемогает плоть моя и сердце мое: Бог твердыня сердца моего и часть моя вовек.
PS|72|27|Ибо вот, удаляющие себя от Тебя гибнут; Ты истребляешь всякого отступающего от Тебя.
PS|72|28|А мне благо приближаться к Богу! На Господа Бога я возложил упование мое, чтобы возвещать все дела Твои.
PS|73|1|Учение Асафа. Для чего, Боже, отринул нас навсегда? возгорелся гнев Твой на овец пажити Твоей?
PS|73|2|Вспомни сонм Твой, [который] Ты стяжал издревле, искупил в жезл достояния Твоего, – эту гору Сион, на которой Ты веселился.
PS|73|3|Подвигни стопы Твои к вековым развалинам: все разрушил враг во святилище.
PS|73|4|Рыкают враги Твои среди собраний Твоих; поставили знаки свои вместо знамений [наших];
PS|73|5|показывали себя подобными поднимающему вверх секиру на сплетшиеся ветви дерева;
PS|73|6|и ныне все резьбы в нем в один раз разрушили секирами и бердышами;
PS|73|7|предали огню святилище Твое; совсем осквернили жилище имени Твоего;
PS|73|8|сказали в сердце своем: "разорим их совсем", – и сожгли все места собраний Божиих на земле.
PS|73|9|Знамений наших мы не видим, нет уже пророка, и нет с нами, кто знал бы, доколе [это будет].
PS|73|10|Доколе, Боже, будет поносить враг? вечно ли будет хулить противник имя Твое?
PS|73|11|Для чего отклоняешь руку Твою и десницу Твою? Из среды недра Твоего порази [их].
PS|73|12|Боже, Царь мой от века, устрояющий спасение посреди земли!
PS|73|13|Ты расторг силою Твоею море, Ты сокрушил головы змиев в воде;
PS|73|14|Ты сокрушил голову левиафана, отдал его в пищу людям пустыни.
PS|73|15|Ты иссек источник и поток, Ты иссушил сильные реки.
PS|73|16|Твой день и Твоя ночь: Ты уготовал светила и солнце;
PS|73|17|Ты установил все пределы земли, лето и зиму Ты учредил.
PS|73|18|Вспомни же: враг поносит Господа, и люди безумные хулят имя Твое.
PS|73|19|Не предай зверям душу горлицы Твоей; собрания убогих Твоих не забудь навсегда.
PS|73|20|Призри на завет Твой; ибо наполнились все мрачные места земли жилищами насилия.
PS|73|21|Да не возвратится угнетенный посрамленным; нищий и убогий да восхвалят имя Твое.
PS|73|22|Восстань, Боже, защити дело Твое, вспомни вседневное поношение Твое от безумного;
PS|73|23|не забудь крика врагов Твоих; шум восстающих против Тебя непрестанно поднимается.
PS|74|1|Начальнику хора. Не погуби. Псалом Асафа. Песнь.
PS|74|2|Славим Тебя, Боже, славим, ибо близко имя Твое; возвещают чудеса Твои.
PS|74|3|"Когда изберу время, Я произведу суд по правде.
PS|74|4|Колеблется земля и все живущие на ней: Я утвержу столпы ее".
PS|74|5|Говорю безумствующим: "не безумствуйте", и нечестивым: "не поднимайте рога,
PS|74|6|не поднимайте высоко рога вашего, [не] говорите жестоковыйно",
PS|74|7|ибо не от востока и не от запада и не от пустыни возвышение,
PS|74|8|но Бог есть судия: одного унижает, а другого возносит;
PS|74|9|ибо чаша в руке Господа, вино кипит в ней, полное смешения, и Он наливает из нее. Даже дрожжи ее будут выжимать и пить все нечестивые земли.
PS|74|10|А я буду возвещать вечно, буду воспевать Бога Иаковлева,
PS|74|11|все роги нечестивых сломлю, и вознесутся роги праведника.
PS|75|1|Начальнику хора. На струнных [орудиях]. Псалом Асафа. Песнь.
PS|75|2|Ведом в Иудее Бог; у Израиля велико имя Его.
PS|75|3|И было в Салиме жилище Его и пребывание Его на Сионе.
PS|75|4|Там сокрушил Он стрелы лука, щит и меч и брань.
PS|75|5|Ты славен, могущественнее гор хищнических.
PS|75|6|Крепкие сердцем стали добычею, уснули сном своим, и не нашли все мужи силы рук своих.
PS|75|7|От прещения Твоего, Боже Иакова, вздремали и колесница и конь.
PS|75|8|Ты страшен, и кто устоит пред лицем Твоим во время гнева Твоего?
PS|75|9|С небес Ты возвестил суд; земля убоялась и утихла,
PS|75|10|когда восстал Бог на суд, чтобы спасти всех угнетенных земли.
PS|75|11|И гнев человеческий обратится во славу Тебе: остаток гнева Ты укротишь.
PS|75|12|Делайте и воздавайте обеты Господу, Богу вашему; все, которые вокруг Него, да принесут дары Страшному:
PS|75|13|Он укрощает дух князей, Он страшен для царей земных.
PS|76|1|Начальнику хора Идифумова. Псалом Асафа.
PS|76|2|Глас мой к Богу, и я буду взывать; глас мой к Богу, и Он услышит меня.
PS|76|3|В день скорби моей ищу Господа; рука моя простерта ночью и не опускается; душа моя отказывается от утешения.
PS|76|4|Вспоминаю о Боге и трепещу; помышляю, и изнемогает дух мой.
PS|76|5|Ты не даешь мне сомкнуть очей моих; я потрясен и не могу говорить.
PS|76|6|Размышляю о днях древних, о летах веков [минувших];
PS|76|7|припоминаю песни мои в ночи, беседую с сердцем моим, и дух мой испытывает:
PS|76|8|неужели навсегда отринул Господь, и не будет более благоволить?
PS|76|9|неужели навсегда престала милость Его, и пресеклось слово Его в род и род?
PS|76|10|неужели Бог забыл миловать? Неужели во гневе затворил щедроты Свои?
PS|76|11|И сказал я: "вот мое горе – изменение десницы Всевышнего".
PS|76|12|Буду вспоминать о делах Господа; буду вспоминать о чудесах Твоих древних;
PS|76|13|буду вникать во все дела Твои, размышлять о великих Твоих деяниях.
PS|76|14|Боже! свят путь Твой. Кто Бог так великий, как Бог [наш]!
PS|76|15|Ты – Бог, творящий чудеса; Ты явил могущество Свое среди народов;
PS|76|16|Ты избавил мышцею народ Твой, сынов Иакова и Иосифа.
PS|76|17|Видели Тебя, Боже, воды, видели Тебя воды и убоялись, и вострепетали бездны.
PS|76|18|Облака изливали воды, тучи издавали гром, и стрелы Твои летали.
PS|76|19|Глас грома Твоего в круге небесном; молнии освещали вселенную; земля содрогалась и тряслась.
PS|76|20|Путь Твой в море, и стезя Твоя в водах великих, и следы Твои неведомы.
PS|76|21|Как стадо, вел Ты народ Твой рукою Моисея и Аарона.
PS|77|1|Учение Асафа. Внимай, народ мой, закону моему, приклоните ухо ваше к словам уст моих.
PS|77|2|Открою уста мои в притче и произнесу гадания из древности.
PS|77|3|Что слышали мы и узнали, и отцы наши рассказали нам,
PS|77|4|не скроем от детей их, возвещая роду грядущему славу Господа, и силу Его, и чудеса Его, которые Он сотворил.
PS|77|5|Он постановил устав в Иакове и положил закон в Израиле, который заповедал отцам нашим возвещать детям их,
PS|77|6|чтобы знал грядущий род, дети, которые родятся, и чтобы они в свое время возвещали своим детям, –
PS|77|7|возлагать надежду свою на Бога и не забывать дел Божиих, и хранить заповеди Его,
PS|77|8|и не быть подобными отцам их, роду упорному и мятежному, неустроенному сердцем и неверному Богу духом своим.
PS|77|9|Сыны Ефремовы, вооруженные, стреляющие из луков, обратились назад в день брани:
PS|77|10|они не сохранили завета Божия и отреклись ходить в законе Его;
PS|77|11|забыли дела Его и чудеса, которые Он явил им.
PS|77|12|Он пред глазами отцов их сотворил чудеса в земле Египетской, на поле Цоан:
PS|77|13|разделил море, и провел их чрез него, и поставил воды стеною;
PS|77|14|и днем вел их облаком, а во всю ночь светом огня;
PS|77|15|рассек камень в пустыне и напоил их, как из великой бездны;
PS|77|16|из скалы извел потоки, и воды потекли, как реки.
PS|77|17|Но они продолжали грешить пред Ним и раздражать Всевышнего в пустыне:
PS|77|18|искушали Бога в сердце своем, требуя пищи по душе своей,
PS|77|19|и говорили против Бога и сказали: "может ли Бог приготовить трапезу в пустыне?"
PS|77|20|Вот, Он ударил в камень, и потекли воды, и полились ручьи. "Может ли Он дать и хлеб, может ли приготовлять мясо народу Своему?"
PS|77|21|Господь услышал и воспламенился гневом, и огонь возгорелся на Иакова, и гнев подвигнулся на Израиля
PS|77|22|за то, что не веровали в Бога и не уповали на спасение Его.
PS|77|23|Он повелел облакам свыше и отверз двери неба,
PS|77|24|и одождил на них манну в пищу, и хлеб небесный дал им.
PS|77|25|Хлеб ангельский ел человек; послал Он им пищу до сытости.
PS|77|26|Он возбудил на небе восточный ветер и навел южный силою Своею
PS|77|27|и, как пыль, одождил на них мясо и, как песок морской, птиц пернатых:
PS|77|28|поверг их среди стана их, около жилищ их, –
PS|77|29|и они ели и пресытились; и желаемое ими дал им.
PS|77|30|Но еще не прошла прихоть их, еще пища была в устах их,
PS|77|31|гнев Божий пришел на них, убил тучных их и юношей Израилевых низложил.
PS|77|32|При всем этом они продолжали грешить и не верили чудесам Его.
PS|77|33|И погубил дни их в суете и лета их в смятении.
PS|77|34|Когда Он убивал их, они искали Его и обращались, и с раннего утра прибегали к Богу,
PS|77|35|и вспоминали, что Бог – их прибежище, и Бог Всевышний – Избавитель их,
PS|77|36|и льстили Ему устами своими и языком своим лгали пред Ним;
PS|77|37|сердце же их было неправо пред Ним, и они не были верны завету Его.
PS|77|38|Но Он, Милостивый, прощал грех и не истреблял их, многократно отвращал гнев Свой и не возбуждал всей ярости Своей:
PS|77|39|Он помнил, что они плоть, дыхание, которое уходит и не возвращается.
PS|77|40|Сколько раз они раздражали Его в пустыне и прогневляли Его в [стране] необитаемой!
PS|77|41|и снова искушали Бога и оскорбляли Святаго Израилева,
PS|77|42|не помнили руки Его, дня, когда Он избавил их от угнетения,
PS|77|43|когда сотворил в Египте знамения Свои и чудеса Свои на поле Цоан;
PS|77|44|и превратил реки их и потоки их в кровь, чтобы они не могли пить;
PS|77|45|послал на них насекомых, чтобы жалили их, и жаб, чтобы губили их;
PS|77|46|земные произрастения их отдал гусенице и труд их – саранче;
PS|77|47|виноград их побил градом и сикоморы их – льдом;
PS|77|48|скот их предал граду и стада их – молниям;
PS|77|49|послал на них пламень гнева Своего, и негодование, и ярость и бедствие, посольство злых ангелов;
PS|77|50|уравнял стезю гневу Своему, не охранял души их от смерти, и скот их предал моровой язве;
PS|77|51|поразил всякого первенца в Египте, начатки сил в шатрах Хамовых;
PS|77|52|и повел народ Свой, как овец, и вел их, как стадо, пустынею;
PS|77|53|вел их безопасно, и они не страшились, а врагов их покрыло море;
PS|77|54|и привел их в область святую Свою, на гору сию, которую стяжала десница Его;
PS|77|55|прогнал от лица их народы и землю их разделил в наследие им, и колена Израилевы поселил в шатрах их.
PS|77|56|Но они еще искушали и огорчали Бога Всевышнего, и уставов Его не сохраняли;
PS|77|57|отступали и изменяли, как отцы их, обращались назад, как неверный лук;
PS|77|58|огорчали Его высотами своими и истуканами своими возбуждали ревность Его.
PS|77|59|Услышал Бог и воспламенился гневом и сильно вознегодовал на Израиля;
PS|77|60|отринул жилище в Силоме, скинию, в которой обитал Он между человеками;
PS|77|61|и отдал в плен крепость Свою и славу Свою в руки врага,
PS|77|62|и предал мечу народ Свой и прогневался на наследие Свое.
PS|77|63|Юношей его поедал огонь, и девицам его не пели брачных песен;
PS|77|64|священники его падали от меча, и вдовы его не плакали.
PS|77|65|Но, как бы от сна, воспрянул Господь, как бы исполин, побежденный вином,
PS|77|66|и поразил врагов его в тыл, вечному сраму предал их;
PS|77|67|и отверг шатер Иосифов и колена Ефремова не избрал,
PS|77|68|а избрал колено Иудино, гору Сион, которую возлюбил.
PS|77|69|И устроил, как небо, святилище Свое и, как землю, утвердил его навек,
PS|77|70|и избрал Давида, раба Своего, и взял его от дворов овчих
PS|77|71|и от доящих привел его пасти народ Свой, Иакова, и наследие Свое, Израиля.
PS|77|72|И он пас их в чистоте сердца своего и руками мудрыми водил их.
PS|78|1|Псалом Асафа. Боже! язычники пришли в наследие Твое, осквернили святый храм Твой, Иерусалим превратили в развалины;
PS|78|2|трупы рабов Твоих отдали на съедение птицам небесным, тела святых Твоих – зверям земным;
PS|78|3|пролили кровь их, как воду, вокруг Иерусалима, и некому было похоронить их.
PS|78|4|Мы сделались посмешищем у соседей наших, поруганием и посрамлением у окружающих нас.
PS|78|5|Доколе, Господи, будешь гневаться непрестанно, будет пылать ревность Твоя, как огонь?
PS|78|6|Пролей гнев Твой на народы, которые не знают Тебя, и на царства, которые имени Твоего не призывают,
PS|78|7|ибо они пожрали Иакова и жилище его опустошили.
PS|78|8|Не помяни нам грехов [наших] предков; скоро да предварят нас щедроты Твои, ибо мы весьма истощены.
PS|78|9|Помоги нам, Боже, Спаситель наш, ради славы имени Твоего; избавь нас и прости нам грехи наши ради имени Твоего.
PS|78|10|Для чего язычникам говорить: "где Бог их?" Да сделается известным между язычниками пред глазами нашими отмщение за пролитую кровь рабов Твоих.
PS|78|11|Да придет пред лице Твое стенание узника; могуществом мышцы Твоей сохрани обреченных на смерть.
PS|78|12|Семикратно возврати соседям нашим в недро их поношение, которым они Тебя, Господи, поносили.
PS|78|13|А мы, народ Твой и Твоей пажити овцы, вечно будем славить Тебя и в род и род возвещать хвалу Тебе.
PS|79|1|Начальнику хора. На музыкальном [орудии] Шошанним–Эдуф. Псалом Асафа.
PS|79|2|Пастырь Израиля! внемли; водящий, как овец, Иосифа, восседающий на Херувимах, яви Себя.
PS|79|3|Пред Ефремом и Вениамином и Манассиею воздвигни силу Твою, и приди спасти нас.
PS|79|4|Боже! восстанови нас; да воссияет лице Твое, и спасемся!
PS|79|5|Господи, Боже сил! доколе будешь гневен к молитвам народа Твоего?
PS|79|6|Ты напитал их хлебом слезным, и напоил их слезами в большой мере,
PS|79|7|положил нас в пререкание соседям нашим, и враги наши издеваются [над нами].
PS|79|8|Боже сил! восстанови нас; да воссияет лице Твое, и спасемся!
PS|79|9|Из Египта перенес Ты виноградную лозу, выгнал народы и посадил ее;
PS|79|10|очистил для нее место, и утвердил корни ее, и она наполнила землю.
PS|79|11|Горы покрылись тенью ее, и ветви ее как кедры Божии;
PS|79|12|она пустила ветви свои до моря и отрасли свои до реки.
PS|79|13|Для чего разрушил Ты ограды ее, так что обрывают ее все, проходящие по пути?
PS|79|14|Лесной вепрь подрывает ее, и полевой зверь объедает ее.
PS|79|15|Боже сил! обратись же, призри с неба, и воззри, и посети виноград сей;
PS|79|16|охрани то, что насадила десница Твоя, и отрасли, которые Ты укрепил Себе.
PS|79|17|Он пожжен огнем, обсечен; от прещения лица Твоего погибнут.
PS|79|18|Да будет рука Твоя над мужем десницы Твоей, над сыном человеческим, которого Ты укрепил Себе,
PS|79|19|и мы не отступим от Тебя; оживи нас, и мы будем призывать имя Твое.
PS|79|20|Господи, Боже сил! восстанови нас; да воссияет лице Твое, и спасемся!
PS|80|1|Начальнику хора. На Гефском орудии. Псалом Асафа.
PS|80|2|Радостно пойте Богу, твердыне нашей; восклицайте Богу Иакова;
PS|80|3|возьмите псалом, дайте тимпан, сладкозвучные гусли с псалтирью;
PS|80|4|трубите в новомесячие трубою, в определенное время, в день праздника нашего;
PS|80|5|ибо это закон для Израиля, устав от Бога Иаковлева.
PS|80|6|Он установил это во свидетельство для Иосифа, когда он вышел из земли Египетской, где услышал звуки языка, которого не знал:
PS|80|7|"Я снял с рамен его тяжести, и руки его освободились от корзин.
PS|80|8|В бедствии ты призвал Меня, и Я избавил тебя; из среды грома Я услышал тебя, при водах Меривы испытал тебя.
PS|80|9|Слушай, народ Мой, и Я буду свидетельствовать тебе: Израиль! о, если бы ты послушал Меня!
PS|80|10|Да не будет у тебя иного бога, и не поклоняйся богу чужеземному.
PS|80|11|Я Господь, Бог твой, изведший тебя из земли Египетской; открой уста твои, и Я наполню их".
PS|80|12|Но народ Мой не слушал гласа Моего, и Израиль не покорялся Мне;
PS|80|13|потому Я оставил их упорству сердца их, пусть ходят по своим помыслам.
PS|80|14|О, если бы народ Мой слушал Меня и Израиль ходил Моими путями!
PS|80|15|Я скоро смирил бы врагов их и обратил бы руку Мою на притеснителей их:
PS|80|16|ненавидящие Господа раболепствовали бы им, а их благоденствие продолжалось бы навсегда;
PS|80|17|Я питал бы их туком пшеницы и насыщал бы их медом из скалы.
PS|81|1|Псалом Асафа. Бог стал в сонме богов; среди богов произнес суд:
PS|81|2|доколе будете вы судить неправедно и оказывать лицеприятие нечестивым?
PS|81|3|Давайте суд бедному и сироте; угнетенному и нищему оказывайте справедливость;
PS|81|4|избавляйте бедного и нищего; исторгайте [его] из руки нечестивых.
PS|81|5|Не знают, не разумеют, во тьме ходят; все основания земли колеблются.
PS|81|6|Я сказал: вы – боги, и сыны Всевышнего – все вы;
PS|81|7|но вы умрете, как человеки, и падете, как всякий из князей.
PS|81|8|Восстань, Боже, суди землю, ибо Ты наследуешь все народы.
PS|82|1|Песнь. Псалом Асафа.
PS|82|2|Боже! Не премолчи, не безмолвствуй и не оставайся в покое, Боже,
PS|82|3|ибо вот, враги Твои шумят, и ненавидящие Тебя подняли голову;
PS|82|4|против народа Твоего составили коварный умысел и совещаются против хранимых Тобою;
PS|82|5|сказали: "пойдем и истребим их из народов, чтобы не вспоминалось более имя Израиля."
PS|82|6|Сговорились единодушно, заключили против Тебя союз:
PS|82|7|селения Едомовы и Измаильтяне, Моав и Агаряне,
PS|82|8|Гевал и Аммон и Амалик, Филистимляне с жителями Тира.
PS|82|9|И Ассур пристал к ним: они стали мышцею для сынов Лотовых.
PS|82|10|Сделай им то же, что Мадиаму, что Сисаре, что Иавину у потока Киссона,
PS|82|11|которые истреблены в Аендоре, сделались навозом для земли.
PS|82|12|Поступи с ними, с князьями их, как с Оривом и Зивом и со всеми вождями их, как с Зевеем и Салманом,
PS|82|13|которые говорили: "возьмем себе во владение селения Божии".
PS|82|14|Боже мой! Да будут они, как пыль в вихре, как солома перед ветром.
PS|82|15|Как огонь сжигает лес, и как пламя опаляет горы,
PS|82|16|так погони их бурею Твоею и вихрем Твоим приведи их в смятение;
PS|82|17|исполни лица их бесчестием, чтобы они взыскали имя Твое, Господи!
PS|82|18|Да постыдятся и смятутся на веки, да посрамятся и погибнут,
PS|82|19|и да познают, что Ты, Которого одного имя Господь, Всевышний над всею землею.
PS|83|1|Начальнику хора. На Гефском [орудии]. Кореевых сынов. Псалом.
PS|83|2|Как вожделенны жилища Твои, Господи сил!
PS|83|3|Истомилась душа моя, желая во дворы Господни; сердце мое и плоть моя восторгаются к Богу живому.
PS|83|4|И птичка находит себе жилье, и ласточка гнездо себе, где положить птенцов своих, у алтарей Твоих, Господи сил, Царь мой и Бог мой!
PS|83|5|Блаженны живущие в доме Твоем: они непрестанно будут восхвалять Тебя.
PS|83|6|Блажен человек, которого сила в Тебе и у которого в сердце стези направлены [к Тебе].
PS|83|7|Проходя долиною плача, они открывают в ней источники, и дождь покрывает ее благословением;
PS|83|8|приходят от силы в силу, являются пред Богом на Сионе.
PS|83|9|Господи, Боже сил! Услышь молитву мою, внемли, Боже Иаковлев!
PS|83|10|Боже, защитник наш! Приникни и призри на лице помазанника Твоего.
PS|83|11|Ибо один день во дворах Твоих лучше тысячи. Желаю лучше быть у порога в доме Божием, нежели жить в шатрах нечестия.
PS|83|12|Ибо Господь Бог есть солнце и щит, Господь дает благодать и славу; ходящих в непорочности Он не лишает благ.
PS|83|13|Господи сил! Блажен человек, уповающий на Тебя!
PS|84|1|Начальнику хора. Кореевых сынов. Псалом.
PS|84|2|Господи! Ты умилосердился к земле Твоей, возвратил плен Иакова;
PS|84|3|простил беззаконие народа Твоего, покрыл все грехи его,
PS|84|4|отъял всю ярость Твою, отвратил лютость гнева Твоего.
PS|84|5|Восстанови нас, Боже спасения нашего, и прекрати негодование Твое на нас.
PS|84|6|Неужели вечно будешь гневаться на нас, прострешь гнев Твой от рода в род?
PS|84|7|Неужели снова не оживишь нас, чтобы народ Твой возрадовался о Тебе?
PS|84|8|Яви нам, Господи, милость Твою, и спасение Твое даруй нам.
PS|84|9|Послушаю, что скажет Господь Бог. Он скажет мир народу Своему и избранным Своим, но да не впадут они снова в безрассудство.
PS|84|10|Так, близко к боящимся Его спасение Его, чтобы обитала слава в земле нашей!
PS|84|11|Милость и истина сретятся, правда и мир облобызаются;
PS|84|12|истина возникнет из земли, и правда приникнет с небес;
PS|84|13|и Господь даст благо, и земля наша даст плод свой;
PS|84|14|правда пойдет пред Ним и поставит на путь стопы свои.
PS|85|1|Молитва Давида. Приклони, Господи, ухо Твое и услышь меня, ибо я беден и нищ.
PS|85|2|Сохрани душу мою, ибо я благоговею пред Тобою; спаси, Боже мой, раба Твоего, уповающего на Тебя.
PS|85|3|Помилуй меня, Господи, ибо к Тебе взываю каждый день.
PS|85|4|Возвесели душу раба Твоего, ибо к Тебе, Господи, возношу душу мою,
PS|85|5|ибо Ты, Господи, благ и милосерд и многомилостив ко всем, призывающим Тебя.
PS|85|6|Услышь, Господи, молитву мою и внемли гласу моления моего.
PS|85|7|В день скорби моей взываю к Тебе, потому что Ты услышишь меня.
PS|85|8|Нет между богами, как Ты, Господи, и нет дел, как Твои.
PS|85|9|Все народы, Тобою сотворенные, приидут и поклонятся пред Тобою, Господи, и прославят имя Твое,
PS|85|10|ибо Ты велик и творишь чудеса, – Ты, Боже, един Ты.
PS|85|11|Наставь меня, Господи, на путь Твой, и буду ходить в истине Твоей; утверди сердце мое в страхе имени Твоего.
PS|85|12|Буду восхвалять Тебя, Господи, Боже мой, всем сердцем моим и славить имя Твое вечно,
PS|85|13|ибо велика милость Твоя ко мне: Ты избавил душу мою от ада преисподнего.
PS|85|14|Боже! гордые восстали на меня, и скопище мятежников ищет души моей: не представляют они Тебя пред собою.
PS|85|15|Но Ты, Господи, Боже щедрый и благосердный, долготерпеливый и многомилостивый и истинный,
PS|85|16|призри на меня и помилуй меня; даруй крепость Твою рабу Твоему, и спаси сына рабы Твоей;
PS|85|17|покажи на мне знамение во благо, да видят ненавидящие меня и устыдятся, потому что Ты, Господи, помог мне и утешил меня.
PS|86|1|Сынов Кореевых. Псалом. Песнь.
PS|86|2|Основание его на горах святых. Господь любит врата Сиона более всех селений Иакова.
PS|86|3|Славное возвещается о тебе, град Божий!
PS|86|4|Упомяну знающим меня о Рааве и Вавилоне; вот Филистимляне и Тир с Ефиопиею, – [скажут]: "такой–то родился там".
PS|86|5|О Сионе же будут говорить: "такой–то и такой–то муж родился в нем, и Сам Всевышний укрепил его".
PS|86|6|Господь в переписи народов напишет: "такой–то родился там".
PS|86|7|И поющие и играющие, – все источники мои в тебе.
PS|87|1|Песнь. Псалом, Сынов Кореевых. Начальнику хора на Махалаф, для пения. Учение Емана Езрахита.
PS|87|2|Господи, Боже спасения моего! днем вопию и ночью пред Тобою:
PS|87|3|да внидет пред лице Твое молитва моя; приклони ухо Твое к молению моему,
PS|87|4|ибо душа моя насытилась бедствиями, и жизнь моя приблизилась к преисподней.
PS|87|5|Я сравнялся с нисходящими в могилу; я стал, как человек без силы,
PS|87|6|между мертвыми брошенный, – как убитые, лежащие во гробе, о которых Ты уже не вспоминаешь и которые от руки Твоей отринуты.
PS|87|7|Ты положил меня в ров преисподний, во мрак, в бездну.
PS|87|8|Отяготела на мне ярость Твоя, и всеми волнами Твоими Ты поразил [меня].
PS|87|9|Ты удалил от меня знакомых моих, сделал меня отвратительным для них; я заключен, и не могу выйти.
PS|87|10|Око мое истомилось от горести: весь день я взывал к Тебе, Господи, простирал к Тебе руки мои.
PS|87|11|Разве над мертвыми Ты сотворишь чудо? Разве мертвые встанут и будут славить Тебя?
PS|87|12|или во гробе будет возвещаема милость Твоя, и истина Твоя – в месте тления?
PS|87|13|разве во мраке познают чудеса Твои, и в земле забвения – правду Твою?
PS|87|14|Но я к Тебе, Господи, взываю, и рано утром молитва моя предваряет Тебя.
PS|87|15|Для чего, Господи, отреваешь душу мою, скрываешь лице Твое от меня?
PS|87|16|Я несчастен и истаеваю с юности; несу ужасы Твои и изнемогаю.
PS|87|17|Надо мною прошла ярость Твоя, устрашения Твои сокрушили меня,
PS|87|18|всякий день окружают меня, как вода: облегают меня все вместе.
PS|87|19|Ты удалил от меня друга и искреннего; знакомых моих не видно.
PS|88|1|Учение Ефама Езрахита.
PS|88|2|Милости [Твои], Господи, буду петь вечно, в род и род возвещать истину Твою устами моими.
PS|88|3|Ибо говорю: навек основана милость, на небесах утвердил Ты истину Твою, [когда сказал]:
PS|88|4|"Я поставил завет с избранным Моим, клялся Давиду, рабу Моему:
PS|88|5|навек утвержу семя твое, в род и род устрою престол твой".
PS|88|6|И небеса прославят чудные дела Твои, Господи, и истину Твою в собрании святых.
PS|88|7|Ибо кто на небесах сравнится с Господом? кто между сынами Божиими уподобится Господу?
PS|88|8|Страшен Бог в великом сонме святых, страшен Он для всех окружающих Его.
PS|88|9|Господи, Боже сил! кто силен, как Ты, Господи? И истина Твоя окрест Тебя.
PS|88|10|Ты владычествуешь над яростью моря: когда воздымаются волны его, Ты укрощаешь их.
PS|88|11|Ты низложил Раава, как пораженного; крепкою мышцею Твоею рассеял врагов Твоих.
PS|88|12|Твои небеса и Твоя земля; вселенную и что наполняет ее, Ты основал.
PS|88|13|Север и юг Ты сотворил; Фавор и Ермон о имени Твоем радуются.
PS|88|14|Крепка мышца Твоя, сильна рука Твоя, высока десница Твоя!
PS|88|15|Правосудие и правота – основание престола Твоего; милость и истина предходят пред лицем Твоим.
PS|88|16|Блажен народ, знающий трубный зов! Они ходят во свете лица Твоего, Господи,
PS|88|17|о имени Твоем радуются весь день и правдою Твоею возносятся,
PS|88|18|ибо Ты украшение силы их, и благоволением Твоим возвышается рог наш.
PS|88|19|От Господа – щит наш, и от Святаго Израилева – царь наш.
PS|88|20|Некогда говорил Ты в видении святому Твоему, и сказал: "Я оказал помощь мужественному, вознес избранного из народа.
PS|88|21|Я обрел Давида, раба Моего, святым елеем Моим помазал его.
PS|88|22|Рука Моя пребудет с ним, и мышца Моя укрепит его.
PS|88|23|Враг не превозможет его, и сын беззакония не притеснит его.
PS|88|24|Сокрушу пред ним врагов его и поражу ненавидящих его.
PS|88|25|И истина Моя и милость Моя с ним, и Моим именем возвысится рог его.
PS|88|26|И положу на море руку его, и на реки – десницу его.
PS|88|27|Он будет звать Меня: Ты отец мой, Бог мой и твердыня спасения моего.
PS|88|28|И Я сделаю его первенцем, превыше царей земли,
PS|88|29|вовек сохраню ему милость Мою, и завет Мой с ним будет верен.
PS|88|30|И продолжу вовек семя его, и престол его – как дни неба.
PS|88|31|Если сыновья его оставят закон Мой и не будут ходить по заповедям Моим;
PS|88|32|если нарушат уставы Мои и повелений Моих не сохранят:
PS|88|33|посещу жезлом беззаконие их, и ударами – неправду их;
PS|88|34|милости же Моей не отниму от него, и не изменю истины Моей.
PS|88|35|Не нарушу завета Моего, и не переменю того, что вышло из уст Моих.
PS|88|36|Однажды Я поклялся святостью Моею: солгу ли Давиду?
PS|88|37|Семя его пребудет вечно, и престол его, как солнце, предо Мною,
PS|88|38|вовек будет тверд, как луна, и верный свидетель на небесах".
PS|88|39|Но [ныне] Ты отринул и презрел, прогневался на помазанника Твоего;
PS|88|40|пренебрег завет с рабом Твоим, поверг на землю венец его;
PS|88|41|разрушил все ограды его, превратил в развалины крепости его.
PS|88|42|Расхищают его все проходящие путем; он сделался посмешищем у соседей своих.
PS|88|43|Ты возвысил десницу противников его, обрадовал всех врагов его;
PS|88|44|Ты обратил назад острие меча его и не укрепил его на брани;
PS|88|45|отнял у него блеск и престол его поверг на землю;
PS|88|46|сократил дни юности его и покрыл его стыдом.
PS|88|47|Доколе, Господи, будешь скрываться непрестанно, будет пылать ярость Твоя, как огонь?
PS|88|48|Вспомни, какой мой век: на какую суету сотворил Ты всех сынов человеческих?
PS|88|49|Кто из людей жил – и не видел смерти, избавил душу свою от руки преисподней?
PS|88|50|Где прежние милости Твои, Господи? Ты клялся Давиду истиною Твоею.
PS|88|51|Вспомни, Господи, поругание рабов Твоих, которое я ношу в недре моем от всех сильных народов;
PS|88|52|как поносят враги Твои, Господи, как бесславят следы помазанника Твоего.
PS|88|53|Благословен Господь вовек! Аминь, аминь.
PS|89|1|Молитва Моисея, человека Божия.
PS|89|2|Господи! Ты нам прибежище в род и род.
PS|89|3|Прежде нежели родились горы, и Ты образовал землю и вселенную, и от века и до века Ты – Бог.
PS|89|4|Ты возвращаешь человека в тление и говоришь: "возвратитесь, сыны человеческие!"
PS|89|5|Ибо пред очами Твоими тысяча лет, как день вчерашний, когда он прошел, и [как] стража в ночи.
PS|89|6|Ты [как] наводнением уносишь их; они – [как] сон, как трава, которая утром вырастает, утром цветет и зеленеет, вечером подсекается и засыхает;
PS|89|7|ибо мы исчезаем от гнева Твоего и от ярости Твоей мы в смятении.
PS|89|8|Ты положил беззакония наши пред Тобою и тайное наше пред светом лица Твоего.
PS|89|9|Все дни наши прошли во гневе Твоем; мы теряем лета наши, как звук.
PS|89|10|Дней лет наших – семьдесят лет, а при большей крепости – восемьдесят лет; и самая лучшая пора их – труд и болезнь, ибо проходят быстро, и мы летим.
PS|89|11|Кто знает силу гнева Твоего, и ярость Твою по мере страха Твоего?
PS|89|12|Научи нас так счислять дни наши, чтобы нам приобрести сердце мудрое.
PS|89|13|Обратись, Господи! Доколе? Умилосердись над рабами Твоими.
PS|89|14|Рано насыти нас милостью Твоею, и мы будем радоваться и веселиться во все дни наши.
PS|89|15|Возвесели нас за дни, [в которые] Ты поражал нас, за лета, [в которые] мы видели бедствие.
PS|89|16|Да явится на рабах Твоих дело Твое и на сынах их слава Твоя;
PS|89|17|и да будет благоволение Господа Бога нашего на нас, и в деле рук наших споспешествуй нам, в деле рук наших споспешествуй.
PS|90|1|Живущий под кровом Всевышнего под сенью Всемогущего покоится,
PS|90|2|говорит Господу: "прибежище мое и защита моя, Бог мой, на Которого я уповаю!"
PS|90|3|Он избавит тебя от сети ловца, от гибельной язвы,
PS|90|4|перьями Своими осенит тебя, и под крыльями Его будешь безопасен; щит и ограждение – истина Его.
PS|90|5|Не убоишься ужасов в ночи, стрелы, летящей днем,
PS|90|6|язвы, ходящей во мраке, заразы, опустошающей в полдень.
PS|90|7|Падут подле тебя тысяча и десять тысяч одесную тебя; но к тебе не приблизится:
PS|90|8|только смотреть будешь очами твоими и видеть возмездие нечестивым.
PS|90|9|Ибо ты [сказал]: "Господь – упование мое"; Всевышнего избрал ты прибежищем твоим;
PS|90|10|не приключится тебе зло, и язва не приблизится к жилищу твоему;
PS|90|11|ибо Ангелам Своим заповедает о тебе – охранять тебя на всех путях твоих:
PS|90|12|на руках понесут тебя, да не преткнешься о камень ногою твоею;
PS|90|13|на аспида и василиска наступишь; попирать будешь льва и дракона.
PS|90|14|"За то, что он возлюбил Меня, избавлю его; защищу его, потому что он познал имя Мое.
PS|90|15|Воззовет ко Мне, и услышу его; с ним Я в скорби; избавлю его и прославлю его,
PS|90|16|долготою дней насыщу его, и явлю ему спасение Мое".
PS|91|1|Псалом. Песнь на день субботний.
PS|91|2|Благо есть славить Господа и петь имени Твоему, Всевышний,
PS|91|3|возвещать утром милость Твою и истину Твою в ночи,
PS|91|4|на десятиструнном и псалтири, с песнью на гуслях.
PS|91|5|Ибо Ты возвеселил меня, Господи, творением Твоим: я восхищаюсь делами рук Твоих.
PS|91|6|Как велики дела Твои, Господи! дивно глубоки помышления Твои!
PS|91|7|Человек несмысленный не знает, и невежда не разумеет того.
PS|91|8|Тогда как нечестивые возникают, как трава, и делающие беззаконие цветут, чтобы исчезнуть на веки, –
PS|91|9|Ты, Господи, высок во веки!
PS|91|10|Ибо вот, враги Твои, Господи, – вот, враги Твои гибнут, и рассыпаются все делающие беззаконие;
PS|91|11|а мой рог Ты возносишь, как рог единорога, и я умащен свежим елеем;
PS|91|12|и око мое смотрит на врагов моих, и уши мои слышат о восстающих на меня злодеях.
PS|91|13|Праведник цветет, как пальма, возвышается подобно кедру на Ливане.
PS|91|14|Насажденные в доме Господнем, они цветут во дворах Бога нашего;
PS|91|15|они и в старости плодовиты, сочны и свежи,
PS|91|16|чтобы возвещать, что праведен Господь, твердыня моя, и нет неправды в Нем.
PS|92|1|Господь царствует; Он облечен величием, облечен Господь могуществом [и] препоясан: потому вселенная тверда, не подвигнется.
PS|92|2|Престол Твой утвержден искони: Ты – от века.
PS|92|3|Возвышают реки, Господи, возвышают реки голос свой, возвышают реки волны свои.
PS|92|4|Но паче шума вод многих, сильных волн морских, силен в вышних Господь.
PS|92|5|Откровения Твои несомненно верны. Дому Твоему, Господи, принадлежит святость на долгие дни.
PS|93|1|Боже отмщений, Господи, Боже отмщений, яви Себя!
PS|93|2|Восстань, Судия земли, воздай возмездие гордым.
PS|93|3|Доколе, Господи, нечестивые, доколе нечестивые торжествовать будут?
PS|93|4|Они изрыгают дерзкие речи; величаются все делающие беззаконие;
PS|93|5|попирают народ Твой, Господи, угнетают наследие Твое;
PS|93|6|вдову и пришельца убивают, и сирот умерщвляют
PS|93|7|и говорят: "не увидит Господь, и не узнает Бог Иаковлев".
PS|93|8|Образумьтесь, бессмысленные люди! когда вы будете умны, невежды?
PS|93|9|Насадивший ухо не услышит ли? и образовавший глаз не увидит ли?
PS|93|10|Вразумляющий народы неужели не обличит, – Тот, Кто учит человека разумению?
PS|93|11|Господь знает мысли человеческие, что они суетны.
PS|93|12|Блажен человек, которого вразумляешь Ты, Господи, и наставляешь законом Твоим,
PS|93|13|чтобы дать ему покой в бедственные дни, доколе нечестивому выроется яма!
PS|93|14|Ибо не отринет Господь народа Своего и не оставит наследия Своего.
PS|93|15|Ибо суд возвратится к правде, и за ним [последуют] все правые сердцем.
PS|93|16|Кто восстанет за меня против злодеев? кто станет за меня против делающих беззаконие?
PS|93|17|Если бы не Господь был мне помощником, вскоре вселилась бы душа моя в [страну] молчания.
PS|93|18|Когда я говорил: "колеблется нога моя", – милость Твоя, Господи, поддерживала меня.
PS|93|19|При умножении скорбей моих в сердце моем, утешения Твои услаждают душу мою.
PS|93|20|Станет ли близ Тебя седалище губителей, умышляющих насилие вопреки закону?
PS|93|21|Толпою устремляются они на душу праведника и осуждают кровь неповинную.
PS|93|22|Но Господь – защита моя, и Бог мой – твердыня убежища моего,
PS|93|23|и обратит на них беззаконие их, и злодейством их истребит их, истребит их Господь Бог наш.
PS|94|1|Приидите, воспоем Господу, воскликнем твердыне спасения нашего;
PS|94|2|предстанем лицу Его со славословием, в песнях воскликнем Ему,
PS|94|3|ибо Господь есть Бог великий и Царь великий над всеми богами.
PS|94|4|В Его руке глубины земли, и вершины гор – Его же;
PS|94|5|Его – море, и Он создал его, и сушу образовали руки Его.
PS|94|6|Приидите, поклонимся и припадем, преклоним колени пред лицем Господа, Творца нашего;
PS|94|7|ибо Он есть Бог наш, и мы – народ паствы Его и овцы руки Его. О, если бы вы ныне послушали гласа Его:
PS|94|8|"не ожесточите сердца вашего, как в Мериве, как в день искушения в пустыне,
PS|94|9|где искушали Меня отцы ваши, испытывали Меня, и видели дело Мое.
PS|94|10|Сорок лет Я был раздражаем родом сим, и сказал: это народ, заблуждающийся сердцем; они не познали путей Моих,
PS|94|11|и потому Я поклялся во гневе Моем, что они не войдут в покой Мой".
PS|95|1|Воспойте Господу песнь новую; воспойте Господу, вся земля;
PS|95|2|пойте Господу, благословляйте имя Его, благовествуйте со дня на день спасение Его;
PS|95|3|возвещайте в народах славу Его, во всех племенах чудеса Его;
PS|95|4|ибо велик Господь и достохвален, страшен Он паче всех богов.
PS|95|5|Ибо все боги народов – идолы, а Господь небеса сотворил.
PS|95|6|Слава и величие пред лицем Его, сила и великолепие во святилище Его.
PS|95|7|Воздайте Господу, племена народов, воздайте Господу славу и честь;
PS|95|8|воздайте Господу славу имени Его, несите дары и идите во дворы Его;
PS|95|9|поклонитесь Господу во благолепии святыни. Трепещи пред лицем Его, вся земля!
PS|95|10|Скажите народам: Господь царствует! потому тверда вселенная, не поколеблется. Он будет судить народы по правде.
PS|95|11|Да веселятся небеса и да торжествует земля; да шумит море и что наполняет его;
PS|95|12|да радуется поле и все, что на нем, и да ликуют все дерева дубравные
PS|95|13|пред лицем Господа; ибо идет, ибо идет судить землю. Он будет судить вселенную по правде, и народы – по истине Своей.
PS|96|1|Господь царствует: да радуется земля; да веселятся многочисленные острова.
PS|96|2|Облако и мрак окрест Его; правда и суд – основание престола Его.
PS|96|3|Пред Ним идет огонь и вокруг попаляет врагов Его.
PS|96|4|Молнии Его освещают вселенную; земля видит и трепещет.
PS|96|5|Горы, как воск, тают от лица Господа, от лица Господа всей земли.
PS|96|6|Небеса возвещают правду Его, и все народы видят славу Его.
PS|96|7|Да постыдятся все служащие истуканам, хвалящиеся идолами. Поклонитесь пред Ним, все боги.
PS|96|8|Слышит Сион и радуется, и веселятся дщери Иудины ради судов Твоих, Господи,
PS|96|9|ибо Ты, Господи, высок над всею землею, превознесен над всеми богами.
PS|96|10|Любящие Господа, ненавидьте зло! Он хранит души святых Своих; из руки нечестивых избавляет их.
PS|96|11|Свет сияет на праведника, и на правых сердцем – веселие.
PS|96|12|Радуйтесь, праведные, о Господе и славьте память святыни Его.
PS|97|1|Псалом Воспойте Господу новую песнь, ибо Он сотворил чудеса. Его десница и святая мышца Его доставили Ему победу.
PS|97|2|Явил Господь спасение Свое, открыл пред очами народов правду Свою.
PS|97|3|Вспомнил Он милость Свою и верность Свою к дому Израилеву. Все концы земли увидели спасение Бога нашего.
PS|97|4|Восклицайте Господу, вся земля; торжествуйте, веселитесь и пойте;
PS|97|5|пойте Господу с гуслями, с гуслями и с гласом псалмопения;
PS|97|6|при звуке труб и рога торжествуйте пред Царем Господом.
PS|97|7|Да шумит море и что наполняет его, вселенная и живущие в ней;
PS|97|8|да рукоплещут реки, да ликуют вместе горы
PS|97|9|пред лицем Господа, ибо Он идет судить землю. Он будет судить вселенную праведно и народы – верно.
PS|98|1|Господь царствует: да трепещут народы! Он восседает на Херувимах: да трясется земля!
PS|98|2|Господь на Сионе велик, и высок Он над всеми народами.
PS|98|3|Да славят великое и страшное имя Твое: свято оно!
PS|98|4|И могущество царя любит суд. Ты утвердил справедливость; суд и правду Ты совершил в Иакове.
PS|98|5|Превозносите Господа, Бога нашего, и поклоняйтесь подножию Его: свято оно!
PS|98|6|Моисей и Аарон между священниками и Самуил между призывающими имя Его взывали к Господу, и Он внимал им.
PS|98|7|В столпе облачном говорил Он к ним; они хранили Его заповеди и устав, который Он дал им.
PS|98|8|Господи, Боже наш! Ты внимал им; Ты был для них Богом прощающим и наказывающим за дела их.
PS|98|9|Превозносите Господа, Бога нашего, и поклоняйтесь на святой горе Его, ибо свят Господь, Бог наш.
PS|99|1|Псалом хвалебный. Воскликните Господу, вся земля!
PS|99|2|Служите Господу с веселием; идите пред лице Его с восклицанием!
PS|99|3|Познайте, что Господь есть Бог, что Он сотворил нас, и мы – Его, Его народ и овцы паствы Его.
PS|99|4|Входите во врата Его со славословием, во дворы Его – с хвалою. Славьте Его, благословляйте имя Его,
PS|99|5|ибо благ Господь: милость Его вовек, и истина Его в род и род.
PS|100|1|Псалом Давида. Милость и суд буду петь; Тебе, Господи, буду петь.
PS|100|2|Буду размышлять о пути непорочном: "когда ты придешь ко мне?" Буду ходить в непорочности моего сердца посреди дома моего.
PS|100|3|Не положу пред очами моими вещи непотребной; дело преступное я ненавижу: не прилепится оно ко мне.
PS|100|4|Сердце развращенное будет удалено от меня; злого я не буду знать.
PS|100|5|Тайно клевещущего на ближнего своего изгоню; гордого очами и надменного сердцем не потерплю.
PS|100|6|Глаза мои на верных земли, чтобы они пребывали при мне; кто ходит путем непорочности, тот будет служить мне.
PS|100|7|Не будет жить в доме моем поступающий коварно; говорящий ложь не останется пред глазами моими.
PS|100|8|С раннего утра буду истреблять всех нечестивцев земли, дабы искоренить из града Господня всех делающих беззаконие.
PS|101|1|Молитва страждущего, когда он унывает и изливает пред Господом печаль свою.
PS|101|2|Господи! услышь молитву мою, и вопль мой да придет к Тебе.
PS|101|3|Не скрывай лица Твоего от меня; в день скорби моей приклони ко мне ухо Твое; в день, [когда воззову к Тебе], скоро услышь меня;
PS|101|4|ибо исчезли, как дым, дни мои, и кости мои обожжены, как головня;
PS|101|5|сердце мое поражено, и иссохло, как трава, так что я забываю есть хлеб мой;
PS|101|6|от голоса стенания моего кости мои прильпнули к плоти моей.
PS|101|7|Я уподобился пеликану в пустыне; я стал как филин на развалинах;
PS|101|8|не сплю и сижу, как одинокая птица на кровле.
PS|101|9|Всякий день поносят меня враги мои, и злобствующие на меня клянут мною.
PS|101|10|Я ем пепел, как хлеб, и питье мое растворяю слезами,
PS|101|11|от гнева Твоего и негодования Твоего, ибо Ты вознес меня и низверг меня.
PS|101|12|Дни мои – как уклоняющаяся тень, и я иссох, как трава.
PS|101|13|Ты же, Господи, вовек пребываешь, и память о Тебе в род и род.
PS|101|14|Ты восстанешь, умилосердишься над Сионом, ибо время помиловать его, – ибо пришло время;
PS|101|15|ибо рабы Твои возлюбили и камни его, и о прахе его жалеют.
PS|101|16|И убоятся народы имени Господня, и все цари земные – славы Твоей.
PS|101|17|Ибо созиждет Господь Сион и явится во славе Своей;
PS|101|18|призрит на молитву беспомощных и не презрит моления их.
PS|101|19|Напишется о сем для рода последующего, и поколение грядущее восхвалит Господа,
PS|101|20|ибо Он приникнул со святой высоты Своей, с небес призрел Господь на землю,
PS|101|21|чтобы услышать стон узников, разрешить сынов смерти,
PS|101|22|дабы возвещали на Сионе имя Господне и хвалу Его – в Иерусалиме,
PS|101|23|когда соберутся народы вместе и царства для служения Господу.
PS|101|24|Изнурил Он на пути силы мои, сократил дни мои.
PS|101|25|Я сказал: Боже мой! не восхити меня в половине дней моих. Твои лета в роды родов.
PS|101|26|В начале Ты, основал землю, и небеса – дело Твоих рук;
PS|101|27|они погибнут, а Ты пребудешь; и все они, как риза, обветшают, и, как одежду, Ты переменишь их, и изменятся;
PS|101|28|но Ты – тот же, и лета Твои не кончатся.
PS|101|29|Сыны рабов Твоих будут жить, и семя их утвердится пред лицем Твоим.
PS|102|1|Псалом Давида. Благослови, душа моя, Господа, и вся внутренность моя – святое имя Его.
PS|102|2|Благослови, душа моя, Господа и не забывай всех благодеяний Его.
PS|102|3|Он прощает все беззакония твои, исцеляет все недуги твои;
PS|102|4|избавляет от могилы жизнь твою, венчает тебя милостью и щедротами;
PS|102|5|насыщает благами желание твое: обновляется, подобно орлу, юность твоя.
PS|102|6|Господь творит правду и суд всем обиженным.
PS|102|7|Он показал пути Свои Моисею, сынам Израилевым – дела Свои.
PS|102|8|Щедр и милостив Господь, долготерпелив и многомилостив:
PS|102|9|не до конца гневается, и не вовек негодует.
PS|102|10|Не по беззакониям нашим сотворил нам, и не по грехам нашим воздал нам:
PS|102|11|ибо как высоко небо над землею, так велика милость [Господа] к боящимся Его;
PS|102|12|как далеко восток от запада, так удалил Он от нас беззакония наши;
PS|102|13|как отец милует сынов, так милует Господь боящихся Его.
PS|102|14|Ибо Он знает состав наш, помнит, что мы – персть.
PS|102|15|Дни человека – как трава; как цвет полевой, так он цветет.
PS|102|16|Пройдет над ним ветер, и нет его, и место его уже не узнает его.
PS|102|17|Милость же Господня от века и до века к боящимся Его,
PS|102|18|и правда Его на сынах сынов, хранящих завет Его и помнящих заповеди Его, чтобы исполнять их.
PS|102|19|Господь на небесах поставил престол Свой, и царство Его всем обладает.
PS|102|20|Благословите Господа, [все] Ангелы Его, крепкие силою, исполняющие слово Его, повинуясь гласу слова Его;
PS|102|21|благословите Господа, все воинства Его, служители Его, исполняющие волю Его;
PS|102|22|благословите Господа, все дела Его, во всех местах владычества Его. Благослови, душа моя, Господа!
PS|103|1|Благослови, душа моя, Господа! Господи, Боже мой! Ты дивно велик, Ты облечен славою и величием;
PS|103|2|Ты одеваешься светом, как ризою, простираешь небеса, как шатер;
PS|103|3|устрояешь над водами горние чертоги Твои, делаешь облака Твоею колесницею, шествуешь на крыльях ветра.
PS|103|4|Ты творишь ангелами Твоими духов, служителями Твоими – огонь пылающий.
PS|103|5|Ты поставил землю на твердых основах: не поколеблется она во веки и веки.
PS|103|6|Бездною, как одеянием, покрыл Ты ее, на горах стоят воды.
PS|103|7|От прещения Твоего бегут они, от гласа грома Твоего быстро уходят;
PS|103|8|восходят на горы, нисходят в долины, на место, которое Ты назначил для них.
PS|103|9|Ты положил предел, которого не перейдут, и не возвратятся покрыть землю.
PS|103|10|Ты послал источники в долины: между горами текут,
PS|103|11|поят всех полевых зверей; дикие ослы утоляют жажду свою.
PS|103|12|При них обитают птицы небесные, из среды ветвей издают голос.
PS|103|13|Ты напояешь горы с высот Твоих, плодами дел Твоих насыщается земля.
PS|103|14|Ты произращаешь траву для скота, и зелень на пользу человека, чтобы произвести из земли пищу,
PS|103|15|и вино, которое веселит сердце человека, и елей, от которого блистает лице его, и хлеб, который укрепляет сердце человека.
PS|103|16|Насыщаются древа Господа, кедры Ливанские, которые Он насадил;
PS|103|17|на них гнездятся птицы: ели – жилище аисту,
PS|103|18|высокие горы – сернам; каменные утесы – убежище зайцам.
PS|103|19|Он сотворил луну для [указания] времен, солнце знает свой запад.
PS|103|20|Ты простираешь тьму и бывает ночь: во время нее бродят все лесные звери;
PS|103|21|львы рыкают о добыче и просят у Бога пищу себе.
PS|103|22|Восходит солнце, [и] они собираются и ложатся в свои логовища;
PS|103|23|выходит человек на дело свое и на работу свою до вечера.
PS|103|24|Как многочисленны дела Твои, Господи! Все соделал Ты премудро; земля полна произведений Твоих.
PS|103|25|Это – море великое и пространное: там пресмыкающиеся, которым нет числа, животные малые с большими;
PS|103|26|там плавают корабли, там этот левиафан, которого Ты сотворил играть в нем.
PS|103|27|Все они от Тебя ожидают, чтобы Ты дал им пищу их в свое время.
PS|103|28|Даешь им – принимают, отверзаешь руку Твою – насыщаются благом;
PS|103|29|скроешь лице Твое – мятутся, отнимешь дух их – умирают и в персть свою возвращаются;
PS|103|30|пошлешь дух Твой – созидаются, и Ты обновляешь лице земли.
PS|103|31|Да будет Господу слава во веки; да веселится Господь о делах Своих!
PS|103|32|Призирает на землю, и она трясется; прикасается к горам, и дымятся.
PS|103|33|Буду петь Господу во [всю] жизнь мою, буду петь Богу моему, доколе есмь.
PS|103|34|Да будет благоприятна Ему песнь моя; буду веселиться о Господе.
PS|103|35|Да исчезнут грешники с земли, и беззаконных да не будет более. Благослови, душа моя, Господа! Аллилуия!
PS|104|1|Славьте Господа; призывайте имя Его; возвещайте в народах дела Его;
PS|104|2|воспойте Ему и пойте Ему; поведайте о всех чудесах Его.
PS|104|3|Хвалитесь именем Его святым; да веселится сердце ищущих Господа.
PS|104|4|Ищите Господа и силы Его, ищите лица Его всегда.
PS|104|5|Воспоминайте чудеса Его, которые сотворил, знамения Его и суды уст Его,
PS|104|6|вы, семя Авраамово, рабы Его, сыны Иакова, избранные Его.
PS|104|7|Он Господь Бог наш: по всей земле суды Его.
PS|104|8|Вечно помнит завет Свой, слово, [которое] заповедал в тысячу родов,
PS|104|9|которое завещал Аврааму, и клятву Свою Исааку,
PS|104|10|и поставил то Иакову в закон и Израилю в завет вечный,
PS|104|11|говоря: "тебе дам землю Ханаанскую в удел наследия вашего".
PS|104|12|Когда их было еще мало числом, очень мало, и они были пришельцами в ней
PS|104|13|и переходили от народа к народу, из царства к иному племени,
PS|104|14|никому не позволял обижать их и возбранял о них царям:
PS|104|15|"не прикасайтесь к помазанным Моим, и пророкам Моим не делайте зла".
PS|104|16|И призвал голод на землю; всякий стебель хлебный истребил.
PS|104|17|Послал пред ними человека: в рабы продан был Иосиф.
PS|104|18|Стеснили оковами ноги его; в железо вошла душа его,
PS|104|19|доколе исполнилось слово Его: слово Господне испытало его.
PS|104|20|Послал царь, и разрешил его владетель народов и освободил его;
PS|104|21|поставил его господином над домом своим и правителем над всем владением своим,
PS|104|22|чтобы он наставлял вельмож его по своей душе и старейшин его учил мудрости.
PS|104|23|Тогда пришел Израиль в Египет, и переселился Иаков в землю Хамову.
PS|104|24|И весьма размножил [Бог] народ Свой и сделал его сильнее врагов его.
PS|104|25|Возбудил в сердце их ненависть против народа Его и ухищрение против рабов Его.
PS|104|26|Послал Моисея, раба Своего, Аарона, которого избрал.
PS|104|27|Они показали между ними слова знамений Его и чудеса [Его] в земле Хамовой.
PS|104|28|Послал тьму и сделал мрак, и не воспротивились слову Его.
PS|104|29|Преложил воду их в кровь, и уморил рыбу их.
PS|104|30|Земля их произвела множество жаб [даже] в спальне царей их.
PS|104|31|Он сказал, и пришли разные насекомые, скнипы во все пределы их.
PS|104|32|Вместо дождя послал на них град, палящий огонь на землю их,
PS|104|33|и побил виноград их и смоковницы их, и сокрушил дерева в пределах их.
PS|104|34|Сказал, и пришла саранча и гусеницы без числа;
PS|104|35|и съели всю траву на земле их, и съели плоды на полях их.
PS|104|36|И поразил всякого первенца в земле их, начатки всей силы их.
PS|104|37|И вывел [Израильтян] с серебром и золотом, и не было в коленах их болящего.
PS|104|38|Обрадовался Египет исшествию их; ибо страх от них напал на него.
PS|104|39|Простер облако в покров [им] и огонь, чтобы светить [им] ночью.
PS|104|40|Просили, и Он послал перепелов, и хлебом небесным насыщал их.
PS|104|41|Разверз камень, и потекли воды, потекли рекою по местам сухим,
PS|104|42|ибо вспомнил Он святое слово Свое к Аврааму, рабу Своему,
PS|104|43|и вывел народ Свой в радости, избранных Своих в веселии,
PS|104|44|и дал им земли народов, и они наследовали труд иноплеменных,
PS|104|45|чтобы соблюдали уставы Его и хранили законы Его. Аллилуия!
PS|105|1|Аллилуия. Славьте Господа, ибо Он благ, ибо вовек милость Его.
PS|105|2|Кто изречет могущество Господа, возвестит все хвалы Его?
PS|105|3|Блаженны хранящие суд и творящие правду во всякое время!
PS|105|4|Вспомни о мне, Господи, в благоволении к народу Твоему; посети меня спасением Твоим,
PS|105|5|дабы мне видеть благоденствие избранных Твоих, веселиться веселием народа Твоего, хвалиться с наследием Твоим.
PS|105|6|Согрешили мы с отцами нашими, совершили беззаконие, соделали неправду.
PS|105|7|Отцы наши в Египте не уразумели чудес Твоих, не помнили множества милостей Твоих, и возмутились у моря, у Чермного моря.
PS|105|8|Но Он спас их ради имени Своего, дабы показать могущество Свое.
PS|105|9|Грозно рек морю Чермному, и оно иссохло; и провел их по безднам, как по суше;
PS|105|10|и спас их от руки ненавидящего и избавил их от руки врага.
PS|105|11|Воды покрыли врагов их, ни одного из них не осталось.
PS|105|12|И поверили они словам Его, [и] воспели хвалу Ему.
PS|105|13|[Но] скоро забыли дела Его, не дождались Его изволения;
PS|105|14|увлеклись похотением в пустыне, и искусили Бога в необитаемой.
PS|105|15|И Он исполнил прошение их, [но] послал язву на души их.
PS|105|16|И позавидовали в стане Моисею [и] Аарону, святому Господню.
PS|105|17|Разверзлась земля, и поглотила Дафана и покрыла скопище Авирона.
PS|105|18|И возгорелся огонь в скопище их, пламень попалил нечестивых.
PS|105|19|Сделали тельца у Хорива и поклонились истукану;
PS|105|20|и променяли славу свою на изображение вола, ядущего траву.
PS|105|21|Забыли Бога, Спасителя своего, совершившего великое в Египте,
PS|105|22|дивное в земле Хамовой, страшное у Чермного моря.
PS|105|23|И хотел истребить их, если бы Моисей, избранный Его, не стал пред Ним в расселине, чтобы отвратить ярость Его, да не погубит [их].
PS|105|24|И презрели они землю желанную, не верили слову Его;
PS|105|25|и роптали в шатрах своих, не слушались гласа Господня.
PS|105|26|И поднял Он руку Свою на них, чтобы низложить их в пустыне,
PS|105|27|низложить племя их в народах и рассеять их по землям.
PS|105|28|Они прилепились к Ваалфегору и ели жертвы бездушным,
PS|105|29|и раздражали [Бога] делами своими, и вторглась к ним язва.
PS|105|30|И восстал Финеес и произвел суд, – и остановилась язва.
PS|105|31|И [это] вменено ему в праведность в роды и роды во веки.
PS|105|32|И прогневали [Бога] у вод Меривы, и Моисей потерпел за них,
PS|105|33|ибо они огорчили дух его, и он погрешил устами своими.
PS|105|34|Не истребили народов, о которых сказал им Господь,
PS|105|35|но смешались с язычниками и научились делам их;
PS|105|36|служили истуканам их, [которые] были для них сетью,
PS|105|37|и приносили сыновей своих и дочерей своих в жертву бесам;
PS|105|38|проливали кровь невинную, кровь сыновей своих и дочерей своих, которых приносили в жертву идолам Ханаанским, – и осквернилась земля кровью;
PS|105|39|оскверняли себя делами своими, блудодействовали поступками своими.
PS|105|40|И воспылал гнев Господа на народ Его, и возгнушался Он наследием Своим
PS|105|41|и предал их в руки язычников, и ненавидящие их стали обладать ими.
PS|105|42|Враги их утесняли их, и они смирялись под рукою их.
PS|105|43|Много раз Он избавлял их; они же раздражали [Его] упорством своим, и были уничижаемы за беззаконие свое.
PS|105|44|Но Он призирал на скорбь их, когда слышал вопль их,
PS|105|45|и вспоминал завет Свой с ними и раскаивался по множеству милости Своей;
PS|105|46|и возбуждал к ним сострадание во всех, пленявших их.
PS|105|47|Спаси нас, Господи, Боже наш, и собери нас от народов, дабы славить святое имя Твое, хвалиться Твоею славою.
PS|105|48|Благословен Господь, Бог Израилев, от века и до века! И да скажет весь народ: аминь! Аллилуия!
PS|106|1|Славьте Господа, ибо Он благ, ибо вовек милость Его!
PS|106|2|Так да скажут избавленные Господом, которых избавил Он от руки врага,
PS|106|3|и собрал от стран, от востока и запада, от севера и моря.
PS|106|4|Они блуждали в пустыне по безлюдному пути и не находили населенного города;
PS|106|5|терпели голод и жажду, душа их истаевала в них.
PS|106|6|Но воззвали к Господу в скорби своей, и Он избавил их от бедствий их,
PS|106|7|и повел их прямым путем, чтобы они шли к населенному городу.
PS|106|8|Да славят Господа за милость Его и за чудные дела Его для сынов человеческих:
PS|106|9|ибо Он насытил душу жаждущую и душу алчущую исполнил благами.
PS|106|10|Они сидели во тьме и тени смертной, окованные скорбью и железом;
PS|106|11|ибо не покорялись словам Божиим и небрегли о воле Всевышнего.
PS|106|12|Он смирил сердце их работами; они преткнулись, и не было помогающего.
PS|106|13|Но воззвали к Господу в скорби своей, и Он спас их от бедствий их;
PS|106|14|вывел их из тьмы и тени смертной, и расторгнул узы их.
PS|106|15|Да славят Господа за милость Его и за чудные дела Его для сынов человеческих:
PS|106|16|ибо Он сокрушил врата медные и вереи железные сломил.
PS|106|17|Безрассудные страдали за беззаконные пути свои и за неправды свои;
PS|106|18|от всякой пищи отвращалась душа их, и они приближались ко вратам смерти.
PS|106|19|Но воззвали к Господу в скорби своей, и Он спас их от бедствий их;
PS|106|20|послал слово Свое и исцелил их, и избавил их от могил их.
PS|106|21|Да славят Господа за милость Его и за чудные дела Его для сынов человеческих!
PS|106|22|Да приносят Ему жертву хвалы и да возвещают о делах Его с пением!
PS|106|23|Отправляющиеся на кораблях в море, производящие дела на больших водах,
PS|106|24|видят дела Господа и чудеса Его в пучине:
PS|106|25|Он речет, – и восстанет бурный ветер и высоко поднимает волны его:
PS|106|26|восходят до небес, нисходят до бездны; душа их истаевает в бедствии;
PS|106|27|они кружатся и шатаются, как пьяные, и вся мудрость их исчезает.
PS|106|28|Но воззвали к Господу в скорби своей, и Он вывел их из бедствия их.
PS|106|29|Он превращает бурю в тишину, и волны умолкают.
PS|106|30|И веселятся, что они утихли, и Он приводит их к желаемой пристани.
PS|106|31|Да славят Господа за милость Его и за чудные дела Его для сынов человеческих!
PS|106|32|Да превозносят Его в собрании народном и да славят Его в сонме старейшин!
PS|106|33|Он превращает реки в пустыню и источники вод – в сушу,
PS|106|34|землю плодородную – в солончатую, за нечестие живущих на ней.
PS|106|35|Он превращает пустыню в озеро, и землю иссохшую – в источники вод;
PS|106|36|и поселяет там алчущих, и они строят город для обитания;
PS|106|37|засевают поля, насаждают виноградники, которые приносят им обильные плоды.
PS|106|38|Он благословляет их, и они весьма размножаются, и скота их не умаляет.
PS|106|39|Уменьшились они и упали от угнетения, бедствия и скорби, –
PS|106|40|он изливает бесчестие на князей и оставляет их блуждать в пустыне, где нет путей.
PS|106|41|Бедного же извлекает из бедствия и умножает род его, как стада овец.
PS|106|42|Праведники видят сие и радуются, а всякое нечестие заграждает уста свои.
PS|106|43|Кто мудр, тот заметит сие и уразумеет милость Господа.
PS|107|1|Песнь. Псалом Давида.
PS|107|2|Готово сердце мое, Боже; буду петь и воспевать во славе моей.
PS|107|3|Воспрянь, псалтирь и гусли! Я встану рано.
PS|107|4|Буду славить Тебя, Господи, между народами; буду воспевать Тебя среди племен,
PS|107|5|ибо превыше небес милость Твоя и до облаков истина Твоя.
PS|107|6|Будь превознесен выше небес, Боже; над всею землею [да] [будет] слава Твоя,
PS|107|7|дабы избавились возлюбленные Твои: спаси десницею Твоею и услышь меня.
PS|107|8|Бог сказал во святилище Своем: "восторжествую, разделю Сихем и долину Сокхоф размерю;
PS|107|9|Мой Галаад, Мой Манассия, Ефрем – крепость главы Моей, Иуда – скипетр Мой,
PS|107|10|Моав – умывальная чаша Моя, на Едома простру сапог Мой, над землею Филистимскою восклицать буду".
PS|107|11|Кто введет меня в укрепленный город? Кто доведет меня до Едома?
PS|107|12|Не Ты ли, Боже, [Который] отринул нас и не выходишь, Боже, с войсками нашими?
PS|107|13|Подай нам помощь в тесноте, ибо защита человеческая суетна.
PS|107|14|С Богом мы окажем силу: Он низложит врагов наших.
PS|108|1|Начальнику хора. Псалом Давида. Боже хвалы моей! не премолчи,
PS|108|2|ибо отверзлись на меня уста нечестивые и уста коварные; говорят со мною языком лживым;
PS|108|3|отвсюду окружают меня словами ненависти, вооружаются против меня без причины;
PS|108|4|за любовь мою они враждуют на меня, а я молюсь;
PS|108|5|воздают мне за добро злом, за любовь мою – ненавистью.
PS|108|6|Поставь над ним нечестивого, и диавол да станет одесную его.
PS|108|7|Когда будет судиться, да выйдет виновным, и молитва его да будет в грех;
PS|108|8|да будут дни его кратки, и достоинство его да возьмет другой;
PS|108|9|дети его да будут сиротами, и жена его – вдовою;
PS|108|10|да скитаются дети его и нищенствуют, и просят [хлеба] из развалин своих;
PS|108|11|да захватит заимодавец все, что есть у него, и чужие да расхитят труд его;
PS|108|12|да не будет сострадающего ему, да не будет милующего сирот его;
PS|108|13|да будет потомство его на погибель, и да изгладится имя их в следующем роде;
PS|108|14|да будет воспомянуто пред Господом беззаконие отцов его, и грех матери его да не изгладится;
PS|108|15|да будут они всегда в очах Господа, и да истребит Он память их на земле,
PS|108|16|за то, что он не думал оказывать милость, но преследовал человека бедного и нищего и сокрушенного сердцем, чтобы умертвить его;
PS|108|17|возлюбил проклятие, – оно и придет на него; не восхотел благословения, – оно и удалится от него;
PS|108|18|да облечется проклятием, как ризою, и да войдет оно, как вода, во внутренность его и, как елей, в кости его;
PS|108|19|да будет оно ему, как одежда, в которую он одевается, и как пояс, которым всегда опоясывается.
PS|108|20|Таково воздаяние от Господа врагам моим и говорящим злое на душу мою!
PS|108|21|Со мною же, Господи, Господи, твори ради имени Твоего, ибо блага милость Твоя; спаси меня,
PS|108|22|ибо я беден и нищ, и сердце мое уязвлено во мне.
PS|108|23|Я исчезаю, как уклоняющаяся тень; гонят меня, как саранчу.
PS|108|24|Колени мои изнемогли от поста, и тело мое лишилось тука.
PS|108|25|Я стал для них посмешищем: увидев меня, кивают головами.
PS|108|26|Помоги мне, Господи, Боже мой, спаси меня по милости Твоей,
PS|108|27|да познают, что это – Твоя рука, и что Ты, Господи, соделал это.
PS|108|28|Они проклинают, а Ты благослови; они восстают, но да будут постыжены; раб же Твой да возрадуется.
PS|108|29|Да облекутся противники мои бесчестьем и, как одеждою, покроются стыдом своим.
PS|108|30|И я громко буду устами моими славить Господа и среди множества прославлять Его,
PS|108|31|ибо Он стоит одесную бедного, чтобы спасти его от судящих душу его.
PS|109|1|Псалом Давида. Сказал Господь Господу моему: седи одесную Меня, доколе положу врагов Твоих в подножие ног Твоих.
PS|109|2|Жезл силы Твоей пошлет Господь с Сиона: господствуй среди врагов Твоих.
PS|109|3|В день силы Твоей народ Твой готов во благолепии святыни; из чрева прежде денницы подобно росе рождение Твое.
PS|109|4|Клялся Господь и не раскается: Ты священник вовек по чину Мелхиседека.
PS|109|5|Господь одесную Тебя. Он в день гнева Своего поразит царей;
PS|109|6|совершит суд над народами, наполнит [землю] трупами, сокрушит голову в земле обширной.
PS|109|7|Из потока на пути будет пить, и потому вознесет главу.
PS|110|1|Аллилуия. Славлю [Тебя], Господи, всем сердцем [моим] в совете праведных и в собрании.
PS|110|2|Велики дела Господни, вожделенны для всех, любящих оные.
PS|110|3|Дело Его – слава и красота, и правда Его пребывает вовек.
PS|110|4|Памятными соделал Он чудеса Свои; милостив и щедр Господь.
PS|110|5|Пищу дает боящимся Его; вечно помнит завет Свой.
PS|110|6|Силу дел Своих явил Он народу Своему, чтобы дать ему наследие язычников.
PS|110|7|Дела рук Его – истина и суд; все заповеди Его верны,
PS|110|8|тверды на веки и веки, основаны на истине и правоте.
PS|110|9|Избавление послал Он народу Своему; заповедал на веки завет Свой. Свято и страшно имя Его!
PS|110|10|Начало мудрости – страх Господень; разум верный у всех, исполняющих [заповеди Его]. Хвала Ему пребудет вовек.
PS|111|1|Аллилуия. Блажен муж, боящийся Господа и крепко любящий заповеди Его.
PS|111|2|Сильно будет на земле семя его; род правых благословится.
PS|111|3|Обилие и богатство в доме его, и правда его пребывает вовек.
PS|111|4|Во тьме восходит свет правым; благ он и милосерд и праведен.
PS|111|5|Добрый человек милует и взаймы дает; он даст твердость словам своим на суде.
PS|111|6|Он вовек не поколеблется; в вечной памяти будет праведник.
PS|111|7|Не убоится худой молвы: сердце его твердо, уповая на Господа.
PS|111|8|Утверждено сердце его: он не убоится, когда посмотрит на врагов своих.
PS|111|9|Он расточил, роздал нищим; правда его пребывает во веки; рог его вознесется во славе.
PS|111|10|Нечестивый увидит [это] и будет досадовать, заскрежещет зубами своими и истает. Желание нечестивых погибнет.
PS|112|1|Аллилуия Хвалите, рабы Господни, хвалите имя Господне.
PS|112|2|Да будет имя Господне благословенно отныне и вовек.
PS|112|3|От восхода солнца до запада [да будет] прославляемо имя Господне.
PS|112|4|Высок над всеми народами Господь; над небесами слава Его.
PS|112|5|Кто, как Господь, Бог наш, Который, обитая на высоте,
PS|112|6|приклоняется, чтобы призирать на небо и на землю;
PS|112|7|из праха поднимает бедного, из брения возвышает нищего,
PS|112|8|чтобы посадить его с князьями, с князьями народа его;
PS|112|9|неплодную вселяет в дом матерью, радующеюся о детях? Аллилуия!
PS|113|1|Когда вышел Израиль из Египта, дом Иакова – из народа иноплеменного,
PS|113|2|Иуда сделался святынею Его, Израиль – владением Его.
PS|113|3|Море увидело и побежало; Иордан обратился назад.
PS|113|4|Горы прыгали, как овны, и холмы, как агнцы.
PS|113|5|Что с тобою, море, что ты побежало, и [с тобою], Иордан, что ты обратился назад?
PS|113|6|Что вы прыгаете, горы, как овны, и вы, холмы, как агнцы?
PS|113|7|Пред лицем Господа трепещи, земля, пред лицем Бога Иаковлева,
PS|113|8|превращающего скалу в озеро воды и камень в источник вод.
PS|113|9|Не нам, Господи, не нам, но имени Твоему дай славу, ради милости Твоей, ради истины Твоей.
PS|113|10|Для чего язычникам говорить: "где же Бог их"?
PS|113|11|Бог наш на небесах; творит все, что хочет.
PS|113|12|А их идолы – серебро и золото, дело рук человеческих.
PS|113|13|Есть у них уста, но не говорят; есть у них глаза, но не видят;
PS|113|14|есть у них уши, но не слышат; есть у них ноздри, но не обоняют;
PS|113|15|есть у них руки, но не осязают; есть у них ноги, но не ходят; и они не издают голоса гортанью своею.
PS|113|16|Подобны им да будут делающие их и все, надеющиеся на них.
PS|113|17|[Дом] Израилев! уповай на Господа: Он наша помощь и щит.
PS|113|18|Дом Ааронов! уповай на Господа: Он наша помощь и щит.
PS|113|19|Боящиеся Господа! уповайте на Господа: Он наша помощь и щит.
PS|113|20|Господь помнит нас, благословляет [нас], благословляет дом Израилев, благословляет дом Ааронов;
PS|113|21|благословляет боящихся Господа, малых с великими.
PS|113|22|Да приложит вам Господь более и более, вам и детям вашим.
PS|113|23|Благословенны вы Господом, сотворившим небо и землю.
PS|113|24|Небо – небо Господу, а землю Он дал сынам человеческим.
PS|113|25|Ни мертвые восхвалят Господа, ни все нисходящие в могилу;
PS|113|26|но мы будем благословлять Господа отныне и вовек. Аллилуия.
PS|114|1|Я радуюсь, что Господь услышал голос мой, моление мое;
PS|114|2|приклонил ко мне ухо Свое, и потому буду призывать Его во [все] дни мои.
PS|114|3|Объяли меня болезни смертные, муки адские постигли меня; я встретил тесноту и скорбь.
PS|114|4|Тогда призвал я имя Господне: Господи! избавь душу мою.
PS|114|5|Милостив Господь и праведен, и милосерд Бог наш.
PS|114|6|Хранит Господь простодушных: я изнемог, и Он помог мне.
PS|114|7|Возвратись, душа моя, в покой твой, ибо Господь облагодетельствовал тебя.
PS|114|8|Ты избавил душу мою от смерти, очи мои от слез и ноги мои от преткновения.
PS|114|9|Буду ходить пред лицем Господним на земле живых.
PS|115|1|Я веровал, и потому говорил: я сильно сокрушен.
PS|115|2|Я сказал в опрометчивости моей: всякий человек ложь.
PS|115|3|Что воздам Господу за все благодеяния Его ко мне?
PS|115|4|Чашу спасения прииму и имя Господне призову.
PS|115|5|Обеты мои воздам Господу пред всем народом Его.
PS|115|6|Дорога в очах Господних смерть святых Его!
PS|115|7|О, Господи! я раб Твой, я раб Твой и сын рабы Твоей; Ты разрешил узы мои.
PS|115|8|Тебе принесу жертву хвалы, и имя Господне призову.
PS|115|9|Обеты мои воздам Господу пред всем народом Его,
PS|115|10|во дворах дома Господня, посреди тебя, Иерусалим! Аллилуия.
PS|116|1|Хвалите Господа, все народы, прославляйте Его, все племена;
PS|116|2|ибо велика милость Его к нам, и истина Господня вовек. Аллилуия.
PS|117|1|Славьте Господа, ибо Он благ, ибо вовек милость Его.
PS|117|2|Да скажет ныне [дом] Израилев: ибо вовек милость Его.
PS|117|3|Да скажет ныне дом Ааронов: ибо вовек милость Его.
PS|117|4|Да скажут ныне боящиеся Господа: ибо вовек милость Его.
PS|117|5|Из тесноты воззвал я к Господу, – и услышал меня, и на пространное место [вывел меня] Господь.
PS|117|6|Господь за меня – не устрашусь: что сделает мне человек?
PS|117|7|Господь мне помощник: буду смотреть на врагов моих.
PS|117|8|Лучше уповать на Господа, нежели надеяться на человека.
PS|117|9|Лучше уповать на Господа, нежели надеяться на князей.
PS|117|10|Все народы окружили меня, но именем Господним я низложил их;
PS|117|11|обступили меня, окружили меня, но именем Господним я низложил их;
PS|117|12|окружили меня, как пчелы, и угасли, как огонь в терне: именем Господним я низложил их.
PS|117|13|Сильно толкнули меня, чтобы я упал, но Господь поддержал меня.
PS|117|14|Господь – сила моя и песнь; Он соделался моим спасением.
PS|117|15|Глас радости и спасения в жилищах праведников: десница Господня творит силу!
PS|117|16|Десница Господня высока, десница Господня творит силу!
PS|117|17|Не умру, но буду жить и возвещать дела Господни.
PS|117|18|Строго наказал меня Господь, но смерти не предал меня.
PS|117|19|Отворите мне врата правды; войду в них, прославлю Господа.
PS|117|20|Вот врата Господа; праведные войдут в них.
PS|117|21|Славлю Тебя, что Ты услышал меня и соделался моим спасением.
PS|117|22|Камень, который отвергли строители, соделался главою угла:
PS|117|23|это – от Господа, и есть дивно в очах наших.
PS|117|24|Сей день сотворил Господь: возрадуемся и возвеселимся в оный!
PS|117|25|О, Господи, спаси же! О, Господи, споспешествуй же!
PS|117|26|Благословен грядущий во имя Господне! Благословляем вас из дома Господня.
PS|117|27|Бог – Господь, и осиял нас; вяжите вервями жертву, [ведите] к рогам жертвенника.
PS|117|28|Ты Бог мой: буду славить Тебя; Ты Бог мой: буду превозносить Тебя.
PS|117|29|Славьте Господа, ибо Он благ, ибо вовек милость Его.
PS|118|1|Блаженны непорочные в пути, ходящие в законе Господнем.
PS|118|2|Блаженны хранящие откровения Его, всем сердцем ищущие Его.
PS|118|3|Они не делают беззакония, ходят путями Его.
PS|118|4|Ты заповедал повеления Твои хранить твердо.
PS|118|5|О, если бы направлялись пути мои к соблюдению уставов Твоих!
PS|118|6|Тогда я не постыдился бы, взирая на все заповеди Твои:
PS|118|7|я славил бы Тебя в правоте сердца, поучаясь судам правды Твоей.
PS|118|8|Буду хранить уставы Твои; не оставляй меня совсем.
PS|118|9|Как юноше содержать в чистоте путь свой? – Хранением себя по слову Твоему.
PS|118|10|Всем сердцем моим ищу Тебя; не дай мне уклониться от заповедей Твоих.
PS|118|11|В сердце моем сокрыл я слово Твое, чтобы не грешить пред Тобою.
PS|118|12|Благословен Ты, Господи! научи меня уставам Твоим.
PS|118|13|Устами моими возвещал я все суды уст Твоих.
PS|118|14|На пути откровений Твоих я радуюсь, как во всяком богатстве.
PS|118|15|О заповедях Твоих размышляю, и взираю на пути Твои.
PS|118|16|Уставами Твоими утешаюсь, не забываю слова Твоего.
PS|118|17|Яви милость рабу Твоему, и буду жить и хранить слово Твое.
PS|118|18|Открой очи мои, и увижу чудеса закона Твоего.
PS|118|19|Странник я на земле; не скрывай от меня заповедей Твоих.
PS|118|20|Истомилась душа моя желанием судов Твоих во всякое время.
PS|118|21|Ты укротил гордых, проклятых, уклоняющихся от заповедей Твоих.
PS|118|22|Сними с меня поношение и посрамление, ибо я храню откровения Твои.
PS|118|23|Князья сидят и сговариваются против меня, а раб Твой размышляет об уставах Твоих.
PS|118|24|Откровения Твои – утешение мое, – советники мои.
PS|118|25|Душа моя повержена в прах; оживи меня по слову Твоему.
PS|118|26|Объявил я пути мои, и Ты услышал меня; научи меня уставам Твоим.
PS|118|27|Дай мне уразуметь путь повелений Твоих, и буду размышлять о чудесах Твоих.
PS|118|28|Душа моя истаевает от скорби: укрепи меня по слову Твоему.
PS|118|29|Удали от меня путь лжи, и закон Твой даруй мне.
PS|118|30|Я избрал путь истины, поставил пред собою суды Твои.
PS|118|31|Я прилепился к откровениям Твоим, Господи; не постыди меня.
PS|118|32|Потеку путем заповедей Твоих, когда Ты расширишь сердце мое.
PS|118|33|Укажи мне, Господи, путь уставов Твоих, и я буду держаться его до конца.
PS|118|34|Вразуми меня, и буду соблюдать закон Твой и хранить его всем сердцем.
PS|118|35|Поставь меня на стезю заповедей Твоих, ибо я возжелал ее.
PS|118|36|Приклони сердце мое к откровениям Твоим, а не к корысти.
PS|118|37|Отврати очи мои, чтобы не видеть суеты; животвори меня на пути Твоем.
PS|118|38|Утверди слово Твое рабу Твоему, ради благоговения пред Тобою.
PS|118|39|Отврати поношение мое, которого я страшусь, ибо суды Твои благи.
PS|118|40|Вот, я возжелал повелений Твоих; животвори меня правдою Твоею.
PS|118|41|Да придут ко мне милости Твои, Господи, спасение Твое по слову Твоему, –
PS|118|42|и я дам ответ поносящему меня, ибо уповаю на слово Твое.
PS|118|43|Не отнимай совсем от уст моих слова истины, ибо я уповаю на суды Твои
PS|118|44|и буду хранить закон Твой всегда, во веки и веки;
PS|118|45|буду ходить свободно, ибо я взыскал повелений Твоих;
PS|118|46|буду говорить об откровениях Твоих пред царями и не постыжусь;
PS|118|47|буду утешаться заповедями Твоими, которые возлюбил;
PS|118|48|руки мои буду простирать к заповедям Твоим, которые возлюбил, и размышлять об уставах Твоих.
PS|118|49|Вспомни слово Твое к рабу Твоему, на которое Ты повелел мне уповать:
PS|118|50|это – утешение в бедствии моем, что слово Твое оживляет меня.
PS|118|51|Гордые крайне ругались надо мною, но я не уклонился от закона Твоего.
PS|118|52|Вспоминал суды Твои, Господи, от века, и утешался.
PS|118|53|Ужас овладевает мною при виде нечестивых, оставляющих закон Твой.
PS|118|54|Уставы Твои были песнями моими на месте странствований моих.
PS|118|55|Ночью вспоминал я имя Твое, Господи, и хранил закон Твой.
PS|118|56|Он стал моим, ибо повеления Твои храню.
PS|118|57|Удел мой, Господи, сказал я, соблюдать слова Твои.
PS|118|58|Молился я Тебе всем сердцем: помилуй меня по слову Твоему.
PS|118|59|Размышлял о путях моих и обращал стопы мои к откровениям Твоим.
PS|118|60|Спешил и не медлил соблюдать заповеди Твои.
PS|118|61|Сети нечестивых окружили меня, но я не забывал закона Твоего.
PS|118|62|В полночь вставал славословить Тебя за праведные суды Твои.
PS|118|63|Общник я всем боящимся Тебя и хранящим повеления Твои.
PS|118|64|Милости Твоей, Господи, полна земля; научи меня уставам Твоим.
PS|118|65|Благо сотворил Ты рабу Твоему, Господи, по слову Твоему.
PS|118|66|Доброму разумению и ведению научи меня, ибо заповедям Твоим я верую.
PS|118|67|Прежде страдания моего я заблуждался; а ныне слово Твое храню.
PS|118|68|Благ и благодетелен Ты, – научи меня уставам Твоим.
PS|118|69|Гордые сплетают на меня ложь; я же всем сердцем буду хранить повеления Твои.
PS|118|70|Ожирело сердце их, как тук; я же законом Твоим утешаюсь.
PS|118|71|Благо мне, что я пострадал, дабы научиться уставам Твоим.
PS|118|72|Закон уст Твоих для меня лучше тысяч золота и серебра.
PS|118|73|Руки Твои сотворили меня и устроили меня; вразуми меня, и научусь заповедям Твоим.
PS|118|74|Боящиеся Тебя увидят меня – и возрадуются, что я уповаю на слово Твое.
PS|118|75|Знаю, Господи, что суды Твои праведны и по справедливости Ты наказал меня.
PS|118|76|Да будет же милость Твоя утешением моим, по слову Твоему к рабу Твоему.
PS|118|77|Да придет ко мне милосердие Твое, и я буду жить; ибо закон Твой – утешение мое.
PS|118|78|Да будут постыжены гордые, ибо безвинно угнетают меня; я размышляю о повелениях Твоих.
PS|118|79|Да обратятся ко мне боящиеся Тебя и знающие откровения Твои.
PS|118|80|Да будет сердце мое непорочно в уставах Твоих, чтобы я не посрамился.
PS|118|81|Истаевает душа моя о спасении Твоем; уповаю на слово Твое.
PS|118|82|Истаевают очи мои о слове Твоем; я говорю: когда Ты утешишь меня?
PS|118|83|Я стал, как мех в дыму, [но] уставов Твоих не забыл.
PS|118|84|Сколько дней раба Твоего? Когда произведешь суд над гонителями моими?
PS|118|85|Яму вырыли мне гордые, вопреки закону Твоему.
PS|118|86|Все заповеди Твои – истина; несправедливо преследуют меня: помоги мне;
PS|118|87|едва не погубили меня на земле, но я не оставил повелений Твоих.
PS|118|88|По милости Твоей оживляй меня, и буду хранить откровения уст Твоих.
PS|118|89|На веки, Господи, слово Твое утверждено на небесах;
PS|118|90|истина Твоя в род и род. Ты поставил землю, и она стоит.
PS|118|91|По определениям Твоим все стоит доныне, ибо все служит Тебе.
PS|118|92|Если бы не закон Твой был утешением моим, погиб бы я в бедствии моем.
PS|118|93|Вовек не забуду повелений Твоих, ибо ими Ты оживляешь меня.
PS|118|94|Твой я, спаси меня; ибо я взыскал повелений Твоих.
PS|118|95|Нечестивые подстерегают меня, чтобы погубить; [а] я углубляюсь в откровения Твои.
PS|118|96|Я видел предел всякого совершенства, [но] Твоя заповедь безмерно обширна.
PS|118|97|Как люблю я закон Твой! весь день размышляю о нем.
PS|118|98|Заповедью Твоею Ты соделал меня мудрее врагов моих, ибо она всегда со мною.
PS|118|99|Я стал разумнее всех учителей моих, ибо размышляю об откровениях Твоих.
PS|118|100|Я сведущ более старцев, ибо повеления Твои храню.
PS|118|101|От всякого злого пути удерживаю ноги мои, чтобы хранить слово Твое;
PS|118|102|от судов Твоих не уклоняюсь, ибо Ты научаешь меня.
PS|118|103|Как сладки гортани моей слова Твои! лучше меда устам моим.
PS|118|104|Повелениями Твоими я вразумлен; потому ненавижу всякий путь лжи.
PS|118|105|Слово Твое – светильник ноге моей и свет стезе моей.
PS|118|106|Я клялся хранить праведные суды Твои, и исполню.
PS|118|107|Сильно угнетен я, Господи; оживи меня по слову Твоему.
PS|118|108|Благоволи же, Господи, принять добровольную жертву уст моих, и судам Твоим научи меня.
PS|118|109|Душа моя непрестанно в руке моей, но закона Твоего не забываю.
PS|118|110|Нечестивые поставили для меня сеть, но я не уклонился от повелений Твоих.
PS|118|111|Откровения Твои я принял, как наследие на веки, ибо они веселие сердца моего.
PS|118|112|Я приклонил сердце мое к исполнению уставов Твоих навек, до конца.
PS|118|113|Вымыслы [человеческие] ненавижу, а закон Твой люблю.
PS|118|114|Ты покров мой и щит мой; на слово Твое уповаю.
PS|118|115|Удалитесь от меня, беззаконные, и буду хранить заповеди Бога моего.
PS|118|116|Укрепи меня по слову Твоему, и буду жить; не посрами меня в надежде моей;
PS|118|117|поддержи меня, и спасусь; и в уставы Твои буду вникать непрестанно.
PS|118|118|Всех, отступающих от уставов Твоих, Ты низлагаешь, ибо ухищрения их – ложь.
PS|118|119|[Как] изгарь, отметаешь Ты всех нечестивых земли; потому я возлюбил откровения Твои.
PS|118|120|Трепещет от страха Твоего плоть моя, и судов Твоих я боюсь.
PS|118|121|Я совершал суд и правду; не предай меня гонителям моим.
PS|118|122|Заступи раба Твоего ко благу [его], чтобы не угнетали меня гордые.
PS|118|123|Истаевают очи мои, ожидая спасения Твоего и слова правды Твоей.
PS|118|124|Сотвори с рабом Твоим по милости Твоей, и уставам Твоим научи меня.
PS|118|125|Я раб Твой: вразуми меня, и познаю откровения Твои.
PS|118|126|Время Господу действовать: закон Твой разорили.
PS|118|127|А я люблю заповеди Твои более золота, и золота чистого.
PS|118|128|Все повеления Твои – все признаю справедливыми; всякий путь лжи ненавижу.
PS|118|129|Дивны откровения Твои; потому хранит их душа моя.
PS|118|130|Откровение слов Твоих просвещает, вразумляет простых.
PS|118|131|Открываю уста мои и вздыхаю, ибо заповедей Твоих жажду.
PS|118|132|Призри на меня и помилуй меня, как поступаешь с любящими имя Твое.
PS|118|133|Утверди стопы мои в слове Твоем и не дай овладеть мною никакому беззаконию;
PS|118|134|избавь меня от угнетения человеческого, и буду хранить повеления Твои;
PS|118|135|осияй раба Твоего светом лица Твоего и научи меня уставам Твоим.
PS|118|136|Из глаз моих текут потоки вод от того, что не хранят закона Твоего.
PS|118|137|Праведен Ты, Господи, и справедливы суды Твои.
PS|118|138|Откровения Твои, которые Ты заповедал, – правда и совершенная истина.
PS|118|139|Ревность моя снедает меня, потому что мои враги забыли слова Твои.
PS|118|140|Слово Твое весьма чисто, и раб Твой возлюбил его.
PS|118|141|Мал я и презрен, [но] повелений Твоих не забываю.
PS|118|142|Правда Твоя – правда вечная, и закон Твой – истина.
PS|118|143|Скорбь и горесть постигли меня; заповеди Твои – утешение мое.
PS|118|144|Правда откровений Твоих вечна: вразуми меня, и буду жить.
PS|118|145|Взываю всем сердцем [моим]: услышь меня, Господи, – и сохраню уставы Твои.
PS|118|146|Призываю Тебя: спаси меня, и буду хранить откровения Твои.
PS|118|147|Предваряю рассвет и взываю; на слово Твое уповаю.
PS|118|148|Очи мои предваряют [утреннюю] стражу, чтобы мне углубляться в слово Твое.
PS|118|149|Услышь голос мой по милости Твоей, Господи; по суду Твоему оживи меня.
PS|118|150|Приблизились замышляющие лукавство; далеки они от закона Твоего.
PS|118|151|Близок Ты, Господи, и все заповеди Твои – истина.
PS|118|152|Издавна узнал я об откровениях Твоих, что Ты утвердил их на веки.
PS|118|153|Воззри на бедствие мое и избавь меня, ибо я не забываю закона Твоего.
PS|118|154|Вступись в дело мое и защити меня; по слову Твоему оживи меня.
PS|118|155|Далеко от нечестивых спасение, ибо они уставов Твоих не ищут.
PS|118|156|Много щедрот Твоих, Господи; по суду Твоему оживи меня.
PS|118|157|Много у меня гонителей и врагов, [но] от откровений Твоих я не удаляюсь.
PS|118|158|Вижу отступников, и сокрушаюсь, ибо они не хранят слова Твоего.
PS|118|159|Зри, как я люблю повеления Твои; по милости Твоей, Господи, оживи меня.
PS|118|160|Основание слова Твоего истинно, и вечен всякий суд правды Твоей.
PS|118|161|Князья гонят меня безвинно, но сердце мое боится слова Твоего.
PS|118|162|Радуюсь я слову Твоему, как получивший великую прибыль.
PS|118|163|Ненавижу ложь и гнушаюсь ею; закон же Твой люблю.
PS|118|164|Семикратно в день прославляю Тебя за суды правды Твоей.
PS|118|165|Велик мир у любящих закон Твой, и нет им преткновения.
PS|118|166|Уповаю на спасение Твое, Господи, и заповеди Твои исполняю.
PS|118|167|Душа моя хранит откровения Твои, и я люблю их крепко.
PS|118|168|Храню повеления Твои и откровения Твои, ибо все пути мои пред Тобою.
PS|118|169|Да приблизится вопль мой пред лице Твое, Господи; по слову Твоему вразуми меня.
PS|118|170|Да придет моление мое пред лице Твое; по слову Твоему избавь меня.
PS|118|171|Уста мои произнесут хвалу, когда Ты научишь меня уставам Твоим.
PS|118|172|Язык мой возгласит слово Твое, ибо все заповеди Твои праведны.
PS|118|173|Да будет рука Твоя в помощь мне, ибо я повеления Твои избрал.
PS|118|174|Жажду спасения Твоего, Господи, и закон Твой – утешение мое.
PS|118|175|Да живет душа моя и славит Тебя, и суды Твои да помогут мне.
PS|118|176|Я заблудился, как овца потерянная: взыщи раба Твоего, ибо я заповедей Твоих не забыл.
PS|119|1|Песнь восхождения. К Господу воззвал я в скорби моей, и Он услышал меня.
PS|119|2|Господи! избавь душу мою от уст лживых, от языка лукавого.
PS|119|3|Что даст тебе и что прибавит тебе язык лукавый?
PS|119|4|Изощренные стрелы сильного, с горящими углями дроковыми.
PS|119|5|Горе мне, что я пребываю у Мосоха, живу у шатров Кидарских.
PS|119|6|Долго жила душа моя с ненавидящими мир.
PS|119|7|Я мирен: но только заговорю, они – к войне.
PS|120|1|Песнь восхождения. Возвожу очи мои к горам, откуда придет помощь моя.
PS|120|2|Помощь моя от Господа, сотворившего небо и землю.
PS|120|3|Не даст Он поколебаться ноге твоей, не воздремлет хранящий тебя;
PS|120|4|не дремлет и не спит хранящий Израиля.
PS|120|5|Господь – хранитель твой; Господь – сень твоя с правой руки твоей.
PS|120|6|Днем солнце не поразит тебя, ни луна ночью.
PS|120|7|Господь сохранит тебя от всякого зла; сохранит душу твою [Господь].
PS|120|8|Господь будет охранять выхождение твое и вхождение твое отныне и вовек.
PS|121|1|Песнь восхождения. Давида. Возрадовался я, когда сказали мне: "пойдем в дом Господень".
PS|121|2|Вот, стоят ноги наши во вратах твоих, Иерусалим, –
PS|121|3|Иерусалим, устроенный как город, слитый в одно,
PS|121|4|куда восходят колена, колена Господни, по закону Израилеву, славить имя Господне.
PS|121|5|Там стоят престолы суда, престолы дома Давидова.
PS|121|6|Просите мира Иерусалиму: да благоденствуют любящие тебя!
PS|121|7|Да будет мир в стенах твоих, благоденствие – в чертогах твоих!
PS|121|8|Ради братьев моих и ближних моих говорю я: "мир тебе!"
PS|121|9|Ради дома Господа, Бога нашего, желаю блага тебе.
PS|122|1|Песнь восхождения. К Тебе возвожу очи мои, Живущий на небесах!
PS|122|2|Вот, как очи рабов [обращены] на руку господ их, как очи рабы – на руку госпожи ее, так очи наши – к Господу, Богу нашему, доколе Он помилует нас.
PS|122|3|Помилуй нас, Господи, помилуй нас, ибо довольно мы насыщены презрением;
PS|122|4|довольно насыщена душа наша поношением от надменных и уничижением от гордых.
PS|123|1|Песнь восхождения. Давида. Если бы не Господь был с нами, – да скажет Израиль, –
PS|123|2|если бы не Господь был с нами, когда восстали на нас люди,
PS|123|3|то живых они поглотили бы нас, когда возгорелась ярость их на нас;
PS|123|4|воды потопили бы нас, поток прошел бы над душею нашею;
PS|123|5|прошли бы над душею нашею воды бурные.
PS|123|6|Благословен Господь, Который не дал нас в добычу зубам их!
PS|123|7|Душа наша избавилась, как птица, из сети ловящих: сеть расторгнута, и мы избавились.
PS|123|8|Помощь наша – в имени Господа, сотворившего небо и землю.
PS|124|1|Песнь восхождения. Давида. Надеющийся на Господа, как гора Сион, не подвигнется: пребывает вовек.
PS|124|2|Горы окрест Иерусалима, а Господь окрест народа Своего отныне и вовек.
PS|124|3|Ибо не оставит [Господь] жезла нечестивых над жребием праведных, дабы праведные не простерли рук своих к беззаконию.
PS|124|4|Благотвори, Господи, добрым и правым в сердцах своих;
PS|124|5|а совращающихся на кривые пути свои да оставит Господь ходить с делающими беззаконие. Мир на Израиля!
PS|125|1|Песнь восхождения. Когда возвращал Господь плен Сиона, мы были как бы видящие во сне:
PS|125|2|тогда уста наши были полны веселья, и язык наш – пения; тогда между народами говорили: "великое сотворил Господь над ними!"
PS|125|3|Великое сотворил Господь над нами: мы радовались.
PS|125|4|Возврати, Господи, пленников наших, как потоки на полдень.
PS|125|5|Сеявшие со слезами будут пожинать с радостью.
PS|125|6|С плачем несущий семена возвратится с радостью, неся снопы свои.
PS|126|1|Песнь восхождения. Соломона. Если Господь не созиждет дома, напрасно трудятся строящие его; если Господь не охранит города, напрасно бодрствует страж.
PS|126|2|Напрасно вы рано встаете, поздно просиживаете, едите хлеб печали, тогда как возлюбленному Своему Он дает сон.
PS|126|3|Вот наследие от Господа: дети; награда от Него – плод чрева.
PS|126|4|Что стрелы в руке сильного, то сыновья молодые.
PS|126|5|Блажен человек, который наполнил ими колчан свой! Не останутся они в стыде, когда будут говорить с врагами в воротах.
PS|127|1|Песнь восхождения. Блажен всякий боящийся Господа, ходящий путями Его!
PS|127|2|Ты будешь есть от трудов рук твоих: блажен ты, и благо тебе!
PS|127|3|Жена твоя, как плодовитая лоза, в доме твоем; сыновья твои, как масличные ветви, вокруг трапезы твоей:
PS|127|4|так благословится человек, боящийся Господа!
PS|127|5|Благословит тебя Господь с Сиона, и увидишь благоденствие Иерусалима во все дни жизни твоей;
PS|127|6|увидишь сыновей у сыновей твоих. Мир на Израиля!
PS|128|1|Песнь восхождения. Много теснили меня от юности моей, да скажет Израиль:
PS|128|2|много теснили меня от юности моей, но не одолели меня.
PS|128|3|На хребте моем орали оратаи, проводили длинные борозды свои.
PS|128|4|Но Господь праведен: Он рассек узы нечестивых.
PS|128|5|Да постыдятся и обратятся назад все ненавидящие Сион!
PS|128|6|Да будут, как трава на кровлях, которая прежде, нежели будет исторгнута, засыхает,
PS|128|7|которою жнец не наполнит руки своей, и вяжущий снопы – горсти своей;
PS|128|8|и проходящие мимо не скажут: "благословение Господне на вас; благословляем вас именем Господним!"
PS|129|1|Песнь восхождения. Из глубины взываю к Тебе, Господи.
PS|129|2|Господи! услышь голос мой. Да будут уши Твои внимательны к голосу молений моих.
PS|129|3|Если Ты, Господи, будешь замечать беззакония, – Господи! кто устоит?
PS|129|4|Но у Тебя прощение, да благоговеют пред Тобою.
PS|129|5|Надеюсь на Господа, надеется душа моя; на слово Его уповаю.
PS|129|6|Душа моя ожидает Господа более, нежели стражи – утра, более, нежели стражи – утра.
PS|129|7|Да уповает Израиль на Господа, ибо у Господа милость и многое у Него избавление,
PS|129|8|и Он избавит Израиля от всех беззаконий его.
PS|130|1|Песнь восхождения. Давида. Господи! не надмевалось сердце мое и не возносились очи мои, и я не входил в великое и для меня недосягаемое.
PS|130|2|Не смирял ли я и не успокаивал ли души моей, как дитяти, отнятого от груди матери? душа моя была во мне, как дитя, отнятое от груди.
PS|130|3|Да уповает Израиль на Господа отныне и вовек.
PS|131|1|Песнь восхождения. Вспомни, Господи, Давида и все сокрушение его:
PS|131|2|как он клялся Господу, давал обет Сильному Иакова:
PS|131|3|"не войду в шатер дома моего, не взойду на ложе мое;
PS|131|4|не дам сна очам моим и веждам моим – дремания,
PS|131|5|доколе не найду места Господу, жилища – Сильному Иакова".
PS|131|6|Вот, мы слышали о нем в Ефрафе, нашли его на полях Иарима.
PS|131|7|Пойдем к жилищу Его, поклонимся подножию ног Его.
PS|131|8|Стань, Господи, на [место] покоя Твоего, – Ты и ковчег могущества Твоего.
PS|131|9|Священники Твои облекутся правдою, и святые Твои возрадуются.
PS|131|10|Ради Давида, раба Твоего, не отврати лица помазанника Твоего.
PS|131|11|Клялся Господь Давиду в истине, и не отречется ее: "от плода чрева твоего посажу на престоле твоем.
PS|131|12|Если сыновья твои будут сохранять завет Мой и откровения Мои, которым Я научу их, то и их сыновья во веки будут сидеть на престоле твоем".
PS|131|13|Ибо избрал Господь Сион, возжелал [его] в жилище Себе.
PS|131|14|"Это покой Мой на веки: здесь вселюсь, ибо Я возжелал его.
PS|131|15|Пищу его благословляя благословлю, нищих его насыщу хлебом;
PS|131|16|священников его облеку во спасение, и святые его радостью возрадуются.
PS|131|17|Там возращу рог Давиду, поставлю светильник помазаннику Моему.
PS|131|18|Врагов его облеку стыдом, а на нем будет сиять венец его".
PS|132|1|Песнь восхождения. Давида. Как хорошо и как приятно жить братьям вместе!
PS|132|2|[Это] – как драгоценный елей на голове, стекающий на бороду, бороду Ааронову, стекающий на края одежды его;
PS|132|3|как роса Ермонская, сходящая на горы Сионские, ибо там заповедал Господь благословение и жизнь на веки.
PS|133|1|Песнь восхождения. Благословите ныне Господа, все рабы Господни, стоящие в доме Господнем, во время ночи.
PS|133|2|Воздвигните руки ваши к святилищу, и благословите Господа.
PS|133|3|Благословит тебя Господь с Сиона, сотворивший небо и землю.
PS|134|1|Аллилуия. Хвалите имя Господне, хвалите, рабы Господни,
PS|134|2|стоящие в доме Господнем, во дворах дома Бога нашего.
PS|134|3|Хвалите Господа, ибо Господь благ; пойте имени Его, ибо это сладостно,
PS|134|4|ибо Господь избрал Себе Иакова, Израиля в собственность Свою.
PS|134|5|Я познал, что велик Господь, и Господь наш превыше всех богов.
PS|134|6|Господь творит все, что хочет, на небесах и на земле, на морях и во всех безднах;
PS|134|7|возводит облака от края земли, творит молнии при дожде, изводит ветер из хранилищ Своих.
PS|134|8|Он поразил первенцев Египта, от человека до скота,
PS|134|9|послал знамения и чудеса среди тебя, Египет, на фараона и на всех рабов его,
PS|134|10|поразил народы многие и истребил царей сильных:
PS|134|11|Сигона, царя Аморрейского, и Ога, царя Васанского, и все царства Ханаанские;
PS|134|12|и отдал землю их в наследие, в наследие Израилю, народу Своему.
PS|134|13|Господи! имя Твое вовек; Господи! память о Тебе в род и род.
PS|134|14|Ибо Господь будет судить народ Свой и над рабами Своими умилосердится.
PS|134|15|Идолы язычников – серебро и золото, дело рук человеческих:
PS|134|16|есть у них уста, но не говорят; есть у них глаза, но не видят;
PS|134|17|есть у них уши, но не слышат, и нет дыхания в устах их.
PS|134|18|Подобны им будут делающие их и всякий, кто надеется на них.
PS|134|19|Дом Израилев! благословите Господа. Дом Ааронов! благословите Господа.
PS|134|20|Дом Левиин! благословите Господа. Боящиеся Господа! благословите Господа.
PS|134|21|Благословен Господь от Сиона, живущий в Иерусалиме! Аллилуия!
PS|135|1|Славьте Господа, ибо Он благ, ибо вовек милость Его.
PS|135|2|Славьте Бога богов, ибо вовек милость Его.
PS|135|3|Славьте Господа господствующих, ибо вовек милость Его;
PS|135|4|Того, Который один творит чудеса великие, ибо вовек милость Его;
PS|135|5|Который сотворил небеса премудро, ибо вовек милость Его;
PS|135|6|утвердил землю на водах, ибо вовек милость Его;
PS|135|7|сотворил светила великие, ибо вовек милость Его;
PS|135|8|солнце – для управления днем, ибо вовек милость Его;
PS|135|9|луну и звезды – для управления ночью, ибо вовек милость Его;
PS|135|10|поразил Египет в первенцах его, ибо вовек милость Его;
PS|135|11|и вывел Израиля из среды его, ибо вовек милость Его;
PS|135|12|рукою крепкою и мышцею простертою, ибо вовек милость Его;
PS|135|13|разделил Чермное море, ибо вовек милость Его;
PS|135|14|и провел Израиля посреди его, ибо вовек милость Его;
PS|135|15|и низверг фараона и войско его в море Чермное, ибо вовек милость Его;
PS|135|16|провел народ Свой чрез пустыню, ибо вовек милость Его;
PS|135|17|поразил царей великих, ибо вовек милость Его;
PS|135|18|и убил царей сильных, ибо вовек милость Его;
PS|135|19|Сигона, царя Аморрейского, ибо вовек милость Его;
PS|135|20|и Ога, царя Васанского, ибо вовек милость Его;
PS|135|21|и отдал землю их в наследие, ибо вовек милость Его;
PS|135|22|в наследие Израилю, рабу Своему, ибо вовек милость Его;
PS|135|23|вспомнил нас в унижении нашем, ибо вовек милость Его;
PS|135|24|и избавил нас от врагов наших, ибо вовек милость Его;
PS|135|25|дает пищу всякой плоти, ибо вовек милость Его.
PS|135|26|Славьте Бога небес, ибо вовек милость Его.
PS|136|1|При реках Вавилона, там сидели мы и плакали, когда вспоминали о Сионе;
PS|136|2|на вербах, посреди его, повесили мы наши арфы.
PS|136|3|Там пленившие нас требовали от нас слов песней, и притеснители наши – веселья: "пропойте нам из песней Сионских".
PS|136|4|Как нам петь песнь Господню на земле чужой?
PS|136|5|Если я забуду тебя, Иерусалим, – забудь меня десница моя;
PS|136|6|прилипни язык мой к гортани моей, если не буду помнить тебя, если не поставлю Иерусалима во главе веселия моего.
PS|136|7|Припомни, Господи, сынам Едомовым день Иерусалима, когда они говорили: "разрушайте, разрушайте до основания его".
PS|136|8|Дочь Вавилона, опустошительница! блажен, кто воздаст тебе за то, что ты сделала нам!
PS|136|9|Блажен, кто возьмет и разобьет младенцев твоих о камень!
PS|137|1|Давида. Славлю Тебя всем сердцем моим, пред богами пою Тебе.
PS|137|2|Поклоняюсь пред святым храмом Твоим и славлю имя Твое за милость Твою и за истину Твою, ибо Ты возвеличил слово Твое превыше всякого имени Твоего.
PS|137|3|В день, когда я воззвал, Ты услышал меня, вселил в душу мою бодрость.
PS|137|4|Прославят Тебя, Господи, все цари земные, когда услышат слова уст Твоих
PS|137|5|и воспоют пути Господни, ибо велика слава Господня.
PS|137|6|Высок Господь: и смиренного видит, и гордого узнает издали.
PS|137|7|Если я пойду посреди напастей, Ты оживишь меня, прострешь на ярость врагов моих руку Твою, и спасет меня десница Твоя.
PS|137|8|Господь совершит за меня! Милость Твоя, Господи, вовек: дело рук Твоих не оставляй.
PS|138|1|Начальнику хора. Псалом Давида. Господи! Ты испытал меня и знаешь.
PS|138|2|Ты знаешь, когда я сажусь и когда встаю; Ты разумеешь помышления мои издали.
PS|138|3|Иду ли я, отдыхаю ли – Ты окружаешь меня, и все пути мои известны Тебе.
PS|138|4|Еще нет слова на языке моем, – Ты, Господи, уже знаешь его совершенно.
PS|138|5|Сзади и спереди Ты объемлешь меня, и полагаешь на мне руку Твою.
PS|138|6|Дивно для меня ведение [Твое], – высоко, не могу постигнуть его!
PS|138|7|Куда пойду от Духа Твоего, и от лица Твоего куда убегу?
PS|138|8|Взойду ли на небо – Ты там; сойду ли в преисподнюю – и там Ты.
PS|138|9|Возьму ли крылья зари и переселюсь на край моря, –
PS|138|10|и там рука Твоя поведет меня, и удержит меня десница Твоя.
PS|138|11|Скажу ли: "может быть, тьма скроет меня, и свет вокруг меня [сделается] ночью";
PS|138|12|но и тьма не затмит от Тебя, и ночь светла, как день: как тьма, так и свет.
PS|138|13|Ибо Ты устроил внутренности мои и соткал меня во чреве матери моей.
PS|138|14|Славлю Тебя, потому что я дивно устроен. Дивны дела Твои, и душа моя вполне сознает это.
PS|138|15|Не сокрыты были от Тебя кости мои, когда я созидаем был в тайне, образуем был во глубине утробы.
PS|138|16|Зародыш мой видели очи Твои; в Твоей книге записаны все дни, для меня назначенные, когда ни одного из них еще не было.
PS|138|17|Как возвышенны для меня помышления Твои, Боже, и как велико число их!
PS|138|18|Стану ли исчислять их, но они многочисленнее песка; когда я пробуждаюсь, я все еще с Тобою.
PS|138|19|О, если бы Ты, Боже, поразил нечестивого! Удалитесь от меня, кровожадные!
PS|138|20|Они говорят против Тебя нечестиво; суетное замышляют враги Твои.
PS|138|21|Мне ли не возненавидеть ненавидящих Тебя, Господи, и не возгнушаться восстающими на Тебя?
PS|138|22|Полною ненавистью ненавижу их: враги они мне.
PS|138|23|Испытай меня, Боже, и узнай сердце мое; испытай меня и узнай помышления мои;
PS|138|24|и зри, не на опасном ли я пути, и направь меня на путь вечный.
PS|139|1|Псалом. Начальнику хора. Псалом Давида.
PS|139|2|Избавь меня, Господи, от человека злого; сохрани меня от притеснителя:
PS|139|3|они злое мыслят в сердце, всякий день ополчаются на брань,
PS|139|4|изощряют язык свой, как змея; яд аспида под устами их.
PS|139|5|Соблюди меня, Господи, от рук нечестивого, сохрани меня от притеснителей, которые замыслили поколебать стопы мои.
PS|139|6|Гордые скрыли силки для меня и петли, раскинули сеть по дороге, тенета разложили для меня.
PS|139|7|Я сказал Господу: Ты Бог мой; услышь, Господи, голос молений моих!
PS|139|8|Господи, Господи, сила спасения моего! Ты покрыл голову мою в день брани.
PS|139|9|Не дай, Господи, желаемого нечестивому; не дай успеха злому замыслу его: они возгордятся.
PS|139|10|Да покроет головы окружающих меня зло собственных уст их.
PS|139|11|Да падут на них горящие угли; да будут они повержены в огонь, в пропасти, так, чтобы не встали.
PS|139|12|Человек злоязычный не утвердится на земле; зло увлечет притеснителя в погибель.
PS|139|13|Знаю, что Господь сотворит суд угнетенным и справедливость бедным.
PS|139|14|Так! праведные будут славить имя Твое; непорочные будут обитать пред лицем Твоим.
PS|140|1|Псалом Давида. Господи! к тебе взываю: поспеши ко мне, внемли голосу моления моего, когда взываю к Тебе.
PS|140|2|Да направится молитва моя, как фимиам, пред лице Твое, воздеяние рук моих – как жертва вечерняя.
PS|140|3|Положи, Господи, охрану устам моим, и огради двери уст моих;
PS|140|4|не дай уклониться сердцу моему к словам лукавым для извинения дел греховных вместе с людьми, делающими беззаконие, и да не вкушу я от сластей их.
PS|140|5|Пусть наказывает меня праведник: это милость; пусть обличает меня: это лучший елей, который не повредит голове моей; но мольбы мои – против злодейств их.
PS|140|6|Вожди их рассыпались по утесам и слышат слова мои, что они кротки.
PS|140|7|Как будто землю рассекают и дробят нас; сыплются кости наши в челюсти преисподней.
PS|140|8|Но к Тебе, Господи, Господи, очи мои; на Тебя уповаю, не отринь души моей!
PS|140|9|Сохрани меня от силков, поставленных для меня, от тенет беззаконников.
PS|140|10|Падут нечестивые в сети свои, а я перейду.
PS|141|1|Учение Давида. Молитва его, когда он был в пещере. Голосом моим к Господу воззвал я, голосом моим к Господу помолился;
PS|141|2|излил пред Ним моление мое; печаль мою открыл Ему.
PS|141|3|Когда изнемогал во мне дух мой, Ты знал стезю мою. На пути, которым я ходил, они скрытно поставили сети для меня.
PS|141|4|Смотрю на правую сторону, и вижу, что никто не признает меня: не стало для меня убежища, никто не заботится о душе моей.
PS|141|5|Я воззвал к Тебе, Господи, я сказал: Ты прибежище мое и часть моя на земле живых.
PS|141|6|Внемли воплю моему, ибо я очень изнемог; избавь меня от гонителей моих, ибо они сильнее меня.
PS|141|7|Выведи из темницы душу мою, чтобы мне славить имя Твое. Вокруг меня соберутся праведные, когда Ты явишь мне благодеяние.
PS|142|1|Псалом Давида. Господи! услышь молитву мою, внемли молению моему по истине Твоей; услышь меня по правде Твоей
PS|142|2|и не входи в суд с рабом Твоим, потому что не оправдается пред Тобой ни один из живущих.
PS|142|3|Враг преследует душу мою, втоптал в землю жизнь мою, принудил меня жить во тьме, как давно умерших, –
PS|142|4|и уныл во мне дух мой, онемело во мне сердце мое.
PS|142|5|Вспоминаю дни древние, размышляю о всех делах Твоих, рассуждаю о делах рук Твоих.
PS|142|6|Простираю к Тебе руки мои; душа моя – к Тебе, как жаждущая земля.
PS|142|7|Скоро услышь меня, Господи: дух мой изнемогает; не скрывай лица Твоего от меня, чтобы я не уподобился нисходящим в могилу.
PS|142|8|Даруй мне рано услышать милость Твою, ибо я на Тебя уповаю. Укажи мне путь, по которому мне идти, ибо к Тебе возношу я душу мою.
PS|142|9|Избавь меня, Господи, от врагов моих; к Тебе прибегаю.
PS|142|10|Научи меня исполнять волю Твою, потому что Ты Бог мой; Дух Твой благий да ведет меня в землю правды.
PS|142|11|Ради имени Твоего, Господи, оживи меня; ради правды Твоей выведи из напасти душу мою.
PS|142|12|И по милости Твоей истреби врагов моих и погуби всех, угнетающих душу мою, ибо я Твой раб.
PS|143|1|Давида. Благословен Господь, твердыня моя, научающий руки мои битве и персты мои брани,
PS|143|2|милость моя и ограждение мое, прибежище мое и Избавитель мой, щит мой, – и я на Него уповаю; Он подчиняет мне народ мой.
PS|143|3|Господи! что есть человек, что Ты знаешь о нем, и сын человеческий, что обращаешь на него внимание?
PS|143|4|Человек подобен дуновению; дни его – как уклоняющаяся тень.
PS|143|5|Господи! Приклони небеса Твои и сойди; коснись гор, и воздымятся;
PS|143|6|блесни молниею и рассей их; пусти стрелы Твои и расстрой их;
PS|143|7|простри с высоты руку Твою, избавь меня и спаси меня от вод многих, от руки сынов иноплеменных,
PS|143|8|которых уста говорят суетное и которых десница – десница лжи.
PS|143|9|Боже! новую песнь воспою Тебе, на десятиструнной псалтири воспою Тебе,
PS|143|10|дарующему спасение царям и избавляющему Давида, раба Твоего, от лютого меча.
PS|143|11|Избавь меня и спаси меня от руки сынов иноплеменных, которых уста говорят суетное и которых десница – десница лжи.
PS|143|12|Да будут сыновья наши, как разросшиеся растения в их молодости; дочери наши – как искусно изваянные столпы в чертогах.
PS|143|13|Да будут житницы наши полны, обильны всяким хлебом; да плодятся овцы наши тысячами и тьмами на пажитях наших;
PS|143|14|[да будут] волы наши тучны; да не будет ни расхищения, ни пропажи, ни воплей на улицах наших.
PS|143|15|Блажен народ, у которого это есть. Блажен народ, у которого Господь есть Бог.
PS|144|1|Хвала Давида. Буду превозносить Тебя, Боже мой, Царь [мой], и благословлять имя Твое во веки и веки.
PS|144|2|Всякий день буду благословлять Тебя и восхвалять имя Твое во веки и веки.
PS|144|3|Велик Господь и достохвален, и величие Его неисследимо.
PS|144|4|Род роду будет восхвалять дела Твои и возвещать о могуществе Твоем.
PS|144|5|А я буду размышлять о высокой славе величия Твоего и о дивных делах Твоих.
PS|144|6|Будут говорить о могуществе страшных дел Твоих, и я буду возвещать о величии Твоем.
PS|144|7|Будут провозглашать память великой благости Твоей и воспевать правду Твою.
PS|144|8|Щедр и милостив Господь, долготерпелив и многомилостив.
PS|144|9|Благ Господь ко всем, и щедроты Его на всех делах Его.
PS|144|10|Да славят Тебя, Господи, все дела Твои, и да благословляют Тебя святые Твои;
PS|144|11|да проповедуют славу царства Твоего, и да повествуют о могуществе Твоем,
PS|144|12|чтобы дать знать сынам человеческим о могуществе Твоем и о славном величии царства Твоего.
PS|144|13|Царство Твое – царство всех веков, и владычество Твое во все роды.
PS|144|14|Господь поддерживает всех падающих и восставляет всех низверженных.
PS|144|15|Очи всех уповают на Тебя, и Ты даешь им пищу их в свое время;
PS|144|16|открываешь руку Твою и насыщаешь все живущее по благоволению.
PS|144|17|Праведен Господь во всех путях Своих и благ во всех делах Своих.
PS|144|18|Близок Господь ко всем призывающим Его, ко всем призывающим Его в истине.
PS|144|19|Желание боящихся Его Он исполняет, вопль их слышит и спасает их.
PS|144|20|Хранит Господь всех любящих Его, а всех нечестивых истребит.
PS|144|21|Уста мои изрекут хвалу Господню, и да благословляет всякая плоть святое имя Его во веки и веки.
PS|145|1|Хвали, душа моя, Господа.
PS|145|2|Буду восхвалять Господа, доколе жив; буду петь Богу моему, доколе есмь.
PS|145|3|Не надейтесь на князей, на сына человеческого, в котором нет спасения.
PS|145|4|Выходит дух его, и он возвращается в землю свою: в тот день исчезают [все] помышления его.
PS|145|5|Блажен, кому помощник Бог Иаковлев, у кого надежда на Господа Бога его,
PS|145|6|сотворившего небо и землю, море и все, что в них, вечно хранящего верность,
PS|145|7|творящего суд обиженным, дающего хлеб алчущим. Господь разрешает узников,
PS|145|8|Господь отверзает очи слепым, Господь восставляет согбенных, Господь любит праведных.
PS|145|9|Господь хранит пришельцев, поддерживает сироту и вдову, а путь нечестивых извращает.
PS|145|10|Господь будет царствовать во веки, Бог твой, Сион, в род и род. Аллилуия.
PS|146|1|Хвалите Господа, ибо благо петь Богу нашему, ибо это сладостно, – хвала подобающая.
PS|146|2|Господь созидает Иерусалим, собирает изгнанников Израиля.
PS|146|3|Он исцеляет сокрушенных сердцем и врачует скорби их;
PS|146|4|исчисляет количество звезд; всех их называет именами их.
PS|146|5|Велик Господь наш и велика крепость [Его], и разум Его неизмерим.
PS|146|6|Смиренных возвышает Господь, а нечестивых унижает до земли.
PS|146|7|Пойте поочередно славословие Господу; пойте Богу нашему на гуслях.
PS|146|8|Он покрывает небо облаками, приготовляет для земли дождь, произращает на горах траву;
PS|146|9|дает скоту пищу его и птенцам ворона, взывающим [к] [Нему].
PS|146|10|Не на силу коня смотрит Он, не к [быстроте] ног человеческих благоволит, –
PS|146|11|благоволит Господь к боящимся Его, к уповающим на милость Его.
PS|147|1|Хвали, Иерусалим, Господа; хвали, Сион, Бога твоего,
PS|147|2|ибо Он укрепляет вереи ворот твоих, благословляет сынов твоих среди тебя;
PS|147|3|утверждает в пределах твоих мир; туком пшеницы насыщает тебя;
PS|147|4|посылает слово Свое на землю; быстро течет слово Его;
PS|147|5|дает снег, как волну; сыплет иней, как пепел;
PS|147|6|бросает град Свой кусками; перед морозом Его кто устоит?
PS|147|7|Пошлет слово Свое, и все растает; подует ветром Своим, и потекут воды.
PS|147|8|Он возвестил слово Свое Иакову, уставы Свои и суды Свои Израилю.
PS|147|9|Не сделал Он того никакому [другому] народу, и судов Его они не знают. Аллилуия.
PS|148|1|Хвалите Господа с небес, хвалите Его в вышних.
PS|148|2|Хвалите Его, все Ангелы Его, хвалите Его, все воинства Его.
PS|148|3|Хвалите Его, солнце и луна, хвалите Его, все звезды света.
PS|148|4|Хвалите Его, небеса небес и воды, которые превыше небес.
PS|148|5|Да хвалят имя Господа, ибо Он повелел, и сотворились;
PS|148|6|поставил их на веки и веки; дал устав, который не прейдет.
PS|148|7|Хвалите Господа от земли, великие рыбы и все бездны,
PS|148|8|огонь и град, снег и туман, бурный ветер, исполняющий слово Его,
PS|148|9|горы и все холмы, дерева плодоносные и все кедры,
PS|148|10|звери и всякий скот, пресмыкающиеся и птицы крылатые,
PS|148|11|цари земные и все народы, князья и все судьи земные,
PS|148|12|юноши и девицы, старцы и отроки
PS|148|13|да хвалят имя Господа, ибо имя Его единого превознесенно, слава Его на земле и на небесах.
PS|148|14|Он возвысил рог народа Своего, славу всех святых Своих, сынов Израилевых, народа, близкого к Нему. Аллилуия.
PS|149|1|Пойте Господу песнь новую; хвала Ему в собрании святых.
PS|149|2|Да веселится Израиль о Создателе своем; сыны Сиона да радуются о Царе своем.
PS|149|3|да хвалят имя Его с ликами, на тимпане и гуслях да поют Ему,
PS|149|4|ибо благоволит Господь к народу Своему, прославляет смиренных спасением.
PS|149|5|Да торжествуют святые во славе, да радуются на ложах своих.
PS|149|6|Да будут славословия Богу в устах их, и меч обоюдоострый в руке их,
PS|149|7|для того, чтобы совершать мщение над народами, наказание над племенами,
PS|149|8|заключать царей их в узы и вельмож их в оковы железные,
PS|149|9|производить над ними суд писанный. Честь сия – всем святым Его. Аллилуия.
PS|150|1|Хвалите Бога во святыне Его, хвалите Его на тверди силы Его.
PS|150|2|Хвалите Его по могуществу Его, хвалите Его по множеству величия Его.
PS|150|3|Хвалите Его со звуком трубным, хвалите Его на псалтири и гуслях.
PS|150|4|Хвалите Его с тимпаном и ликами, хвалите Его на струнах и органе.
PS|150|5|Хвалите Его на звучных кимвалах, хвалите Его на кимвалах громогласных.
PS|150|6|Все дышащее да хвалит Господа! Аллилуия.
