2PET|1|1|耶穌基督的僕人和使徒 西門．彼得 寫信給那因我們的上帝和 救主耶穌基督的義，與我們同得一樣寶貴信心的人。
2PET|1|2|願恩惠、平安 ，因你們認識上帝和我們的主耶穌，多多加給你們！
2PET|1|3|上帝的神能已把一切關乎生命和虔敬的事賜給我們，因我們認識那用自己榮耀和美德召我們的上帝。
2PET|1|4|因此，他已把又寶貴又極大的應許賜給我們，使我們既脫離世上從情慾來的敗壞，就得分享上帝的本性。
2PET|1|5|正因這緣故，你們要分外地努力。有了信心，又要加上德行；有了德行，又要加上知識；
2PET|1|6|有了知識，又要加上節制；有了節制，又要加上忍耐；有了忍耐，又要加上虔敬；
2PET|1|7|有了虔敬，又要加上愛弟兄的心；有了愛弟兄的心，又要加上愛眾人的心。
2PET|1|8|你們有了這幾樣，再繼續增長，就必使你們在認識我們的主耶穌基督上，不至於懶散和不結果子了。
2PET|1|9|沒有這幾樣的人就是瞎眼，是短視，忘了他過去的罪已經得了潔淨。
2PET|1|10|所以，弟兄們，要更加努力，使你們的蒙召和被選堅定不移。你們實行這幾樣，就永不失腳。
2PET|1|11|這樣，必叫你們豐豐富富地得以進入我們主－救主耶穌基督永遠的國度。
2PET|1|12|雖然你們已經知道這些事，並且在你們已有的真道上得到堅固，我還是要常常提醒你們這些事。
2PET|1|13|我認為趁我還在這帳棚的時候，應該激發你們的記憶，
2PET|1|14|因為知道我脫離這帳棚的時候快到了，正如我們的主耶穌基督所指示我的。
2PET|1|15|我也要盡心竭力，使你們在我去世以後時常記念這些事。
2PET|1|16|我們從前把我們主耶穌基督的大能和他來臨的事告訴你們，並不是隨從一些捏造出來的無稽傳說，我們是曾經親眼見過他的威榮的人。
2PET|1|17|他從父上帝得尊貴榮耀的時候，從至高無上的榮耀有聲音出來，對他說：「這是我的愛子，我所喜悅的。」
2PET|1|18|我們同他在聖山的時候，親自聽見這聲音從天上出來。
2PET|1|19|我們有先知更確實的信息，你們要好好地留意這信息，如同留意照耀在暗處的明燈，直等到天亮，晨星在你們心裏升起的時候。
2PET|1|20|第一要緊的，你們要知道，經上所有的預言是不可隨私意解釋的，
2PET|1|21|因為預言從來沒有出於人意的，而是人被聖靈感動說出上帝的話來。
2PET|2|1|從前在民間有假先知起來；同樣，將來在你們中間也會有假教師，偷偷地引進使人滅亡的異端。他們甚至不認買他們的主人，自取迅速滅亡。
2PET|2|2|許多人會隨從他們淫蕩的行為，以致真理之道因他們的緣故被毀謗。
2PET|2|3|他們因貪婪，要用捏造的言語在你們身上取得利益。他們的懲罰，自古以來並不遲延；他們的滅亡也必迅速來到。
2PET|2|4|既然上帝沒有寬容犯了罪的天使，反而把他們丟在地獄裏，囚禁在幽暗中等候審判；
2PET|2|5|既然上帝也沒有寬容上古的世界，曾叫洪水臨到那不敬虔的世界，只保護了報公義信息的 挪亞 一家八口；
2PET|2|6|既然上帝判決了 所多瑪 和 蛾摩拉 ，將二城傾覆 ，焚燒成灰，作為後世不敬虔人的鑒戒，
2PET|2|7|只搭救了那常為惡人的淫蕩憂傷的義人 羅得 —
2PET|2|8|因為那義人住在他們當中，他正義的心因天天看見和聽見他們不法的事而傷痛；
2PET|2|9|那麼，主知道搭救敬虔的人脫離試煉，把不義的人留在懲罰之下等候審判的日子，
2PET|2|10|尤其那些隨從肉體、放縱污穢的情慾、藐視主的權威的人更是如此。 他們膽大任性，無懼地毀謗眾尊榮者；
2PET|2|11|就是天使，雖然力量權能更大，在對他們宣告從主來的審判的時候還不用毀謗的話 。
2PET|2|12|但這些人好像沒有理性的牲畜，生來就是要被捉拿宰殺的。他們毀謗自己所不知道的事，正在敗壞人的時候，自己也遭遇敗壞，
2PET|2|13|為所行的不義受不義的工錢。他們喜愛白晝狂歡，他們已被玷污，又有瑕疵，正與你們一同歡宴，以自己的詭詐為樂。
2PET|2|14|他們滿眼是淫色，是止不住的罪，引誘心不堅定的人，心中習慣了貪婪，正是被詛咒的種類。
2PET|2|15|他們離棄了正路，走入歧途，隨從 比珥 的兒子 巴蘭 的路； 巴蘭 就是那貪愛不義的工錢的人，
2PET|2|16|他卻為自己的過犯受了責備，而那不能說話的驢以人的聲音阻止了先知的狂妄。
2PET|2|17|這些人是無水的泉源，是狂風催逼的霧氣，有漆黑的幽暗為他們存留。
2PET|2|18|他們說虛妄誇大的話，用肉體的情慾和淫蕩的事引誘那些剛脫離錯謬生活的人。
2PET|2|19|他們應許人自由，自己卻作了腐敗的奴隸，因為人被誰制伏就是誰的奴隸。
2PET|2|20|倘若他們因認識我們的主和救主耶穌基督而得以脫離世上的污穢，後來又被污穢纏住，被制伏，他們末後的景況就比先前更不好了。
2PET|2|21|他們知道義路，竟背棄了傳授給他們那神聖的誡命，倒不如不知道為妙。
2PET|2|22|俗語說得好，這話正印證在他們身上了： 「狗轉過來吃自己所吐的；」 又說： 「豬洗淨了，又回到爛泥裏打滾。」
2PET|3|1|親愛的，我現在寫給你們的是第二封信。在這兩封信裏，我都提醒你們，激發你們真誠的心，
2PET|3|2|要你們記得聖先知預先所說的話和主—救主的命令，就是使徒所傳給你們的。
2PET|3|3|第一要緊的，你們要知道，在末世必有好譏誚的人隨從自己的私慾出來譏誚，
2PET|3|4|說：「他要來臨的應許在哪裏呢？因為從列祖長眠以來，萬物與起初創造的時候仍是一樣啊！」
2PET|3|5|他們故意忘記這事，就是從太古憑上帝的話有了天，並由水而出和藉著水而成的地；
2PET|3|6|藉著水，當時的世界被水淹沒而消滅了。
2PET|3|7|但現在的天地還是憑著上帝的話存留，直留到不敬虔之人受審判遭沉淪的日子，用火焚燒。
2PET|3|8|親愛的，有一件事你們不可忘記，就是：主看一日如千年，千年如一日。
2PET|3|9|主沒有遲延他的應許，就如有人以為他是遲延，其實他是寬容你們，不願一人沉淪，而是人人都來悔改。
2PET|3|10|但主的日子要像賊一樣來到；那日，天必在轟然一聲中消失，天體都要被烈火熔化，地和地上的萬物都要燒盡 。
2PET|3|11|既然這一切都要如此消失，你們 處世為人必須聖潔敬虔，
2PET|3|12|等候並催促上帝的日子來到。因為在那日，天要被火燒而消滅，天體都要被烈火熔化。
2PET|3|13|但照他的應許，我們等候新天新地，其中有正義常住。
2PET|3|14|所以，親愛的，既然你們等候這些事，就要竭力使自己沒有玷污，無可指責，在主前和睦；
2PET|3|15|並且要以我們主的容忍作為你們得救的機會，就如我們所親愛的弟兄 保羅 ，照著所賜給他的智慧寫信給你們。
2PET|3|16|他一切的信上都談到這事。信中有些難明白的，那無學問、不堅定的人加以曲解，如曲解別的經書一樣，自取滅亡。
2PET|3|17|所以，親愛的，既然你們預先知道這事，就當防備，免得被惡人的錯謬誘惑，從自己穩定的立場上墜落。
2PET|3|18|你們倒要在我們的主和救主耶穌基督的恩典和知識上有長進。願榮耀歸給他，從今直到永遠之日。阿們！
