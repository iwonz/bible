JOSH|1|1|et factum est ut post mortem Mosi servi Domini loqueretur Dominus ad Iosue filium Nun ministrum Mosi et diceret ei
JOSH|1|2|Moses servus meus mortuus est surge et transi Iordanem istum tu et omnis populus tecum in terram quam ego dabo filiis Israhel
JOSH|1|3|omnem locum quem calcaverit vestigium pedis vestri vobis tradam sicut locutus sum Mosi
JOSH|1|4|a deserto et Libano usque ad fluvium magnum Eufraten omnis terra Hettheorum usque ad mare Magnum contra solis occasum erit terminus vester
JOSH|1|5|nullus vobis poterit resistere cunctis diebus vitae tuae sicut fui cum Mose ero et tecum non dimittam nec derelinquam te
JOSH|1|6|confortare et esto robustus tu enim sorte divides populo huic terram pro qua iuravi patribus suis ut traderem eam illis
JOSH|1|7|confortare igitur et esto robustus valde ut custodias et facias omnem legem quam praecepit tibi Moses servus meus ne declines ab ea ad dextram vel ad sinistram ut intellegas cuncta quae agis
JOSH|1|8|non recedat volumen legis huius de ore tuo sed meditaberis in eo diebus ac noctibus ut custodias et facias omnia quae scripta sunt in eo tunc diriges viam tuam et intelleges eam
JOSH|1|9|ecce praecipio tibi confortare et esto robustus noli metuere et noli timere quoniam tecum est Dominus Deus tuus in omnibus ad quaecumque perrexeris
JOSH|1|10|praecepitque Iosue principibus populi dicens transite per medium castrorum et imperate populo ac dicite
JOSH|1|11|praeparate vobis cibaria quoniam post diem tertium transibitis Iordanem et intrabitis ad possidendam terram quam Dominus Deus vester daturus est vobis
JOSH|1|12|Rubenitis quoque et Gadditis et dimidiae tribui Manasse ait
JOSH|1|13|mementote sermonis quem praecepit vobis Moses famulus Domini dicens Dominus Deus vester dedit vobis requiem et omnem terram
JOSH|1|14|uxores vestrae et filii ac iumenta manebunt in terra quam tradidit vobis Moses trans Iordanem vos autem transite armati ante fratres vestros omnes fortes manu et pugnate pro eis
JOSH|1|15|donec det requiem Dominus fratribus vestris sicut et vobis dedit et possideant ipsi quoque terram quam Dominus Deus vester daturus est eis et sic revertemini in terram possessionis vestrae et habitabitis in ea quam vobis dedit Moses famulus Domini trans Iordanem contra solis ortum
JOSH|1|16|responderuntque ad Iosue atque dixerunt omnia quae praecepisti nobis faciemus et quocumque miseris ibimus
JOSH|1|17|sicut oboedivimus in cunctis Mosi ita oboediemus et tibi tantum sit Dominus Deus tecum sicut fuit cum Mose
JOSH|1|18|qui contradixerit ori tuo et non oboedierit cunctis sermonibus quos praeceperis ei moriatur tu tantum confortare et viriliter age
JOSH|2|1|misit ergo Iosue filius Nun de Setthim duos viros exploratores abscondito et dixit eis ite et considerate terram urbemque Hiericho qui pergentes ingressi sunt domum mulieris meretricis nomine Raab et quieverunt apud eam
JOSH|2|2|nuntiatumque est regi Hiericho et dictum ecce viri ingressi sunt huc per noctem de filiis Israhel ut explorarent terram
JOSH|2|3|misitque rex Hiericho ad Raab dicens educ viros qui venerunt ad te et ingressi sunt domum tuam exploratores quippe sunt et omnem terram considerare venerunt
JOSH|2|4|tollensque mulier viros abscondit et ait fateor venerunt ad me sed nesciebam unde essent
JOSH|2|5|cumque porta clauderetur in tenebris et illi pariter exierunt nescio quo abierunt persequimini cito et conprehendetis eos
JOSH|2|6|ipsa autem fecit ascendere viros in solarium domus suae operuitque eos lini stipula quae ibi erat
JOSH|2|7|hii autem qui missi fuerant secuti sunt eos per viam quae ducit ad vadum Iordanis illisque egressis statim porta clausa est
JOSH|2|8|necdum obdormierant qui latebant et ecce mulier ascendit ad eos et ait
JOSH|2|9|novi quod tradiderit Dominus vobis terram etenim inruit in nos terror vester et elanguerunt omnes habitatores terrae
JOSH|2|10|audivimus quod siccaverit Dominus aquas maris Rubri ad vestrum introitum quando egressi estis ex Aegypto et quae feceritis duobus Amorreorum regibus qui erant trans Iordanem Seon et Og quos interfecistis
JOSH|2|11|et haec audientes pertimuimus et elanguit cor nostrum nec remansit in nobis spiritus ad introitum vestrum Dominus enim Deus vester ipse est Deus in caelo sursum et in terra deorsum
JOSH|2|12|nunc ergo iurate mihi per Dominum ut quomodo ego feci vobiscum misericordiam ita et vos faciatis cum domo patris mei detisque mihi signum verum
JOSH|2|13|et salvetis patrem meum et matrem fratres ac sorores meas et omnia quae eorum sunt et eruatis animas nostras de morte
JOSH|2|14|qui responderunt ei anima nostra sit pro vobis in mortem si tamen non prodideris nos cumque tradiderit nobis Dominus terram faciemus in te misericordiam et veritatem
JOSH|2|15|dimisit ergo eos per funem de fenestra domus enim eius herebat muro
JOSH|2|16|dixitque ad eos ad montana conscendite ne forte occurrant vobis revertentes ibique latete diebus tribus donec redeant et sic ibitis per viam vestram
JOSH|2|17|qui dixerunt ad eam innoxii erimus a iuramento hoc quo adiurasti nos
JOSH|2|18|si ingredientibus nobis terram signum fuerit funiculus iste coccineus et ligaveris eum in fenestra per quam nos dimisisti et patrem tuum ac matrem fratresque et omnem cognationem tuam congregaveris in domum tuam
JOSH|2|19|qui ostium domus tuae egressus fuerit sanguis ipsius erit in caput eius et nos erimus alieni cunctorum autem sanguis qui tecum fuerint in domo redundabit in caput nostrum si eos aliquis tetigerit
JOSH|2|20|quod si nos prodere volueris et sermonem istum proferre in medium erimus mundi ab hoc iuramento quo adiurasti nos
JOSH|2|21|et illa respondit sicut locuti estis ita fiat dimittensque eos ut pergerent adpendit funiculum coccineum in fenestra
JOSH|2|22|illi vero ambulantes pervenerunt ad montana et manserunt ibi tres dies donec reverterentur qui fuerant persecuti quaerentes enim per omnem viam non reppererunt eos
JOSH|2|23|quibus urbem ingressis reversi sunt et descenderunt exploratores de monte et Iordane transmisso venerunt ad Iosue filium Nun narraveruntque ei omnia quae acciderant sibi
JOSH|2|24|atque dixerunt tradidit Dominus in manus nostras omnem terram hanc et timore prostrati sunt cuncti habitatores eius
JOSH|3|1|igitur Iosue de nocte consurgens movit castra egredientesque de Setthim venerunt ad Iordanem ipse et omnes filii Israhel et morati sunt ibi per tres dies
JOSH|3|2|quibus evolutis transierunt praecones per castrorum medium
JOSH|3|3|et clamare coeperunt quando videritis arcam foederis Domini Dei vestri et sacerdotes stirpis leviticae portantes eam vos quoque consurgite et sequimini praecedentes
JOSH|3|4|sitque inter vos et arcam spatium cubitorum duum milium ut procul videre possitis et nosse per quam viam ingrediamini quia prius non ambulastis per eam et cavete ne adpropinquetis ad arcam
JOSH|3|5|dixitque Iosue ad populum sanctificamini cras enim faciet Dominus inter vos mirabilia
JOSH|3|6|et ait ad sacerdotes tollite arcam foederis et praecedite populum qui iussa conplentes tulerunt et ambulaverunt ante eos
JOSH|3|7|dixitque Dominus ad Iosue hodie incipiam exaltare te coram omni Israhel ut sciant quod sicut cum Mosi fui ita et tecum sim
JOSH|3|8|tu autem praecipe sacerdotibus qui portant arcam foederis et dic eis cum ingressi fueritis partem aquae Iordanis state in ea
JOSH|3|9|dixitque Iosue ad filios Israhel accedite huc et audite verba Domini Dei vestri
JOSH|3|10|et rursum in hoc inquit scietis quod Dominus Deus vivens in medio vestri est et disperdat in conspectu vestro Chananeum Hettheum Eveum et Ferezeum Gergeseum quoque et Amorreum et Iebuseum
JOSH|3|11|ecce arca foederis Domini omnis terrae antecedet vos per Iordanem
JOSH|3|12|parate duodecim viros de tribubus Israhel singulos per singulas tribus
JOSH|3|13|et cum posuerint vestigia pedum suorum sacerdotes qui portant arcam Domini Dei universae terrae in aquis Iordanis aquae quae inferiores sunt decurrent atque deficient quae autem desuper veniunt in una mole consistent
JOSH|3|14|igitur egressus est populus de tabernaculis suis ut transirent Iordanem et sacerdotes qui portabant arcam foederis pergebant ante eum
JOSH|3|15|ingressisque eis Iordanem et pedibus eorum tinctis in parte aquae cum Iordanis autem ripas alvei sui tempore messis impleret
JOSH|3|16|steterunt aquae descendentes in uno loco et instar montis intumescentes apparebant procul ab urbe quae vocatur Adom usque ad locum Sarthan quae autem inferiores erant in mare Solitudinis quod nunc vocatur Mortuum descenderunt usquequo omnino deficerent
JOSH|3|17|populus autem incedebat contra Iordanem et sacerdotes qui portabant arcam foederis Domini stabant super siccam humum in medio Iordanis accincti omnisque populus per arentem alveum transiebat
JOSH|4|1|quibus transgressis dixit Dominus ad Iosue
JOSH|4|2|elige duodecim viros singulos per singulas tribus
JOSH|4|3|et praecipe eis ut tollant de medio Iordanis alveo ubi steterunt sacerdotum pedes duodecim durissimos lapides quos ponetis in loco castrorum ubi fixeritis hac nocte tentoria
JOSH|4|4|vocavitque Iosue duodecim viros quos elegerat de filiis Israhel singulos de tribubus singulis
JOSH|4|5|et ait ad eos ite ante arcam Domini Dei vestri ad Iordanis medium et portate singuli singulos lapides in umeris vestris iuxta numerum filiorum Israhel
JOSH|4|6|ut sit signum inter vos et quando interrogaverint vos filii vestri cras dicentes quid sibi volunt isti lapides
JOSH|4|7|respondebitis eis defecerunt aquae Iordanis ante arcam foederis Domini cum transiret eum idcirco positi sunt lapides isti in monumentum filiorum Israhel usque in aeternum
JOSH|4|8|fecerunt ergo filii Israhel sicut eis praecepit Iosue portantes de medio Iordanis alveo duodecim lapides ut ei Dominus imperarat iuxta numerum filiorum Israhel usque ad locum in quo castrametati sunt ibique posuerunt eos
JOSH|4|9|alios quoque duodecim lapides posuit Iosue in medio Iordanis alveo ubi steterunt sacerdotes qui portabant arcam foederis et sunt ibi usque in praesentem diem
JOSH|4|10|sacerdotes autem qui portabant arcam stabant in Iordanis medio donec omnia conplerentur quae Iosue ut loqueretur ad populum praeceperat Dominus et dixerat ei Moses festinavitque populus et transiit
JOSH|4|11|cumque transissent omnes transivit et arca Domini sacerdotesque pergebant ante populum
JOSH|4|12|filii quoque Ruben et Gad et dimidiae tribus Manasse armati praecedebant filios Israhel sicut eis praeceperat Moses
JOSH|4|13|et quadraginta pugnatorum milia per turmas et cuneos incedebant per plana atque campestria urbis Hiericho
JOSH|4|14|in illo die magnificavit Dominus Iosue coram omni Israhel ut timerent eum sicut timuerant Mosen dum adviveret
JOSH|4|15|dixitque ad eum
JOSH|4|16|praecipe sacerdotibus qui portant arcam foederis ut ascendant de Iordane
JOSH|4|17|qui praecepit eis dicens ascendite de Iordane
JOSH|4|18|cumque ascendissent portantes arcam foederis Domini et siccam humum calcare coepissent reversae sunt aquae in alveum suum et fluebant sicut ante consueverant
JOSH|4|19|populus autem ascendit de Iordane decimo mensis primi die et castrametati sunt in Galgalis contra orientalem plagam urbis Hiericho
JOSH|4|20|duodecim quoque lapides quos de Iordanis alveo sumpserant posuit Iosue in Galgalis
JOSH|4|21|et dixit ad filios Israhel quando interrogaverint filii vestri cras patres suos et dixerint eis quid sibi volunt isti lapides
JOSH|4|22|docebitis eos atque dicetis per arentem alveum transivit Israhel Iordanem istum
JOSH|4|23|siccante Domino Deo vestro aquas eius in conspectu vestro donec transiretis
JOSH|4|24|sicut fecerat prius in mari Rubro quod siccavit donec transiremus
JOSH|4|25|ut discant omnes terrarum populi fortissimam Domini manum et ut vos timeatis Dominum Deum vestrum omni tempore
JOSH|5|1|postquam ergo audierunt omnes reges Amorreorum qui habitabant trans Iordanem ad occidentalem plagam et cuncti reges Chanaan qui propinqua possidebant Magno mari loca quod siccasset Dominus fluenta Iordanis coram filiis Israhel donec transirent dissolutum est cor eorum et non remansit in eis spiritus timentium introitum filiorum Israhel
JOSH|5|2|eo tempore ait Dominus ad Iosue fac tibi cultros lapideos et circumcide secundo filios Israhel
JOSH|5|3|fecit quod iusserat Dominus et circumcidit filios Israhel in colle Praeputiorum
JOSH|5|4|haec autem causa est secundae circumcisionis omnis populus qui egressus est ex Aegypto generis masculini universi bellatores viri mortui sunt in deserto per longissimos viae circuitus
JOSH|5|5|qui omnes circumcisi erant populus autem qui natus est in deserto
JOSH|5|6|per quadraginta annos itineris latissimae solitudinis incircumcisus fuit donec consumerentur qui non audierant vocem Domini et quibus ante iuraverat ut ostenderet eis terram lacte et melle manantem
JOSH|5|7|horum filii in locum successerunt patrum et circumcisi sunt ab Iosue quia sicut nati fuerant in praeputio erant nec eos in via aliquis circumciderat
JOSH|5|8|postquam autem omnes circumcisi sunt manserunt in eodem castrorum loco donec sanarentur
JOSH|5|9|dixitque Dominus ad Iosue hodie abstuli obprobrium Aegypti a vobis vocatumque est nomen loci illius Galgala usque in praesentem diem
JOSH|5|10|manseruntque filii Israhel in Galgalis et fecerunt phase quartadecima die mensis ad vesperum in campestribus Hiericho
JOSH|5|11|et comederunt de frugibus terrae die altero azymos panes et pulentam eiusdem anni
JOSH|5|12|defecitque manna postquam comederunt de frugibus terrae nec usi sunt ultra illo cibo filii Israhel sed comederunt de frugibus praesentis anni terrae Chanaan
JOSH|5|13|cum autem esset Iosue in agro urbis Hiericho levavit oculos et vidit virum stantem contra se et evaginatum tenentem gladium perrexitque ad eum et ait noster es an adversariorum
JOSH|5|14|qui respondit nequaquam sed sum princeps exercitus Domini et nunc venio
JOSH|5|15|cecidit Iosue pronus in terram et adorans ait quid dominus meus loquitur ad servum suum
JOSH|5|16|solve inquit calciamentum de pedibus tuis locus enim in quo stas sanctus est fecitque Iosue ut sibi fuerat imperatum
JOSH|6|1|Hiericho autem clausa erat atque munita timore filiorum Israhel et nullus egredi audebat aut ingredi
JOSH|6|2|dixitque Dominus ad Iosue ecce dedi in manus tuas Hiericho et regem eius omnesque fortes viros
JOSH|6|3|circuite urbem cuncti bellatores semel per diem sic facietis sex diebus
JOSH|6|4|septimo autem die sacerdotes tollant septem bucinas quarum usus est in iobeleo et praecedant arcam foederis septiesque circuibitis civitatem et sacerdotes clangent bucinis
JOSH|6|5|cumque insonuerit vox tubae longior atque concisior et in auribus vestris increpuerit conclamabit omnis populus vociferatione maxima et muri funditus corruent civitatis ingredienturque singuli per locum contra quem steterint
JOSH|6|6|vocavit ergo Iosue filius Nun sacerdotes et dixit ad eos tollite arcam foederis et septem alii sacerdotes tollant septem iobeleorum bucinas et incedant ante arcam Domini
JOSH|6|7|ad populum quoque ait vadite et circuite civitatem armati praecedentes arcam Domini
JOSH|6|8|cumque Iosue verba finisset et septem sacerdotes septem bucinis clangerent ante arcam foederis Domini
JOSH|6|9|omnisque praecederet armatus exercitus reliquum vulgus arcam sequebatur ac bucinis omnia concrepabant
JOSH|6|10|praeceperat autem Iosue populo dicens non clamabitis nec audietur vox vestra neque ullus sermo ex ore vestro egredietur donec veniat dies in quo dicam vobis clamate et vociferamini
JOSH|6|11|circuivit ergo arca Domini civitatem semel per diem et reversa in castra mansit ibi
JOSH|6|12|igitur Iosue de nocte consurgente tulerunt sacerdotes arcam Domini
JOSH|6|13|et septem ex eis septem bucinas quarum in iobeleis usus est praecedebantque arcam Domini ambulantes atque clangentes et armatus populus ibat ante eos vulgus autem reliquum sequebatur arcam et bucinis personabat
JOSH|6|14|circumieruntque civitatem secundo die semel et reversi sunt in castra sic fecerunt sex diebus
JOSH|6|15|die autem septimo diluculo consurgentes circumierunt urbem sicut dispositum erat septies
JOSH|6|16|cumque septimo circuitu clangerent bucinis sacerdotes dixit Iosue ad omnem Israhel vociferamini tradidit enim vobis Dominus civitatem
JOSH|6|17|sitque civitas haec anathema et omnia quae in ea sunt Domino sola Raab meretrix vivat cum universis qui cum ea in domo sunt abscondit enim nuntios quos direximus
JOSH|6|18|vos autem cavete ne de his quae praecepta sunt quippiam contingatis et sitis praevaricationis rei et omnia castra Israhel sub peccato sint atque turbentur
JOSH|6|19|quicquid autem auri et argenti fuerit et vasorum aeneorum ac ferri Domino consecretur repositum in thesauris eius
JOSH|6|20|igitur omni vociferante populo et clangentibus tubis postquam in aures multitudinis vox sonitusque increpuit muri ilico corruerunt et ascendit unusquisque per locum qui contra se erat ceperuntque civitatem
JOSH|6|21|et interfecerunt omnia quae erant in ea a viro usque ad mulierem ab infante usque ad senem boves quoque et oves et asinos in ore gladii percusserunt
JOSH|6|22|duobus autem viris qui exploratores missi fuerant dixit Iosue ingredimini domum mulieris meretricis et producite eam omniaque quae illius sunt sicut illi iuramento firmastis
JOSH|6|23|ingressique iuvenes eduxerunt Raab et parentes eius fratres quoque et cunctam supellectilem ac cognationem illius et extra castra Israhel manere fecerunt
JOSH|6|24|urbem autem et omnia quae in ea sunt succenderunt absque argento et auro et vasis aeneis ac ferro quae in aerarium Domini consecrarunt
JOSH|6|25|Raab vero meretricem et domum patris eius atque omnia quae habebat fecit Iosue vivere et habitaverunt in medio Israhel usque in praesentem diem eo quod absconderit nuntios quos miserat ut explorarent Hiericho in tempore illo inprecatus est Iosue dicens
JOSH|6|26|maledictus vir coram Domino qui suscitaverit et aedificaverit civitatem Hiericho in primogenito suo fundamenta illius iaciat et in novissimo liberorum ponat portas eius
JOSH|6|27|fuit ergo Dominus cum Iosue et nomen eius in omni terra vulgatum est
JOSH|7|1|filii autem Israhel praevaricati sunt mandatum et usurpaverunt de anathemate nam Achan filius Charmi filii Zabdi filii Zare de tribu Iuda tulit aliquid de anathemate iratusque est Dominus contra filios Israhel
JOSH|7|2|cumque mitteret Iosue de Hiericho viros contra Ahi quae est iuxta Bethaven ad orientalem plagam oppidi Bethel dixit eis ascendite et explorate terram qui praecepta conplentes exploraverunt Ahi
JOSH|7|3|et reversi dixerunt ei non ascendat omnis populus sed duo vel tria milia virorum pergant et deleant civitatem quare omnis populus frustra vexatur contra hostes paucissimos
JOSH|7|4|ascenderunt ergo tria milia pugnatores qui statim terga vertentes
JOSH|7|5|percussi sunt a viris urbis Ahi et corruerunt ex eis triginta et sex homines persecutique sunt eos adversarii de porta usque Sabarim et ceciderunt per prona fugientes pertimuitque cor populi et instar aquae liquefactum est
JOSH|7|6|Iosue vero scidit vestimenta sua et cecidit pronus in terram coram arca Domini usque ad vesperum tam ipse quam omnes senes Israhel miseruntque pulverem super capita sua
JOSH|7|7|et dixit Iosue heu Domine Deus quid voluisti transducere populum istum Iordanem fluvium ut traderes nos in manus Amorrei et perderes utinam ut coepimus mansissemus trans Iordanem
JOSH|7|8|mi Domine Deus quid dicam videns Israhelem hostibus suis terga vertentem
JOSH|7|9|audient Chananei et omnes habitatores terrae ac pariter conglobati circumdabunt nos atque delebunt nomen nostrum de terra et quid facies magno nomini tuo
JOSH|7|10|dixitque Dominus ad Iosue surge cur iaces pronus in terra
JOSH|7|11|peccavit Israhel et praevaricatus est pactum meum tuleruntque de anathemate et furati sunt atque mentiti et absconderunt inter vasa sua
JOSH|7|12|nec poterit Israhel stare ante hostes suos eosque fugiet quia pollutus est anathemate non ero ultra vobiscum donec conteratis eum qui huius sceleris reus est
JOSH|7|13|surge sanctifica populum et dic eis sanctificamini in crastinum haec enim dicit Dominus Deus Israhel anathema in medio tui est Israhel non poteris stare coram hostibus tuis donec deleatur ex te qui hoc contaminatus est scelere
JOSH|7|14|accedetisque mane singuli per tribus vestras et quamcumque tribum sors invenerit accedet per cognationes suas et cognatio per domos domusque per viros
JOSH|7|15|et quicumque ille in hoc facinore fuerit deprehensus conburetur igni cum omni substantia sua quoniam praevaricatus est pactum Domini et fecit nefas in Israhel
JOSH|7|16|surgens itaque Iosue mane adplicavit Israhel per tribus suas et inventa est tribus Iuda
JOSH|7|17|quae cum iuxta familias suas esset oblata inventa est familia Zarai illam quoque per viros offerens repperit Zabdi
JOSH|7|18|cuius domum in singulos dividens viros invenit Achan filium Charmi filii Zabdi filii Zare de tribu Iuda
JOSH|7|19|et ait ad Achan fili mi da gloriam Domino Deo Israhel et confitere atque indica mihi quid feceris ne abscondas
JOSH|7|20|responditque Achan Iosue et dixit ei vere ego peccavi Domino Deo Israhel et sic et sic feci
JOSH|7|21|vidi enim inter spolia pallium coccineum valde bonum et ducentos siclos argenti regulamque auream quinquaginta siclorum et concupiscens abstuli et abscondi in terra contra medium tabernaculi mei argentumque fossa humo operui
JOSH|7|22|misit ergo Iosue ministros qui currentes ad tabernaculum illius reppererunt cuncta abscondita in eodem loco et argentum simul
JOSH|7|23|auferentesque de tentorio tulerunt ea ad Iosue et ad omnes filios Israhel proieceruntque ante Dominum
JOSH|7|24|tollens itaque Iosue Achan filium Zare argentumque et pallium et auream regulam filiosque eius et filias boves et asinos et oves ipsumque tabernaculum et cunctam supellectilem et omnis Israhel cum eo duxerunt eos ad vallem Achor
JOSH|7|25|ubi dixit Iosue quia turbasti nos exturbet te Dominus in die hac lapidavitque eum omnis Israhel et cuncta quae illius erant igne consumpta sunt
JOSH|7|26|congregaverunt quoque super eum acervum magnum lapidum qui permanet usque in praesentem diem et aversus est furor Domini ab eis vocatumque est nomen loci illius vallis Achor usque hodie
JOSH|8|1|dixit autem Dominus ad Iosue ne timeas neque formides tolle tecum omnem multitudinem pugnatorum et consurgens ascende in oppidum Ahi ecce tradidi in manu tua regem eius et populum urbemque et terram
JOSH|8|2|faciesque urbi Ahi et regi eius sicut fecisti Hiericho et regi illius praedam vero et omnia animantia diripietis vobis pone insidias urbi post eam
JOSH|8|3|surrexitque Iosue et omnis exercitus bellatorum cum eo ut ascenderent in Ahi et electa triginta milia virorum fortium misit nocte
JOSH|8|4|praecepitque eis dicens ponite insidias post civitatem nec longius recedatis et eritis omnes parati
JOSH|8|5|ego autem et reliqua multitudo quae mecum est accedemus ex adverso contra urbem cumque exierint contra nos sicut ante fecimus fugiemus et terga vertemus
JOSH|8|6|donec persequentes ab urbe longius protrahantur putabunt enim fugere nos sicut prius
JOSH|8|7|nobis ergo fugientibus et illis sequentibus consurgetis de insidiis et vastabitis civitatem tradetque eam Dominus Deus vester in manus vestras
JOSH|8|8|cumque ceperitis succendite eam sic omnia facietis ut iussi
JOSH|8|9|dimisitque eos et perrexerunt ad insidiarum locum sederuntque inter Bethel et Ahi ad occidentalem plagam urbis Ahi Iosue autem nocte illa in medio mansit populi
JOSH|8|10|surgensque diluculo recensuit socios et ascendit cum senioribus in fronte exercitus vallatus auxilio pugnatorum
JOSH|8|11|cumque venissent et ascendissent ex adverso civitatis steterunt ad septentrionalem urbis plagam inter quam et eos vallis media erat
JOSH|8|12|quinque milia autem viros elegerat et posuerat in insidiis inter Bethaven et Ahi ex occidentali parte eiusdem civitatis
JOSH|8|13|omnis vero reliquus exercitus ad aquilonem aciem dirigebat ita ut novissimi multitudinis occidentalem plagam urbis adtingerent abiit ergo Iosue nocte illa et stetit in vallis medio
JOSH|8|14|quod cum vidisset rex Ahi festinavit mane et egressus est cum omni exercitu civitatis direxitque aciem contra desertum ignorans quod post tergum laterent insidiae
JOSH|8|15|Iosue vero et omnis Israhel cesserunt loco simulantes metum et fugientes per viam solitudinis
JOSH|8|16|at illi vociferantes pariter et se mutuo cohortantes persecuti sunt eos cumque recessissent a civitate
JOSH|8|17|et ne unus quidem in urbe Ahi et Bethel remansisset qui non persequeretur Israhel sicut eruperant aperta oppida relinquentes
JOSH|8|18|dixit Dominus ad Iosue leva clypeum qui in manu tua est contra urbem Ahi quoniam tibi tradam eam
JOSH|8|19|cumque elevasset clypeum ex adverso civitatis insidiae quae latebant surrexerunt confestim et pergentes ad civitatem ceperunt et succenderunt eam
JOSH|8|20|viri autem civitatis qui persequebantur Iosue respicientes et videntes fumum urbis ad caelum usque conscendere non potuerunt ultra huc illucque diffugere praesertim cum hii qui simulaverant fugam et tendebant ad solitudinem contra persequentes fortissime restitissent
JOSH|8|21|vidensque Iosue et omnis Israhel quod capta esset civitas et fumus urbis ascenderet reversus percussit viros Ahi
JOSH|8|22|siquidem et illi qui ceperant et succenderant civitatem egressi ex urbe contra suos medios hostium ferire coeperunt cum ergo ex utraque parte adversarii caederentur ita ut nullus de tanta multitudine salvaretur
JOSH|8|23|regem quoque urbis Ahi adprehendere viventem et obtulerunt Iosue
JOSH|8|24|igitur omnibus interfectis qui Israhelem ad deserta tendentem fuerant persecuti et in eodem loco gladio corruentibus reversi filii Israhel percusserunt civitatem
JOSH|8|25|erant autem qui in eo die conciderant a viro usque ad mulierem duodecim milia hominum omnes urbis Ahi
JOSH|8|26|Iosue vero non contraxit manum quam in sublime porrexerat tenens clypeum donec interficerentur omnes habitatores Ahi
JOSH|8|27|iumenta autem et praedam civitatis diviserunt sibi filii Israhel sicut praeceperat Dominus Iosue
JOSH|8|28|qui succendit urbem et fecit eam tumulum sempiternum
JOSH|8|29|regem quoque eius suspendit in patibulo usque ad vesperum et solis occasum praecepitque et deposuerunt cadaver eius de cruce proieceruntque in ipso introitu civitatis congesto super eum magno acervo lapidum qui permanet usque in praesentem diem
JOSH|8|30|tunc aedificavit Iosue altare Domino Deo Israhel in monte Hebal
JOSH|8|31|sicut praeceperat Moses famulus Domini filiis Israhel et scriptum est in volumine legis Mosi altare de lapidibus inpolitis quos ferrum non tetigit et obtulit super eo holocausta Domino immolavitque pacificas victimas
JOSH|8|32|et scripsit super lapides deuteronomium legis Mosi quod ille digesserat coram filiis Israhel
JOSH|8|33|omnis autem populus et maiores natu ducesque ac iudices stabant ex utraque parte arcae in conspectu sacerdotum qui portabant arcam foederis Domini ut advena ita et indigena media eorum pars iuxta montem Garizim et media iuxta montem Hebal sicut praeceperat Moses famulus Domini et primum quidem benedixit populo Israhel
JOSH|8|34|post haec legit omnia verba benedictionis et maledictionis et cuncta quae scripta erant in legis volumine
JOSH|8|35|nihil ex his quae Moses iusserat reliquit intactum sed universa replicavit coram omni multitudine Israhel mulieribus ac parvulis et advenis qui inter eos morabantur
JOSH|9|1|quibus auditis cuncti reges trans Iordanem qui versabantur in montanis et in campestribus in maritimis ac litore maris Magni hii quoque qui habitabant iuxta Libanum Hettheus et Amorreus et Chananeus Ferezeus et Eveus et Iebuseus
JOSH|9|2|congregati sunt pariter ut pugnarent contra Iosue et Israhel uno animo eademque sententia
JOSH|9|3|at hii qui habitabant in Gabaon audientes cuncta quae fecerat Iosue Hiericho et Ahi
JOSH|9|4|et callide cogitantes tulerunt sibi cibaria saccos veteres asinis inponentes et utres vinarios scissos atque consutos
JOSH|9|5|calciamentaque perantiqua quae ad indicium vetustatis pittaciis consuta erant induti veteribus vestimentis panes quoque quos portabant ob viaticum duri erant et in frusta comminuti
JOSH|9|6|perrexeruntque ad Iosue qui tunc morabatur in castris Galgalae et dixerunt ei atque omni simul Israheli de terra longinqua venimus pacem vobiscum facere cupientes responderuntque viri Israhel ad eos atque dixerunt
JOSH|9|7|ne forsitan in terra quae nobis sorte debetur habitetis et non possimus foedus inire vobiscum
JOSH|9|8|at illi ad Iosue servi inquiunt tui sumus quibus Iosue quinam ait estis et unde venistis
JOSH|9|9|responderunt de terra longinqua valde venerunt servi tui in nomine Domini Dei tui audivimus enim famam potentiae eius cuncta quae fecit in Aegypto
JOSH|9|10|et duobus Amorreorum regibus trans Iordanem Seon regi Esebon et Og regi Basan qui erat in Astharoth
JOSH|9|11|dixeruntque nobis seniores et omnes habitatores terrae nostrae tollite in manibus cibaria ob longissimam viam et occurrite eis ac dicite servi vestri sumus foedus inite nobiscum
JOSH|9|12|en panes quando egressi sumus de domibus nostris ut veniremus ad vos calidos sumpsimus nunc sicci facti sunt et vetustate nimia comminuti
JOSH|9|13|utres vini novos implevimus nunc rupti sunt et soluti vestes et calciamenta quibus induimur et quae habemus in pedibus ob longitudinem largioris viae trita sunt et paene consumpta
JOSH|9|14|susceperunt igitur de cibariis eorum et os Domini non interrogaverunt
JOSH|9|15|fecitque Iosue cum eis pacem et inito foedere pollicitus est quod non occiderentur principes quoque multitudinis iuraverunt eis
JOSH|9|16|post dies autem tres initi foederis audierunt quod in vicino habitarent et inter eos futuri essent
JOSH|9|17|moveruntque castra filii Israhel et venerunt in civitates eorum die tertio quarum haec vocabula sunt Gabaon et Caphira et Beroth et Cariathiarim
JOSH|9|18|et non percusserunt eos eo quod iurassent eis principes multitudinis in nomine Domini Dei Israhel murmuravit itaque omne vulgus contra principes
JOSH|9|19|qui responderunt eis iuravimus illis in nomine Domini Dei Israhel et idcirco non possumus eos contingere
JOSH|9|20|sed hoc faciemus eis reserventur quidem ut vivant ne contra nos ira Domini concitetur si peieraverimus
JOSH|9|21|sed sic vivant ut in usus universae multitudinis ligna caedant aquasque conportent quibus haec loquentibus
JOSH|9|22|vocavit Gabaonitas Iosue et dixit eis cur nos decipere fraude voluistis ut diceretis procul valde habitamus a vobis cum in medio nostri sitis
JOSH|9|23|itaque sub maledictione eritis et non deficiet de stirpe vestra ligna caedens aquasque conportans in domum Dei mei
JOSH|9|24|qui responderunt nuntiatum est nobis servis tuis quae promisisset Dominus Deus tuus Mosi servo suo ut traderet vobis omnem terram et disperderet cunctos habitatores eius timuimus igitur valde et providimus animabus nostris vestro terrore conpulsi et hoc consilium inivimus
JOSH|9|25|nunc autem in manu tua sumus quod tibi bonum et rectum videtur fac nobis
JOSH|9|26|fecit ergo Iosue ut dixerat et liberavit eos de manibus filiorum Israhel ut non occiderentur
JOSH|9|27|decrevitque in illo die esse eos in ministerium cuncti populi et altaris Domini caedentes ligna et aquas conportantes usque in praesens tempus in loco quem Dominus elegisset
JOSH|10|1|quae cum audisset Adonisedec rex Hierusalem quod scilicet cepisset Iosue Ahi et subvertisset eam sicut enim fecerat Hiericho et regi eius sic fecit Ahi et regi illius et quod transfugissent Gabaonitae ad Israhel et essent foederati eorum
JOSH|10|2|timuit valde urbs enim magna erat Gabaon et una regalium civitatum et maior oppido Ahi omnesque bellatores eius fortissimi
JOSH|10|3|misit ergo Adonisedec rex Hierusalem ad Oham regem Hebron et ad Pharam regem Hieremoth ad Iaphie quoque regem Lachis et ad Dabir regem Eglon dicens
JOSH|10|4|ascendite ad me et ferte praesidium ut expugnemus Gabaon quare transfugerit ad Iosue et filios Israhel
JOSH|10|5|congregati igitur ascenderunt quinque reges Amorreorum rex Hierusalem rex Hebron rex Hieremoth rex Lachis rex Eglon simul cum exercitibus suis et castrametati sunt circa Gabaon obpugnantes eam
JOSH|10|6|habitatores autem Gabaon urbis obsessae miserunt ad Iosue qui tunc morabatur in castris apud Galgalam et dixerunt ei ne retrahas manus tuas ab auxilio servorum tuorum ascende cito et libera nos ferque praesidium convenerunt enim adversum nos omnes reges Amorreorum qui habitant in montanis
JOSH|10|7|ascenditque Iosue de Galgalis et omnis exercitus bellatorum cum eo viri fortissimi
JOSH|10|8|dixitque Dominus ad Iosue ne timeas eos in manus enim tuas tradidi illos nullus tibi ex eis resistere poterit
JOSH|10|9|inruit itaque Iosue super eos repente tota ascendens nocte de Galgalis
JOSH|10|10|et conturbavit eos Dominus a facie Israhel contrivitque plaga magna in Gabaon ac persecutus est per viam ascensus Bethoron et percussit usque Azeca et Maceda
JOSH|10|11|cumque fugerent filios Israhel et essent in descensu Bethoron Dominus misit super eos lapides magnos de caelo usque Azeca et mortui sunt multo plures lapidibus grandinis quam quos gladio percusserant filii Israhel
JOSH|10|12|tunc locutus est Iosue Domino in die qua tradidit Amorreum in conspectu filiorum Israhel dixitque coram eis sol contra Gabaon ne movearis et luna contra vallem Ahialon
JOSH|10|13|steteruntque sol et luna donec ulcisceretur se gens de inimicis suis nonne scriptum est hoc in libro Iustorum stetit itaque sol in medio caeli et non festinavit occumbere spatio unius diei
JOSH|10|14|non fuit ante et postea tam longa dies oboediente Domino voci hominis et pugnante pro Israhel
JOSH|10|15|reversusque est Iosue cum omni Israhel in castra Galgalae
JOSH|10|16|fugerant enim quinque reges et se absconderant in spelunca urbis Maceda
JOSH|10|17|nuntiatumque est Iosue quod inventi essent quinque reges latentes in spelunca Maceda
JOSH|10|18|qui praecepit sociis et ait volvite saxa ingentia ad os speluncae et ponite viros industrios qui clausos custodiant
JOSH|10|19|vos autem nolite stare sed persequimini hostes et extremos quosque fugientium caedite ne dimittatis eos urbium suarum intrare praesidia quos tradidit Dominus Deus in manus vestras
JOSH|10|20|caesis igitur adversariis plaga magna et usque ad internicionem paene consumptis hii qui Israhel effugere potuerunt ingressi sunt civitates munitas
JOSH|10|21|reversusque est omnis exercitus ad Iosue in Maceda ubi tunc erant castra sani et integro numero nullusque contra filios Israhel muttire ausus est
JOSH|10|22|praecepitque Iosue dicens aperite os speluncae et producite ad me quinque reges qui in ea latitant
JOSH|10|23|fecerunt ministri ut sibi fuerat imperatum et eduxerunt ad eum quinque reges de spelunca regem Hierusalem regem Hebron regem Hieremoth regem Lachis regem Eglon
JOSH|10|24|cumque educti essent ad eum vocavit omnes viros Israhel et ait ad principes exercitus qui secum erant ite et ponite pedes super colla regum istorum qui cum perrexissent et subiectorum pedibus colla calcarent
JOSH|10|25|rursum ait ad eos nolite timere nec paveatis confortamini et estote robusti sic enim faciet Dominus cunctis hostibus vestris adversum quos dimicatis
JOSH|10|26|percussitque Iosue et interfecit eos atque suspendit super quinque stipites fueruntque suspensi usque ad vesperum
JOSH|10|27|cumque occumberet sol praecepit sociis ut deponerent eos de patibulis qui depositos proiecerunt in speluncam in qua latuerant et posuerunt super os eius saxa ingentia quae permanent usque in praesens
JOSH|10|28|eodem die Macedam quoque cepit Iosue et percussit in ore gladii regemque illius interfecit et omnes habitatores eius non dimisit in ea saltim parvas reliquias fecitque regi Maceda sicut fecerat regi Hiericho
JOSH|10|29|transivit cum omni Israhel de Maceda in Lebna et pugnabat contra eam
JOSH|10|30|quam tradidit Dominus cum rege suo in manu Israhel percusseruntque urbem in ore gladii et omnes habitatores eius non dimiserunt in ea ullas reliquias feceruntque regi Lebna sicut fecerant regi Hiericho
JOSH|10|31|de Lebna transivit in Lachis et exercitu per gyrum disposito obpugnabat eam
JOSH|10|32|tradiditque Dominus Lachis in manu Israhel et cepit eam die altero atque percussit in ore gladii omnemque animam quae fuerat in ea sicut fecerat Lebna
JOSH|10|33|eo tempore ascendit Hiram rex Gazer ut auxiliaretur Lachis quem percussit Iosue cum omni populo eius usque ad internicionem
JOSH|10|34|transivitque de Lachis in Eglon et circumdedit
JOSH|10|35|atque expugnavit eam eadem die percussitque in ore gladii omnes animas quae erant in ea iuxta omnia quae fecerat Lachis
JOSH|10|36|ascendit quoque cum omni Israhele de Eglon in Hebron et pugnavit contra eam
JOSH|10|37|cepitque et percussit in ore gladii regem quoque eius et omnia oppida regionis illius universasque animas quae in ea fuerant commoratae non reliquit in ea ullas reliquias sicut fecerat Eglon sic fecit et Hebron cuncta quae in ea repperit consumens gladio
JOSH|10|38|inde reversus in Dabir
JOSH|10|39|cepit eam atque vastavit
JOSH|10|40|regem quoque eius et omnia per circuitum oppida percussit in ore gladii non dimisit in ea ullas reliquias sicut fecerat Hebron et Lebna et regibus earum sic fecit Dabir et regi illius
JOSH|10|41|percussit itaque Iosue omnem terram montanam et meridianam atque campestrem et Asedoth cum regibus suis non dimisit in ea ullas reliquias sed omne quod spirare poterat interfecit sicut praeceperat ei Dominus Deus Israhel
JOSH|10|42|a Cadesbarne usque Gazam omnem terram Gosen usque Gabaon
JOSH|10|43|universos reges et regiones eorum uno cepit impetu atque vastavit Dominus enim Deus Israhel pugnabat pro eo
JOSH|10|44|reversusque est cum omni Israhele ad locum castrorum in Galgala
JOSH|11|1|quae cum audisset Iabin rex Asor misit ad Iobab regem Madon et ad regem Someron atque ad regem Acsaph
JOSH|11|2|ad reges quoque aquilonis qui habitabant in montanis et in planitie contra meridiem Cheneroth in campestribus quoque et in regionibus Dor iuxta mare
JOSH|11|3|Chananeumque ab oriente et occidente et Amorreum atque Hettheum ac Ferezeum et Iebuseum in montanis Eveum quoque qui habitabat ad radices Hermon in terra Masphe
JOSH|11|4|egressique sunt omnes cum turmis suis populus multus nimis sicut harena quae est in litore maris equi quoque et currus inmensae multitudinis
JOSH|11|5|conveneruntque omnes reges isti in unum ad aquas Merom ut pugnarent contra Israhel
JOSH|11|6|dixitque Dominus ad Iosue ne timeas eos cras enim hac eadem hora ego tradam omnes istos vulnerandos in conspectu Israhel equos eorum subnervabis et currus igne conbures
JOSH|11|7|venitque Iosue et omnis exercitus cum eo adversum illos ad aquas Merom subito et inruerunt super eos
JOSH|11|8|tradiditque illos Dominus in manu Israhel qui percusserunt eos et persecuti sunt usque ad Sidonem magnam et aquas Maserefoth campumque Masphe qui est ad orientalem illius partem ita percussit omnes ut nullas dimitteret ex eis reliquias
JOSH|11|9|fecit sicut praeceperat ei Dominus equos eorum subnervavit currusque conbusit
JOSH|11|10|reversusque statim cepit Asor et regem eius percussit gladio Asor enim antiquitus inter omnia regna haec principatum tenebat
JOSH|11|11|percussitque omnes animas quae ibidem morabantur non dimisit in ea ullas reliquias sed usque ad internicionem universa vastavit ipsamque urbem permisit incendio
JOSH|11|12|et omnes per circuitum civitates regesque earum cepit percussit atque delevit sicut praeceperat ei Moses famulus Domini
JOSH|11|13|absque urbibus quae erant in collibus et in tumulis sitae ceteras succendit Israhel unam tantum Asor munitissimam flamma consumpsit
JOSH|11|14|omnemque praedam istarum urbium ac iumenta diviserunt sibi filii Israhel cunctis hominibus interfectis
JOSH|11|15|sicut praeceperat Dominus Mosi servo suo ita praecepit Moses Iosue et ille universa conplevit non praeteriit de universis mandatis ne unum quidem verbum quod iusserat Dominus Mosi
JOSH|11|16|cepit itaque Iosue omnem terram montanam et meridianam terramque Gosen et planitiem et occidentalem plagam montemque Israhel et campestria eius
JOSH|11|17|et partem montis quae ascendit Seir usque Baalgad per planitiem Libani subter montem Hermon omnes reges eorum cepit percussit occidit
JOSH|11|18|multo tempore pugnavit Iosue contra reges istos
JOSH|11|19|non fuit civitas quae se non traderet filiis Israhel praeter Eveum qui habitabat in Gabaon omnes bellando cepit
JOSH|11|20|Domini enim sententiae fuerat ut indurarentur corda eorum et pugnarent contra Israhel et caderent et non mererentur ullam clementiam ac perirent sicut praeceperat Dominus Mosi
JOSH|11|21|in tempore illo venit Iosue et interfecit Enacim de montanis Hebron et Dabir et Anab et de omni monte Iuda et Israhel urbesque eorum delevit
JOSH|11|22|non reliquit ullum de stirpe Enacim in terra filiorum Israhel absque civitatibus Gaza et Geth et Azoto in quibus solis relicti sunt
JOSH|11|23|cepit ergo Iosue omnem terram sicut locutus est Dominus ad Mosen et tradidit eam in possessionem filiis Israhel secundum partes et tribus suas quievitque terra a proeliis
JOSH|12|1|hii sunt reges quos percusserunt filii Israhel et possederunt terram eorum trans Iordanem ad solis ortum a torrente Arnon usque ad montem Hermon et omnem orientalem plagam quae respicit solitudinem
JOSH|12|2|Seon rex Amorreorum qui habitavit in Esebon dominatus est ab Aroer quae sita est super ripam torrentis Arnon et mediae partis in valle dimidiique Galaad usque ad torrentem Iaboc qui est terminus filiorum Ammon
JOSH|12|3|et a solitudine usque ad mare Cheneroth contra orientem et usque ad mare Deserti quod est mare Salsissimum ad orientalem plagam per viam quae ducit Bethesimoth et ab australi parte quae subiacent Asedothphasga
JOSH|12|4|terminus Og regis Basan de reliquiis Rafaim qui habitavit in Astharoth et in Edrain et dominatus est in monte Hermon et in Salacha atque in universa Basan usque ad terminos
JOSH|12|5|Gesuri et Machathi et dimidiae partis Galaad terminos Seon regis Esebon
JOSH|12|6|Moses famulus Domini et filii Israhel percusserunt eos tradiditque terram eorum Moses in possessionem Rubenitis et Gadditis et dimidiae tribui Manasse
JOSH|12|7|hii sunt reges terrae quos percussit Iosue et filii Israhel trans Iordanem ad occidentalem plagam a Baalgad in campo Libani usque ad montem cuius pars ascendit in Seir tradiditque eam Iosue in possessionem tribubus Israhel singulis partes suas
JOSH|12|8|tam in montanis quam in planis atque campestribus in Aseroth et solitudine ac meridie Hettheus fuit et Amorreus Chananeus et Ferezeus Eveus et Iebuseus
JOSH|12|9|rex Hiericho unus rex Ahi quae est ex latere Bethel unus
JOSH|12|10|rex Hierusalem unus rex Hebron unus
JOSH|12|11|rex Hierimoth unus rex Lachis unus
JOSH|12|12|rex Eglon unus rex Gazer unus
JOSH|12|13|rex Dabir unus rex Gader unus
JOSH|12|14|rex Herma unus rex Hered unus
JOSH|12|15|rex Lebna unus rex Odollam unus
JOSH|12|16|rex Maceda unus rex Bethel unus
JOSH|12|17|rex Thaffua unus rex Afer unus
JOSH|12|18|rex Afec unus rex Saron unus
JOSH|12|19|rex Madon unus rex Asor unus
JOSH|12|20|rex Someron unus rex Acsaph unus
JOSH|12|21|rex Thenach unus rex Mageddo unus
JOSH|12|22|rex Cades unus rex Iachanaem Chermeli unus
JOSH|12|23|rex Dor et provinciae Dor unus rex gentium Galgal unus
JOSH|12|24|rex Thersa unus omnes reges triginta et unus
JOSH|13|1|Iosue senex provectaeque aetatis erat et dixit Dominus ad eum senuisti et longevus es terraque latissima derelicta est quae necdum est sorte divisa
JOSH|13|2|omnis videlicet Galilea Philisthim et universa Gesuri
JOSH|13|3|a fluvio turbido qui inrigat Aegyptum usque ad terminos Accaron contra aquilonem terra Chanaan quae in quinque regulos Philisthim dividitur Gazeos Azotios Ascalonitas Gettheos et Accaronitas
JOSH|13|4|ad meridiem vero sunt Evei omnis terra Chanaan et Maara Sidoniorum usque Afeca et terminos Amorrei
JOSH|13|5|eiusque confinia Libani quoque regio contra orientem a Baalgad sub monte Hermon donec ingrediaris Emath
JOSH|13|6|omnium qui habitant in monte a Libano usque ad aquas Masrefoth universique Sidonii ego sum qui delebo eos a facie filiorum Israhel veniat ergo in parte hereditatis Israhel sicut praecepi tibi
JOSH|13|7|et nunc divide terram in possessionem novem tribubus et dimidiae tribui Manasse
JOSH|13|8|cum qua Ruben et Gad possederunt terram quam tradidit eis Moses famulus Domini trans fluenta Iordanis ad orientalem plagam
JOSH|13|9|ab Aroer quae sita est in ripa torrentis Arnon et in vallis medio universaque campestria Medaba usque Dibon
JOSH|13|10|et cunctas civitates Seon regis Amorrei qui regnavit in Esebon usque ad terminos filiorum Ammon
JOSH|13|11|et Galaad ac terminum Gesuri et Machathi omnemque montem Hermon et universam Basan usque Saleca
JOSH|13|12|omne regnum Og in Basan qui regnavit in Astharoth et Edraim ipse fuit de reliquiis Rafaim percussitque eos Moses atque delevit
JOSH|13|13|nolueruntque disperdere filii Israhel Gesuri et Machathi et habitaverunt in medio Israhel usque in praesentem diem
JOSH|13|14|tribui autem Levi non dedit possessionem sed sacrificia et victimae Domini Dei Israhel ipsa est eius hereditas sicut locutus est illi
JOSH|13|15|dedit ergo Moses possessionem tribui filiorum Ruben iuxta cognationes suas
JOSH|13|16|fuitque terminus eorum ab Aroer quae sita est in ripa torrentis Arnon et in valle eiusdem torrentis media universam planitiem quae ducit Medaba
JOSH|13|17|et Esebon cunctosque viculos earum qui sunt in campestribus Dibon quoque et Bamothbaal et oppidum Baalmaon
JOSH|13|18|Iessa et Cedmoth et Mepheeth
JOSH|13|19|Cariathaim et Sebama et Sarathasar in monte convallis
JOSH|13|20|Bethpheor et Asedothphasga et Bethaisimoth
JOSH|13|21|omnes urbes campestres universaque regna Seon regis Amorrei qui regnavit in Esebon quem percussit Moses cum principibus Madian Eveum et Recem et Sur et Ur et Rabee duces Seon habitatores terrae
JOSH|13|22|et Balaam filium Beor ariolum occiderunt filii Israhel gladio cum ceteris interfectis
JOSH|13|23|factusque est terminus filiorum Ruben Iordanis fluvius haec est possessio Rubenitarum per cognationes suas urbium et viculorum
JOSH|13|24|deditque Moses tribui Gad et filiis eius per cognationes suas possessionem cuius haec divisio est
JOSH|13|25|terminus Iazer et omnes civitates Galaad dimidiamque partem terrae filiorum Ammon usque ad Aroer quae est contra Rabba
JOSH|13|26|et ab Esebon usque Ramoth Masphe et Batanim et a Manaim usque ad terminos Dabir
JOSH|13|27|in valle quoque Betharaam et Bethnemra et Soccoth et Saphon reliquam partem regni Seon regis Esebon huius quoque Iordanis finis est usque ad extremam partem maris Chenereth trans Iordanem ad orientalem plagam
JOSH|13|28|haec est possessio filiorum Gad per familias suas civitates et villae earum
JOSH|13|29|dedit et dimidiae tribui Manasse filiisque eius iuxta cognationes suas possessionem
JOSH|13|30|cuius hoc principium est a Manaim universam Basan et cuncta regna Og regis Basan omnesque vicos Air qui sunt in Basan sexaginta oppida
JOSH|13|31|et dimidiam partem Galaad Astharoth et Edrai urbes regni Og in Basan filiis Machir filii Manasse dimidiae parti filiorum Machir iuxta cognationes suas
JOSH|13|32|hanc possessionem divisit Moses in campestribus Moab trans Iordanem contra Hiericho ad orientalem plagam
JOSH|13|33|tribui autem Levi non dedit possessionem quoniam Dominus Deus Israhel ipse est possessio eius ut locutus est illi
JOSH|14|1|hoc est quod possederunt filii Israhel in terra Chanaan quam dederunt eis Eleazar sacerdos et Iosue filius Nun et principes familiarum per tribus Israhel
JOSH|14|2|sorte omnia dividentes sicut praeceperat Dominus in manu Mosi novem tribubus et dimidiae tribui
JOSH|14|3|duabus enim tribubus et dimidiae dederat Moses trans Iordanem possessionem absque Levitis qui nihil terrae acceperunt inter fratres suos
JOSH|14|4|sed in eorum successerant locum filii Ioseph in duas divisi tribus Manasse et Ephraim nec acceperunt Levitae aliam in terra partem nisi urbes ad habitandum et suburbana earum ad alenda iumenta et pecora sua
JOSH|14|5|sicut praecepit Dominus Mosi ita fecerunt filii Israhel et diviserunt terram
JOSH|14|6|accesserunt itaque filii Iuda ad Iosue in Galgala locutusque est ad eum Chaleb filius Iepphonne Cenezeus nosti quid locutus sit Dominus ad Mosen hominem Dei de me et te in Cadesbarne
JOSH|14|7|quadraginta annorum eram quando me misit Moses famulus Domini de Cadesbarne ut considerarem terram nuntiavique ei quod mihi verum videbatur
JOSH|14|8|fratres autem mei qui ascenderant mecum dissolverunt cor populi et nihilominus ego secutus sum Dominum Deum meum
JOSH|14|9|iuravitque Moses in die illo dicens terram quam calcavit pes tuus erit possessio tua et filiorum tuorum in aeternum quia secutus es Dominum Deum meum
JOSH|14|10|concessit ergo Dominus vitam mihi sicut pollicitus est usque in praesentem diem quadraginta et quinque anni sunt ex quo locutus est Dominus verbum istud ad Mosen quando ambulabat Israhel per solitudinem hodie octoginta quinque annorum sum
JOSH|14|11|sic valens ut eo valebam tempore quando ad explorandum missus sum illius in me temporis fortitudo usque hodie perseverat tam ad bellandum quam ad gradiendum
JOSH|14|12|da ergo mihi montem istum quem pollicitus est Dominus te quoque audiente in quo Enacim sunt et urbes magnae atque munitae si forte sit Dominus mecum et potuero delere eos sicut promisit mihi
JOSH|14|13|benedixitque ei Iosue et tradidit Hebron in possessionem
JOSH|14|14|atque ex eo fuit Hebron Chaleb filio Iepphonne Cenezeo usque in praesentem diem quia secutus est Dominum Deum Israhel
JOSH|14|15|nomen Hebron antea vocabatur Cariatharbe Adam maximus ibi inter Enacim situs est et terra cessavit a proeliis
JOSH|15|1|igitur sors filiorum Iudae per cognationes suas ista fuit a termino Edom desertum Sin contra meridiem et usque ad extremam partem australis plagae
JOSH|15|2|initium eius a summitate maris Salsissimi et a lingua eius quae respicit meridiem
JOSH|15|3|egrediturque contra ascensum Scorpionis et pertransit in Sina ascenditque in Cadesbarne et pervenit in Esrom ascendens Addara et circumiens Caricaa
JOSH|15|4|atque inde pertransiens in Asemona et perveniens ad torrentem Aegypti eruntque termini eius mare Magnum hic erit finis meridianae plagae
JOSH|15|5|ab oriente vero erit initium mare Salsissimum usque ad extrema Iordanis et ea quae respiciunt aquilonem a lingua maris usque ad eundem Iordanem fluvium
JOSH|15|6|ascenditque terminus in Bethagla et transit ab aquilone in Betharaba ascendens ad lapidem Boem filii Ruben
JOSH|15|7|et tendens usque ad terminos Debera de valle Achor contra aquilonem respiciens Galgala quae est ex adverso ascensionis Adommim ab australi parte torrentis transitque aquas quae vocantur fons Solis et erunt exitus eius ad fontem Rogel
JOSH|15|8|ascenditque per convallem filii Ennom ex latere Iebusei ad meridiem haec est Hierusalem et inde se erigens ad verticem montis qui est contra Gehennom ad occidentem in summitate vallis Rafaim contra aquilonem
JOSH|15|9|pertransitque a vertice montis usque ad fontem aquae Nepthoa et pervenit usque ad vicos montis Ephron inclinaturque in Bala quae est Cariathiarim id est urbs Silvarum
JOSH|15|10|et circuit de Bala contra occidentem usque ad montem Seir transitque iuxta latus montis Iarim ad aquilonem in Cheslon et descendit in Bethsames transitque in Thamna
JOSH|15|11|et pervenit contra aquilonem partis Accaron ex latere inclinaturque Sechrona et transit montem Baala pervenitque in Iebnehel et maris Magni contra occidentem fine concluditur
JOSH|15|12|hii sunt termini filiorum Iuda per circuitum in cognationibus suis
JOSH|15|13|Chaleb vero filio Iepphonne dedit partem in medio filiorum Iuda sicut praeceperat ei Dominus Cariatharbe patris Enach ipsa est Hebron
JOSH|15|14|delevitque ex ea Chaleb tres filios Enach Sesai et Ahiman et Tholmai de stirpe Enach
JOSH|15|15|atque inde conscendens venit ad habitatores Dabir quae prius vocabatur Cariathsepher id est civitas Litterarum
JOSH|15|16|dixitque Chaleb qui percusserit Cariathsepher et ceperit eam dabo illi Axam filiam meam uxorem
JOSH|15|17|cepitque eam Othonihel filius Cenez frater Chaleb iunior deditque ei Axam filiam suam uxorem
JOSH|15|18|quae cum pergerent simul suasit viro ut peteret a patre suo agrum suspiravitque ut sedebat in asino cui Chaleb quid habes inquit
JOSH|15|19|at illa respondit da mihi benedictionem terram australem et arentem dedisti mihi iunge et inriguam dedit itaque ei Chaleb inriguum superius et inferius
JOSH|15|20|haec est possessio tribus filiorum Iuda per cognationes suas
JOSH|15|21|erantque civitates ab extremis partibus filiorum Iuda iuxta terminos Edom a meridie Cabsehel et Eder et Iagur
JOSH|15|22|et Cina et Dimona Adeda
JOSH|15|23|et Cedes et Asor Iethnan
JOSH|15|24|Zif et Thelem Baloth
JOSH|15|25|et Asor nova et Cariothesrom haec est Asor
JOSH|15|26|Aman Same et Molada
JOSH|15|27|et Asergadda et Asemon Bethfeleth
JOSH|15|28|et Asersual et Bersabee et Baziothia
JOSH|15|29|Bala et Hiim Esem
JOSH|15|30|et Heltholad Exiil et Harma
JOSH|15|31|Siceleg et Medemena et Sensenna
JOSH|15|32|Lebaoth et Selim et Aenremmon omnes civitates viginti novem et villae earum
JOSH|15|33|in campestribus vero Esthaul et Saraa et Asena
JOSH|15|34|et Azanoe et Aengannim Thaffua et Aenaim
JOSH|15|35|et Hierimoth Adulam Soccho et Azeca
JOSH|15|36|et Saraim Adithaim et Gedera et Giderothaim urbes quattuordecim et villae earum
JOSH|15|37|Sanan et Adesa et Magdalgad
JOSH|15|38|Delean et Mesfa et Iecthel
JOSH|15|39|Lachis et Bascath et Aglon
JOSH|15|40|Thebbon et Lehemas et Chethlis
JOSH|15|41|et Gideroth Bethdagon et Neema et Maceda civitates sedecim et villae earum
JOSH|15|42|Labana et Aether et Asan
JOSH|15|43|Ieptha et Esna et Nesib
JOSH|15|44|Ceila et Achzib et Maresa civitates novem et villae earum
JOSH|15|45|Accaron cum vicis et villulis suis
JOSH|15|46|ab Accaron usque ad mare omnia quae vergunt ad Azotum et viculos eius
JOSH|15|47|Azotus cum vicis et villulis suis Gaza cum viculis et villulis suis usque ad torrentem Aegypti mare Magnum terminus eius
JOSH|15|48|et in monte Samir et Iether et Soccho
JOSH|15|49|et Edenna Cariathsenna haec est Dabir
JOSH|15|50|Anab et Isthemo et Anim
JOSH|15|51|Gosen et Olon et Gilo civitates undecim et villae earum
JOSH|15|52|Arab et Roma et Esaan
JOSH|15|53|Ianum et Bethafua et Afeca
JOSH|15|54|Ammatha et Cariatharbe haec est Hebron et Sior civitates novem et villae earum
JOSH|15|55|Maon et Chermel et Zif et Iotae
JOSH|15|56|Iezrehel et Iucadam et Zanoe
JOSH|15|57|Accaim Gebaa et Thamna civitates decem et villae earum
JOSH|15|58|Alul et Bethsur et Gedor
JOSH|15|59|Mareth et Bethanoth et Elthecen civitates sex et villae earum
JOSH|15|60|Cariathbaal haec est Cariathiarim urbs Silvarum et Arebba civitates duae et villae earum
JOSH|15|61|in deserto Betharaba Meddin et Schacha
JOSH|15|62|Anepsan et civitas Salis et Engaddi civitates sex et villae earum
JOSH|15|63|Iebuseum autem habitatorem Hierusalem non potuerunt filii Iuda delere habitavitque Iebuseus cum filiis Iuda in Hierusalem usque in praesentem diem
JOSH|16|1|cecidit quoque sors filiorum Ioseph ab Iordane contra Hiericho et aquas eius ab oriente solitudo quae ascendit de Hiericho ad montana Bethel
JOSH|16|2|et egreditur de Bethel Luzam transitque terminum Archiatharoth
JOSH|16|3|et descendit ad occidentem iuxta terminum Ieflethi usque ad terminos Bethoron inferioris et Gazer finiunturque regiones eius mari Magno
JOSH|16|4|possederuntque filii Ioseph Manasse et Ephraim
JOSH|16|5|et factus est terminus filiorum Ephraim per cognationes suas et possessio eorum contra orientem Atharothaddar usque Bethoron superiorem
JOSH|16|6|egrediunturque confinia in mare Machmethath vero aquilonem respicit et circuit terminus contra orientem in Thanathselo et pertransit ab oriente Ianoe
JOSH|16|7|descenditque de Ianoe in Atharoth et Noaratha et pervenit in Hiericho et egreditur ad Iordanem
JOSH|16|8|de Taffua pertransitque contra mare in valle Harundineti suntque egressus eius in mare Salsissimum haec est possessio tribus filiorum Ephraim per familias suas
JOSH|16|9|urbesque quae separatae sunt filiis Ephraim in medio possessionis filiorum Manasse et villae earum
JOSH|16|10|et non interfecerunt filii Ephraim Chananeum qui habitabat in Gazer habitavitque Chananeus in medio Ephraim usque in diem hanc tributarius
JOSH|17|1|cecidit autem sors tribui Manasse ipse est enim primogenitus Ioseph Machir primogenito Manasse patri Galaad qui fuit vir pugnator habuitque possessionem Galaad et Basan
JOSH|17|2|et reliquis filiorum Manasse iuxta familias suas filiis Abiezer et filiis Elech et filiis Esrihel et filiis Sechem et filiis Epher et filiis Semida isti sunt filii Manasse filii Ioseph mares per cognationes suas
JOSH|17|3|Salphaad vero filio Epher filii Galaad filii Machir filii Manasse non erant filii sed solae filiae quarum ista sunt nomina Maala et Noa Egla et Melcha et Thersa
JOSH|17|4|veneruntque in conspectu Eleazari sacerdotis et Iosue filii Nun et principum dicentes Dominus praecepit per manum Mosi ut daretur nobis possessio in medio fratrum nostrorum deditque eis iuxta imperium Domini possessionem in medio fratrum patris earum
JOSH|17|5|et ceciderunt funiculi Manasse decem absque terra Galaad et Basan trans Iordanem
JOSH|17|6|filiae enim Manasse possederunt hereditatem in medio filiorum eius terra autem Galaad cecidit in sortem filiorum Manasse qui reliqui erant
JOSH|17|7|fuitque terminus Manasse ab Aser Machmathath quae respicit Sychem et egreditur ad dextram iuxta habitatores fontis Taffuae
JOSH|17|8|etenim in sorte Manasse ceciderat terra Taffuae quae est iuxta terminos Manasse filiorum Ephraim
JOSH|17|9|descenditque terminus vallis Harundineti in meridiem torrentis civitatum Ephraim quae in medio sunt urbium Manasse terminus Manasse ab aquilone torrentis et exitus eius pergit ad mare
JOSH|17|10|ita ut ab austro sit possessio Ephraim et ab aquilone Manasse et utramque claudat mare et coniungantur sibi in tribu Aser ab aquilone et in tribu Isachar ab oriente
JOSH|17|11|fuitque hereditas Manasse in Isachar et in Aser Bethsan et viculi eius et Ieblaam cum villulis suis et habitatores Dor cum oppidis suis habitatores quoque Hendor cum villulis suis similiterque habitatores Thanach cum villulis suis et habitatores Mageddo cum viculis suis et tertia pars urbis Nofeth
JOSH|17|12|nec potuerunt filii Manasse has subvertere civitates sed coepit Chananeus habitare in terra ista
JOSH|17|13|postquam autem convaluerunt filii Israhel subiecerunt Chananeos et fecerunt sibi tributarios nec interfecerunt eos
JOSH|17|14|locutique sunt filii Ioseph ad Iosue atque dixerunt quare dedisti mihi possessionem sortis et funiculi unius cum sim tantae multitudinis et benedixerit mihi Dominus
JOSH|17|15|ad quos Iosue ait si populus multus es ascende in silvam et succide tibi spatia in terra Ferezei et Rafaim quia angusta est tibi possessio montis Ephraim
JOSH|17|16|cui responderunt filii Ioseph non poterimus ad montana conscendere cum ferreis curribus utantur Chananei qui habitant in terra campestri in qua sitae sunt Bethsan cum viculis suis et Iezrahel mediam possidens vallem
JOSH|17|17|dixitque Iosue ad domum Ioseph Ephraim et Manasse populus multus es et magnae fortitudinis non habebis sortem unam
JOSH|17|18|sed transibis ad montem et succides tibi atque purgabis ad habitandum spatia et poteris ultra procedere cum subverteris Chananeum quem dicis ferreos habere currus et esse fortissimum
JOSH|18|1|congregatique sunt omnes filii Israhel in Silo ibique fixerunt tabernaculum testimonii et fuit eis terra subiecta
JOSH|18|2|remanserant autem filiorum Israhel septem tribus quae necdum acceperant possessiones suas
JOSH|18|3|ad quos Iosue ait usquequo marcetis ignavia et non intratis ad possidendam terram quam Dominus Deus patrum vestrorum dedit vobis
JOSH|18|4|eligite de singulis tribubus ternos viros ut mittam eos et pergant atque circumeant terram et describant eam iuxta numerum uniuscuiusque multitudinis referantque ad me quod descripserint
JOSH|18|5|dividite vobis terram in septem partes Iudas sit in terminis suis ab australi plaga et domus Ioseph ab aquilone
JOSH|18|6|mediam inter hos terram in septem partes describite et huc venietis ad me ut coram Domino Deo vestro mittam vobis hic sortem
JOSH|18|7|quia non est inter vos pars Levitarum sed sacerdotium Domini est eorum hereditas Gad autem et Ruben et dimidia tribus Manasse iam acceperant possessiones suas trans Iordanem ad orientalem plagam quas dedit eis Moses famulus Domini
JOSH|18|8|cumque surrexissent viri ut pergerent ad describendam terram praecepit eis Iosue dicens circuite terram et describite eam ac revertimini ad me ut hic coram Domino Deo in Silo mittam vobis sortem
JOSH|18|9|itaque perrexerunt et lustrantes eam in septem partes diviserunt scribentes in volumine reversique sunt ad Iosue in castra Silo
JOSH|18|10|qui misit sortes coram Domino in Silo divisitque terram filiis Israhel in septem partes
JOSH|18|11|et ascendit sors prima filiorum Beniamin per familias suas ut possiderent terram inter filios Iuda et filios Ioseph
JOSH|18|12|fuitque terminus eorum contra aquilonem ab Iordane pergens iuxta latus Hiericho septentrionalis plagae et inde contra occidentem ad montana conscendens et perveniens in solitudinem Bethaven
JOSH|18|13|atque pertransiens iuxta Luzam ad meridiem ipsa est Bethel descenditque in Atharothaddar in montem qui est ad meridiem Bethoron inferioris
JOSH|18|14|et inclinatur circumiens contra mare a meridie montis qui respicit Bethoron contra africum suntque exitus eius in Cariathbaal quae vocatur et Cariathiarim urbem filiorum Iuda haec est plaga contra mare et occidentem
JOSH|18|15|a meridie autem ex parte Cariathiarim egreditur terminus contra mare et pervenit usque ad fontem aquarum Nepthoa
JOSH|18|16|descenditque in partem montis qui respicit vallem filiorum Ennom et est contra septentrionalem plagam in extrema parte vallis Rafaim descenditque Gehennom id est vallis Ennom iuxta latus Iebusei ad austrum et pervenit ad fontem Rogel
JOSH|18|17|transiens ad aquilonem et egrediens ad Aensemes id est fontem Solis
JOSH|18|18|et pertransit usque ad tumulos qui sunt e regione ascensus Adommim descenditque ad Abenboen id est lapidem Boen filii Ruben et pertransit ex latere aquilonis ad campestria descenditque in planitiem
JOSH|18|19|et praetergreditur contra aquilonem Bethagla suntque exitus eius contra linguam maris Salsissimi ab aquilone in fine Iordanis ad australem plagam
JOSH|18|20|qui est terminus illius ab oriente haec est possessio filiorum Beniamin per terminos suos in circuitu et familias singulas
JOSH|18|21|fueruntque civitates eius Hiericho et Bethagla et vallis Casis
JOSH|18|22|Betharaba et Semaraim et Bethel
JOSH|18|23|Avim et Affara et Ofra
JOSH|18|24|villa Emona et Ofni et Gabee civitates duodecim et villae earum
JOSH|18|25|Gabaon et Rama et Beroth
JOSH|18|26|et Mesfe Cafera et Ammosa
JOSH|18|27|et Recem Iarafel et Tharala
JOSH|18|28|et Sela Eleph et Iebus quae est Hierusalem Gabaath et Cariath civitates quattuordecim et villae earum haec est possessio filiorum Beniamin iuxta familias suas
JOSH|19|1|et egressa est sors secunda filiorum Symeon per cognationes suas fuitque hereditas
JOSH|19|2|eorum in medio possessionis filiorum Iuda Bersabee et Sabee et Molada
JOSH|19|3|et Asersual Bala et Asem
JOSH|19|4|et Heltholath Bethul Arma
JOSH|19|5|et Seceleg et Bethmarchaboth Asersusa
JOSH|19|6|et Bethlebaoth et Saroen civitates tredecim et villae earum
JOSH|19|7|Ahin et Remmon et Athar et Asan civitates quattuor et villae earum
JOSH|19|8|omnes viculi per circuitum urbium istarum usque ad Balaath Berrameth contra australem plagam haec est hereditas filiorum Symeon iuxta cognationes suas
JOSH|19|9|in funiculo et possessione filiorum Iuda quia maior erat et idcirco possederunt filii Symeon in medio hereditatis eorum
JOSH|19|10|cecidit quoque sors tertia filiorum Zabulon per cognationes suas et factus est terminus possessionis eorum usque Sarith
JOSH|19|11|ascenditque de mari et Medala ac pervenit in Debbaseth usque ad torrentem qui est contra Iecennam
JOSH|19|12|et revertitur de Sarith contra orientem in fines Ceseleththabor et egreditur ad Dabereth ascenditque contra Iafie
JOSH|19|13|et inde pertransit ad orientalem plagam Getthefer Etthacasin et egreditur in Remmon Ampthar et Noa
JOSH|19|14|et circuit ad aquilonem et Nathon suntque egressus eius vallis Iepthahel
JOSH|19|15|et Catheth et Nehalal et Semron et Iedala et Bethleem civitates duodecim et villae earum
JOSH|19|16|haec est hereditas tribus filiorum Zabulon per cognationes suas urbes et viculi earum
JOSH|19|17|Isachar egressa est sors quarta per cognationes suas
JOSH|19|18|fuitque eius hereditas Hiezrahel et Chasaloth et Sunem
JOSH|19|19|et Afaraim Seon et Anaarath
JOSH|19|20|et Rabbith et Cesion Abes
JOSH|19|21|et Rameth et Engannim et Enadda et Bethfeses
JOSH|19|22|et pervenit terminus usque Thabor et Seesima et Bethsemes eruntque exitus eius Iordanes civitates sedecim et villae earum
JOSH|19|23|haec est possessio filiorum Isachar per cognationes suas urbes et viculi earum
JOSH|19|24|cecidit sors quinta tribui filiorum Aser per cognationes suas
JOSH|19|25|fuitque terminus eorum Alchath et Oali et Beten et Axab
JOSH|19|26|Elmelech et Amaad et Messal et pervenit usque ad Carmelum maris et Siorlabanath
JOSH|19|27|ac revertitur contra orientem Bethdagon et pertransit usque Zabulon et vallem Iepthahel contra aquilonem in Bethemech et Neihel egrediturque ad levam Chabul
JOSH|19|28|et Achran et Roob et Amon et Canae usque ad Sidonem magnam
JOSH|19|29|revertiturque in Orma usque ad civitatem munitissimam Tyrum et usque Osa eruntque exitus eius in mare de funiculo Acziba
JOSH|19|30|et Amma et Afec et Roob civitates viginti duae et villae earum
JOSH|19|31|haec est possessio filiorum Aser per cognationes suas urbes et viculi earum
JOSH|19|32|filiorum Nepthalim sexta pars cecidit per familias suas
JOSH|19|33|et coepit terminus de Heleb et Helon in Sananim et Adami quae est Neceb et Iebnahel usque Lecum et egressus eorum usque ad Iordanem
JOSH|19|34|revertiturque terminus contra occidentem in Aznoththabor atque inde egreditur in Ucoca et pertransit in Zabulon contra meridiem et in Aser contra occidentem et in Iuda ad Iordanem contra ortum solis
JOSH|19|35|civitates munitissimae Aseddim Ser et Ammath et Recchath Chenereth
JOSH|19|36|et Edema et Arama Asor
JOSH|19|37|et Cedes et Edrai Nasor
JOSH|19|38|et Ieron et Magdalel Horem et Bethanath et Bethsemes civitates decem et novem et villae earum
JOSH|19|39|haec est possessio tribus filiorum Nepthali per cognationes suas urbes et viculi earum
JOSH|19|40|tribui filiorum Dan per familias suas egressa est sors septima
JOSH|19|41|et fuit terminus possessionis eius Saraa et Esthaol et Ahirsemes id est civitas Solis
JOSH|19|42|Selebin et Ahialon et Iethela
JOSH|19|43|Helon et Themna et Acron
JOSH|19|44|Helthecen et Gebthon et Baalath
JOSH|19|45|Iud et Benebarach et Gethremmon
JOSH|19|46|aquae Hiercon et Areccon cum termino qui respicit Ioppen
JOSH|19|47|et ipso fine concluditur ascenderuntque filii Dan et pugnaverunt contra Lesem ceperuntque eam et percusserunt in ore gladii ac possederunt et habitaverunt in ea vocantes nomen eius Lesemdan ex nomine Dan patris sui
JOSH|19|48|haec est possessio tribus filiorum Dan per cognationes suas urbes et viculi earum
JOSH|19|49|cumque conplesset terram sorte dividere singulis per tribus suas dederunt filii Israhel possessionem Iosue filio Nun in medio sui
JOSH|19|50|iuxta praeceptum Domini urbem quam postulavit Thamnathseraa in monte Ephraim et aedificavit civitatem habitavitque in ea
JOSH|19|51|hae sunt possessiones quas sorte diviserunt Eleazar sacerdos et Iosue filius Nun et principes familiarum ac tribuum filiorum Israhel in Silo coram Domino ad ostium tabernaculi testimonii partitique sunt terram
JOSH|20|1|et locutus est Dominus ad Iosue dicens loquere filiis Israhel et dic eis
JOSH|20|2|separate urbes fugitivorum de quibus locutus sum ad vos per manum Mosi
JOSH|20|3|ut confugiat ad eas quicumque animam percusserit nescius et possit evadere iram proximi qui ultor est sanguinis
JOSH|20|4|cum ad unam harum confugerit civitatum stabitque ante portam civitatis et loquetur senioribus urbis illius ea quae se conprobent innocentem sicque suscipient eum et dabunt ei locum ad habitandum
JOSH|20|5|cumque ultor sanguinis eum fuerit persecutus non tradent in manus eius quia ignorans percussit proximum eius nec ante biduum triduumve eius probatur inimicus
JOSH|20|6|et habitabit in civitate illa donec stet ante iudicium causam reddens facti sui et moriatur sacerdos magnus qui fuerit in illo tempore tunc revertetur homicida et ingredietur civitatem et domum suam de qua fugerat
JOSH|20|7|decreveruntque Cedes in Galilea montis Nepthali et Sychem in monte Ephraim et Cariatharbe ipsa est Hebron in monte Iuda
JOSH|20|8|et trans Iordanem contra orientalem plagam Hiericho statuerunt Bosor quae sita est in campestri solitudine de tribu Ruben et Ramoth in Galaad de tribu Gad et Gaulon in Basan de tribu Manasse
JOSH|20|9|hae civitates constitutae sunt cunctis filiis Israhel et advenis qui habitant inter eos ut fugeret ad eas qui animam nescius percussisset et non moreretur in manu proximi effusum sanguinem vindicare cupientis donec staret ante populum expositurus causam suam
JOSH|21|1|accesseruntque principes familiarum Levi ad Eleazar sacerdotem et Iosue filium Nun et ad duces cognationum per singulas tribus filiorum Israhel
JOSH|21|2|locutique sunt ad eos in Silo terrae Chanaan atque dixerunt Dominus praecepit per manum Mosi ut darentur nobis urbes ad habitandum et suburbana earum ad alenda iumenta
JOSH|21|3|dederuntque filii Israhel de possessionibus suis iuxta imperium Domini civitates et suburbana earum
JOSH|21|4|egressaque est sors in familiam Caath filiorum Aaron sacerdotis de tribubus Iuda et Symeon et Beniamin civitates tredecim
JOSH|21|5|et reliquis filiorum Caath id est Levitis qui superflui erant de tribubus Ephraim et Dan et dimidia tribu Manasse civitates decem
JOSH|21|6|porro filiis Gerson egressa est sors ut acciperent de tribubus Isachar et Aser et Nepthalim dimidiaque tribu Manasse in Basan civitates numero tredecim
JOSH|21|7|et filiis Merari per cognationes suas de tribubus Ruben et Gad et Zabulon urbes duodecim
JOSH|21|8|dederuntque filii Israhel Levitis civitates et suburbana earum sicut praecepit Dominus per manum Mosi singulis sorte tribuentes
JOSH|21|9|de tribubus filiorum Iuda et Symeon dedit Iosue civitates quarum ista sunt nomina
JOSH|21|10|filiis Aaron per familias Caath levitici generis prima enim sors illis egressa est
JOSH|21|11|Cariatharbe patris Enach quae vocatur Hebron in monte Iuda et suburbana eius per circuitum
JOSH|21|12|agros vero et villas eius dederat Chaleb filio Iepphonne ad possidendum
JOSH|21|13|dedit ergo filiis Aaron sacerdotis Hebron confugii civitatem ac suburbana eius et Lebnam cum suburbanis suis
JOSH|21|14|et Iether et Isthimon
JOSH|21|15|et Helon Dabir
JOSH|21|16|et Ahin et Iethan et Bethsemes cum suburbanis suis civitates novem de tribubus ut dictum est duabus
JOSH|21|17|de tribu autem filiorum Beniamin Gabaon et Gabee
JOSH|21|18|et Anathoth et Almon cum suburbanis suis civitates quattuor
JOSH|21|19|omnes simul civitates filiorum Aaron sacerdotis tredecim cum suburbanis suis
JOSH|21|20|reliquis vero per familias filiorum Caath levitici generis haec est data possessio
JOSH|21|21|de tribu Ephraim urbs confugii Sychem cum suburbanis suis in monte Ephraim et Gazer
JOSH|21|22|et Cebsain et Bethoron cum suburbanis suis civitates quattuor
JOSH|21|23|de tribu quoque Dan Elthece et Gebbethon
JOSH|21|24|et Ahialon et Gethremmon cum suburbanis suis civitates quattuor
JOSH|21|25|porro de dimidia tribu Manasse Thanach et Gethremmon cum suburbanis suis civitates duae
JOSH|21|26|omnes civitates decem et suburbana earum datae sunt filiis Caath inferioris gradus
JOSH|21|27|filiis quoque Gerson levitici generis dedit de dimidia tribu Manasse confugii civitatem Gaulon in Basan et Bosram cum suburbanis suis civitates duas
JOSH|21|28|porro de tribu Isachar Cesion et Dabereth
JOSH|21|29|et Iaramoth et Engannim cum suburbanis suis civitates quattuor
JOSH|21|30|de tribu autem Aser Masal et Abdon
JOSH|21|31|et Elacoth et Roob cum suburbanis suis civitates quattuor
JOSH|21|32|de tribu quoque Nepthali civitatem confugii Cedes in Galilea et Ammothdor et Charthan cum suburbanis suis civitates tres
JOSH|21|33|omnes urbes familiarum Gerson tredecim cum suburbanis suis
JOSH|21|34|filiis autem Merari Levitis inferioris gradus per familias suas data est de tribu Zabulon Iechenam et Chartha
JOSH|21|35|et Damna et Nalol civitates quattuor cum suburbanis suis
JOSH|21|36|de tribu quoque Ruben ciuitates confugii Bosor in solitudine et Cedson et Misor et Ocho ciuitates quattuor cum suburbanis suis]
JOSH|21|37|et de tribu Gad civitates confugii Ramoth in Galaad et Manaim et Esebon et Iazer civitates quattuor cum suburbanis suis
JOSH|21|38|omnes urbes filiorum Merari per familias et cognationes suas duodecim
JOSH|21|39|itaque universae civitates Levitarum in medio possessionis filiorum Israhel fuerunt quadraginta octo
JOSH|21|40|cum suburbanis suis singulae per familias distributae
JOSH|21|41|deditque Dominus Israheli omnem terram quam traditurum se patribus eorum iuraverat et possederunt illam atque habitaverunt in ea
JOSH|21|42|dataque est ab eo pax in omnes per circuitum nationes nullusque eis hostium resistere ausus est sed cuncti in eorum dicionem redacti sunt
JOSH|21|43|ne unum quidem verbum quod illis praestaturum se esse promiserat irritum fuit sed rebus expleta sunt omnia
JOSH|22|1|eodem tempore vocavit Iosue Rubenitas et Gadditas et dimidiam tribum Manasse
JOSH|22|2|dixitque ad eos fecistis omnia quae vobis praecepit Moses famulus Domini mihi quoque in omnibus oboedistis
JOSH|22|3|nec reliquistis fratres vestros longo tempore usque in praesentem diem custodientes imperium Domini Dei vestri
JOSH|22|4|quia igitur dedit Dominus Deus vester fratribus vestris quietem ac pacem sicut pollicitus est revertimini et ite in tabernacula vestra et in terram possessionis quam tradidit vobis Moses famulus Domini trans Iordanem
JOSH|22|5|ita dumtaxat ut custodiatis adtente et opere conpleatis mandatum et legem quam praecepit vobis Moses servus Domini ut diligatis Dominum Deum vestrum et ambuletis in omnibus viis eius et observetis mandata illius adhereatisque ei ac serviatis in omni corde et in omni anima vestra
JOSH|22|6|benedixitque eis Iosue et dimisit eos qui reversi sunt in tabernacula sua
JOSH|22|7|tribui autem Manasse mediae possessionem Moses dederat in Basan et idcirco mediae quae superfuit dedit Iosue sortem inter ceteros fratres suos trans Iordanem ad occidentalem eius plagam cumque dimitteret eos in tabernacula sua et benedixisset illis
JOSH|22|8|dixit ad eos in multa substantia atque divitiis revertimini ad sedes vestras cum argento et auro aere ac ferro et veste multiplici dividite praedam hostium cum fratribus vestris
JOSH|22|9|reversique sunt et abierunt filii Ruben et filii Gad et dimidia tribus Manasse a filiis Israhel de Silo quae sita est in Chanaan ut intrarent Galaad terram possessionis suae quam obtinuerant iuxta imperium Domini in manu Mosi
JOSH|22|10|cumque venissent ad tumulos Iordanis in terra Chanaan aedificaverunt iuxta Iordanem altare infinitae magnitudinis
JOSH|22|11|quod cum audissent filii Israhel et ad eos certi nuntii detulissent aedificasse filios Ruben et Gad et dimidiae tribus Manasse altare in terra Chanaan super Iordanis tumulos contra filios Israhel
JOSH|22|12|convenerunt omnes in Silo ut ascenderent et dimicarent contra eos
JOSH|22|13|et interim miserunt ad illos in terram Galaad Finees filium Eleazar sacerdotem
JOSH|22|14|et decem principes cum eo singulos de tribubus singulis
JOSH|22|15|qui venerunt ad filios Ruben et Gad et dimidiae tribus Manasse in terram Galaad dixeruntque ad eos
JOSH|22|16|haec mandat omnis populus Domini quae est ista transgressio cur reliquistis Dominum Deum Israhel aedificantes altare sacrilegum et a cultu illius recedentes
JOSH|22|17|an parum vobis est quod peccastis in Beelphegor et usque in praesentem diem macula huius sceleris in nobis permanet multique de populo corruerunt
JOSH|22|18|et vos hodie reliquistis Dominum et cras in universum Israhel eius ira desaeviet
JOSH|22|19|quod si putatis inmundam esse terram possessionis vestrae transite ad terram in qua tabernaculum Domini est et habitate inter nos tantum ut a Domino et a nostro consortio non recedatis aedificato altari praeter altare Domini Dei vestri
JOSH|22|20|nonne Achan filius Zare praeteriit mandatum Domini et super omnem populum Israhel ira eius incubuit et ille erat unus homo atque utinam solus perisset in scelere suo
JOSH|22|21|responderuntque filii Ruben et Gad et dimidiae tribus Manasse principibus legationis Israhel
JOSH|22|22|fortissimus Deus Dominus fortissimus Deus Dominus ipse novit et Israhel simul intelleget si praevaricationis animo hoc altare construximus non custodiat nos sed puniat in praesenti
JOSH|22|23|et si ea mente fecimus ut holocausta et sacrificium et pacificas victimas super eo inponeremus ipse quaerat et iudicet
JOSH|22|24|et non ea magis cogitatione atque tractatu ut diceremus cras dicent filii vestri filiis nostris quid vobis et Domino Deo Israhel
JOSH|22|25|terminum posuit Dominus inter nos et vos o filii Ruben et filii Gad Iordanem fluvium et idcirco partem non habetis in Domino et per hanc occasionem avertent filii vestri filios nostros a timore Domini putavimus itaque melius
JOSH|22|26|et diximus extruamus nobis altare non in holocausta neque ad victimas offerendas
JOSH|22|27|sed in testimonium inter nos et vos et subolem nostram vestramque progeniem ut serviamus Domino et iuris nostri sit offerre holocausta et victimas et pacificas hostias et nequaquam dicant cras filii vestri filiis nostris non est vobis pars in Domino
JOSH|22|28|quod si voluerint dicere respondebunt eis ecce altare Domini quod fecerunt patres nostri non in holocausta neque in sacrificium sed in testimonium vestrum ac nostrum
JOSH|22|29|absit a nobis hoc scelus ut recedamus a Domino et eius vestigia relinquamus extructo altari ad holocausta et sacrificia et victimas offerendas praeter altare Domini Dei nostri quod extructum est ante tabernaculum eius
JOSH|22|30|quibus auditis Finees sacerdos et principes legationis Israhel qui erant cum eo placati sunt et verba filiorum Ruben et Gad et dimidiae tribus Manasse libentissime susceperunt
JOSH|22|31|dixitque Finees filius Eleazari sacerdos ad eos nunc scimus quod nobiscum sit Dominus quoniam alieni estis a praevaricatione hac et liberastis filios Israhel de manu Domini
JOSH|22|32|reversusque est cum principibus a filiis Ruben et Gad de terra Galaad finium Chanaan ad filios Israhel et rettulit eis
JOSH|22|33|placuitque sermo cunctis audientibus et laudaverunt Deum filii Israhel et nequaquam ultra dixerunt ut ascenderent contra eos atque pugnarent et delerent terram possessionis eorum
JOSH|22|34|vocaveruntque filii Ruben et filii Gad altare quod extruxerant Testimonium nostrum quod Dominus ipse sit Deus
JOSH|23|1|evoluto autem multo tempore postquam pacem Dominus dederat Israheli subiectis in gyro nationibus universis et Iosue iam longevo et persenilis aetatis
JOSH|23|2|vocavit Iosue omnem Israhelem maioresque natu et principes ac duces et magistros dixitque ad eos ego senui et progressioris aetatis sum
JOSH|23|3|vosque cernitis omnia quae fecerit Dominus Deus vester cunctis per circuitum nationibus quomodo pro vobis ipse pugnaverit
JOSH|23|4|et nunc quia vobis sorte divisit omnem terram ab orientali parte Iordanis usque ad mare Magnum multaeque adhuc supersunt nationes
JOSH|23|5|Dominus Deus vester disperdet eas et auferet a facie vestra et possidebitis terram sicut vobis pollicitus est
JOSH|23|6|tantum confortamini et estote solliciti ut custodiatis cuncta quae scripta sunt in volumine legis Mosi et non declinetis ab eis nec ad dextram nec ad sinistram
JOSH|23|7|ne postquam intraveritis ad gentes quae inter vos futurae sunt iuretis in nomine deorum earum et serviatis eis et adoretis illos
JOSH|23|8|sed adhereatis Domino Deo vestro quod fecistis usque in diem hanc
JOSH|23|9|et tunc auferet Dominus in conspectu vestro gentes magnas et robustissimas et nullus vobis resistere poterit
JOSH|23|10|unus e vobis persequetur hostium mille viros quia Dominus Deus vester pro vobis ipse pugnabit sicut pollicitus est
JOSH|23|11|hoc tantum diligentissime praecavete ut diligatis Dominum Deum vestrum
JOSH|23|12|quod si volueritis gentium harum quae inter vos habitant erroribus adherere et cum eis miscere conubia atque amicitias copulare
JOSH|23|13|iam nunc scitote quod Dominus Deus vester non eas deleat ante faciem vestram sed sint vobis in foveam ac laqueum et offendiculum ex latere vestro et sudes in oculis vestris donec vos auferat atque disperdat de terra hac optima quam tradidit vobis
JOSH|23|14|en ego hodie ingrediar viam universae terrae et toto animo cognoscetis quod de omnibus verbis quae se Dominus praestaturum nobis esse pollicitus est unum non praeterierit in cassum
JOSH|23|15|sicut ergo implevit opere quod promisit et prospera cuncta venerunt sic adducet super vos quicquid malorum comminatus est donec vos auferat atque disperdat de terra hac optima quam tradidit vobis
JOSH|23|16|eo quod praeterieritis pactum Domini Dei vestri quod pepigit vobiscum et servieritis diis alienis et adoraveritis eos cito atque velociter consurget in vos furor Domini et auferemini de terra hac optima quam tradidit vobis
JOSH|24|1|congregavitque Iosue omnes tribus Israhel in Sychem et vocavit maiores natu ac principes et iudices et magistros steteruntque in conspectu Domini
JOSH|24|2|et ad populum sic locutus est haec dicit Dominus Deus Israhel trans fluvium habitaverunt patres vestri ab initio Thare pater Abraham et Nahor servieruntque diis alienis
JOSH|24|3|tuli ergo patrem vestrum Abraham de Mesopotamiae finibus et adduxi eum in terram Chanaan multiplicavique semen eius
JOSH|24|4|et dedi ei Isaac illique rursum dedi Iacob et Esau e quibus Esau dedi montem Seir ad possidendum Iacob vero et filii eius descenderunt in Aegyptum
JOSH|24|5|misique Mosen et Aaron et percussi Aegyptum multis signis atque portentis
JOSH|24|6|eduxique vos et patres vestros de Aegypto et venistis ad mare persecutique sunt Aegyptii patres vestros cum curribus et equitatu usque ad mare Rubrum
JOSH|24|7|clamaverunt autem ad Dominum filii Israhel qui posuit tenebras inter vos et Aegyptios et adduxit super eos mare et operuit illos viderunt oculi vestri cuncta quae in Aegypto fecerim et habitastis in solitudine multo tempore
JOSH|24|8|et introduxi vos ad terram Amorrei qui habitabat trans Iordanem cumque pugnarent contra vos tradidi eos in manus vestras et possedistis terram eorum atque interfecistis illos
JOSH|24|9|surrexit autem Balac filius Sepphor rex Moab et pugnavit contra Israhelem misitque et vocavit Balaam filium Beor ut malediceret vobis
JOSH|24|10|et ego nolui audire eum sed e contrario per illum benedixi vobis et liberavi vos de manu eius
JOSH|24|11|transistisque Iordanem et venistis ad Hiericho pugnaveruntque contra vos viri civitatis eius Amorreus et Ferezeus et Chananeus et Hettheus et Gergeseus et Eveus et Iebuseus et tradidi illos in manus vestras
JOSH|24|12|misique ante vos crabrones et eieci eos de locis suis duos reges Amorreorum non in gladio et arcu tuo
JOSH|24|13|dedique vobis terram in qua non laborastis et urbes quas non aedificastis ut habitaretis in eis vineas et oliveta quae non plantastis
JOSH|24|14|nunc ergo timete Dominum et servite ei perfecto corde atque verissimo et auferte deos quibus servierunt patres vestri in Mesopotamia et in Aegypto ac servite Domino
JOSH|24|15|sin autem malum vobis videtur ut Domino serviatis optio vobis datur eligite hodie quod placet cui potissimum servire debeatis utrum diis quibus servierunt patres vestri in Mesopotamia an diis Amorreorum in quorum terra habitatis ego autem et domus mea serviemus Domino
JOSH|24|16|responditque populus et ait absit a nobis ut relinquamus Dominum et serviamus diis alienis
JOSH|24|17|Dominus Deus noster ipse eduxit nos et patres nostros de terra Aegypti de domo servitutis fecitque videntibus nobis signa ingentia et custodivit nos in omni via per quam ambulavimus et in cunctis populis per quos transivimus
JOSH|24|18|et eiecit universas gentes Amorreum habitatorem terrae quam nos intravimus serviemus igitur Domino quia ipse est Deus noster
JOSH|24|19|dixitque Iosue ad populum non poteritis servire Domino Deus enim sanctus et fortis aemulator est nec ignoscet sceleribus vestris atque peccatis
JOSH|24|20|si dimiseritis Dominum et servieritis diis alienis convertet se et adfliget vos atque subvertet postquam vobis praestiterit bona
JOSH|24|21|dixitque populus ad Iosue nequaquam ita ut loqueris erit sed Domino serviemus
JOSH|24|22|et Iosue ad populum testes inquit vos estis quia ipsi elegeritis vobis Dominum ut serviatis ei responderuntque testes
JOSH|24|23|nunc ergo ait auferte deos alienos de medio vestrum et inclinate corda vestra ad Dominum Deum Israhel
JOSH|24|24|dixitque populus ad Iosue Domino Deo nostro serviemus oboedientes praeceptis eius
JOSH|24|25|percussit igitur Iosue in die illo foedus et proposuit populo praecepta atque iudicia in Sychem
JOSH|24|26|scripsitque omnia verba haec in volumine legis Dei et tulit lapidem pergrandem posuitque eum subter quercum quae erat in sanctuario Domini
JOSH|24|27|et dixit ad omnem populum en lapis iste erit vobis in testimonium quod audierit omnia verba Domini quae locutus est vobis ne forte postea negare velitis et mentiri Domino Deo vestro
JOSH|24|28|dimisitque populum singulos in possessionem suam
JOSH|24|29|et post haec mortuus est Iosue filius Nun servus Domini centum decem annorum
JOSH|24|30|sepelieruntque eum in finibus possessionis suae in Thamnathsare quae sita est in monte Ephraim a septentrionali parte montis Gaas
JOSH|24|31|servivitque Israhel Domino cunctis diebus Iosue et seniorum qui longo vixerunt tempore post Iosue et qui noverant omnia opera Domini quae fecerat in Israhel
JOSH|24|32|ossa quoque Ioseph quae tulerant filii Israhel de Aegypto sepelierunt in Sychem in parte agri quem emerat Iacob a filiis Emmor patris Sychem centum novellis ovibus et fuit in possessione filiorum Ioseph
JOSH|24|33|Eleazar quoque filius Aaron mortuus est et sepelierunt eum in Gaab Finees filii eius quae data est ei in monte Ephraim
