NUM|1|1|以色列 人出 埃及 地後第二年二月初一，耶和華在 西奈 曠野，在會幕中吩咐 摩西 說：
NUM|1|2|「你要按宗族、父家、人名的數目計算 以色列 全會眾，數點所有的男丁。
NUM|1|3|以色列 中凡二十歲以上能出去打仗的，你和 亞倫 要按照他們的隊伍數點。
NUM|1|4|每支派要有一個人，就是父家的家長跟你們一起。
NUM|1|5|這是幫助你們的人的名字： 屬 呂便 的， 示丟珥 的兒子 以利蓿 ；
NUM|1|6|屬 西緬 的， 蘇利沙代 的兒子 示路蔑 ；
NUM|1|7|屬 猶大 的， 亞米拿達 的兒子 拿順 ；
NUM|1|8|屬 以薩迦 的， 蘇押 的兒子 拿坦業 ；
NUM|1|9|屬 西布倫 的， 希倫 的兒子 以利押 ；
NUM|1|10|約瑟 子孫、屬 以法蓮 的， 亞米忽 的兒子 以利沙瑪 ；屬 瑪拿西 的， 比大蓿 的兒子 迦瑪列 ；
NUM|1|11|屬 便雅憫 的， 基多尼 的兒子 亞比但 ；
NUM|1|12|屬 但 的， 亞米沙代 的兒子 亞希以謝 ；
NUM|1|13|屬 亞設 的， 俄蘭 的兒子 帕結 ；
NUM|1|14|屬 迦得 的， 丟珥 的兒子 以利雅薩 ；
NUM|1|15|屬 拿弗他利 的， 以南 的兒子 亞希拉 。」
NUM|1|16|這些是從會眾中選出來的父系支派的領袖，是 以色列 部隊的官長。
NUM|1|17|於是， 摩西 和 亞倫 帶著這些按名指定的人，
NUM|1|18|在二月初一召集全會眾。會眾就照他們的宗族、父家、人名的數目，登記二十歲以上的人口。
NUM|1|19|耶和華怎樣吩咐 摩西 ，他就照樣在 西奈 的曠野數點他們。
NUM|1|20|以色列 的長子， 呂便 子孫的後代，照著宗族、父家、人名的數目，他們的人口凡二十歲以上能出去打仗的男丁，
NUM|1|21|呂便 支派被數的共有四萬六千五百名。
NUM|1|22|西緬 子孫的後代，照著宗族、父家、被數 人名的數目，他們的人口凡二十歲以上能出去打仗的男丁，
NUM|1|23|西緬 支派被數的共有五萬九千三百名。
NUM|1|24|迦得 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|25|迦得 支派被數的共有四萬五千六百五十名。
NUM|1|26|猶大 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|27|猶大 支派被數的共有七萬四千六百名。
NUM|1|28|以薩迦 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|29|以薩迦 支派被數的共有五萬四千四百名。
NUM|1|30|西布倫 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|31|西布倫 支派被數的共有五萬七千四百名。
NUM|1|32|約瑟 子孫屬 以法蓮 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|33|以法蓮 支派被數的共有四萬零五百名。
NUM|1|34|瑪拿西 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|35|瑪拿西 支派被數的共有三萬二千二百名。
NUM|1|36|便雅憫 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|37|便雅憫 支派被數的共有三萬五千四百名。
NUM|1|38|但 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|39|但 支派被數的共有六萬二千七百名。
NUM|1|40|亞設 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|41|亞設 支派被數的共有四萬一千五百名。
NUM|1|42|拿弗他利 子孫的後代，照著宗族、父家、人名的數目，凡二十歲以上能出去打仗的，
NUM|1|43|拿弗他利 支派被數的共有五萬三千四百名。
NUM|1|44|這些就是被數點的，是 摩西 、 亞倫 和 以色列 十二個領袖所數點的；每一個領袖代表他們的父家。
NUM|1|45|以色列 人被數點的總數， 以色列 中照著父家，凡二十歲以上能出去打仗的，
NUM|1|46|他們被數點的總數是六十萬三千五百五十名。
NUM|1|47|利未 人卻沒有按照父系支派數在其中。
NUM|1|48|耶和華吩咐 摩西 說：
NUM|1|49|「惟獨 利未 支派你不可數點，也不可在 以色列 人中計算他們的人口。
NUM|1|50|你要派 利未 人管理法櫃的帳幕和其中一切的器具，以及屬帳幕的一切。他們要抬帳幕和其中一切的器具，並要辦理帳幕的事務，在帳幕的四圍安營。
NUM|1|51|帳幕將往前行的時候， 利未 人要拆卸；將駐紮的時候， 利未 人要支搭帳幕。近前來的外人必被處死。
NUM|1|52|以色列 人要按照各自的隊伍安營，各歸本營，各歸本旗。
NUM|1|53|但 利未 人要在法櫃帳幕的四圍安營，免得憤怒臨到 以色列 會眾； 利未 人要負責看守法櫃的帳幕。」
NUM|1|54|以色列 人就這樣做了。凡耶和華所吩咐 摩西 的，他們都照樣做了。
NUM|2|1|耶和華吩咐 摩西 和 亞倫 說：
NUM|2|2|「 以色列 人各人要在自己的旗幟下，按照自己父家的旗號安營，對著會幕的四圍安營。
NUM|2|3|「在東邊，向日出的方向， 猶大 營按照他們的隊伍，在它的旗幟下安營。 猶大 人的領袖是 亞米拿達 的兒子 拿順 ，
NUM|2|4|他的軍隊被數的有七萬四千六百名。
NUM|2|5|在他旁邊安營的是 以薩迦 支派。 以薩迦 人的領袖是 蘇押 的兒子 拿坦業 ，
NUM|2|6|他的軍隊被數的有五萬四千四百名。
NUM|2|7|還有 西布倫 支派， 西布倫 人的領袖是 希倫 的兒子 以利押 ，
NUM|2|8|他的軍隊被數的有五萬七千四百名。
NUM|2|9|凡屬 猶大 營，照他們隊伍被數的共有十八萬六千四百名；他們要作第一隊往前行。
NUM|2|10|「在南邊，按照他們的隊伍是 呂便 營的旗幟。 呂便 人的領袖是 示丟珥 的兒子 以利蓿 ，
NUM|2|11|他的軍隊被數的有四萬六千五百名。
NUM|2|12|在他旁邊安營的是 西緬 支派。 西緬 人的領袖是 蘇利沙代 的兒子 示路蔑 ，
NUM|2|13|他的軍隊被數的有五萬九千三百名。
NUM|2|14|還有 迦得 支派， 迦得 人的領袖是 丟珥 的兒子 以利雅薩 ，
NUM|2|15|他的軍隊被數的有四萬五千六百五十名。
NUM|2|16|凡屬 呂便 營，照他們隊伍被數的共有十五萬一千四百五十名；他們要作第二隊往前行。
NUM|2|17|「會幕與 利未 營在諸營中間往前行。他們怎樣安營就怎樣往前行，各按本位，各歸本旗。
NUM|2|18|「在西邊，按照他們的隊伍是 以法蓮 營的旗幟。 以法蓮 人的領袖是 亞米忽 的兒子 以利沙瑪 ，
NUM|2|19|他的軍隊被數的有四萬零五百名。
NUM|2|20|在他旁邊的是 瑪拿西 支派。 瑪拿西 人的領袖是 比大蓿 的兒子 迦瑪列 ，
NUM|2|21|他的軍隊被數的有三萬二千二百名。
NUM|2|22|還有 便雅憫 支派， 便雅憫 人的領袖是 基多尼 的兒子 亞比但 ，
NUM|2|23|他的軍隊被數的有三萬五千四百名。
NUM|2|24|凡屬 以法蓮 營，照他們隊伍被數的共有十萬八千一百名；他們要作第三隊往前行。
NUM|2|25|「在北邊，按照他們的隊伍是 但 營的旗幟。 但 人的領袖是 亞米沙代 的兒子 亞希以謝 ，
NUM|2|26|他的軍隊被數的有六萬二千七百名。
NUM|2|27|在他旁邊安營的是 亞設 支派。 亞設 人的領袖是 俄蘭 的兒子 帕結 ，
NUM|2|28|他的軍隊被數的有四萬一千五百名。
NUM|2|29|還有 拿弗他利 支派， 拿弗他利 人的領袖是 以南 的兒子 亞希拉 ，
NUM|2|30|他的軍隊被數的有五萬三千四百名。
NUM|2|31|凡屬 但 營被數的共有十五萬七千六百名；他們隨著自己的旗幟行在最後。」
NUM|2|32|以上是 以色列 人按照各自的父家被數的，在諸營中按照各自的隊伍被數的，共有六十萬三千五百五十名。
NUM|2|33|但 利未 人沒有數在 以色列 人中，正如耶和華所吩咐 摩西 的。
NUM|2|34|以色列 人就照著耶和華所吩咐 摩西 的做了，在各自的旗幟下安營，隨著各自的宗族、父家起行。
NUM|3|1|耶和華在 西奈山 與 摩西 說話的日子， 亞倫 和 摩西 的後代如下：
NUM|3|2|這些是 亞倫 兒子的名字，長子 拿答 ，及 亞比戶 、 以利亞撒 、 以他瑪 。
NUM|3|3|這些是 亞倫 兒子的名字，都是受膏的祭司，是 摩西 授聖職使他們擔任祭司職分的。
NUM|3|4|拿答 、 亞比戶 在 西奈 的曠野向耶和華獻上凡火的時候，死在耶和華面前。他們沒有兒子。 以利亞撒 和 以他瑪 在他們的父親 亞倫 面前擔任祭司的職分。
NUM|3|5|耶和華吩咐 摩西 說：
NUM|3|6|「你要帶 利未 支派近前來，站在 亞倫 祭司面前伺候他。
NUM|3|7|他們要替他，又替全會眾，在會幕前執行任務，辦理帳幕的事。
NUM|3|8|他們要看守會幕一切的器具，為 以色列 人執行任務，辦理帳幕的事。
NUM|3|9|你要把 利未 人給 亞倫 和他的兒子；他們是從 以色列 人中選出來完全給他的。
NUM|3|10|你要指派 亞倫 和他的兒子謹守祭司的職分；近前來的外人必被處死。」
NUM|3|11|耶和華吩咐 摩西 說：
NUM|3|12|「看哪，我從 以色列 人中選了 利未 人，代替 以色列 人中所有頭胎的長子； 利未 人要歸我。
NUM|3|13|因為凡頭生的是我的；我在 埃及 地擊殺所有頭生的那日，就把 以色列 中所有頭生的，無論是人或牲畜，都分別為聖歸我；他們定要屬我。我是耶和華。」
NUM|3|14|耶和華在 西奈 的曠野吩咐 摩西 說：
NUM|3|15|「你要照父家、宗族計算 利未 人。凡一個月以上的男子都要數點。」
NUM|3|16|於是 摩西 遵照耶和華的吩咐，按所指示的數點他們。
NUM|3|17|利未 兒子的名字是 革順 、 哥轄 、 米拉利 。
NUM|3|18|按照宗族， 革順 兒子的名字是 立尼 、 示每 。
NUM|3|19|按照宗族， 哥轄 的兒子是 暗蘭 、 以斯哈 、 希伯倫 、 烏薛 。
NUM|3|20|按照宗族， 米拉利 的兒子是 抹利 、 母示 。按照父家，這些都是 利未 人的宗族。
NUM|3|21|屬 革順 的有 立尼 族、 示每 族，他們是 革順 人的宗族。
NUM|3|22|他們被數的，一個月以上所有男子的數目共有七千五百名。
NUM|3|23|這 革順 人的宗族要在西邊，在帳幕後面安營。
NUM|3|24|革順 人父家的領袖是 拉伊勒 的兒子 以利雅薩 。
NUM|3|25|革順 的子孫在會幕中要看守的是帳幕、罩棚、罩棚的蓋、會幕的門簾、
NUM|3|26|帳幕和祭壇周圍院子的帷幔和門簾，以及所有需用的繩子。
NUM|3|27|屬 哥轄 的有 暗蘭 族、 以斯哈 族、 希伯倫 族、 烏薛 族，他們是 哥轄 人的宗族。
NUM|3|28|一個月以上所有男子的數目共有八千六百 名；他們負責看守聖所。
NUM|3|29|哥轄 子孫的宗族要在帳幕的南邊安營。
NUM|3|30|哥轄 人父家宗族的領袖是 烏薛 的兒子 以利撒反 。
NUM|3|31|他們要看守的是約櫃、供桌、燈臺、祭壇、香壇、祭司在聖所內用的器皿、簾子，與一切相關事奉的物件。
NUM|3|32|亞倫 祭司的兒子 以利亞撒 是 利未 人眾領袖的主管，他要監督那些負責看守聖所的人。
NUM|3|33|屬 米拉利 的有 抹利 族、 母示 族，他們是 米拉利 的宗族。
NUM|3|34|他們被數的，一個月以上所有男子的數目共有六千二百名。
NUM|3|35|米拉利 宗族的領袖是 亞比亥 的兒子 蘇列 ，他們要在帳幕的北邊安營。
NUM|3|36|米拉利 子孫的職分是看守帳幕的豎板、橫木、柱子、帶卯眼的座和一切的器具，就是一切相關事奉的物件，
NUM|3|37|以及院子四圍的柱子、其上帶卯眼的座、橛子和繩子。
NUM|3|38|在帳幕前東邊，向日出的方向，安營的是 摩西 、 亞倫 和 亞倫 的兒子。他們負責看守聖所，是為 以色列 人看守的。近前來的外人必被處死。
NUM|3|39|凡被數的 利未 人，就是 摩西 、 亞倫 照耶和華所指示、按宗族所數的，一個月以上所有的男子共有二萬二千名。
NUM|3|40|耶和華對 摩西 說：「你要數點 以色列 人中凡一個月以上頭生的男子，登記他們的名字。
NUM|3|41|我是耶和華。你要揀選 利未 人歸我，代替所有頭生的 以色列 人，也取 利未 人的牲畜代替 以色列 人所有頭生的牲畜。」
NUM|3|42|摩西 就遵照耶和華所吩咐的，把所有 以色列 人頭生的都數點了。
NUM|3|43|按人名的數目，凡一個月以上頭生的男子共有二萬二千二百七十三名。
NUM|3|44|耶和華吩咐 摩西 說：
NUM|3|45|「你要揀選 利未 人代替所有頭生的 以色列 人，也要取 利未 人的牲畜代替 以色列 人的牲畜。 利未 人要歸我，我是耶和華。
NUM|3|46|以色列 人頭生的男子比 利未 人多了二百七十三名，必須把他們贖出來；
NUM|3|47|按照人丁，照聖所的舍客勒，每人當付五舍客勒，一舍客勒是二十季拉。
NUM|3|48|你要把這些多出來的人的贖銀交給 亞倫 和他的兒子。」
NUM|3|49|於是 摩西 從那被 利未 人所贖以外多出來的人取了贖銀。
NUM|3|50|從頭生的 以色列 人所取的銀子，按照聖所的舍客勒，共計一千三百六十五舍客勒。
NUM|3|51|摩西 遵照耶和華指示的話，把贖銀交給 亞倫 和他的兒子，正如耶和華所吩咐的。
NUM|4|1|耶和華吩咐 摩西 和 亞倫 說：
NUM|4|2|「你要照宗族、父家計算 利未 人中 哥轄 子孫的人口，
NUM|4|3|就是從三十歲到五十歲，凡前來任職，在會幕裏事奉的人。
NUM|4|4|這是 哥轄 子孫在會幕裏有關至聖之物的職責。
NUM|4|5|「拔營的時候， 亞倫 和他兒子要進去，把遮掩的幔子取下，用它來遮蓋法櫃，
NUM|4|6|又用精美皮料蓋在上面，鋪上純藍色的布，再把槓穿上。
NUM|4|7|他們要用藍色的布鋪在供餅的桌上，將盤、碟，以及澆酒祭的杯和壺擺在上面；經常供的餅也要留在桌上。
NUM|4|8|他們要在這些東西的上面鋪上朱紅色的布，把精美皮料蓋在上面，再把槓穿上。
NUM|4|9|他們要用藍色的布遮蓋供職用的燈臺、燈臺上的燈盞、燈剪、燈盤，以及所有盛油的器皿；
NUM|4|10|又要用精美皮料把燈臺和燈臺的一切器具包好，放在抬架上。
NUM|4|11|他們要用藍色的布鋪在金壇上，用精美皮料蓋在上面，再把槓穿上。
NUM|4|12|要用藍色的布把聖所供職用的一切器具包好，再用精美皮料蓋在上面，放在抬架上。
NUM|4|13|他們要清理祭壇上的灰，用紫色的布鋪在壇上；
NUM|4|14|又要把供職用的一切器具，就是祭壇一切的器具，火盆、肉叉、鏟子和盤子，都擺在壇上，鋪上精美皮料，再把槓穿上。
NUM|4|15|「拔營的時候， 亞倫 和他兒子把聖所和聖所一切的器具蓋好之後， 哥轄 的子孫才好來抬，免得他們摸聖物而死；這是 哥轄 子孫在會幕裏所當抬的。
NUM|4|16|「祭司 亞倫 的兒子 以利亞撒 所要照管的是點燈的油和香料，以及常獻的素祭和膏油。他要照管整個帳幕和其中所有的，以及聖所和聖所的器具。」
NUM|4|17|耶和華吩咐 摩西 和 亞倫 說：
NUM|4|18|「你們不可使 哥轄 人宗族的這一支從 利未 人中剪除。
NUM|4|19|他們挨近至聖之物的時候，要向他們這樣做，使他們存活，不致死亡； 亞倫 和他的兒子要進去，分派各人當做的，當抬的。
NUM|4|20|但是他們不可進去觀看聖所的拆卸 ，免得死亡。」
NUM|4|21|耶和華吩咐 摩西 說：
NUM|4|22|「你要照父家、宗族計算 革順 子孫的人口；
NUM|4|23|從三十歲到五十歲，凡前來任職，在會幕裏事奉的，都要數點。
NUM|4|24|這是 革順 人宗族的職責，要做的事，要抬的東西如下：
NUM|4|25|他們要抬帳幕的幔子、會幕和會幕的蓋、外層精美皮料的蓋、會幕的門簾、
NUM|4|26|帳幕和祭壇周圍院子的帷幔和門簾、繩子，以及所有需用的器具；一切與這些東西相關的事務，他們要盡職。
NUM|4|27|革順 人的子孫一切的事奉，就是所當抬的，所當做的，都要遵照 亞倫 和他兒子的指示；他們所當抬的，你們要派他們負責。
NUM|4|28|這是 革順 人子孫的宗族在會幕裏的事奉；他們要在 亞倫 祭司的兒子 以他瑪 的手下盡職。」
NUM|4|29|「至於 米拉利 的子孫，你要照宗族、父家數點他們；
NUM|4|30|從三十歲到五十歲，凡前來任職，在會幕裏事奉的，你都要數點。
NUM|4|31|這是他們在會幕裏的事奉，他們負責要抬的是帳幕的豎板、橫木、柱子和帶卯眼的座，
NUM|4|32|院子四圍的柱子和其上帶卯眼的座、橛子、繩子和一切的器具，與一切相關事奉的物件。你們要按名指定他們要抬的器具。
NUM|4|33|這是 米拉利 子孫的宗族在會幕裏的事奉，都在 亞倫 祭司的兒子 以他瑪 的手下。」
NUM|4|34|摩西 、 亞倫 和會眾的領袖按照宗族、父家數點 哥轄 人的子孫；
NUM|4|35|從三十歲到五十歲，凡前來任職，在會幕裏事奉的，
NUM|4|36|按照宗族被數的共有二千七百五十名。
NUM|4|37|這是所有在會幕裏事奉的 哥轄 人宗族中被數的，是 摩西 和 亞倫 遵照耶和華藉 摩西 所指示數點的。
NUM|4|38|革順 子孫被數的，按照宗族、父家，
NUM|4|39|從三十歲到五十歲，凡前來任職，在會幕裏事奉的，
NUM|4|40|按照宗族、父家被數的共有二千六百三十名。
NUM|4|41|這是所有在會幕裏事奉的 革順 子孫宗族中被數的，是 摩西 和 亞倫 遵照耶和華的指示所數點的。
NUM|4|42|米拉利 子孫宗族被數的，按照宗族、父家，
NUM|4|43|從三十歲到五十歲，凡前來任職，在會幕裏事奉的，
NUM|4|44|按照宗族被數的共有三千二百名。
NUM|4|45|這是 米拉利 子孫宗族中被數的，是 摩西 和 亞倫 遵照耶和華藉 摩西 所指示數點的。
NUM|4|46|摩西 、 亞倫 和 以色列 領袖按照宗族、父家數點 利未 人，
NUM|4|47|從三十歲到五十歲，凡前來任職，在會幕裏事奉，做抬物之工的，
NUM|4|48|他們被數的共有八千五百八十名。
NUM|4|49|按照耶和華藉 摩西 所指示的來分派，各人都有自己所做的事、所抬的物；他們就這樣被數點，正如耶和華所吩咐 摩西 的。
NUM|5|1|耶和華吩咐 摩西 說：
NUM|5|2|「你要吩咐 以色列 人，把一切患痲瘋 的、患漏症的和因屍體而不潔淨的，都送到營外去。
NUM|5|3|無論男女你都要送，把他們送到營外，免得他們玷污了他們的營，這是我住在他們中間的地方。」
NUM|5|4|以色列 人就照樣做，把他們送到營外去。耶和華怎樣吩咐 摩西 ， 以色列 人就照樣做了。
NUM|5|5|耶和華吩咐 摩西 說：
NUM|5|6|「你要吩咐 以色列 人：無論男女，若犯了人所常犯的任何罪 ，以致干犯耶和華，那人就有了罪。
NUM|5|7|他要承認所犯的罪，將所虧負人的如數賠償，另外再加五分之一，交給所虧負的人。
NUM|5|8|那人若沒有至親可接受所賠償的，所賠償的就要歸耶和華，交給祭司；另外還要獻一隻贖罪的公羊為他贖罪。
NUM|5|9|以色列 人一切的聖物中，所奉給祭司的一切禮物都要歸給祭司。
NUM|5|10|各人自己的聖物歸自己，給祭司的要歸給祭司。」
NUM|5|11|耶和華吩咐 摩西 說：
NUM|5|12|「你要吩咐 以色列 人，對他們說：若任何人的妻子背離婦道，對丈夫不貞，
NUM|5|13|有人與她同寢交合，這事瞞過她的丈夫，沒有被發現；她玷污自己，沒有證人指控她，也沒有被捉住；
NUM|5|14|丈夫若生了疑忌的心，對妻子起了疑忌，認為她玷污自己；或是丈夫生了疑忌的心，對妻子起了疑忌，雖然她沒有玷污自己，
NUM|5|15|這人要帶妻子到祭司那裏，同時為她帶十分之一伊法大麥麵粉作供物。不可澆上油，也不可加乳香，因為這是疑忌的素祭，是紀念的素祭，使人記得罪孽。
NUM|5|16|「祭司要使那婦人近前來，站在耶和華面前。
NUM|5|17|祭司要把聖水盛在瓦器裏，從帳幕的地上取些塵土，放在水中。
NUM|5|18|祭司要帶那婦人站在耶和華面前，使她蓬頭散髮，再把紀念的素祭，就是疑忌的素祭，放在她的手掌，祭司手裏捧著致詛咒的苦水。
NUM|5|19|祭司要叫婦人起誓，對她說：『若沒有人與你同寢，若你未曾背著丈夫做污穢的事，你就能免去這致詛咒的苦水。
NUM|5|20|但你背著丈夫，玷污自己，跟丈夫以外的人同寢。』
NUM|5|21|祭司叫婦人賭咒起誓，祭司對她說：『當耶和華使你大腿萎縮，肚腹腫脹時，願耶和華使你在你百姓中成為詛咒和咒罵；
NUM|5|22|願這致詛咒的水進入你體內，使你肚腹腫脹，大腿萎縮。』婦人要說：『阿們，阿們。』
NUM|5|23|「祭司要把這詛咒寫在冊上，然後用苦水塗去，
NUM|5|24|又叫婦人喝這致詛咒的苦水，這詛咒的水要進入她裏面，令她痛苦。
NUM|5|25|祭司要從婦人手中取那疑忌的素祭，把素祭在耶和華面前搖一搖，拿到祭壇前；
NUM|5|26|又要從素祭中取出一把，作為紀念，燒在壇上，然後叫婦人喝這水。
NUM|5|27|祭司叫她喝了以後，她若玷污自己，確實對丈夫不貞，這致詛咒的水必進入她裏面，令她痛苦，她的肚腹就要腫脹起來，大腿萎縮；這婦人就在她百姓中成為詛咒。
NUM|5|28|這婦人若沒有玷污自己，是貞潔的，就要免受這災，並且能夠生育。
NUM|5|29|「這是疑忌的條例。妻子背離丈夫玷污自己，
NUM|5|30|或是丈夫生了疑忌的心，對妻子起了疑忌，祭司要使那婦人站在耶和華面前，在她身上照這條例而行。
NUM|5|31|男人可免罪責；女人必須擔當自己的罪孽。」
NUM|6|1|耶和華吩咐 摩西 說：
NUM|6|2|「你要吩咐 以色列 人，對他們說：無論男女，若許了特別的願，就是拿細耳人的願，願意離俗歸耶和華，
NUM|6|3|他就要遠離清酒烈酒，也不可喝任何清酒烈酒做的醋；不可喝任何葡萄汁，也不可吃鮮葡萄和乾葡萄。
NUM|6|4|在一切離俗的日子，任何葡萄樹上所結的，甚至果核和果皮，都不可吃。
NUM|6|5|「在他一切許願離俗的日子，不可用剃刀剃頭。在離俗歸耶和華的日子未滿之前，他要成為聖，要任由頭上的髮綹生長。
NUM|6|6|在他一切離俗歸耶和華的日子，不可挨近死屍。
NUM|6|7|即使他的父母或兄弟姊妹死了，他也不可因他們使自己不潔淨，因為他頭上有離俗歸上帝的記號 。
NUM|6|8|在他一切離俗的日子，他是歸耶和華為聖的。
NUM|6|9|「若在他旁邊忽然有人死了，因而玷污了他離俗的頭，他要在第七日，得潔淨的日子剃頭。
NUM|6|10|第八日，他要把兩隻斑鳩或兩隻雛鴿帶到會幕門口，交給祭司。
NUM|6|11|祭司要獻一隻作贖罪祭，一隻作燔祭，為他贖因屍體而有的罪，並要在當日使他的頭分別為聖。
NUM|6|12|他要另選離俗歸耶和華的日子，牽一隻一歲的小公羊來作贖愆祭。先前的那段日子算為無效，因為他在離俗期間被玷污了。
NUM|6|13|「拿細耳人的條例是這樣的：離俗的日子滿了，祭司要領他到會幕門口，
NUM|6|14|他要將供物獻給耶和華，就是一隻沒有殘疾的一歲小公羊作燔祭，一隻沒有殘疾的一歲小母羊作贖罪祭，和一隻沒有殘疾的公綿羊作平安祭，
NUM|6|15|一籃用油調和的無酵細麵餅和抹了油的無酵薄餅，以及同獻的素祭和澆酒祭。
NUM|6|16|祭司要來到耶和華面前，獻上那人的贖罪祭和燔祭。
NUM|6|17|祭司要把公綿羊和那籃無酵餅獻給耶和華作平安祭，又要獻上同獻的素祭和澆酒祭。
NUM|6|18|拿細耳人要在會幕門口剃離俗的頭，把離俗頭上的髮放在平安祭下的火上。
NUM|6|19|他剃了離俗的頭以後，祭司要取那煮好的公綿羊的一條前腿，連同籃子裏的一塊無酵餅和一塊無酵薄餅，放在他手掌上。
NUM|6|20|祭司要拿這些在耶和華面前搖一搖，作為搖祭；這和所搖的胸、所舉的腿一樣是聖物，是歸給祭司的。然後拿細耳人才可以喝酒。
NUM|6|21|「這是拿細耳人許願的條例，除了他手頭財力所及之外，他要為離俗獻供物給耶和華。他怎樣許願，就當照離俗的條例做。」
NUM|6|22|耶和華吩咐 摩西 說：
NUM|6|23|「你要吩咐 亞倫 和他兒子說：你們要這樣為 以色列 人祝福，對他們說：
NUM|6|24|『願耶和華賜福給你，保護你。
NUM|6|25|願耶和華使他的臉光照你，賜恩給你。
NUM|6|26|願耶和華向你仰臉，賜你平安。』
NUM|6|27|「他們要如此奉我的名為 以色列 人祝福；我也要賜福給他們。」
NUM|7|1|摩西 豎立帳幕後，就用膏抹了帳幕，使它分別為聖，又用膏抹其中的一切器具，以及祭壇和壇上的一切器具，使它們分別為聖。
NUM|7|2|以色列 的領袖，各父家的家長，都前來奉獻。他們是各支派的領袖，管理那些被數的人。
NUM|7|3|他們把自己的供物送到耶和華面前，就是六輛篷車和十二頭公牛。每兩個領袖奉獻一輛車，每個領袖奉獻一頭牛。他們把這些都帶到帳幕前。
NUM|7|4|耶和華對 摩西 說：
NUM|7|5|「你要從他們收下這些，作為會幕事奉的用途，照著 利未 人所事奉的交給他們各人。」
NUM|7|6|於是 摩西 收了車和牛，交給 利未 人。
NUM|7|7|他把兩輛車和四頭牛，照著 革順 子孫所事奉的交給他們，
NUM|7|8|又把四輛車和八頭牛，照著 米拉利 子孫所事奉的交給他們。他們都在 亞倫 祭司的兒子 以他瑪 的手下。
NUM|7|9|但沒有交給 哥轄 子孫任何東西，因為他們所事奉的是聖物，必須抬在肩頭上。
NUM|7|10|用膏抹祭壇的那一天，眾領袖前來為獻壇奉獻；眾領袖都在祭壇前獻供物。
NUM|7|11|耶和華對 摩西 說：「眾領袖為獻壇奉獻供物，每天要有一個領袖前來奉獻。」
NUM|7|12|第一天獻供物的是 猶大 支派的 亞米拿達 的兒子 拿順 。
NUM|7|13|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|14|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|15|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|16|一隻公山羊作贖罪祭；
NUM|7|17|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 亞米拿達 的兒子 拿順 的供物。
NUM|7|18|第二天來獻的是 以薩迦 的領袖， 蘇押 的兒子 拿坦業 。
NUM|7|19|他獻為供物的是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|20|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|21|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|22|一隻公山羊作贖罪祭；
NUM|7|23|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 蘇押 的兒子 拿坦業 的供物。
NUM|7|24|第三天是 西布倫 子孫的領袖， 希倫 的兒子 以利押 。
NUM|7|25|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|26|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|27|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|28|一隻公山羊作贖罪祭；
NUM|7|29|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 希倫 的兒子 以利押 的供物。
NUM|7|30|第四天是 呂便 子孫的領袖， 示丟珥 的兒子 以利蓿 。
NUM|7|31|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|32|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|33|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|34|一隻公山羊作贖罪祭；
NUM|7|35|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 示丟珥 的兒子 以利蓿 的供物。
NUM|7|36|第五天是 西緬 子孫的領袖， 蘇利沙代 的兒子 示路蔑 。
NUM|7|37|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|38|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|39|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|40|一隻公山羊作贖罪祭；
NUM|7|41|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 蘇利沙代 的兒子 示路蔑 的供物。
NUM|7|42|第六天是 迦得 子孫的領袖， 丟珥 的兒子 以利雅薩 。
NUM|7|43|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|44|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|45|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|46|一隻公山羊作贖罪祭；
NUM|7|47|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 丟珥 的兒子 以利雅薩 的供物。
NUM|7|48|第七天是 以法蓮 子孫的領袖， 亞米忽 的兒子 以利沙瑪 。
NUM|7|49|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|50|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|51|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|52|一隻公山羊作贖罪祭；
NUM|7|53|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 亞米忽 的兒子 以利沙瑪 的供物。
NUM|7|54|第八天是 瑪拿西 子孫的領袖， 比大蓿 的兒子 迦瑪列 。
NUM|7|55|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|56|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|57|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|58|一隻公山羊作贖罪祭；
NUM|7|59|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 比大蓿 的兒子 迦瑪列 的供物。
NUM|7|60|第九天是 便雅憫 子孫的領袖， 基多尼 的兒子 亞比但 。
NUM|7|61|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|62|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|63|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|64|一隻公山羊作贖罪祭；
NUM|7|65|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 基多尼 的兒子 亞比但 的供物。
NUM|7|66|第十天是 但 子孫的領袖， 亞米沙代 的兒子 亞希以謝 。
NUM|7|67|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|68|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|69|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|70|一隻公山羊作贖罪祭；
NUM|7|71|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 亞米沙代 的兒子 亞希以謝 的供物。
NUM|7|72|第十一天是 亞設 子孫的領袖， 俄蘭 的兒子 帕結 。
NUM|7|73|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|74|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|75|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|76|一隻公山羊作贖罪祭；
NUM|7|77|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 俄蘭 的兒子 帕結 的供物。
NUM|7|78|第十二天是 拿弗他利 子孫的領袖， 以南 兒子 亞希拉 。
NUM|7|79|他的供物是：一個重一百三十舍客勒的銀盤，一個重七十舍客勒的銀碗，都是按照聖所的舍客勒，裏面盛滿了調油的細麵作素祭；
NUM|7|80|一個重十舍客勒的金碟子，盛滿了香；
NUM|7|81|一頭公牛犢、一隻公綿羊、一隻一歲的小公羊作燔祭；
NUM|7|82|一隻公山羊作贖罪祭；
NUM|7|83|兩頭公牛、五隻公綿羊、五隻公山羊、五隻一歲的小公羊作平安祭。這是 以南 的兒子 亞希拉 的供物。
NUM|7|84|用膏抹祭壇的那一天， 以色列 的眾領袖為獻壇所獻的是：銀盤十二個、銀碗十二個、金碟子十二個；
NUM|7|85|一個銀盤重一百三十，一個碗七十。一切器皿的銀子，按照聖所的舍客勒共二千四百舍客勒。
NUM|7|86|十二個金碟子盛滿了香，按照聖所的舍客勒，一個碟子重十舍客勒，所有碟子的金子共一百二十舍客勒。
NUM|7|87|作燔祭的共有公牛十二頭、公羊十二隻、一歲的小公羊十二隻，和同獻的素祭，以及作贖罪祭的公山羊十二隻；
NUM|7|88|作平安祭的共有公牛二十四頭、公綿羊六十隻、公山羊六十隻、一歲的小公羊六十隻。這就是用膏抹壇之後，為獻壇的奉獻。
NUM|7|89|摩西 進會幕要與耶和華說話的時候，聽見法櫃的櫃蓋以上二基路伯中間有對他說話的聲音。耶和華向他說話。
NUM|8|1|耶和華吩咐 摩西 說：
NUM|8|2|「你要吩咐 亞倫 ，對他說：點燈的時候，七盞燈都要照亮燈臺前面。」
NUM|8|3|亞倫 就照樣做了；他點燈，照亮了燈臺前面，正如耶和華所吩咐 摩西 的。
NUM|8|4|燈臺是這樣造的：燈臺是用金子錘出來的，連座帶花都是錘出來的。 摩西 照著耶和華所指示的樣式造了燈臺。
NUM|8|5|耶和華吩咐 摩西 說：
NUM|8|6|「你要從 以色列 人中選出 利未 人來，潔淨他們。
NUM|8|7|你要這樣做來潔淨他們：要用潔淨的水彈在他們身上，又叫他們用剃刀剃刮全身，洗淨衣服，潔淨自己。
NUM|8|8|然後他們要取一頭公牛犢，以及同獻的素祭，就是調油的細麵。你要另取一頭公牛犢作贖罪祭。
NUM|8|9|你要帶 利未 人到會幕前，並且要召集 以色列 全會眾。
NUM|8|10|你要把 利未 人帶到耶和華面前， 以色列 人要為 利未 人按手。
NUM|8|11|亞倫 要從 以色列 人中將 利未 人奉獻 在耶和華面前，作為搖祭，使他們事奉耶和華。
NUM|8|12|利未 人要按手在那兩頭牛的頭上；你要將一頭作贖罪祭，一頭作燔祭，獻給耶和華，為 利未 人贖罪。
NUM|8|13|你也要使 利未 人站在 亞倫 和他兒子面前，將他們奉獻給耶和華，作為搖祭。
NUM|8|14|「你從 以色列 人中將 利未 人分別出來， 利未 人就歸我了。
NUM|8|15|你潔淨了 利未 人，奉獻他們作為搖祭之後，他們就可以進會幕事奉。
NUM|8|16|因為他們是從 以色列 人中全然獻給我的；我選他們歸我，代替 以色列 人中所有頭胎的長子。
NUM|8|17|因為 以色列 人中凡頭生的，無論是人或牲畜，都是我的。我在 埃及 地擊殺所有頭生的那日，已將他們分別為聖歸我。
NUM|8|18|我選 利未 人代替 以色列 人中所有頭生的。
NUM|8|19|我從 以色列 人中將 利未 人給 亞倫 和他的兒子作為賞賜，在會幕中為 以色列 人事奉，又為 以色列 人贖罪，免得 以色列 人因挨近聖所而遭受災禍。」
NUM|8|20|摩西 、 亞倫 和 以色列 全會眾就向 利未 人這樣做。關於 利未 人，凡耶和華怎樣吩咐 摩西 ， 以色列 人就向他們照樣做了。
NUM|8|21|於是 利未 人從罪中潔淨自己，洗淨衣服。 亞倫 將他們奉獻在耶和華面前，作為搖祭，又為他們贖罪，潔淨他們。
NUM|8|22|然後 利未 人進去，在 亞倫 和他兒子面前，在會幕中事奉。關於 利未 人，耶和華怎樣吩咐 摩西 ，他們就向 利未 人照樣做了。
NUM|8|23|耶和華吩咐 摩西 說：
NUM|8|24|「這是有關 利未 人的：二十五歲以上的人都要前來任職，在會幕裏事奉。
NUM|8|25|到了五十歲，他們就要從事奉的工作中退休，不再事奉，
NUM|8|26|只可在會幕裏輔助他們的弟兄盡責，他們自己不再事奉了。關於 利未 人的職責，你要向他們這樣做。」
NUM|9|1|以色列 人出 埃及 地以後，第二年正月，耶和華在 西奈 的曠野吩咐 摩西 說：
NUM|9|2|「 以色列 人應當在所定的日期守逾越節。
NUM|9|3|你們要在本月十四日黃昏的時候 ，在所定的日期守這節，按照一切的律例典章守節。」
NUM|9|4|於是 摩西 吩咐 以色列 人守逾越節。
NUM|9|5|正月十四日黃昏的時候，他們就在 西奈 的曠野守逾越節。凡耶和華所吩咐 摩西 的， 以色列 人都照樣做了。
NUM|9|6|有幾個人因屍體成了不潔淨，不能在那日守逾越節。當天他們到 摩西 、 亞倫 面前。
NUM|9|7|那些人對他說：「我們因屍體而不潔淨，為何禁止我們，不能和 以色列 人在所定的日期獻供物給耶和華呢？」
NUM|9|8|摩西 對他們說：「你們稍等，讓我去聽耶和華對你們有甚麼吩咐。」
NUM|9|9|耶和華吩咐 摩西 說：
NUM|9|10|「你要吩咐 以色列 人說：你們和你們後代中，若有人因屍體成了不潔淨，或出外遠行，仍然要向耶和華守逾越節，
NUM|9|11|他們就要在二月十四日黃昏的時候守節，要吃羔羊，以及無酵餅和苦菜。
NUM|9|12|他們不可留一點食物到早晨；羔羊的骨頭一根也不可折斷。他們要照逾越節的一切律例守這節。
NUM|9|13|但潔淨又不出外遠行的人若不守逾越節，那人要從百姓中剪除，因為他沒有在所定的日期獻供物給耶和華，必須擔當自己的罪。
NUM|9|14|若有寄居在你們那裏的外人要向耶和華守逾越節，他要照逾越節的律例和典章做。無論是寄居的或是本地人，都用同樣的律例。」
NUM|9|15|立起帳幕的那日，有雲彩遮蓋帳幕，就是法櫃的帳幕；從晚上到早晨，雲彩在帳幕上，形狀如火。
NUM|9|16|經常都是這樣：雲彩遮蓋帳幕，夜間雲彩形狀如火。
NUM|9|17|雲彩幾時從帳幕上升， 以色列 人就幾時起行；雲彩在哪裏停住， 以色列 人就在哪裏安營。
NUM|9|18|以色列 人遵照耶和華的指示起行，也遵照耶和華的指示安營。雲彩在帳幕上停留多久，他們就留在營裏多久。
NUM|9|19|雲彩在帳幕上停留許多日子， 以色列 人就遵照耶和華的吩咐不起行。
NUM|9|20|有時雲彩在帳幕上只停了幾天，他們就遵照耶和華的指示留在營裏，也遵照耶和華的指示起行。
NUM|9|21|有時雲彩從晚上留到早晨；早晨雲彩上升，他們就起行。無論是白天是黑夜，當雲彩上升的時候，他們就要起行。
NUM|9|22|雲彩停留在帳幕上，無論是兩天，一個月，或更長的日子， 以色列 人就留在營裏不起行；但雲彩一上升，他們就起行。
NUM|9|23|他們遵照耶和華的指示安營，也遵照耶和華的指示起行。他們遵守耶和華的吩咐，是耶和華藉 摩西 所指示的話。
NUM|10|1|耶和華吩咐 摩西 說：
NUM|10|2|「你要用銀子做兩枝號筒，把它們錘出來，給你用來召集會眾，拔營起行。
NUM|10|3|吹號的時候，全會眾要到你那裏，聚集在會幕的門口。
NUM|10|4|若只吹一枝，眾領袖，就是 以色列 部隊的官長，要到你那裏聚集。
NUM|10|5|你們大聲吹號的時候，東邊安營的要起行。
NUM|10|6|第二次大聲吹號的時候，南邊安營的要起行。起行的時候，要大聲吹號；
NUM|10|7|但召集會眾的時候，你們要吹號，卻不要吹出大聲。
NUM|10|8|亞倫 子孫作祭司的要吹這號筒，作為你們世世代代永遠的定例。
NUM|10|9|當你們在自己的土地上，與欺壓你們的敵人打仗時，要用號筒吹出大聲。你們就在耶和華－你們的上帝面前得蒙記念，也必蒙拯救脫離仇敵。
NUM|10|10|在快樂的日子，節期和初一，獻燔祭與平安祭的時候，你們要吹號筒，在你們的上帝面前作為紀念。我是耶和華－你們的上帝。」
NUM|10|11|第二年二月二十日，雲彩從法櫃的帳幕上升。
NUM|10|12|以色列 人離開 西奈 的曠野，一段一段地往前行，雲彩停在 巴蘭 的曠野。
NUM|10|13|他們遵照耶和華藉 摩西 所指示的，初次往前行。
NUM|10|14|按照隊伍首先起行的是 猶大 營旗幟下的人，帶隊的是 亞米拿達 的兒子 拿順 。
NUM|10|15|以薩迦 支派帶隊的是 蘇押 的兒子 拿坦業 。
NUM|10|16|西布倫 支派帶隊的是 希倫 的兒子 以利押 。
NUM|10|17|帳幕拆卸了， 革順 的子孫和 米拉利 的子孫就抬著帳幕往前行。
NUM|10|18|按照隊伍往前行的是 呂便 營旗幟下的人，帶隊的是 示丟珥 的兒子 以利蓿 。
NUM|10|19|西緬 支派帶隊的是 蘇利沙代 的兒子 示路蔑 。
NUM|10|20|迦得 支派帶隊的是 丟珥 的兒子 以利雅薩 。
NUM|10|21|哥轄 人抬著聖物往前行。他們未到以前，帳幕已經立好了。
NUM|10|22|按照隊伍往前行的是 以法蓮 營旗幟下的人，帶隊的是 亞米忽 的兒子 以利沙瑪 。
NUM|10|23|瑪拿西 支派帶隊的是 比大蓿 的兒子 迦瑪列 。
NUM|10|24|便雅憫 支派帶隊的是 基多尼 的兒子 亞比但 。
NUM|10|25|作全營後衛，按隊伍往前行的是 但 營旗幟下的人，帶隊的是 亞米沙代 的兒子 亞希以謝 。
NUM|10|26|亞設 支派帶隊的是 俄蘭 的兒子 帕結 。
NUM|10|27|拿弗他利 支派帶隊的是 以南 的兒子 亞希拉 。
NUM|10|28|以色列 人就這樣按著隊伍往前行。
NUM|10|29|摩西 對他岳父 ， 米甸 人 流珥 的兒子 何巴 說：「我們要往前行，到耶和華所說的地方；他曾說：『我要將這地賜給你們。』現在請你和我們同去，我們必善待你，因為耶和華已經應許賜福氣給 以色列 人。」
NUM|10|30|何巴 對他說：「我不去，我要回本地本族去。」
NUM|10|31|摩西 說：「請你不要離開我們，因為你知道我們要在曠野安營，你可以當我們的眼目。
NUM|10|32|你若和我們同去，將來耶和華以甚麼福氣恩待我們，我們也必這樣善待你。」
NUM|10|33|以色列 人離開耶和華的山，往前行了三天的路程。耶和華的約櫃在前面行了三天的路程，為他們尋找安歇的地方。
NUM|10|34|他們拔營往前行，日間有耶和華的雲彩在他們上面。
NUM|10|35|約櫃往前行的時候， 摩西 說： 「耶和華啊，求你興起！ 願你的仇敵潰散！ 願恨你的人從你面前逃跑！」
NUM|10|36|約櫃停住的時候，他說： 「 以色列 千萬人的耶和華啊，求你回來 ！」
NUM|11|1|百姓發怨言，惡言傳達到耶和華的耳中。耶和華聽見了就怒氣發作，耶和華的火在他們中間焚燒，燒燬營的外圍。
NUM|11|2|百姓向 摩西 哀求， 摩西 祈求耶和華，火就熄了。
NUM|11|3|那地方就叫做 他備拉 ，因為耶和華的火曾在他們中間焚燒。
NUM|11|4|他們中間的閒雜人動了貪慾的心； 以色列 人又再哭著說：「誰給我們肉吃呢？
NUM|11|5|我們記得在 埃及 的時候，不花錢就可以吃魚，還有黃瓜、西瓜、韭菜、蔥、蒜。
NUM|11|6|現在我們的精力枯乾了。除了這嗎哪以外，在我們眼前甚麼都沒有。」
NUM|11|7|嗎哪好像芫荽子，看上去如同樹脂的樣子。
NUM|11|8|百姓四處走動撿取嗎哪，把它用磨磨碎或用臼搗成粉，在鍋中煮了做成餅，滋味好像油烤餅的滋味。
NUM|11|9|夜間露水降在營中，嗎哪也隨著降下。
NUM|11|10|摩西 聽見百姓家家戶戶在帳棚門口哀哭。因此， 耶和華的怒氣大大發作， 摩西 看了也不高興。
NUM|11|11|摩西 對耶和華說：「你為何苦待僕人？我為何不在你眼前蒙恩，竟把這眾百姓的擔子加在我身上呢？
NUM|11|12|這眾百姓豈是我懷的胎，豈是我生下來的呢？你竟對我說：『把他們抱在懷裏，如養育之父抱著吃奶的嬰孩，一直抱到你起誓應許給他們祖宗的土地去。』
NUM|11|13|我從哪裏拿肉給這眾百姓吃呢？他們都向我哭著說：『給我們肉吃！』
NUM|11|14|我不能獨自帶領這眾百姓，這對我太沉重了。
NUM|11|15|如果你這樣待我，倒不如立刻把我殺了吧！我若在你眼前蒙恩，求你不要讓我再受這樣的苦。」
NUM|11|16|耶和華對 摩西 說：「你要從 以色列 的長老中為我召集七十個人，就是你所認識，作百姓的長老和官長的，領他們到會幕，使他們和你一同站在那裏。
NUM|11|17|我要在那裏降臨，與你說話，把降給你的靈分給他們。他們就和你分擔帶領百姓的擔子，免得你獨自承擔。
NUM|11|18|你要對百姓說：『你們要為了明天使自己分別為聖，你們將有肉吃。因你們哭著說：誰給我們肉吃呢？我們在 埃及 多麼好！這聲音傳到了耶和華的耳中，所以他必給你們肉吃。
NUM|11|19|你們不只吃一天、兩天、五天、十天、二十天，
NUM|11|20|而是整整一個月，直到肉從你們的鼻孔噴出來，使你們厭惡。因為你們厭棄那住在你們中間的耶和華，在他面前哭著說：我們為何出 埃及 呢？』」
NUM|11|21|摩西 說：「跟我在一起的百姓，步行的男人就有六十萬，你還說：『我要把肉賜給他們，使他們可以整整吃一個月。』
NUM|11|22|難道宰了羊群牛群，就夠給他們嗎？或者把海中所有的魚都捕來，就夠給他們嗎？」
NUM|11|23|耶和華對 摩西 說：「耶和華的膀臂 豈是縮短了嗎？現在你要看我的話向你應驗不應驗。」
NUM|11|24|摩西 出去，把耶和華的話告訴百姓，並從百姓的長老中召集七十個人來，叫他們站在會幕的四圍。
NUM|11|25|耶和華在雲中降臨，對 摩西 說話，把降給他的靈分給那七十個長老。靈停在他們身上的時候，他們就說預言，以後卻沒有再說了。
NUM|11|26|但有兩個人仍在營裏，一個名叫 伊利達 ，一個名叫 米達 。他們本是在那些登記的人中，卻沒有到會幕那裏去。靈停在他們身上，他們就在營裏說預言。
NUM|11|27|有一個年輕人跑來告訴 摩西 說：「 伊利達 和 米達 在營裏說預言。」
NUM|11|28|嫩 的兒子 約書亞 ，年輕時就作 摩西 的助手 ，說：「請我主 摩西 禁止他們。」
NUM|11|29|摩西 對他說：「你為我的緣故嫉妒嗎？惟願耶和華的百姓都是先知，願耶和華把他的靈降在他們身上！」
NUM|11|30|於是， 摩西 回到營裏去， 以色列 的長老也回去了。
NUM|11|31|有一陣風從耶和華那裏颳起，把鵪鶉從海上颳來，散落在營地和周圍；一邊約有一天的路程，另一邊也約有一天的路程，離地面約有二肘。
NUM|11|32|百姓起來，整天整夜，甚至次日一整天，都在捕捉鵪鶉。每人至少捉到十賀梅珥，各自擺在營的四圍。
NUM|11|33|但肉在他們牙間還未咀嚼時，耶和華的怒氣向百姓發作，用極重的災禍擊殺百姓。
NUM|11|34|那地方就叫 基博羅‧哈他瓦 ，因為他們在那裏埋葬了貪慾的百姓。
NUM|11|35|百姓從 基博羅‧哈他瓦 起程，到 哈洗錄 ，就住在 哈洗錄 。
NUM|12|1|摩西 娶了 古實 女子為妻。 米利暗 和 亞倫 因他娶了 古實 女子就批評他，
NUM|12|2|他們說：「難道耶和華只與 摩西 說話嗎？他不也與我們說話嗎？」耶和華聽見了。
NUM|12|3|摩西 為人極其謙和，勝過地面上的任何人。
NUM|12|4|忽然，耶和華對 摩西 、 亞倫 和 米利暗 說：「你們三個人都出來，到會幕這裏。」他們三個人就出來了。
NUM|12|5|耶和華在雲柱中降臨，停在會幕門口，叫 亞倫 和 米利暗 。二人就出來，
NUM|12|6|耶和華說：「你們要聽我的話：你們中間若有先知，我－耶和華必在異象中向他顯現，在夢中與他說話；
NUM|12|7|但我的僕人 摩西 不是這樣，他在我全家是盡忠的。
NUM|12|8|我與他面對面說話，清清楚楚，不用謎語，他甚至看見我的形像。你們為何批評我的僕人 摩西 而不懼怕呢？」
NUM|12|9|耶和華向他們怒氣發作，就離開了。
NUM|12|10|當雲彩從帳幕上離開時，看哪， 米利暗 長了痲瘋，像雪那麼白。 亞倫 轉向 米利暗 ，看哪，她長了痲瘋。
NUM|12|11|亞倫 對 摩西 說：「我主啊，求你不要因我們愚昧，因我們犯罪，就將這罪加在我們身上。
NUM|12|12|求你不要使她像那一出母腹、肉已侵蝕了一半的死胎。」
NUM|12|13|於是 摩西 哀求耶和華說：「上帝啊，求你醫治她！」
NUM|12|14|耶和華對 摩西 說：「她父親若吐唾沫在她臉上，她豈不蒙羞七天嗎？現在要把她隔離在營外七天，然後才領她回來。」
NUM|12|15|於是 米利暗 被隔離在營外七天；百姓沒有起程，直等到 米利暗 回來。
NUM|12|16|以後百姓從 哈洗錄 起行，來到 巴蘭 的曠野安營。
NUM|13|1|耶和華吩咐 摩西 說：
NUM|13|2|「你要派人去窺探我所賜給 以色列 人的 迦南 地；每個父系支派要派一個人，是他們中間的族長。」
NUM|13|3|摩西 就遵照耶和華的指示，從 巴蘭 曠野差派他們去；他們都是 以色列 人中的領袖。
NUM|13|4|這是他們的名字： 屬 呂便 支派的， 撒刻 的兒子 沙母亞 。
NUM|13|5|屬 西緬 支派的， 何利 的兒子 沙法 。
NUM|13|6|屬 猶大 支派的， 耶孚尼 的兒子 迦勒 。
NUM|13|7|屬 以薩迦 支派的， 約色 的兒子 以迦 。
NUM|13|8|屬 以法蓮 支派的， 嫩 的兒子 何西阿 。
NUM|13|9|屬 便雅憫 支派的， 拉孚 的兒子 帕提 。
NUM|13|10|屬 西布倫 支派的， 梭底 的兒子 迦疊 。
NUM|13|11|屬 約瑟 支派，就是 瑪拿西 支派的， 穌西 的兒子 迦底 。
NUM|13|12|屬 但 支派的， 基瑪利 的兒子 亞米利 。
NUM|13|13|屬 亞設 支派的， 米迦勒 的兒子 西帖 。
NUM|13|14|屬 拿弗他利 支派的， 縛西 的兒子 拿比 。
NUM|13|15|屬 迦得 支派的， 瑪基 的兒子 臼利 。
NUM|13|16|這些是 摩西 差派去窺探那地之人的名字。 摩西 叫 嫩 的兒子 何西阿 為 約書亞 。
NUM|13|17|摩西 差派他們去窺探 迦南 地，對他們說：「你們上到 尼革夫 那裏，上到山區去，
NUM|13|18|看看那地如何：住那裏的百姓是強是弱，是多是少，
NUM|13|19|他們所住的地是好是壞，所住的城鎮是營地還是堡壘，
NUM|13|20|那地是肥沃還是貧瘠，當中有樹木沒有。你們要放膽，把那地的果子帶些回來。」那時正是葡萄初熟的季節。
NUM|13|21|他們上去窺探那地，從 尋 的曠野到 利合 ，直到 哈馬口 。
NUM|13|22|他們從 尼革夫 上去，到了 希伯崙 。在那裏有 亞衲 族的 亞希幔 人、 示篩 人和 撻買 人。 希伯崙 的建造比 埃及 的 瑣安 早七年。
NUM|13|23|他們到了 以實各谷 ，從那裏砍下葡萄樹枝，上面有一掛葡萄，兩個人用槓抬著，又帶了一些石榴和無花果。
NUM|13|24|以色列 人從那裏砍下一掛葡萄，所以那地方就叫 以實各谷 。
NUM|13|25|他們窺探那地四十天之後，就回來了。
NUM|13|26|他們來到 巴蘭 曠野的 加低斯 ， 摩西 、 亞倫 ，以及 以色列 全會眾那裏，向他們和全會眾報告，又把那地的果子給他們看。
NUM|13|27|他們告訴 摩西 說：「我們到了你派我們去的那地，果然是流奶與蜜之地；這就是那地的果子。
NUM|13|28|但是住那地的百姓很強悍，城鎮又大又堅固，我們也在那裏看見了 亞衲 族人。
NUM|13|29|亞瑪力 人住在 尼革夫 ； 赫 人、 耶布斯 人和 亞摩利 人住在山區； 迦南 人住在沿海一帶和 約旦河 旁。」
NUM|13|30|迦勒 在 摩西 面前安撫百姓，說：「我們立刻上去得那地吧！我們必能征服它。」
NUM|13|31|但那些和他同去的人卻說：「我們不能上去攻打那些百姓，因為他們比我們強大。」
NUM|13|32|於是探子中有人向 以色列 人散佈有關所窺探之地的謠言，說：「我們所走過、所窺探之地是吞沒居民之地，並且我們在那裏所看見的百姓都身材高大。
NUM|13|33|我們在那裏看見巨人，就是巨人中的 亞衲 族人。我們在自己眼中像蚱蜢一樣，而在他們眼中，我們也確是這樣。」
NUM|14|1|全會眾大聲喧嚷，那夜百姓哭號。
NUM|14|2|以色列 眾人向 摩西 和 亞倫 發怨言，全會眾對他們說：「我們寧願死在 埃及 地，寧願死在這曠野！
NUM|14|3|耶和華為甚麼要把我們領到那地，讓我們倒在刀下呢？我們的妻子和孩子必成為擄物。我們回 埃及 去豈不更好嗎？」
NUM|14|4|他們彼此說：「我們不如選一個領袖，回 埃及 去吧！」
NUM|14|5|摩西 和 亞倫 在 以色列 全會眾面前臉伏於地。
NUM|14|6|窺探那地的人中， 嫩 的兒子 約書亞 和 耶孚尼 的兒子 迦勒 撕裂衣服，
NUM|14|7|對 以色列 全會眾說：「我們所走過、所窺探之地是極美之地。
NUM|14|8|耶和華若喜愛我們，就必領我們進入那地，把這流奶與蜜之地賜給我們。
NUM|14|9|但你們不可背叛耶和華，也不要怕那地的百姓，因為他們是我們的食物。保護他們的已經離開他們，耶和華卻與我們同在。不要怕他們！」
NUM|14|10|當全會眾正說著要拿石頭打死他們的時候，耶和華的榮光在會幕中向 以色列 眾人顯現。
NUM|14|11|耶和華對 摩西 說：「這百姓藐視我要到幾時呢？我在他們中間行了這一切神蹟，他們還不信我要到幾時呢？
NUM|14|12|我要用瘟疫擊殺他們，使他們不得承受那地。我要使你成為大國，比他們強大。」
NUM|14|13|摩西 對耶和華說：「 埃及 人必聽見，因你曾施展大能，領這百姓從他們中間出來。
NUM|14|14|埃及 人要告訴這地的居民，他們已經聽見你─耶和華是在這百姓中間，因為你─耶和華面對面 顯示自己，你的雲彩停在他們以上。你日間在雲柱中，夜間在火柱中，在他們的前面行。
NUM|14|15|你若把這百姓殺了，好像殺一個人那樣，那聽見你名聲的列國必說：
NUM|14|16|『耶和華因為不能把這百姓領進他向他們起誓應許之地，所以在曠野把他們殺了。』
NUM|14|17|現在求主顯出大能，照你說過的話說：
NUM|14|18|『耶和華不輕易發怒， 且有豐盛的慈愛。 他赦免罪孽和過犯， 萬不以有罪的為無罪， 必懲罰人的罪， 從父到子，直到三、四代。』
NUM|14|19|求你照你的大慈愛赦免這百姓的罪孽，好像你從 埃及 到如今饒恕這百姓一樣。」
NUM|14|20|耶和華說：「我照著你的話赦免他們。
NUM|14|21|然而，我指著我的永生與遍地充滿了耶和華的榮耀起誓：
NUM|14|22|這些人雖然都看過我的榮耀和我在 埃及 與曠野所行的神蹟，仍然這十次試探我，不聽從我的話，
NUM|14|23|他們絕不能看見我向他們祖宗所起誓應許之地；凡藐視我的，一個也不得看見。
NUM|14|24|惟獨我的僕人 迦勒 ，因他另有一個心志，專心跟從我，我要領他進入他所去過的那地；他的後裔必得那地為業。
NUM|14|25|亞瑪力 人和 迦南 人住在谷中，明天你們要轉回去，沿著 紅海 的路往曠野去。」
NUM|14|26|耶和華對 摩西 和 亞倫 說：
NUM|14|27|「這邪惡的會眾向我發怨言要到幾時呢？ 以色列 人向我發的怨言，我都聽見了。
NUM|14|28|你要告訴他們，耶和華說：『我指著我的永生起誓，我必照你們在我耳中所說的待你們。
NUM|14|29|你們的屍體必倒在這曠野中。你們中間被數點，凡二十歲以上向我發怨言的，
NUM|14|30|必不得進我所起誓應許給你們居住的那地。惟有 耶孚尼 的兒子 迦勒 和 嫩 的兒子 約書亞 才能進去。
NUM|14|31|你們的孩子，就是你們說要成為擄物的，我必領他們進去，他們就得知你們所厭棄的那地。
NUM|14|32|至於你們，你們的屍體必倒在這曠野中；
NUM|14|33|你們的兒女必在曠野遊牧四十年，擔當你們不信的罪 ，直到你們的屍體在曠野消滅為止。
NUM|14|34|按你們窺探那地的四十日，一年抵一日，你們要擔當你們的罪孽四十年，你們就知道我疏遠你們了。』
NUM|14|35|我－耶和華說過，我必這樣對待這一切聚集對抗我的邪惡會眾。他們必在這曠野中消滅，死在這裏。」
NUM|14|36|摩西 所差派去窺探那地的人回來，散佈有關那地的謠言，使全會眾向 摩西 發怨言，
NUM|14|37|這些散佈謠言的人都遭受瘟疫，死在耶和華面前。
NUM|14|38|窺探那地的人中，惟有 嫩 的兒子 約書亞 和 耶孚尼 的兒子 迦勒 得以存活。
NUM|14|39|摩西 把這些話告訴 以色列 眾人，他們都極其悲哀。
NUM|14|40|他們清晨起來，上到山頂，說：「看哪，我們要上到耶和華所說的地方；因為我們犯了罪。」
NUM|14|41|摩西 說：「你們為何要這樣違背耶和華的指示呢？這事必不能順利。
NUM|14|42|不要上去，因為耶和華不在你們中間，恐怕你們在仇敵面前被擊敗。
NUM|14|43|亞瑪力 人和 迦南 人都在你們面前，你們必倒在刀下。因為你們背離不跟從耶和華，耶和華必不與你們同在。」
NUM|14|44|他們卻擅自上到山頂。但耶和華的約櫃和 摩西 都沒有離開營地。
NUM|14|45|於是 亞瑪力 人和住在那山區的 迦南 人下來，擊敗他們，追擊他們直到 何珥瑪 。
NUM|15|1|耶和華吩咐 摩西 說：
NUM|15|2|「你要吩咐 以色列 人，對他們說：你們到了我所賜給你們居住的地，
NUM|15|3|你們要從牛群羊群中取牲畜獻給耶和華為火祭，無論是燔祭或祭物，為要還所許特別的願或甘心祭，或節期的祭，作為獻給耶和華的馨香之祭，
NUM|15|4|那獻供物的要將十分之一伊法細麵和四分之一欣油調和作素祭，獻給耶和華。
NUM|15|5|無論是燔祭或祭物，要為每隻小綿羊預備四分之一欣酒作澆酒祭。
NUM|15|6|要為每隻公綿羊預備十分之二伊法細麵，和三分之一欣油調和作素祭，
NUM|15|7|又用三分之一欣酒作澆酒祭，獻給耶和華為馨香之祭。
NUM|15|8|你預備公牛獻給耶和華作燔祭或祭物，為要還所許特別的願，或平安祭，
NUM|15|9|就要把十分之三伊法細麵和半欣油調和作素祭，和公牛一同獻上，
NUM|15|10|又用半欣酒作澆酒祭，獻給耶和華為馨香的火祭。
NUM|15|11|「獻公牛、或公綿羊、或小綿羊、或小山羊，每隻都要這樣處理；
NUM|15|12|無論你們所獻的數目多少，照著數目每隻都要這樣處理。
NUM|15|13|凡本地人將馨香的火祭獻給耶和華，都要照樣處理。
NUM|15|14|若有外人寄居在你們那裏，或有人世世代代住在你們中間，願意將馨香的火祭獻給耶和華，你們怎樣處理，他也要照樣處理。
NUM|15|15|至於會眾，無論是你們或寄居的外人都要遵守同一條例；這是你們世世代代永遠的定例。在耶和華面前，你們怎樣，寄居的也要怎樣。
NUM|15|16|你們和寄居在你們那裏的外人要遵守同一律法，同一典章。」
NUM|15|17|耶和華吩咐 摩西 說：
NUM|15|18|「你要吩咐 以色列 人，對他們說：你們到了我領你們進去的那地，
NUM|15|19|吃那地的糧食時，要把舉祭獻給耶和華。
NUM|15|20|你們要用初熟的麥子磨麵，做成餅當舉祭獻上。你們要舉上，如同舉禾場的舉祭。
NUM|15|21|你們世世代代要用初熟的麥子磨麵，當舉祭獻給耶和華。
NUM|15|22|「你們若犯了錯，不遵守耶和華所吩咐 摩西 的這一切命令，
NUM|15|23|就是耶和華藉 摩西 一切所命令你們的，從耶和華命令的那日直到你們的世世代代，
NUM|15|24|會眾因沒有察覺而犯了無心之過，全會眾就要將一頭公牛犢作燔祭，遵照典章把素祭和澆酒祭一同獻給耶和華為馨香的祭，又要獻一隻公山羊作贖罪祭。
NUM|15|25|祭司要為 以色列 全會眾贖罪，他們就必蒙赦免，因為這是無心之過。他們要因自己的無心之過，把供物，就是向耶和華當獻的火祭和贖罪祭，帶到耶和華面前。
NUM|15|26|以色列 全會眾和寄居在他們中間的外人就必蒙赦免，因為這是眾百姓的無心之過。
NUM|15|27|「若有一個人無意中犯了罪，他就要獻一隻一歲的母山羊作贖罪祭。
NUM|15|28|這誤犯罪的人因無意中犯了罪，祭司要在耶和華面前為他贖罪，他就必蒙赦免。
NUM|15|29|以色列 中的本地人和寄居在他們中間的外人，若無意中犯了罪，都要遵守同一律法。
NUM|15|30|但那故意犯罪的人，無論是本地人是寄居的，褻瀆了耶和華，這人必從百姓中剪除。
NUM|15|31|因為他藐視耶和華的話，違背耶和華的命令，這人一定要剪除；他的罪孽要歸到自己身上。」
NUM|15|32|以色列 人還在曠野的時候，發現有一個人在安息日撿柴。
NUM|15|33|發現他撿柴的人把他帶到 摩西 、 亞倫 以及全會眾那裏。
NUM|15|34|他們把他收押在監裏，因為還不知道要怎樣懲罰他。
NUM|15|35|耶和華吩咐 摩西 說：「這人應當處死；全會眾要在營外用石頭打死他。」
NUM|15|36|於是全會眾把他帶到營外，用石頭打死他，是照耶和華所吩咐 摩西 的。
NUM|15|37|耶和華對 摩西 說：
NUM|15|38|「你吩咐 以色列 人，對他們說，他們世世代代要在衣服邊上縫繸子，並在邊上的繸子釘一條藍色帶子。
NUM|15|39|你們要佩帶這繸子，好叫你們看見它就記起耶和華一切的命令，並且遵行，不隨從自己內心和眼目的情慾而跟著行淫。
NUM|15|40|這樣，你們就必記得並遵行我一切的命令，成為聖，歸你們的上帝。
NUM|15|41|「我是耶和華－你們的上帝，曾把你們從 埃及 地領出來，要作你們的上帝。我是耶和華－你們的上帝。」
NUM|16|1|利未 的曾孫， 哥轄 的孫子， 以斯哈 的兒子 可拉 ，連同 呂便 子孫中 以利押 的兒子 大坍 和 亞比蘭 ，與 比勒 的兒子 安 ，帶了
NUM|16|2|以色列 人中的二百五十個領袖，就是有名望、從會眾中選出來的人，在 摩西 面前一同起來，
NUM|16|3|聚集攻擊 摩西 、 亞倫 ，說：「你們太過分了！全會眾人人都成為聖，耶和華也在他們中間。你們為甚麼抬高自己，在耶和華的會眾之上呢？」
NUM|16|4|摩西 聽見就臉伏於地，
NUM|16|5|對 可拉 和他所有同夥的人說：「到了早晨，耶和華必指示誰是屬他的，誰是成為聖的，就准許誰親近他。他要叫自己所揀選的人親近他。
NUM|16|6|可拉 和你所有同夥的人哪，你們要這樣做：要拿著香爐，
NUM|16|7|明天在耶和華面前把火盛在爐中，把香放在上面。耶和華揀選誰，誰就成為聖。 利未 的子孫哪，你們太過分了！」
NUM|16|8|摩西 又對 可拉 說：「 利未 的子孫，聽吧！
NUM|16|9|以色列 的上帝將你們從 以色列 會眾中分別出來，使你們親近他，在耶和華的帳幕中事奉，並且站在會眾面前替他們供職。這對你們豈是小事嗎？
NUM|16|10|耶和華已經准許你和你所有的弟兄，就是 利未 的子孫，一同親近他，你們還要求祭司的職分嗎？
NUM|16|11|所以，你和你所有同夥的人聚集是在攻擊耶和華。 亞倫 算甚麼，你們竟向他發怨言？」
NUM|16|12|摩西 派人去叫 以利押 的兒子 大坍 和 亞比蘭 。他們卻說：「我們不上去！
NUM|16|13|你把我們從流奶與蜜之地領出來，讓我們死在曠野，這豈是小事？你還要自立為王管轄我們嗎？
NUM|16|14|你根本沒有領我們到流奶與蜜之地，也沒有給我們田地和葡萄園作為產業。難道你想要挖這些人的眼睛嗎？我們不上去！」
NUM|16|15|摩西 非常生氣，就對耶和華說：「求你不要接受他們的供物。我並沒有奪過他們一匹驢，也沒有害過他們中任何一個人。」
NUM|16|16|摩西 對 可拉 說：「明天，你和你所有同夥的人，以及 亞倫 ，都要站在耶和華面前。
NUM|16|17|你們各人要拿一個香爐，把香放在上面，各人帶香爐到耶和華面前，共二百五十個；你和 亞倫 也各拿自己的香爐。」
NUM|16|18|於是他們各人拿一個香爐，盛著火，加上香，和 摩西 、 亞倫 一同站在會幕的門口。
NUM|16|19|可拉 召集全會眾到會幕門口攻擊 摩西 和 亞倫 。這時，耶和華的榮光向全會眾顯現。
NUM|16|20|耶和華吩咐 摩西 和 亞倫 說：
NUM|16|21|「你們離開這會眾，我好立刻把他們滅絕。」
NUM|16|22|摩西 、 亞倫 臉伏於地，說：「上帝，賜萬人氣息的上帝啊，一人犯罪，你就要向全會眾發怒嗎？」
NUM|16|23|耶和華吩咐 摩西 說：
NUM|16|24|「你吩咐會眾說：『你們遠離 可拉 、 大坍 和 亞比蘭 帳棚的周圍。』」
NUM|16|25|摩西 起來，到 大坍 、 亞比蘭 那裏去； 以色列 的長老也都跟著他去。
NUM|16|26|他吩咐會眾說：「你們離開這些惡人的帳棚吧！不可碰他們的任何東西，免得你們因他們一切的罪而消滅。」
NUM|16|27|於是會眾遠離了 可拉 、 大坍 和 亞比蘭 的帳棚。 大坍 和 亞比蘭 帶著妻子、兒女和小孩子出來，站在自己的帳棚門口。
NUM|16|28|摩西 說：「因這件事，你們就必知道這一切事是耶和華差派我做的，並非出於我的心意。
NUM|16|29|這些人的死若和世人無異，或者他們所遭遇的和其他人相同，那麼耶和華就不曾差派我了。
NUM|16|30|但是，倘若耶和華創作一件新事，使地開了裂口，把他們和一切屬他們的都吞下去，叫他們活活墜落陰間，你們就知道是這些人藐視了耶和華。」
NUM|16|31|摩西 剛說完這些話，他們腳下的地就裂開，
NUM|16|32|地開了裂口，把他們和他們的家眷，以及一切屬 可拉 的人和財物，都吞了下去。
NUM|16|33|他們和一切屬他們的，都活活墜落陰間；地在他們上面又合攏起來，他們就從會眾中滅亡了。
NUM|16|34|在他們四圍的 以色列 眾人聽見他們的叫聲，就都逃跑，說：「恐怕地也要把我們吞下去了！」
NUM|16|35|有火從耶和華那裏出來，吞滅了那上香的二百五十人。
NUM|16|36|耶和華吩咐 摩西 說：
NUM|16|37|「你要對 亞倫 祭司的兒子 以利亞撒 說，把香爐從火中移開，再把炭火撒在別處，因為這些香爐是分別為聖的。
NUM|16|38|要把那些犯罪自喪己命之人的香爐錘成薄片，用以包祭壇；因為這些本是他們在耶和華面前獻過，分別為聖的，可以給 以色列 人作記號。」
NUM|16|39|於是 以利亞撒 祭司把被燒死的人所獻的銅香爐拿來；它們被錘出來，用以包壇，
NUM|16|40|給 以色列 人作紀念，為要叫 亞倫 子孫之外的人不得近前來，在耶和華面前燒香，免得他和 可拉 與同他一夥的人一樣，正如耶和華藉 摩西 所吩咐的。
NUM|16|41|第二天， 以色列 全會眾都向 摩西 、 亞倫 發怨言說：「你們殺了耶和華的百姓了。」
NUM|16|42|會眾聚集攻擊 摩西 、 亞倫 的時候， 摩西 和 亞倫 轉向會幕，看哪，雲彩遮蓋會幕，耶和華的榮光顯現。
NUM|16|43|摩西 、 亞倫 就來到會幕前。
NUM|16|44|耶和華吩咐 摩西 說：
NUM|16|45|「你們離開這會眾，我好立刻把他們滅絕。」他們二人就臉伏於地。
NUM|16|46|摩西 對 亞倫 說：「拿你的香爐，把祭壇的火盛在裏面，加上香，趕快帶到會眾那裏，為他們贖罪。因為有憤怒從耶和華面前發出，瘟疫已經開始了。」
NUM|16|47|亞倫 照 摩西 所說的拿了香爐，跑到會眾中。看哪，瘟疫已經在百姓中開始了。他就加上香，為百姓贖罪。
NUM|16|48|他站在活人和死人之間，瘟疫就止住了。
NUM|16|49|除了因 可拉 事件死的以外，遭瘟疫死的共有一萬四千七百人。
NUM|16|50|亞倫 回到會幕門口 ，到 摩西 那裏，瘟疫已經止住了。
NUM|17|1|耶和華吩咐 摩西 說：
NUM|17|2|「你要吩咐 以色列 人，從他們當中取杖，每父家一根；從他們所有的領袖，按著父家，共取十二根。你要把各人的名字寫在他的杖上，
NUM|17|3|並要把 亞倫 的名字寫在 利未 的杖上，因為各父家的家長都有一根杖。
NUM|17|4|你要把這些杖放在會幕裏法櫃前，我與你們 相會的地方。
NUM|17|5|我所揀選的人，他的杖必發芽。我就平息了 以色列 人向你們所發的怨言，不再達到我這裏。」
NUM|17|6|於是， 摩西 吩咐 以色列 人，他們的眾領袖就把杖給他，一個領袖一根杖，按照父家一個領袖一根杖，共有十二根； 亞倫 的杖也在其中。
NUM|17|7|摩西 把這些杖放在耶和華面前，在法櫃的帳幕裏。
NUM|17|8|第二天， 摩西 進到法櫃的帳幕去，看哪， 利未 族 亞倫 的杖已經發芽，長了花苞，開了花，也結出熟的杏子！
NUM|17|9|摩西 把所有的杖從耶和華面前拿出來，給 以色列 眾人看。他們都看見了，各領袖就把自己的杖拿去。
NUM|17|10|耶和華吩咐 摩西 說：「把 亞倫 的杖放回法櫃前，給這些背叛之子留作記號。你就可以平息他們向我所發的怨言，他們也不會死亡。」
NUM|17|11|摩西 就照樣做了；耶和華怎樣吩咐他，他就照樣做。
NUM|17|12|以色列 人對 摩西 說：「看哪，我們死啦！我們滅亡啦！我們全都滅亡啦！
NUM|17|13|凡挨近耶和華帳幕的，就必死亡。我們都要消滅而死嗎？」
NUM|18|1|耶和華對 亞倫 說：「你和你的兒子，以及你父家的人，要一同擔當干犯聖所的罪孽；你和你的兒子也要擔當干犯祭司職分的罪孽。
NUM|18|2|你也要帶你弟兄 利未 人，就是你父系支派的人前來，與你聯合，服事你。你和你的兒子要一起在法櫃的帳幕前；
NUM|18|3|他們要遵守你的吩咐，負責看守整個帳幕，只是不可挨近聖所的器具和祭壇，免得他們和你們都死亡。
NUM|18|4|他們要與你聯合，負責看守會幕和帳幕一切的事；只是外人不可挨近你們。
NUM|18|5|你們要負責看守聖所和祭壇，免得憤怒再臨到 以色列 人。
NUM|18|6|看哪，我已從 以色列 人中選了你們的弟兄 利未 人，交給你們為賞賜，歸給耶和華，為要在會幕裏事奉。
NUM|18|7|你和你的兒子要謹守祭司的職分，負責一切關於祭壇和幔子內的事。我把祭司的職分賜給你們，作為賞賜好事奉我；凡挨近的外人必被處死。」
NUM|18|8|耶和華吩咐 亞倫 說：「看哪，我已將歸我的舉祭，就是 以色列 人一切分別為聖之物，交給你照管；我把受膏的份賜給你和你的子孫，作為永遠當得的份。
NUM|18|9|這是至聖供物中所給你的，一切獻給我為至聖的素祭、贖罪祭、贖愆祭，其中所有不被火燒的供物，都要歸你和你的子孫。
NUM|18|10|你要把它當作至聖之物吃 ；凡男丁都可以吃。你要以這祭物為聖。
NUM|18|11|這也是你的， 以色列 人所獻的舉祭和搖祭，我已賜給你和你的兒女，作為永遠當得的份；你家中任何潔淨的人都可以吃。
NUM|18|12|凡最好的新油、最好的新酒和五穀，就是 以色列 人獻給耶和華的初熟之物，我都賜給你。
NUM|18|13|凡他們從地上所帶來給耶和華的初熟之物也都要歸給你。你家中任何潔淨的人都可以吃。
NUM|18|14|以色列 中一切永獻的都必歸給你。
NUM|18|15|他們所有奉給耶和華的，無論是人是牲畜，凡頭胎的，都要歸給你；但是人的長子，一定要贖出來。不潔淨牲畜中頭生的，也要贖出來。
NUM|18|16|其中一個月以上所當贖的，要照你的估價，按聖所的舍客勒，付五舍客勒銀子將他贖回，一舍客勒是二十季拉。
NUM|18|17|但是頭生的牛，或頭生的綿羊，或頭生的山羊，卻不可贖，因為牠們都是聖的。要把牠們的血灑在祭壇上，把牠們的脂肪焚燒，當作馨香的火祭獻給耶和華。
NUM|18|18|牠們的肉必歸你，像被搖的胸、被舉的右腿歸你一樣。
NUM|18|19|凡 以色列 人所獻給耶和華聖物中的舉祭，我都賜給你和你的兒女，作為永遠當得的份。這要成為你和你的後裔在耶和華面前永遠的鹽 約。
NUM|18|20|耶和華對 亞倫 說：「你在 以色列 人的境內不可有產業，在他們中間也不可有份。在 以色列 人中，我是你的份，你的產業。
NUM|18|21|「至於 利未 的子孫，看哪，我已賜給他們 以色列 所有出產的十分之一為業，作為他們在會幕中事奉的酬勞。
NUM|18|22|以色列 人不可再挨近會幕，免得他們擔當罪而死。
NUM|18|23|惟獨 利未 人要在會幕中事奉，他們要擔當罪孽，作為你們世世代代永遠的定例。他們在 以色列 人中不可有產業；
NUM|18|24|因為 以色列 人出產的十分之一，就是獻給耶和華為舉祭的，我已賜給 利未 人為業。所以我對他們說，他們不可在 以色列 人中有產業。」
NUM|18|25|耶和華吩咐 摩西 說：
NUM|18|26|「你要吩咐 利未 人，對他們說：你們從 以色列 人中所取的十分之一，就是我給你們為業的，要從這十分之一中取十分之一，作為獻給耶和華的舉祭。
NUM|18|27|這可算為你們的舉祭，如同禾場上的穀，酒池中盛滿的酒。
NUM|18|28|這樣，從 以色列 人中所收取所有的十分之一，你們要從其中取舉祭獻給耶和華；你們要把獻給耶和華的舉祭歸給 亞倫 祭司。
NUM|18|29|你們要將給你們一切禮物中最好的，就是分別為聖的，獻給耶和華為舉祭。
NUM|18|30|你要對 利未 人說：當你們把其中最好的獻上為舉祭之後，這剩下的就算是你們禾場上的農作物，酒池中的酒。
NUM|18|31|你們和你們的家人可以在任何地方吃；這本是你們的賞賜，是你們在會幕裏事奉的酬勞。
NUM|18|32|當你們把其中最好的獻上為舉祭，就不致於因它擔當罪。你們不可玷污 以色列 人的聖物，免得死亡。」
NUM|19|1|耶和華吩咐 摩西 和 亞倫 說：
NUM|19|2|「耶和華所吩咐的律法中，其中一條律例這樣說：要吩咐 以色列 人，把一頭健康、沒有殘疾、未曾負軛的紅母牛牽到你這裏來，
NUM|19|3|交給 以利亞撒 祭司。他要把牛牽到營外，人就在他面前把牛宰了。
NUM|19|4|以利亞撒 祭司要用指頭蘸這牛的血，向會幕前面彈七次。
NUM|19|5|人要在他眼前焚燒這母牛，牛的皮、肉、血和糞都要焚燒。
NUM|19|6|祭司要把香柏木、牛膝草和朱紅色紗都丟在焚燒牛的火中。
NUM|19|7|祭司要洗衣服，用水洗身，然後才可以進營；祭司必不潔淨到晚上。
NUM|19|8|焚燒牛的人也要用水洗衣服，用水洗身，必不潔淨到晚上。
NUM|19|9|一個潔淨的人要收母牛的灰，存放在營外潔淨的地方，為 以色列 會眾留作除污穢的水之用。這是為除罪用的。
NUM|19|10|收取母牛灰的人要洗衣服，必不潔淨到晚上。這要成為 以色列 人和寄居在他們中間的外人永遠的定例。
NUM|19|11|「摸了任何人死屍的，必不潔淨七天。
NUM|19|12|那人要在第三天和第七天潔淨自己，他就潔淨了。若他不在第三天和第七天潔淨自己，他就不潔淨了。
NUM|19|13|凡摸了死屍，就是死了的人的屍體，又不潔淨自己的，就玷污了耶和華的帳幕，這人必從 以色列 中剪除；因為那除污穢的水沒有灑在他身上，他就不潔淨，污穢還在他身上。
NUM|19|14|「若有人死在帳棚裏，條例是這樣：凡進那帳棚的，和所有在帳棚裏的人，都必不潔淨七天。
NUM|19|15|凡敞開的，沒有用繩子紮好蓋子的器皿，也不潔淨。
NUM|19|16|任何人在田野裏摸了被刀殺的，或自然死的，或人的骨頭，或墳墓，就必不潔淨七天。
NUM|19|17|要為這不潔淨的人拿一些燒好的除罪灰放在器皿裏，倒上清水。
NUM|19|18|一個潔淨的人要拿牛膝草蘸在這水中，把水彈在帳棚上，和一切器皿以及帳棚內的人身上，又要彈在那摸了骨頭，或摸了被殺的或自然死的，或摸了墳墓的人身上。
NUM|19|19|那潔淨的人要在第三天和第七天把水彈在不潔淨的人身上，在第七天潔淨那人。那人要洗衣服，用水洗澡，到晚上就潔淨了。
NUM|19|20|但任何不潔淨的人，他若不潔淨自己，那人要從會中剪除，因為他玷污了耶和華的聖所，除污穢的水沒有灑在他身上，他是不潔淨的。
NUM|19|21|這要成為你們永遠的定例。此外，那彈除污穢水的人也要洗衣服。凡碰除污穢水的，必不潔淨到晚上。
NUM|19|22|不潔淨的人所摸的任何東西都不潔淨；摸了這東西的人必不潔淨到晚上。」
NUM|20|1|正月間， 以色列 全會眾到了 尋 的曠野；百姓住在 加低斯 。 米利暗 死在那裏，也葬在那裏。
NUM|20|2|會眾沒有水，就聚集反對 摩西 和 亞倫 。
NUM|20|3|百姓與 摩西 爭鬧，說：「我們恨不得與我們的弟兄一同死在耶和華面前。
NUM|20|4|你們為甚麼領耶和華的會眾到這曠野，使我們和我們的牲畜都死在這裏呢？
NUM|20|5|你們為甚麼領我們從 埃及 上來，把我們帶到這壞的地方呢？這地方不能撒種，沒有無花果樹、葡萄樹、石榴樹，也沒有水喝。」
NUM|20|6|摩西 、 亞倫 離開會眾面前，到會幕的門口，臉伏於地；耶和華的榮光向他們顯現。
NUM|20|7|耶和華吩咐 摩西 說：
NUM|20|8|「你拿著杖去，和你的哥哥 亞倫 召集會眾，在他們眼前吩咐磐石湧出水來，水就會從磐石流出，給會眾和他們的牲畜喝。」
NUM|20|9|於是 摩西 遵照耶和華所吩咐他的，從耶和華面前拿了杖去。
NUM|20|10|摩西 和 亞倫 召集會眾到磐石前。 摩西 對他們說：「聽著，你們這些悖逆的人！我們要叫這磐石流出水來給你們嗎？」
NUM|20|11|摩西 舉起手來，用杖擊打磐石兩下，就有許多水流出來，會眾和他們的牲畜都喝了。
NUM|20|12|但是耶和華對 摩西 、 亞倫 說：「因為你們不信我，沒有在 以色列 人眼前尊我為聖，所以你們必不能領這會眾進入我所要賜給他們的地去。」
NUM|20|13|這就是 米利巴 水，因 以色列 人與耶和華爭鬧，耶和華在他們面前顯為聖。
NUM|20|14|摩西 從 加低斯 差遣使者到 以東 王那裏，說：「你的弟兄 以色列 這樣說：『你知道我們所遭遇的一切困難。
NUM|20|15|我們的祖先曾下到 埃及 ，我們也在 埃及 住了很多年。然而， 埃及 人卻惡待我們和我們的祖先。
NUM|20|16|我們哀求耶和華，他垂聽了我們的聲音，差遣使者把我們從 埃及 領出來。看哪，我們到了你邊界的 加低斯城 。
NUM|20|17|求你讓我們穿越你的地。我們不走田間和葡萄園，也不喝井裏的水。我們只走王的大路，不偏左右，直到過了你的邊界。』」
NUM|20|18|但是， 以東 對他說：「你不可從我這裏穿越！否則，我要帶刀出去攻擊你。」
NUM|20|19|以色列 人對他說：「我們只上大道。如果我和我的牲畜喝了你的水，我必付錢給你。我不求別的事，只求讓我步行過去。」
NUM|20|20|以東 說：「你不可經過！」他就率領一大群軍隊，以強硬的手出來攻擊 以色列 。
NUM|20|21|這樣， 以東 不肯讓 以色列 穿越他的境內， 以色列 就轉去，離開他了。
NUM|20|22|以色列 全會眾從 加低斯 起行，到了 何珥山 。
NUM|20|23|耶和華在 以東 地邊界的 何珥山 對 摩西 、 亞倫 說：
NUM|20|24|「 亞倫 要歸到他祖先 那裏。他必不得進入我所賜給 以色列 人的地，因為你們在 米利巴 水的事上違背了我的指示。
NUM|20|25|你要帶 亞倫 和他的兒子 以利亞撒 上 何珥山 ，
NUM|20|26|把 亞倫 的聖衣脫下，給他的兒子 以利亞撒 穿上。 亞倫 必歸去，死在那裏。」
NUM|20|27|摩西 就遵照耶和華的吩咐去做，他們在全會眾的眼前上了 何珥山 。
NUM|20|28|摩西 把 亞倫 的聖衣脫下，給他的兒子 以利亞撒 穿上， 亞倫 就死在山頂那裏。於是， 摩西 和 以利亞撒 下了山。
NUM|20|29|全會眾見 亞倫 死了， 以色列 全家就為 亞倫 舉哀三十天。
NUM|21|1|住 尼革夫 的 迦南 人的 亞拉得 王，聽說 以色列 從 亞他林 路來，就和 以色列 交戰，擄去他們一些人。
NUM|21|2|以色列 向耶和華許願說：「你若把這百姓真的交在我手中，我就把他們的城鎮徹底毀滅。」
NUM|21|3|耶和華垂聽了 以色列 的聲音，把 迦南 人交出來。 以色列 就把 迦南 人和他們的城鎮徹底毀滅。因此，那地方名叫 何珥瑪 。
NUM|21|4|他們從 何珥山 起行，繞過 以東 地往 紅海 那條路走。在路上，百姓心中煩躁。
NUM|21|5|百姓向上帝和 摩西 發怨言，說：「你們為甚麼把我們從 埃及 領上來 ，使我們死在曠野呢？這裏沒有糧食，沒有水，我們厭惡這淡而無味的食物。」
NUM|21|6|耶和華派火蛇進入百姓當中去咬他們，於是 以色列 中死了許多百姓。
NUM|21|7|百姓到 摩西 那裏，說：「我們有罪了，因為我們向耶和華和你發怨言。求你向耶和華禱告，叫蛇離開我們。」於是 摩西 為百姓禱告。
NUM|21|8|耶和華對 摩西 說：「你要造一條火蛇，掛在杆子上。凡被咬的，一望這蛇就必存活。」
NUM|21|9|摩西 就造了一條銅蛇，掛在杆子上。凡被蛇咬的，一望這銅蛇就活了。
NUM|21|10|以色列 人起行，安營在 阿伯 。
NUM|21|11|又從 阿伯 起行，安營在 以耶‧亞巴琳 ，在 摩押 對面的曠野，向日出的方向。
NUM|21|12|又從那裏起行，安營在 撒烈谷 。
NUM|21|13|從那裏再起行，安營在 亞嫩河 的另一邊。這 亞嫩河 在曠野，從 亞摩利 人的境內流出來； 亞嫩河 是 摩押 的邊界，在 摩押 和 亞摩利 人之間。
NUM|21|14|所以《耶和華的戰記》中提到： 「 蘇法 的 哇哈伯 ， 亞嫩河 谷，
NUM|21|15|以及 亞珥 地區眾河床的斜坡， 都靠近 摩押 的邊境。」
NUM|21|16|以色列 人從那裏起行，到了 比珥 。從前耶和華對 摩西 說：「召集百姓，我要給他們水」，說的就是這井。
NUM|21|17|當時， 以色列 人唱這首歌： 「井啊，湧出水來！ 你們要向它歌唱！
NUM|21|18|這井是領袖用權杖所挖， 是百姓中的貴族用手杖所掘。」 以色列 人從曠野往 瑪他拿 去，
NUM|21|19|從 瑪他拿 到 拿哈列 ，從 拿哈列 到 巴末 ，
NUM|21|20|從 巴末 到 摩押 地的谷，又到那可以瞭望曠野的 毗斯迦山 頂。
NUM|21|21|以色列 差遣使者到 亞摩利 人的王 西宏 那裏，說：
NUM|21|22|「求你讓我們穿越你的地；我們不岔進田間和葡萄園，也不喝井裏的水，只走王的大道，直到過了你的邊界。」
NUM|21|23|但 西宏 不讓 以色列 人穿越他的境內，就召集他的眾百姓出到曠野，要攻擊 以色列 ，到了 雅雜 與 以色列 交戰。
NUM|21|24|以色列 人用刀殺了他，佔領了他的地，從 亞嫩河 到 雅博河 ，直到 亞捫 人的邊界，因為 亞捫 人的邊防堅固。
NUM|21|25|以色列 人奪取這裏所有的城鎮，就住在 亞摩利 人的城鎮中，包括 希實本 和所屬的一切鄉鎮 。
NUM|21|26|希實本 是 亞摩利 王 西宏 的首都； 西宏 曾與先前的 摩押 王交戰，從他手中奪取了他所有的地，直到 亞嫩河 。
NUM|21|27|所以那些作詩歌的說： 你們到 希實本 來吧； 願 西宏 的城被修造建立。
NUM|21|28|因為有火從 希實本 發出， 有火焰從 西宏 的城冒出， 燒燬了 摩押 的 亞珥 ， 亞嫩河 丘壇的主 。
NUM|21|29|摩押 啊，你有禍了！ 基抹 的百姓啊，你們滅亡了！ 基抹 的男子逃亡， 女子被擄， 交給了 亞摩利 王 西宏 。
NUM|21|30|我們射了他們； 希實本 直到 底本 盡都毀滅 。 我們劫掠，直到 挪法 ； 這 挪法 直延到 米底巴 。
NUM|21|31|這樣， 以色列 人就住在 亞摩利 人的地。
NUM|21|32|摩西 差派人去窺探 雅謝 ； 以色列 人佔領了 雅謝 附近的鄉村，趕出那裏的 亞摩利 人。
NUM|21|33|後來， 以色列 人轉回，往上 巴珊 的路去。 巴珊 王 噩 率領他的眾百姓出來，在 以得來 與他們交戰。
NUM|21|34|耶和華對 摩西 說：「不要怕他！因為我已將他和他的眾百姓，以及他的地都交在你手中。你要待他如同待住在 希實本 的 亞摩利 王 西宏 一樣。」
NUM|21|35|於是他們殺了 巴珊 王和他的眾子，以及他的眾百姓，沒有留下一個倖存者，並且佔領了他的地。
NUM|22|1|以色列 人起行，在 摩押 平原， 約旦河 東，對著 耶利哥 安營。
NUM|22|2|西撥 的兒子 巴勒 看見 以色列 向 亞摩利 人所做的一切。
NUM|22|3|摩押 因 以色列 百姓這麼多，非常懼怕。 摩押 因 以色列 人的緣故就憂懼。
NUM|22|4|摩押 對 米甸 的長老說：「現在這群人要舔盡我們四圍的一切，好像牛舔盡田間的草一樣。」 那時， 西撥 的兒子 巴勒 作 摩押 王。
NUM|22|5|他派使者往 大河 附近的 毗奪 去，到 比珥 的兒子 巴蘭 的家鄉 ，召 巴蘭 來，說：「看哪，有一群百姓從 埃及 出來；看哪，他們遮滿地面，住在我的對面。
NUM|22|6|現在請你來，為我詛咒這百姓，因為他們比我強大，或許我能打敗他們，把他們趕出此地。因為我知道，你為誰祝福，誰就得福；你詛咒誰，誰就受詛咒。」
NUM|22|7|摩押 的長老和 米甸 的長老手裏拿著占卜的禮金到 巴蘭 那裏，將 巴勒 的話告訴他。
NUM|22|8|巴蘭 對他們說：「今晚你們在這裏過夜，我必照著耶和華向我說的話給你們答覆。」 摩押 的官員就在 巴蘭 那裏住下。
NUM|22|9|上帝臨到 巴蘭 那裏，說：「你這裏的這些人是誰？」
NUM|22|10|巴蘭 對上帝說：「 摩押 王 西撥 的兒子 巴勒 送信給我：
NUM|22|11|『看哪，從 埃及 出來的百姓遮滿了地面，現在請你來，為我詛咒他們，或許我能打敗他們，把他們趕走。』」
NUM|22|12|上帝對 巴蘭 說：「你不可跟他們去，也不可詛咒這百姓，因為他們是蒙福的。」
NUM|22|13|巴蘭 早晨起來，對 巴勒 的官員說：「你們回本地去吧，因為耶和華不允許我和你們一起去。」
NUM|22|14|摩押 的官員就起來，到 巴勒 那裏，說：「 巴蘭 不肯和我們一起來。」
NUM|22|15|巴勒 又差遣比這些更多，更尊貴的官員。
NUM|22|16|他們來到 巴蘭 那裏，對他說：「 西撥 的兒子 巴勒 這樣說：『請你不要再推辭到我這裏來！
NUM|22|17|我必使你得極大的尊榮，無論你向我要甚麼，我都給你。只求你來為我詛咒這百姓。』」
NUM|22|18|巴蘭 回答 巴勒 的臣僕說：「 巴勒 就是將他滿屋的金銀給我，我也不能做任何大小的事，違背耶和華－我上帝的指示。
NUM|22|19|現在請你們今晚也在這裏住下，我好知道耶和華還要對我說甚麼。」
NUM|22|20|上帝在夜裏臨到 巴蘭 那裏，說：「這些人若來求你，你就起來跟他們去吧，只是你必須照著我對你說的話去做。」
NUM|22|21|巴蘭 早晨起來，備了驢，就和 摩押 的官員一同去了。
NUM|22|22|上帝因他去就怒氣發作；耶和華的使者站在路中間敵對他。他騎著驢，有兩個僕人跟隨他。
NUM|22|23|驢看見耶和華的使者站在路中間，手裏有拔出來的刀，就離開了路，岔入田間。 巴蘭 就打驢，要牠回到路上。
NUM|22|24|耶和華的使者站在葡萄園的窄路上，這邊有牆，那邊也有牆。
NUM|22|25|驢看見耶和華的使者，就往牆擠去，把 巴蘭 的腳擠到牆上； 巴蘭 再打驢。
NUM|22|26|耶和華的使者又往前去，站在狹窄的地方，那裏左右都無路可轉。
NUM|22|27|驢看見耶和華的使者，就伏在 巴蘭 底下。 巴蘭 怒氣發作，用杖打驢。
NUM|22|28|耶和華使驢開口，對 巴蘭 說：「我向你做了甚麼，你竟打我這三次呢？」
NUM|22|29|巴蘭 對驢說：「因為你戲弄我，我恨不得手中有刀，現在就把你殺了。」
NUM|22|30|驢對 巴蘭 說：「我不是你從小直到今天所騎的驢嗎？我平時有這樣待過你嗎？」 巴蘭 說：「沒有。」
NUM|22|31|耶和華使 巴蘭 的眼目明亮，他看見耶和華的使者站在路中間，手裏有拔出來的刀； 巴蘭 就低頭俯伏下拜。
NUM|22|32|耶和華的使者對他說：「你為甚麼這三次打你的驢呢？看哪，我出來敵對你，因為這路在我面前已經偏離了。
NUM|22|33|驢看見我就從我面前迴避了這三次；驢若沒有迴避我，我早把你殺了，留牠存活。」
NUM|22|34|巴蘭 對耶和華的使者說：「我有罪了。我不知道你站在路中間阻擋我；現在你若看為不好，我就回去。」
NUM|22|35|耶和華的使者對 巴蘭 說：「你和這些人去吧！你只要說我對你說的話。」於是 巴蘭 和 巴勒 的官員一同去了。
NUM|22|36|巴勒 聽見 巴蘭 來了，就到 摩押 的城 去迎接他；這城是在邊界的 亞嫩河 旁。
NUM|22|37|巴勒 對 巴蘭 說：「我不是急切地派人到你那裏去召你嗎？你為何不到我這裏來呢？我豈不能使你得尊榮嗎？」
NUM|22|38|巴蘭 對 巴勒 說：「看哪，我已經到你這裏來了！現在我豈能擅自說甚麼呢？上帝將甚麼話放在我口中，我就說甚麼。」
NUM|22|39|巴蘭 和 巴勒 同去，來到 基列‧胡瑣 。
NUM|22|40|巴勒 宰了牛羊為祭物，送給 巴蘭 和陪伴他的官員。
NUM|22|41|到了早晨， 巴勒 領 巴蘭 到 巴末‧巴力 ，從那裏可以看到一部分 以色列 的百姓。
NUM|23|1|巴蘭 對 巴勒 說：「你要在這裏為我築七座壇，又要在這裏為我預備七頭公牛，七隻公羊。」
NUM|23|2|巴勒 照 巴蘭 的話做了。 巴勒 和 巴蘭 在每座壇上獻一頭公牛，一隻公羊。
NUM|23|3|巴蘭 對 巴勒 說：「你站在你的燔祭旁邊，我要往前去，或許耶和華會向我顯現。他指示我甚麼事，我必告訴你。」於是 巴蘭 上到一個光禿的高地。
NUM|23|4|上帝向 巴蘭 顯現。 巴蘭 對他說：「我預備了七座壇，在每座壇上獻了一頭公牛，一隻公羊。」
NUM|23|5|耶和華把話放在 巴蘭 口中，說：「你回到 巴勒 那裏，要這樣說。」
NUM|23|6|他就回到 巴勒 那裏，看哪， 巴勒 和 摩押 的眾官員站在燔祭旁邊。
NUM|23|7|巴蘭 唱起詩歌說： 「 巴勒 領我出 亞蘭 ， 摩押 王領我出東方的山脈： 『來啊，為我詛咒 雅各 ； 來啊，怒罵 以色列 。』
NUM|23|8|上帝沒有詛咒的， 我焉能詛咒？ 耶和華沒有怒罵的， 我豈能怒罵？
NUM|23|9|我從磐石的巔峰看到他， 我從山丘望見他。 看哪，這是獨居的民， 不算在列國中。
NUM|23|10|誰能數點 雅各 的塵土？ 誰能計算 以色列 的塵沙 ？ 我願如正直人之死而死； 我願如正直人之終而終。」
NUM|23|11|巴勒 對 巴蘭 說：「你向我做的是甚麼呢？我帶你來詛咒我的仇敵，看哪，你竟為他們祝福。」
NUM|23|12|他回答說：「耶和華放在我口中的話，我豈能不謹慎地說呢？」
NUM|23|13|巴勒 對他說：「請你跟我到別的地方，在那裏可以看見他們。你只能看見他們的一部分，卻不能看見全部。請你在那裏為我詛咒他們。」
NUM|23|14|於是 巴勒 領 巴蘭 到了 瑣腓 的田野，上了 毗斯迦山 頂 ，築了七座壇，在每座壇上獻一頭公牛，一隻公羊。
NUM|23|15|巴蘭 對 巴勒 說：「你站在你的燔祭旁邊，我要到那邊去看看。」
NUM|23|16|耶和華向 巴蘭 顯現，把話放在他口中，說：「你回到 巴勒 那裏，要這樣說。」
NUM|23|17|他回到 巴勒 那裏，看哪， 巴勒 站在燔祭旁邊， 摩押 的官員也和他在一起。 巴勒 對他說：「耶和華說了甚麼呢？」
NUM|23|18|巴蘭 唱起詩歌說： 「 巴勒 啊，起來，聽； 西撥 的兒子啊，側耳聽我。
NUM|23|19|上帝非人，必不致說謊， 也非人子，必不致後悔。 他說了豈不照著做呢？ 他發了言豈不實現呢？
NUM|23|20|看哪，我奉命祝福； 上帝賜福，我不能扭轉。
NUM|23|21|他未見 雅各 中有災難 ， 也未見 以色列 中有禍患 。 耶和華－他的上帝和他同在； 在他中間有歡呼王的聲音。
NUM|23|22|上帝領他們出 埃及 ， 為 以色列 有如野牛的角。
NUM|23|23|絕沒有法術可以傷 雅各 ， 沒有占卜可以害 以色列 。 現在，人論及 雅各 ，論及 以色列 必說： 『上帝成就了何等的事啊！』
NUM|23|24|看哪，這百姓興起如母獅， 挺身像公獅， 未曾吃獵物， 未曾喝被殺者的血， 絕不躺臥。」
NUM|23|25|巴勒 對 巴蘭 說：「你一點也不要詛咒他們，一點也不要為他們祝福！」
NUM|23|26|巴蘭 回答 巴勒 說：「我不是告訴過你：『凡耶和華所說的，我必須遵行』嗎？」
NUM|23|27|巴勒 對 巴蘭 說：「來，我領你到別的地方，或許上帝喜歡你在那裏為我詛咒他們。」
NUM|23|28|巴勒 就領 巴蘭 到那可瞭望曠野的 毗珥山 頂。
NUM|23|29|巴蘭 對 巴勒 說：「你要在這裏為我築七座壇，又要在這裏為我預備七頭公牛，七隻公羊。」
NUM|23|30|巴勒 就照 巴蘭 的話做，在每座壇上獻一頭公牛，一隻公羊。
NUM|24|1|巴蘭 見耶和華喜歡賜福給 以色列 ，就不像前兩次去求法術，卻面向曠野。
NUM|24|2|巴蘭 舉目，看見 以色列 人照著支派紮營。上帝的靈就臨到他身上，
NUM|24|3|他唱起詩歌說： 「 比珥 的兒子 巴蘭 說， 眼目關閉 的人說，
NUM|24|4|聽見上帝的言語， 得見全能者的異象， 俯伏著，眼睛卻睜開的人說：
NUM|24|5|雅各 啊，你的帳棚何等華美！ 以色列 啊，你的帳幕何其華麗！
NUM|24|6|如連綿的山谷， 如河畔的園子， 如耶和華栽種的沉香樹， 又如水邊的香柏木。
NUM|24|7|水要從他的桶裏流出， 種子要撒在多水之處。 他的王必超越 亞甲 ， 他的國必要振興。
NUM|24|8|上帝領他出 埃及 ， 為他有如野牛的角。 他要吞滅那敵對他的國， 壓碎他們的骨頭， 用箭射透他們。
NUM|24|9|他蹲如公獅， 臥如母獅， 誰敢惹他？ 凡為你祝福的，願他蒙福； 凡詛咒你的，願他受詛咒。」
NUM|24|10|巴勒 向 巴蘭 怒氣發作，就緊握拳頭 。 巴勒 對 巴蘭 說：「我召你來詛咒我的仇敵，看哪，你竟然這三次為他們祝福。
NUM|24|11|如今你趕快回本地去吧！我想使你大得尊榮，看哪，耶和華卻阻止你得尊榮。」
NUM|24|12|巴蘭 對 巴勒 說：「我不是對你所差遣到我那裏的使者說：
NUM|24|13|『 巴勒 就是把他滿屋的金銀給我，我也不能違背耶和華的指示，隨自己的心意做好做歹。耶和華說甚麼，我就說甚麼。』
NUM|24|14|現在，看哪，我要回到我的百姓那裏。來，讓我告訴你這百姓日後要怎樣對待你的百姓。」
NUM|24|15|他就唱起詩歌說： 「 比珥 的兒子 巴蘭 說， 眼目關閉的人說，
NUM|24|16|聽見上帝的言語， 明白至高者的知識， 看見全能者的異象， 俯伏著，眼睛卻睜開的人說：
NUM|24|17|我看見他，卻不在現時； 我望見他，卻不在近處。 有星出於 雅各 ， 有杖從 以色列 興起， 必打破 摩押 的額頭， 必毀壞所有的 塞特 人 。
NUM|24|18|以東 將成為產業， 西珥 將成為它敵人的產業 ； 但 以色列 卻要得勝。
NUM|24|19|有一位出於 雅各 的，必掌大權， 他要除滅城中的倖存者。」
NUM|24|20|巴蘭 看見 亞瑪力 人，就唱起詩歌說： 「 亞瑪力 是諸國之首， 但它終必永遠沉淪 。」
NUM|24|21|巴蘭 看見 基尼 人，就唱起詩歌說： 「你的住處堅固； 你的巢窩造在巖石中。
NUM|24|22|然而 基尼 族 必被吞滅， 直到何時 亞述 把你擄去？ 」
NUM|24|23|巴蘭 又唱起詩歌說： 「哀哉！若上帝做這事， 誰能存活呢？
NUM|24|24|有船隻 從 基提 邊界來到， 要壓制 亞述 ， 要壓制 希伯 ； 他也必永遠沉淪 。」
NUM|24|25|於是 巴蘭 起來，回本地去； 巴勒 也回他的路去了。
NUM|25|1|以色列 人住在 什亭 ，百姓開始與 摩押 女子行淫。
NUM|25|2|這些女子請百姓一同為她們的神明獻祭，百姓吃了祭物，跪拜她們的神明。
NUM|25|3|以色列 與 巴力‧毗珥 聯合，耶和華的怒氣就向 以色列 發作。
NUM|25|4|耶和華對 摩西 說：「拿下百姓中所有的領袖，對著太陽把他們懸掛在我面前，使我向 以色列 所發的怒氣可以平息。」
NUM|25|5|於是 摩西 對 以色列 的審判官說：「你們的人若有與 巴力‧毗珥 聯合的，你們各人就要把他們殺了。」
NUM|25|6|摩西 和 以色列 全會眾在會幕門口哭泣的時候，看哪，有一個 以色列 人，在他們眼前帶著一個 米甸 女子，到他弟兄那裏。
NUM|25|7|亞倫 祭司的孫子， 以利亞撒 的兒子 非尼哈 看見了，就從會眾中起來，手裏拿著槍，
NUM|25|8|跟這 以色列 人進入帳棚，刺穿了二人，就是 以色列 人和那女子的肚腹。這樣， 以色列 人遭受的瘟疫就停止了。
NUM|25|9|遭瘟疫死的，有二萬四千人。
NUM|25|10|耶和華吩咐 摩西 說：
NUM|25|11|「 亞倫 祭司的孫子， 以利亞撒 的兒子 非尼哈 ，使我的憤怒轉離 以色列 人，因為在他們中間，他以我的妒忌為他的妒忌，使我不在妒忌中毀滅 以色列 人。
NUM|25|12|因此，你要說：『看哪，我將我平安的約賜給他。
NUM|25|13|這是他和他的後裔永遠當祭司職任的約，因他為了上帝而妒忌，他為 以色列 人贖罪。』」
NUM|25|14|那與 米甸 女子一起被殺的 以色列 人，名叫 心利 ，是 撒路 的兒子，是 西緬 一個父家的領袖。
NUM|25|15|那被殺的 米甸 女子，名叫 哥斯比 ，是 蘇珥 的女兒； 蘇珥 是 米甸 一個父家的領袖。
NUM|25|16|耶和華吩咐 摩西 說：
NUM|25|17|「你要苦害 米甸 人，擊殺他們；
NUM|25|18|因為他們用詭計苦害你們，在 毗珥 的事上和他們的姊妹， 米甸 領袖的女兒 哥斯比 的事上，欺騙了你們；在瘟疫的日子，這女子因 毗珥 的事件被殺了。」
NUM|26|1|瘟疫過了之後，耶和華對 摩西 和 亞倫 祭司的兒子 以利亞撒 說：
NUM|26|2|「你們要將 以色列 全會眾，按他們的父家，凡二十歲以上能出去為 以色列 打仗的，計算總數。」
NUM|26|3|摩西 和 以利亞撒 祭司在 摩押 平原與 耶利哥 相對的 約旦河 邊吩咐他們說：
NUM|26|4|「計算你們中間從二十歲以上的人數。」正如耶和華所吩咐 摩西 的。 從 埃及 地出來的 以色列 人如下：
NUM|26|5|以色列 的長子是 呂便 。 呂便 的眾子：屬 哈諾 的，有 哈諾 族；屬 法路 的，有 法路 族；
NUM|26|6|屬 希斯倫 的，有 希斯倫 族；屬 迦米 的，有 迦米 族。
NUM|26|7|這就是 呂便 的各族；被數的共有四萬三千七百三十名。
NUM|26|8|法路 的兒子是 以利押 。
NUM|26|9|以利押 的兒子是 尼母利 、 大坍 、 亞比蘭 。這 大坍 、 亞比蘭 ，就是從會中選出來，當 可拉 一夥的人向耶和華爭鬧的時候，一起向 摩西 、 亞倫 爭鬧的；
NUM|26|10|地開了裂口，吞了他們和 可拉 ， 可拉 一夥的人也一同死亡。當時火吞滅了二百五十個人；他們就成為鑑戒。
NUM|26|11|然而 可拉 的眾子沒有死亡。
NUM|26|12|按著宗族， 西緬 的眾子：屬 尼母利 的，有 尼母利 族；屬 雅憫 的，有 雅憫 族；屬 雅斤 的，有 雅斤 族；
NUM|26|13|屬 謝拉 的，有 謝拉 族；屬 掃羅 的，有 掃羅 族。
NUM|26|14|這就是 西緬 的各族，共有二萬二千二百名。
NUM|26|15|按著宗族， 迦得 的眾子：屬 洗分 的，有 洗分 族；屬 哈基 的，有 哈基 族；屬 書尼 的，有 書尼 族；
NUM|26|16|屬 阿斯尼 的，有 阿斯尼 族；屬 以利 的，有 以利 族；
NUM|26|17|屬 亞律 的，有 亞律 族；屬 亞列利 的，有 亞列利 族。
NUM|26|18|這就是 迦得 子孫的各族；他們被數的共有四萬零五百名。
NUM|26|19|猶大 的兒子是 珥 和 俄南 。 珥 和 俄南 死在 迦南 地。
NUM|26|20|按著宗族， 猶大 的眾子：屬 示拉 的，有 示拉 族；屬 法勒斯 的，有 法勒斯 族；屬 謝拉 的，有 謝拉 族。
NUM|26|21|法勒斯 的眾子：屬 希斯崙 的，有 希斯崙 族；屬 哈母勒 的，有 哈母勒 族。
NUM|26|22|這就是 猶大 的各族；他們被數的共有七萬六千五百名。
NUM|26|23|按著宗族， 以薩迦 的眾子：屬 陀拉 的，有 陀拉 族；屬 普瓦 的，有 普瓦 族；
NUM|26|24|屬 雅述 的，有 雅述 族；屬 伸崙 的，有 伸崙 族。
NUM|26|25|這就是 以薩迦 的各族；他們被數的共有六萬四千三百名。
NUM|26|26|按著宗族， 西布倫 的眾子：屬 西烈 的，有 西烈 族；屬 以倫 的，有 以倫 族；屬 雅利 的，有 雅利 族。
NUM|26|27|這就是 西布倫 的各族；他們被數的共有六萬零五百名。
NUM|26|28|按著宗族， 約瑟 的兒子有 瑪拿西 、 以法蓮 。
NUM|26|29|瑪拿西 的眾子：屬 瑪吉 的，有 瑪吉 族； 瑪吉 生 基列 ；屬 基列 的，有 基列 族。
NUM|26|30|這就是 基列 的眾子：屬 伊以謝 的，有 伊以謝 族；屬 希勒 的，有 希勒 族；
NUM|26|31|屬 亞斯烈 的，有 亞斯烈 族；屬 示劍 的，有 示劍 族；
NUM|26|32|屬 示米大 的，有 示米大 族；屬 希弗 的，有 希弗 族。
NUM|26|33|希弗 的兒子 西羅非哈 沒有兒子，只有女兒。 西羅非哈 的女兒的名字是 瑪拉 、 挪阿 、 曷拉 、 密迦 、 得撒 。
NUM|26|34|這就是 瑪拿西 的各族；他們被數的共有五萬二千七百名。
NUM|26|35|這就是按著宗族， 以法蓮 的眾子：屬 書提拉 的，有 書提拉 族；屬 比結 的，有 比結 族；屬 他罕 的，有 他罕 族。
NUM|26|36|這就是 書提拉 的眾子：屬 以蘭 的，有 以蘭 族。
NUM|26|37|這就是 以法蓮 子孫的各族；他們被數的共有三萬二千五百名。按著宗族，以上這些都是 約瑟 的子孫。
NUM|26|38|按著宗族， 便雅憫 的眾子：屬 比拉 的，有 比拉 族；屬 亞實別 的，有 亞實別 族；屬 亞希蘭 的，有 亞希蘭 族；
NUM|26|39|屬 書反 的，有 書反 族；屬 戶反 的，有 戶反 族。
NUM|26|40|比拉 的兒子是 亞勒 、 乃幔 ；屬 亞勒 的 ，有 亞勒 族；屬 乃幔 的，有 乃幔 族。
NUM|26|41|按著宗族，這就是 便雅憫 的子孫；他們被數的共有四萬五千六百名。
NUM|26|42|這就是按著宗族， 但 的眾子：屬 書含 的，有 書含 族。按著宗族，這就是 但 的各族。
NUM|26|43|按照他們被數的， 書含 全宗族共有六萬四千四百名。
NUM|26|44|按著宗族， 亞設 的眾子：屬 音拿 的，有 音拿 族；屬 亦施韋 的，有 亦施韋 族；屬 比利亞 的，有 比利亞 族。
NUM|26|45|比利亞 的眾子：屬 希別 的，有 希別 族；屬 瑪結 的，有 瑪結 族。
NUM|26|46|亞設 的女兒名叫 西拉 。
NUM|26|47|這就是 亞設 子孫的各族；他們被數的共有五萬三千四百名。
NUM|26|48|按著宗族， 拿弗他利 的眾子：屬 雅薛 的，有 雅薛 族；屬 沽尼 的，有 沽尼 族；
NUM|26|49|屬 耶色 的，有 耶色 族；屬 示冷 的，有 示冷 族。
NUM|26|50|按著宗族，這就是 拿弗他利 的各族；他們被數的共有四萬五千四百名。
NUM|26|51|這就是 以色列 人中被數的，共有六十萬零一千七百三十名。
NUM|26|52|耶和華吩咐 摩西 說：
NUM|26|53|「你要按著人名的數目，將地分給這些人為產業。
NUM|26|54|人多的要多給他們產業，人少的要少給他們產業；各照被數的人數分配產業。
NUM|26|55|此外，要以抽籤來分地，按著父系各支派的名字承受產業。
NUM|26|56|要根據抽籤，看人數的多寡，給他們分配產業。」
NUM|26|57|這就是按著宗族，被數的 利未 人：屬 革順 的，有 革順 族；屬 哥轄 的，有 哥轄 族；屬 米拉利 的，有 米拉利 族。
NUM|26|58|這就是 利未 的宗族： 立尼 族、 希伯倫 族、 瑪利 族、 母示 族、 可拉 族。 哥轄 生 暗蘭 。
NUM|26|59|暗蘭 的妻子名叫 約基別 ，是 利未 的女兒，是 利未 在 埃及 所生的。她給 暗蘭 生了 亞倫 、 摩西 ，和他們的姊姊 米利暗 。
NUM|26|60|亞倫 生 拿答 、 亞比戶 、 以利亞撒 、 以他瑪 。
NUM|26|61|拿答 、 亞比戶 在耶和華面前獻凡火的時候死了。
NUM|26|62|利未 人中，凡一個月以上所有被數的男子，共有二萬三千名。他們沒有數在 以色列 人中；因為在 以色列 人中，沒有分給他們產業。
NUM|26|63|這些是 摩西 和 以利亞撒 祭司所數的；他們在 摩押 平原與 耶利哥 相對的 約旦河 邊數點 以色列 人。
NUM|26|64|這些被數的人中，沒有一個是 摩西 和 亞倫 祭司先前在 西奈 曠野所數的 以色列 人，
NUM|26|65|因為耶和華論到他們說：「他們必死在曠野。」所以，除了 耶孚尼 的兒子 迦勒 和 嫩 的兒子 約書亞 以外，他們一個也沒有存留。
NUM|27|1|約瑟 的兒子 瑪拿西 的宗族中，有 瑪拿西 的玄孫， 瑪吉 的曾孫， 基列 的孫子， 希弗 的兒子 西羅非哈 的女兒，名叫 瑪拉 、 挪阿 、 曷拉 、 密迦 、 得撒 。她們前來，
NUM|27|2|站在會幕門口，在 摩西 和 以利亞撒 祭司，以及眾領袖與全會眾面前，說：
NUM|27|3|「我們的父親死在曠野。他沒有與 可拉 同夥聚集攻擊耶和華，是在自己的罪中死的；他沒有兒子。
NUM|27|4|為甚麼因我們的父親沒有兒子就把他的名從他族中除掉呢？求你們在我們父親的兄弟中分給我們產業。」
NUM|27|5|於是， 摩西 將她們的案件呈到耶和華面前。
NUM|27|6|耶和華對 摩西 說：
NUM|27|7|「 西羅非哈 的女兒說得有理。你定要在她們父親的兄弟中，把地分給她們為業，把她們父親的產業傳給她們。
NUM|27|8|你也要吩咐 以色列 人說：『人死了，若沒有兒子，就要把他的產業傳給他的女兒。
NUM|27|9|他若沒有女兒，就要把他的產業給他的兄弟。
NUM|27|10|他若沒有兄弟，就要把他的產業給他父親的兄弟。
NUM|27|11|他父親若沒有兄弟，就要把他的產業給他族中最近的親屬繼承為業。』」這要作 以色列 人的律例典章，是照耶和華所吩咐 摩西 的。
NUM|27|12|耶和華對 摩西 說：「你上這 亞巴琳山脈 ，看我所賜給 以色列 人的地。
NUM|27|13|看了以後，你也必歸到你祖先 那裏，像你哥哥 亞倫 歸去一樣。
NUM|27|14|因為你們在 尋 的曠野，當會眾爭鬧的時候，違背了我的命令，在取水之事上沒有在會眾眼前尊我為聖。」這水就是 尋 的曠野中， 加低斯 的 米利巴 水。
NUM|27|15|摩西 對耶和華說：
NUM|27|16|「願耶和華，賜萬人氣息的上帝，立一個人治理會眾，
NUM|27|17|可以在他們面前出入，引導他們進出，免得耶和華的會眾如同沒有牧人的羊群一般。」
NUM|27|18|耶和華對 摩西 說：「 嫩 的兒子 約書亞 是一個有聖靈的人；你要領他來，為他按手，
NUM|27|19|使他站在 以利亞撒 祭司和全會眾面前，在他們眼前委派他，
NUM|27|20|又將你的尊榮給他一些，好使 以色列 全會眾都聽從他。
NUM|27|21|他要站在 以利亞撒 祭司面前； 以利亞撒 要憑烏陵的判斷，在耶和華面前為他求問。他和 以色列 全會眾都要照 以利亞撒 的指示出入。」
NUM|27|22|於是 摩西 照耶和華所吩咐他的，將 約書亞 領來，使他站在 以利亞撒 祭司和全會眾面前，
NUM|27|23|為他按手，委派他，是照耶和華藉 摩西 所說的。
NUM|28|1|耶和華吩咐 摩西 說：
NUM|28|2|「你要吩咐 以色列 人說：『你們要按時把我的供物，就是獻給我作馨香火祭的食物，獻給我。』
NUM|28|3|要對他們說：『這是當獻給耶和華的火祭：每天兩隻沒有殘疾一歲的小公羊，作為經常獻的燔祭。
NUM|28|4|早晨獻第一隻小公羊，黃昏獻第二隻小公羊；
NUM|28|5|又用十分之一伊法細麵和四分之一欣搗成的油，調和作為素祭。
NUM|28|6|這是在 西奈山 上規定為經常獻的燔祭，是獻給耶和華為馨香的火祭。
NUM|28|7|為每隻小公羊，要有四分之一欣的澆酒祭；在聖所中，你要將醇酒獻給耶和華作澆酒祭。
NUM|28|8|黃昏你獻第二隻小公羊，要照早晨的素祭和同獻的澆酒祭獻上，作為馨香的火祭，獻給耶和華。』」
NUM|28|9|「在安息日，要獻兩隻沒有殘疾，一歲的小公羊、十分之二伊法調了油的細麵為素祭，和同獻的澆酒祭。
NUM|28|10|除了經常獻的燔祭和同獻的澆酒祭之外，這是每一個安息日當獻的燔祭。」
NUM|28|11|「每月初一，要將兩頭公牛犢、一隻公綿羊、七隻沒有殘疾一歲的小公羊，獻給耶和華為燔祭。
NUM|28|12|為每頭公牛，要用十分之三伊法調了油的細麵作為素祭；為那隻公綿羊，要用十分之二伊法調了油的細麵作為素祭；
NUM|28|13|為每隻小公羊，要用十分之一伊法調了油的細麵作為素祭。這是馨香的燔祭，是獻給耶和華的火祭。
NUM|28|14|每頭公牛要有半欣的澆酒祭，每隻公綿羊三分之一欣的澆酒祭，每隻小公羊四分之一欣的澆酒祭。這是一年之中每月初一當獻的燔祭。
NUM|28|15|除了經常獻的燔祭和同獻的澆酒祭之外，又要將一隻公山羊，獻給耶和華為贖罪祭。」
NUM|28|16|「正月十四日是向耶和華守的逾越節。
NUM|28|17|這月十五日是節期，要吃無酵餅七日。
NUM|28|18|第一日要有聖會，任何勞動的工都不可做。
NUM|28|19|要把火祭，就是兩頭公牛犢，一隻公綿羊、七隻一歲的小公羊，都要沒有殘疾的，獻給耶和華為燔祭。
NUM|28|20|要同時獻調了油的細麵為素祭：每頭公牛要獻十分之三伊法；每隻公綿羊要獻十分之二伊法；
NUM|28|21|為那七隻小公羊，每隻要獻十分之一伊法。
NUM|28|22|此外，要獻一隻公山羊作贖罪祭，為你們贖罪。
NUM|28|23|除了早晨經常獻的燔祭之外，你們也要獻這些祭。
NUM|28|24|一連七天，在經常獻的燔祭和同獻的澆酒祭之外，每天要這樣把馨香火祭的食物獻給耶和華。
NUM|28|25|第七日要有聖會，任何勞動的工都不可做。」
NUM|28|26|「七七初熟節，就是你們獻初熟穀物給耶和華為素祭的那一天，要宣告聖會；任何勞動的工都不可做。
NUM|28|27|要將兩頭公牛犢，一隻公綿羊，七隻一歲的小公羊，作為馨香的燔祭獻給耶和華。
NUM|28|28|要同時獻調了油的細麵為素祭：每頭公牛要獻十分之三伊法；每隻公綿羊要獻十分之二伊法；
NUM|28|29|為那七隻小公羊，每隻要獻十分之一伊法。
NUM|28|30|此外，要獻一隻公山羊為你們贖罪。
NUM|28|31|除了經常獻的燔祭和同獻的素祭，你們也要獻上這些沒有殘疾的，和同獻的澆酒祭。」
NUM|29|1|「七月初一，你們當有聖會；任何勞動的工都不可做，是你們當守為吹角的日子。
NUM|29|2|你們要將一頭公牛犢、一隻公綿羊、七隻一歲的小公羊，都是沒有殘疾的，獻給耶和華為馨香的燔祭。
NUM|29|3|要同時獻調了油的細麵為素祭：每頭公牛要獻十分之三伊法；每隻公綿羊要獻十分之二伊法；
NUM|29|4|為那七隻小公羊，每隻要獻十分之一伊法。
NUM|29|5|此外，要獻一隻公山羊作贖罪祭，為你們贖罪。
NUM|29|6|除了初一的燔祭和同獻的素祭、經常獻的燔祭與同獻的素祭，以及同獻的澆酒祭以外，這些都照例作為馨香的火祭獻給耶和華。」
NUM|29|7|「七月初十，你們當有聖會；要刻苦己心，任何工都不可做。
NUM|29|8|要將一頭公牛犢、一隻公綿羊、七隻一歲的小公羊，都是沒有殘疾的，獻給耶和華為馨香的燔祭。
NUM|29|9|要同時獻調了油的細麵為素祭：每頭公牛要獻十分之三伊法；每隻公綿羊要獻十分之二伊法；
NUM|29|10|為那七隻小公羊，每隻要獻十分之一伊法。
NUM|29|11|又要獻一隻公山羊為贖罪祭。這是在贖罪祭和經常獻的燔祭，以及同獻的素祭和澆酒祭以外所獻的。」
NUM|29|12|「七月十五日，你們當有聖會；任何勞動的工都不可做，要向耶和華守節七天。
NUM|29|13|要將十三頭公牛犢、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，獻上作火祭，是獻給耶和華馨香的燔祭。
NUM|29|14|要同時獻調了油的細麵為素祭：為那十三頭公牛犢，每頭要獻十分之三伊法；為那兩隻公綿羊，每隻要獻十分之二伊法；
NUM|29|15|為那十四隻小公羊，每隻要獻十分之一伊法。
NUM|29|16|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|17|「第二日要獻十二頭公牛犢、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，
NUM|29|18|並為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|19|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|20|「第三日要獻十一頭公牛、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，
NUM|29|21|並為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|22|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|23|「第四日要獻十頭公牛、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，
NUM|29|24|並為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|25|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|26|「第五日要獻九頭公牛、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，
NUM|29|27|並為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|28|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|29|「第六日要獻八頭公牛、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，
NUM|29|30|並為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|31|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|32|「第七日要獻七頭公牛、兩隻公綿羊、十四隻一歲的小公羊，都是沒有殘疾的，
NUM|29|33|並為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|34|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|35|「第八日你們當有嚴肅會；任何勞動的工都不可做；
NUM|29|36|要將一頭公牛、一隻公綿羊、七隻一歲的小公羊，都是沒有殘疾的，獻上作火祭，是獻給耶和華馨香的燔祭。
NUM|29|37|要為公牛、公綿羊和小公羊，按數照例奉獻同獻的素祭和澆酒祭。
NUM|29|38|又要獻一隻公山羊為贖罪祭。這是在經常獻的燔祭、同獻的素祭和澆酒祭以外所獻的。
NUM|29|39|「這些祭要在你們的節期獻給耶和華，都是在所許的願和甘心獻的以外所獻的，作為你們的燔祭、素祭、澆酒祭和平安祭。」
NUM|29|40|於是， 摩西 照耶和華所吩咐他的一切話告訴 以色列 人。
NUM|30|1|摩西 對 以色列 各支派的領袖說：「這是耶和華所吩咐的話：
NUM|30|2|人若向耶和華許願或起誓，要約束自己，就不可食言，必須照口中所出的一切話去做。
NUM|30|3|女子年輕，還在父家的時候，若向耶和華許願，要約束自己，
NUM|30|4|她父親聽見她所許的願和約束自己的話，卻向她默默不言，她所許的願和約束自己的話就都有效。
NUM|30|5|但是，若她父親在聽見的日子不允許她一切所許的願和約束自己的話，這就不算為有效；耶和華也必赦免她，因為她的父親不允許。
NUM|30|6|她若已出嫁，有願在身，或口中出了約束自己的冒失話，
NUM|30|7|她丈夫聽見了，卻在聽見的日子向她默默不言，她所許的願和約束自己的話就都有效。
NUM|30|8|但是，若她丈夫在聽見的日子不允許，丈夫就廢了她所許的願和口中所出約束自己的冒失話；耶和華也必赦免她。
NUM|30|9|寡婦或被休的婦人所許的願，她所有約束自己的話，都是有效的。
NUM|30|10|她若在丈夫家裏許了願或起了誓，要約束自己，
NUM|30|11|丈夫聽見了，卻向她默默不言，沒有不允許，她所許的願和約束自己的話就都有效。
NUM|30|12|她丈夫聽見的日子，若把這些全廢了，她口中一切所許的願或約束自己的話就不算為有效。她丈夫已把這些都廢了，耶和華也必赦免她。
NUM|30|13|凡她所許的願和刻苦約束自己所起的誓，丈夫可以堅立，也可以廢去。
NUM|30|14|倘若她丈夫天天向她默默不言，這就算是堅立她一切所許的願或約束自己的話；因為丈夫在聽見的日子向她默默不言，就算是堅立了這些話。
NUM|30|15|但她丈夫聽見了，以後若再廢了這些話，就要擔當婦人的罪孽。」
NUM|30|16|這是關於丈夫待妻子，父親待女兒，女兒年輕還在父家，耶和華所吩咐 摩西 的條例。
NUM|31|1|耶和華吩咐 摩西 說：
NUM|31|2|「你要為 以色列 人向 米甸 人報仇，然後歸到你祖先 那裏。」
NUM|31|3|摩西 吩咐百姓說：「要在你們中間叫人帶兵器去攻擊 米甸 ，為耶和華向 米甸 報仇。
NUM|31|4|從 以色列 眾支派中，每支派要派一千人去打仗。」
NUM|31|5|於是從 以色列 千萬人中，每支派徵召一千人，一共一萬二千名，帶著兵器預備打仗。
NUM|31|6|摩西 派他們去打仗，每支派一千人；又派 以利亞撒 祭司的兒子 非尼哈 同去； 非尼哈 手裏拿著聖所的器皿和吹號的號筒。
NUM|31|7|他們遵照耶和華所吩咐 摩西 的，與 米甸 打仗，殺了所有的男丁。
NUM|31|8|在所殺的人中，他們殺了 米甸 的王，就是 以未 、 利金 、 蘇珥 、 戶珥 、 利巴 五個 米甸 的王，又用刀殺了 比珥 的兒子 巴蘭 。
NUM|31|9|以色列 人擄了 米甸 的婦女和孩童，搶奪他們一切的牲畜、牛羊和所有的財物，
NUM|31|10|又用火焚燒了他們所住的一切城鎮和所有的營寨。
NUM|31|11|以色列 人把一切擄物和掠物，連人和牲畜都帶走，
NUM|31|12|將俘虜、掠物、擄物帶到 摩押 平原，在 約旦河 邊與 耶利哥 相對的營地，交給 摩西 和 以利亞撒 祭司，以及 以色列 的會眾。
NUM|31|13|摩西 和 以利亞撒 祭司，以及會眾中所有的領袖，都出營迎接他們。
NUM|31|14|摩西 向打仗回來的軍官，就是千夫長和百夫長發怒。
NUM|31|15|摩西 對他們說：「你們要讓這所有的婦女活著嗎？
NUM|31|16|看哪，正是這些婦女，因 巴蘭 的話，在 毗珥 的事上導致 以色列 人背叛耶和華，以致耶和華的會眾遭遇瘟疫。
NUM|31|17|現在，你們要殺所有的男孩，也要把所有曾與男人同房共寢的女子都殺了。
NUM|31|18|但那些未曾與男人同房共寢的女孩，你們可以讓她們存活。
NUM|31|19|你們和你們所擄來的人，要住在營外七天；凡殺了人的，和一切摸了屍體的，要在第三日和第七日潔淨自己。
NUM|31|20|你們也要潔淨一切的衣服，以及用皮革、山羊毛和木頭做的任何東西。」
NUM|31|21|以利亞撒 祭司對打仗回來的士兵說：「耶和華所吩咐 摩西 律法中的條例是這樣：
NUM|31|22|金、銀、銅、鐵、錫、鉛，
NUM|31|23|凡能耐火的，你們要使它經過火，它就潔淨，然而還要用除污穢的水來潔淨它；凡不能耐火的，你們要使它經過水。
NUM|31|24|第七日，你們要洗衣服，才為潔淨，然後可以進營。」
NUM|31|25|耶和華對 摩西 說：
NUM|31|26|「你和 以利亞撒 祭司，以及會眾的各父系家長，要計算所擄掠的人和牲畜的總數。
NUM|31|27|要把所擄掠的分成兩半：一半給那出去打仗的精兵，一半給全會眾。
NUM|31|28|再從那出去打仗的戰士所得的人、牛、驢、羊中，每五百取一，獻給耶和華為貢物。
NUM|31|29|要從他們那一半中取出這些，交給 以利亞撒 祭司，作為耶和華的舉祭。
NUM|31|30|又要從 以色列 人的那一半中，就是從人、牛、驢、羊，各樣牲畜中，每五十取一，交給照管耶和華帳幕的 利未 人。」
NUM|31|31|於是 摩西 和 以利亞撒 祭司遵照耶和華所吩咐 摩西 的做了。
NUM|31|32|除了士兵所奪的財物以外，所擄來的有羊六十七萬五千隻，
NUM|31|33|牛七萬二千頭，
NUM|31|34|驢六萬一千匹；
NUM|31|35|至於人，就是未曾與男人同房共寢的女子，總共三萬二千名。
NUM|31|36|出去打仗之人的那分，就是他們所得的一半，共計羊三十三萬七千五百隻，
NUM|31|37|其中歸耶和華為貢物的羊，六百七十五隻；
NUM|31|38|牛三萬六千頭，其中歸耶和華為貢物的七十二頭；
NUM|31|39|驢三萬零五百匹，其中歸耶和華為貢物的六十一匹；
NUM|31|40|人一萬六千名，其中歸耶和華的三十二名。
NUM|31|41|摩西 把貢物，就是歸給耶和華的舉祭，交給 以利亞撒 祭司，是照耶和華所吩咐 摩西 的。
NUM|31|42|以色列 人所得的另一半，是 摩西 從打仗的人取來分給他們的。
NUM|31|43|會眾的這一半有羊三十三萬七千五百隻，
NUM|31|44|牛三萬六千頭，
NUM|31|45|驢三萬零五百匹，
NUM|31|46|人一萬六千名。
NUM|31|47|無論是人或牲畜， 摩西 都每五十取一，交給照管耶和華帳幕的 利未 人，是照耶和華所吩咐 摩西 的。
NUM|31|48|帶領眾軍隊的軍官，就是千夫長、百夫長，進到 摩西 那裏，
NUM|31|49|對他說：「你的僕人已經計算屬下戰士的總數，一個也沒有少。
NUM|31|50|如今我們把各人所得的金器，就是腳鏈子、手鐲、打印的戒指、耳環、項鏈，都送給耶和華為供物，好在耶和華面前為我們贖罪。」
NUM|31|51|摩西 和 以利亞撒 祭司就收了他們的金子，就是各樣的首飾。
NUM|31|52|千夫長、百夫長所獻給耶和華為舉祭的金子共有一萬六千七百五十舍客勒。
NUM|31|53|打仗的人都把自己所掠奪的各自留下。
NUM|31|54|摩西 和 以利亞撒 祭司收了千夫長、百夫長的金子，就帶進會幕，好使 以色列 人在耶和華面前蒙記念。
NUM|32|1|呂便 子孫和 迦得 子孫的牲畜極其眾多。他們看到 雅謝 地和 基列 地；看哪，這是可牧放牲畜的地方。
NUM|32|2|呂便 子孫和 迦得 子孫就到 摩西 和 以利亞撒 祭司，以及會眾的領袖那裏，說：
NUM|32|3|「 亞他錄 、 底本 、 雅謝 、 寧拉 、 希實本 、 以利亞利 、 示班 、 尼波 、 比穩 ，
NUM|32|4|就是耶和華在 以色列 會眾面前所攻取之地，是可牧放牲畜之地，而你的僕人也有牲畜。」
NUM|32|5|又說：「我們若在你眼前蒙恩，求你把這地給我們為業；不要領我們過 約旦河 。」
NUM|32|6|摩西 對 迦得 子孫和 呂便 子孫說：「難道你們的弟兄去打仗，你們卻留在這裏嗎？
NUM|32|7|你們為甚麼使 以色列 人灰心，不渡過去，進入耶和華所賜給他們的那地呢？
NUM|32|8|我從 加低斯‧巴尼亞 派你們的父執之輩去窺探那地時，他們就曾這樣做過。
NUM|32|9|他們上到 以實各谷 ，窺探了那地之後，竟然使 以色列 人灰心，不願進入耶和華所賜給他們的地。
NUM|32|10|當日，耶和華的怒氣發作，起誓說：
NUM|32|11|『凡從 埃及 上來二十歲以上的人，斷不得看見我對 亞伯拉罕 、 以撒 、 雅各 起誓應許之地，因為他們沒有專心跟從我；
NUM|32|12|惟有 基尼洗 族 耶孚尼 的兒子 迦勒 ，還有 嫩 的兒子 約書亞 可以看見，因為他們專心跟從耶和華。』
NUM|32|13|耶和華的怒氣向 以色列 發作，使他們在曠野飄流四十年，直到在耶和華眼前作惡的那一代都消滅了。
NUM|32|14|看哪，你們這一夥罪人，竟然接續你們父執之輩，再增加耶和華對 以色列 所發的怒氣。
NUM|32|15|你們若轉離不跟從他，他要再把 以色列 人撇在曠野；這樣，你們就使這眾百姓滅亡了。」
NUM|32|16|他們挨近 摩西 ，說：「我們要在這裏為牲畜築圈，為孩童建城。
NUM|32|17|我們自己卻要帶兵器，急速行在 以色列 人的前面，領他們直到他們的地方。我們的孩童可以留在堅固的城內，躲避當地的居民。
NUM|32|18|我們必不回自己的家，直等到 以色列 人各自承受了自己的產業。
NUM|32|19|我們不和他們在 約旦河 那邊分產業，因為我們的產業是在 約旦河 的東邊。」
NUM|32|20|摩西 對他們說：「你們若要這麼做，若要在耶和華面前帶著兵器出去打仗，
NUM|32|21|你們中間所有帶兵器的人都要在耶和華面前過 約旦河 ，直到耶和華把仇敵從他面前趕出去。
NUM|32|22|那地在耶和華面前被征服以後，你們方可回來。這樣，你們向耶和華和 以色列 才算為無罪，這地也必在耶和華面前歸你們為業。
NUM|32|23|倘若你們不這樣做，看哪，你們就得罪了耶和華，當知道你們的罪必找上你們。
NUM|32|24|如今你們可以為孩童建城，為羊群築圈，但你們口所講出來的話，必須實踐。」
NUM|32|25|迦得 子孫和 呂便 子孫對 摩西 說：「你的僕人們必照我主所吩咐的去做。
NUM|32|26|我們的孩子、妻子、牛羊和所有的牲畜都要留在 基列 的各城。
NUM|32|27|但你的僕人，凡能帶兵器上戰場的，都要照我主所說的話，在耶和華面前渡過去打仗。」
NUM|32|28|於是， 摩西 為他們吩咐 以利亞撒 祭司和 嫩 的兒子 約書亞 ，以及 以色列 人各支派父系的領袖。
NUM|32|29|摩西 對他們說：「 迦得 子孫和 呂便 子孫，凡帶兵器在耶和華面前去打仗的，若與你們一同渡過 約旦河 ，那地被你們征服以後，你們就要把 基列 地給他們為業。
NUM|32|30|倘若他們不帶兵器與你們一同渡過去，他們就要在 迦南 地你們中間得產業。」
NUM|32|31|迦得 子孫和 呂便 子孫回答說：「耶和華怎樣吩咐僕人，我們就必照樣做。
NUM|32|32|我們自己必帶著兵器，在耶和華面前渡過去，進入 迦南 地，好使我們在 約旦河 這邊得到我們的產業。」
NUM|32|33|摩西 把 亞摩利 王 西宏 的國和 巴珊 王 噩 的國，就是他們的國土和周圍的城鎮，都給了 迦得 子孫和 呂便 子孫，以及 約瑟 的兒子 瑪拿西 半個支派。
NUM|32|34|迦得 子孫建造了 底本 、 亞他錄 、 亞羅珥 、
NUM|32|35|亞他錄‧朔反 、 雅謝 、 約比哈 、
NUM|32|36|伯‧寧拉 、 伯‧哈蘭 ，都是堅固城，並築有羊圈。
NUM|32|37|呂便 子孫建造了 希實本 、 以利亞利 、 基列亭 、
NUM|32|38|尼波 、 巴力‧免 （名字是改了的）、 西比瑪 ；他們給建造的城另起別名。
NUM|32|39|瑪拿西 的兒子 瑪吉 的子孫往 基列 去，佔了那地，趕出那裏的 亞摩利 人。
NUM|32|40|摩西 把 基列 賜給 瑪拿西 的兒子 瑪吉 ，他就住在那裏。
NUM|32|41|瑪拿西 的子孫 睚珥 佔了 基列 的城鎮，就稱這些城鎮為 哈倭特‧睚珥 。
NUM|32|42|挪巴 佔了 基納 和 基納 的鄉鎮，就照自己的名字稱 基納 為 挪巴 。
NUM|33|1|這是 以色列 人按著隊伍，在 摩西 、 亞倫 的手下，出 埃及 地的行程。
NUM|33|2|摩西 遵照耶和華的指示記錄他們每段行程的起點，這些行程的起點如下：
NUM|33|3|第一個月，就是正月十五日，逾越的第二天，他們從 蘭塞 起行，在所有 埃及 人的眼前抬起頭 來出去了。
NUM|33|4|那時， 埃及 人正埋葬他們的長子，就是耶和華在他們中間所擊殺的；耶和華也懲治了他們的眾神明。
NUM|33|5|以色列 人從 蘭塞 起行，安營在 疏割 。
NUM|33|6|從 疏割 起行，安營在曠野邊上的 以倘 。
NUM|33|7|從 以倘 起行，轉向 巴力‧洗分 對面的 比‧哈希錄 ，安營在 密奪 。
NUM|33|8|從 比‧哈希錄 起行，經過海，進入曠野，在 以倘 的曠野走了三天的路程，就安營在 瑪拉 。
NUM|33|9|從 瑪拉 起行，來到 以琳 ， 以琳 有十二股水泉，七十棵棕樹，就安營在那裏。
NUM|33|10|從 以琳 起行，安營在 紅海 邊。
NUM|33|11|從 紅海 邊起行，安營在 汛 的曠野。
NUM|33|12|從 汛 的曠野起行，安營在 脫加 。
NUM|33|13|從 脫加 起行，安營在 亞錄 。
NUM|33|14|從 亞錄 起行，安營在 利非訂 ；在那裏，百姓沒有水喝。
NUM|33|15|從 利非訂 起行，安營在 西奈 的曠野。
NUM|33|16|從 西奈 的曠野起行，安營在 基博羅‧哈他瓦 。
NUM|33|17|從 基博羅‧哈他瓦 起行，安營在 哈洗錄 。
NUM|33|18|從 哈洗錄 起行，安營在 利提瑪 。
NUM|33|19|從 利提瑪 起行，安營在 臨門‧帕烈 。
NUM|33|20|從 臨門‧帕烈 起行，安營在 立拿 。
NUM|33|21|從 立拿 起行，安營在 勒撒 。
NUM|33|22|從 勒撒 起行，安營在 基希拉他 。
NUM|33|23|從 基希拉他 起行，安營在 沙斐山 。
NUM|33|24|從 沙斐山 起行，安營在 哈拉大 。
NUM|33|25|從 哈拉大 起行，安營在 瑪吉希錄 。
NUM|33|26|從 瑪吉希錄 起行，安營在 他哈 。
NUM|33|27|從 他哈 起行，安營在 他拉 。
NUM|33|28|從 他拉 起行，安營在 密加 。
NUM|33|29|從 密加 起行，安營在 哈摩拿 。
NUM|33|30|從 哈摩拿 起行，安營在 摩西錄 。
NUM|33|31|從 摩西錄 起行，安營在 比尼‧亞干 。
NUM|33|32|從 比尼‧亞干 起行，安營在 曷‧哈及甲 。
NUM|33|33|從 曷‧哈及甲 起行，安營在 約巴他 。
NUM|33|34|從 約巴他 起行，安營在 阿博拿 。
NUM|33|35|從 阿博拿 起行，安營在 以旬‧迦別 。
NUM|33|36|從 以旬‧迦別 起行，安營在 尋 的曠野，就是 加低斯 。
NUM|33|37|從 加低斯 起行，安營在 以東 地邊界的 何珥山 。
NUM|33|38|以色列 人出 埃及 地後四十年，五月初一， 亞倫 祭司遵照耶和華的指示，上 何珥山 ，死在那裏。
NUM|33|39|亞倫 死在 何珥山 的時候一百二十三歲。
NUM|33|40|住在 迦南 地 尼革夫 的 迦南 人 亞拉得 王聽說 以色列 人來了。
NUM|33|41|以色列 人從 何珥山 起行，安營在 撒摩拿 。
NUM|33|42|從 撒摩拿 起行，安營在 普嫩 。
NUM|33|43|從 普嫩 起行，安營在 阿伯 。
NUM|33|44|從 阿伯 起行，安營在 摩押 境內的 以耶‧亞巴琳 。
NUM|33|45|從 以耶‧亞巴琳 起行，安營在 底本‧迦得 。
NUM|33|46|從 底本‧迦得 起行，安營在 亞門‧低比拉太音 。
NUM|33|47|從 亞門‧低比拉太音 起行，安營在 尼波 前面的 亞巴琳山脈 。
NUM|33|48|從 亞巴琳山脈 起行，安營在 約旦河 邊， 耶利哥 對面的 摩押 平原。
NUM|33|49|他們在 摩押 平原，沿著 約旦河 安營，從 伯‧耶施末 直到 亞伯‧什亭 。
NUM|33|50|耶和華在 約旦河 邊， 耶利哥 對面的 摩押 平原吩咐 摩西 說：
NUM|33|51|「你要吩咐 以色列 人說：你們過 約旦河 進 迦南 地的時候，
NUM|33|52|要從你們面前趕出那地所有的居民，摧毀他們一切的石像和鑄成的偶像，也要拆毀他們一切的丘壇。
NUM|33|53|你們要佔領那地，住在那裏，因我已把那地賜給你們為業。
NUM|33|54|你們要按照宗族抽籤，承受土地：人多的要多給他們產業；人少的要少給他們產業。抽到何地給何人，那地就屬於他。你們要按照父系的支派承受產業。
NUM|33|55|倘若你們不把那地的居民從你們面前趕出去，那留下的居民就必成為你們眼中的刺，肋下的荊棘，也必在你們所住的地上擾亂你們；
NUM|33|56|我想要怎樣待他們，也必照樣待你們。」
NUM|34|1|耶和華吩咐 摩西 說：
NUM|34|2|「你要吩咐 以色列 人，對他們說：你們到了 迦南 地，這就是歸你們為業的地， 迦南 地和它四周的邊界：
NUM|34|3|你們的南邊是從 尋 的曠野起，沿著 以東 的邊界；南邊的地界從 鹽海 東邊開始，
NUM|34|4|繞過 亞克拉濱 斜坡的南邊，經過 尋 ，直通到 加低斯‧巴尼亞 的南邊，又通到 哈薩‧亞達 ，經過 押們 ，
NUM|34|5|從 押們 轉向 埃及 溪谷，直通到海。
NUM|34|6|「你們西邊的地界要以 大海 為邊界；這就是你們西邊的地界。
NUM|34|7|「你們北邊的地界要從 大海 開始劃界，直到 何珥山 ，
NUM|34|8|從 何珥山 劃到 哈馬口 ，直通到 西達達 ，
NUM|34|9|又通到 西斐崙 ，直達 哈薩‧以難 。這就是你們北邊的地界。
NUM|34|10|「東邊的地界，你們要從 哈薩‧以難 開始劃界，直到 示番 ，
NUM|34|11|這地界要從 示番 下到 亞延 東邊的 利比拉 ，這地界要下延到 基尼烈海 的東邊，
NUM|34|12|這地界又下到 約旦河 ，直通到 鹽海 。這就是你們的地和它四圍的邊界。」
NUM|34|13|摩西 吩咐 以色列 人說：「這就是耶和華吩咐抽籤給九個半支派承受為業的地。
NUM|34|14|因為 呂便 子孫的支派按著父家、 迦得 子孫的支派按著父家，和 瑪拿西 半個支派已經得到了他們的產業：
NUM|34|15|這兩個半支派已經在 耶利哥 對面， 約旦河 東邊，向日出的方向承受了產業。」
NUM|34|16|耶和華吩咐 摩西 說：
NUM|34|17|「這是為你們分地為業的人的名字： 以利亞撒 祭司和 嫩 的兒子 約書亞 。
NUM|34|18|你要從每個支派中選一個領袖來分配產業。
NUM|34|19|這些人的名字如下： 猶大 支派， 耶孚尼 的兒子 迦勒 。
NUM|34|20|西緬 子孫的支派， 亞米忽 的兒子 示母利 。
NUM|34|21|便雅憫 支派， 基斯倫 的兒子 以利達 。
NUM|34|22|但 子孫支派的領袖， 約利 的兒子 布基 。
NUM|34|23|約瑟 的子孫， 瑪拿西 子孫支派的領袖： 以弗 的兒子 漢尼業 。
NUM|34|24|以法蓮 子孫支派的領袖： 拾弗但 的兒子 基摩利 。
NUM|34|25|西布倫 子孫支派的領袖： 帕納 的兒子 以利撒番 。
NUM|34|26|以薩迦 子孫支派的領袖： 阿散 的兒子 帕鐵 。
NUM|34|27|亞設 子孫支派的領袖： 示羅米 的兒子 亞希忽 。
NUM|34|28|拿弗他利 子孫支派的領袖： 亞米忽 的兒子 比大黑 。」
NUM|34|29|這些就是耶和華所吩咐，在 迦南 地為 以色列 人分產業的人。
NUM|35|1|耶和華在 約旦河 邊， 耶利哥 對面的 摩押 平原吩咐 摩西 說：
NUM|35|2|「你吩咐 以色列 人，要從所得為業的地中把一些城給 利未 人居住，也要把這些城四圍的郊野給 利未 人。
NUM|35|3|這些城鎮要歸他們居住，郊外可以給他們牧放牛羊、牲畜和所有的動物。
NUM|35|4|你們給 利未 人城的郊外，要從城牆量起，四圍往外量一千肘。
NUM|35|5|你們要往東量二千肘，往南量二千肘，往西量二千肘，往北量二千肘為邊界，以城為中心；這城鎮的郊外要歸給他們。」
NUM|35|6|「你們給 利未 人的城鎮中，要設立六座逃城，讓誤殺人的可以逃到那裏。此外還要給他們四十二座城。
NUM|35|7|所以，給 利未 人的城一共有四十八座，連同城的郊外都給他們。
NUM|35|8|從 以色列 人所得的產業中給 利未 人的這些城鎮，多的要多給，少的要少給；各支派要按照所承受為業之地的多少把城鎮給 利未 人。」
NUM|35|9|耶和華吩咐 摩西 說：
NUM|35|10|「你要吩咐 以色列 人，對他們說：你們過了 約旦河 ，進入 迦南 地，
NUM|35|11|要指定幾座城，作為你們的逃城，使誤殺人的可以逃到那裏。
NUM|35|12|這些城要作為逃避報仇者的城，使誤殺人的不至於死，等他站在會眾面前受審判。
NUM|35|13|「你們指定的城，是要作你們的六座逃城。
NUM|35|14|約旦河 東指定三座， 迦南 地也指定三座，作為逃城。
NUM|35|15|這六座城要給 以色列 人和他們中間的外人，以及寄居者，作為逃城，讓誤殺人的可以逃到那裏。
NUM|35|16|「倘若人用鐵器打死人，他是故意殺人的；故意殺人的必被處死。
NUM|35|17|若用手中可以致命的石頭打死人，他是故意殺人的；故意殺人的必被處死。
NUM|35|18|若用手中可以致命的木器打死人，他是故意殺人的；故意殺人的必被處死。
NUM|35|19|報血仇者可以親自殺死那故意殺人的；他一找到兇手，就可以殺死他。
NUM|35|20|人若因怨恨把人推倒，或埋伏等著丟東西砸人，以至於死，
NUM|35|21|或因仇恨用手打死人，打人的必被處死，他是故意殺人的；報血仇者一遇見兇手就可以殺死他。
NUM|35|22|「人若不是出於仇恨，把人推倒，或不是埋伏等著丟東西砸人，
NUM|35|23|或是在不注意的時候，用可以致命的石頭扔在人身上，以至於死，彼此沒有仇恨，也無意害對方，
NUM|35|24|會眾就要照著這些典章，在殺人者和報血仇者中間審判。
NUM|35|25|會眾要救這誤殺人的脫離報血仇者的手，送他回到他曾逃入的逃城那裏。他要住在城中，直到受聖膏的大祭司去世。
NUM|35|26|但誤殺人的，無論甚麼時候，若離開了他所逃入的逃城邊界，
NUM|35|27|報血仇者在逃城邊界外遇見他，把兇手殺了，報血仇者就沒有流人血之罪。
NUM|35|28|因為誤殺人的應該住在逃城裏，直到大祭司去世。大祭司去世以後，誤殺人的才可以回到他所得為業之地。
NUM|35|29|在你們一切的住處，這些都要作為你們世世代代的律例典章。
NUM|35|30|「無論誰殺了人，必須憑幾個證人的口，才可把那故意殺人的處死；只憑一個證人，不足以判人死。
NUM|35|31|那犯死罪的殺人犯，你們不可收贖價來代替他的命；他必須被處死。
NUM|35|32|那逃到逃城的人，你們不可向他收贖價，使他在大祭司未死以先回本地居住。
NUM|35|33|這樣，你們就不會污穢所住之地，因為血能使地污穢；若有血流在地上，除非流那殺人者的血，否則那地就不得潔淨。
NUM|35|34|你們不可玷污所住之地，就是我住在當中的地，因為我－耶和華住在 以色列 人中間。」
NUM|36|1|約瑟 子孫的宗族， 瑪拿西 的孫子， 瑪吉 的兒子 基列 ，他父系宗族的領袖來到 摩西 和作領袖的 以色列 眾父系家長面前，說：
NUM|36|2|「耶和華曾吩咐我主抽籤分地給 以色列 人為業，我主也遵照耶和華的吩咐，把我們兄弟 西羅非哈 的產業給他的女兒。
NUM|36|3|她們若嫁給 以色列 別個支派的人，必拿走我們祖宗所遺留的產業，加在她們丈夫支派的產業上。這樣，我們抽籤所得的產業就要減少了。
NUM|36|4|到了 以色列 人的禧年，她們的產業就必加在她們丈夫支派的產業上。這樣，我們祖宗支派的產業就要減少了。」
NUM|36|5|摩西 照耶和華的指示吩咐 以色列 人說：「 約瑟 子孫支派的人說得有理。
NUM|36|6|關於 西羅非哈 的女兒們，這是耶和華吩咐的話說：『她們可以隨意嫁人，只是必須嫁給同宗，她們父親支派的人。
NUM|36|7|這樣， 以色列 人的產業就不會從這支派轉到另一個支派，因為 以色列 人要各自守住祖宗支派的產業。
NUM|36|8|凡在 以色列 支派中得了產業的女兒，必須嫁給同宗，她們父親支派的人，好使 以色列 人各自承受他們祖宗的產業。
NUM|36|9|產業不可從一個支派轉到另一個支派，因為 以色列 支派的人要各自守住自己的產業。』」
NUM|36|10|耶和華怎樣吩咐 摩西 ， 西羅非哈 的女兒就照樣做。
NUM|36|11|西羅非哈 的女兒 瑪拉 、 得撒 、 曷拉 、 密迦 、 挪阿 都嫁給她們叔伯的兒子。
NUM|36|12|她們嫁給了 約瑟 兒子 瑪拿西 子孫宗族的人；她們的產業保留在同宗，她們父親的支派中。
NUM|36|13|這是耶和華在 約旦河 邊， 耶利哥 對面的 摩押 平原，藉著 摩西 吩咐 以色列 人的命令和典章。
