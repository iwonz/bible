MAL|1|1|onus verbi Domini ad Israhel in manu Malachi
MAL|1|2|dilexi vos dicit Dominus et dixistis in quo dilexisti nos nonne frater erat Esau Iacob dicit Dominus et dilexi Iacob
MAL|1|3|Esau autem odio habui et posui montes eius in solitudinem et hereditatem eius in dracones deserti
MAL|1|4|quod si dixerit Idumea destructi sumus sed revertentes aedificabimus quae deserta sunt haec dicit Dominus exercituum isti aedificabunt et ego destruam et vocabuntur Termini impietatis et Populus cui iratus est Dominus usque in aeternum
MAL|1|5|et oculi vestri videbunt et vos dicetis magnificetur Dominus super terminum Israhel
MAL|1|6|filius honorat patrem et servus dominum suum si ergo pater ego sum ubi est honor meus et si dominus ego sum ubi est timor meus dicit Dominus exercituum ad vos o sacerdotes qui despicitis nomen meum et dixistis in quo despeximus nomen tuum
MAL|1|7|offertis super altare meum panem pollutum et dicitis in quo polluimus te in eo quod dicitis mensa Domini despecta est
MAL|1|8|si offeratis caecum ad immolandum nonne malum est et si offeratis claudum et languidum nonne malum est offer illud duci tuo si placuerit ei aut si susceperit faciem tuam dicit Dominus exercituum
MAL|1|9|et nunc deprecamini vultum Dei ut misereatur vestri de manu enim vestra factum est hoc si quo modo suscipiat facies vestras dicit Dominus exercituum
MAL|1|10|quis est in vobis qui claudat ostia et incendat altare meum gratuito non est mihi voluntas in vobis dicit Dominus exercituum et munus non suscipiam de manu vestra
MAL|1|11|ab ortu enim solis usque ad occasum magnum est nomen meum in gentibus et in omni loco sacrificatur et offertur nomini meo oblatio munda quia magnum nomen meum in gentibus dicit Dominus exercituum
MAL|1|12|et vos polluistis illud in eo quod dicitis mensa Domini contaminata est et quod superponitur contemptibile est cum igni qui illud devorat
MAL|1|13|et dixistis ecce de labore et exsuflastis illud dicit Dominus exercituum et intulistis de rapinis claudum et languidum et intulistis munus numquid suscipiam illud de manu vestra dicit Dominus
MAL|1|14|maledictus dolosus qui habet in grege suo masculum et votum faciens immolat debile Domino quia rex magnus ego dicit Dominus exercituum et nomen meum horribile in gentibus
MAL|2|1|et nunc ad vos mandatum hoc o sacerdotes
MAL|2|2|si nolueritis audire et si nolueritis ponere super cor ut detis gloriam nomini meo ait Dominus exercituum mittam in vos egestatem et maledicam benedictionibus vestris et maledicam illis quoniam non posuistis super cor
MAL|2|3|ecce ego proiciam vobis brachium et dispergam super vultum vestrum stercus sollemnitatum vestrarum et adsumet vos secum
MAL|2|4|et scietis quia misi ad vos mandatum istud ut esset pactum meum cum Levi dicit Dominus exercituum
MAL|2|5|pactum meum fuit cum eo vitae et pacis et dedi ei timorem et timuit me et a facie nominis mei pavebat
MAL|2|6|lex veritatis fuit in ore eius et iniquitas non est inventa in labiis eius in pace et in aequitate ambulavit mecum et multos avertit ab iniquitate
MAL|2|7|labia enim sacerdotis custodient scientiam et legem requirent ex ore eius quia angelus Domini exercituum est
MAL|2|8|vos autem recessistis de via et scandalizastis plurimos in lege irritum fecistis pactum Levi dicit Dominus exercituum
MAL|2|9|propter quod et ego dedi vos contemptibiles et humiles omnibus populis sicut non servastis vias meas et accepistis faciem in lege
MAL|2|10|numquid non pater unus omnium nostrum numquid non Deus unus creavit nos quare ergo despicit unusquisque nostrum fratrem suum violans pactum patrum nostrorum
MAL|2|11|transgressus est Iuda et abominatio facta est in Israhel et in Hierusalem quia contaminavit Iudas sanctificationem Domini quam dilexit et habuit filiam dei alieni
MAL|2|12|disperdat Dominus virum qui fecerit hoc magistrum et discipulum de tabernaculis Iacob et offerentem munus Domino exercituum
MAL|2|13|et hoc rursum fecistis operiebatis lacrimis altare Domini fletu et mugitu ita ut ultra non respiciam ad sacrificium nec accipiam placabile quid de manu vestra
MAL|2|14|et dixistis quam ob causam quia Dominus testificatus est inter te et uxorem pubertatis tuae quam tu despexisti et haec particeps tua et uxor foederis tui
MAL|2|15|nonne unus fecit et residuum spiritus eius est et quid unus quaerit nisi semen Dei custodite ergo spiritum vestrum et uxorem adulescentiae tuae noli despicere
MAL|2|16|cum odio habueris dimitte dicit Dominus Deus Israhel operiet autem iniquitas vestimentum eius dicit Dominus exercituum custodite spiritum vestrum et nolite despicere
MAL|2|17|laborare fecistis Dominum in sermonibus vestris et dixistis in quo eum fecimus laborare in eo cum diceretis omnis qui facit malum bonus est in conspectu Domini et tales ei placent aut certe ubi est Deus iudicii
MAL|3|1|ecce ego mittam angelum meum et praeparabit viam ante faciem meam et statim veniet ad templum suum dominator quem vos quaeritis et angelus testamenti quem vos vultis ecce venit dicit Dominus exercituum
MAL|3|2|et quis poterit cogitare diem adventus eius et quis stabit ad videndum eum ipse enim quasi ignis conflans et quasi herba fullonum
MAL|3|3|et sedebit conflans et emundans argentum et purgabit filios Levi et colabit eos quasi aurum et quasi argentum et erunt Domino offerentes sacrificia in iustitia
MAL|3|4|et placebit Domino sacrificium Iuda et Hierusalem sicut dies saeculi et sicut anni antiqui
MAL|3|5|et accedam ad vos in iudicio et ero testis velox maleficis et adulteris et periuris et qui calumniantur mercedem mercennarii viduas et pupillos et opprimunt peregrinum nec timuerunt me dicit Dominus exercituum
MAL|3|6|ego enim Dominus et non mutor et vos filii Iacob non estis consumpti
MAL|3|7|a diebus enim patrum vestrorum recessistis a legitimis meis et non custodistis revertimini ad me et revertar ad vos dicit Dominus exercituum et dixistis in quo revertemur
MAL|3|8|si adfiget homo Deum quia vos configitis me et dixistis in quo confiximus te in decimis et in primitivis
MAL|3|9|et in penuria vos maledicti estis et me vos configitis gens tota
MAL|3|10|inferte omnem decimam in horreum et sit cibus in domo mea et probate me super hoc dicit Dominus si non aperuero vobis cataractas caeli et effudero vobis benedictionem usque ad abundantiam
MAL|3|11|et increpabo pro vobis devorantem et non corrumpet fructum terrae vestrae nec erit sterilis vinea in agro dicit Dominus exercituum
MAL|3|12|et beatos vos dicent omnes gentes eritis enim vos terra desiderabilis dicit Dominus exercituum
MAL|3|13|invaluerunt super me verba vestra dicit Dominus
MAL|3|14|et dixistis quid locuti sumus contra te dixistis vanus est qui servit Deo et quod emolumentum quia custodivimus praecepta eius et quia ambulavimus tristes coram Domino exercituum
MAL|3|15|ergo nunc beatos dicimus arrogantes siquidem aedificati sunt facientes impietatem et temptaverunt Deum et salvi facti sunt
MAL|3|16|tunc locuti sunt timentes Deum unusquisque cum proximo suo et adtendit Dominus et audivit et scriptus est liber monumenti coram eo timentibus Dominum et cogitantibus nomen eius
MAL|3|17|et erunt mihi ait Dominus exercituum in die qua ego facio in peculium et parcam eis sicut parcit vir filio suo servienti sibi
MAL|3|18|et convertemini et videbitis quid sit inter iustum et impium et inter servientem Deo et non servientem ei
MAL|4|1|ecce enim dies veniet succensa quasi caminus et erunt omnes superbi et omnes facientes impietatem stipula et inflammabit eos dies veniens dicit Dominus exercituum quae non relinquet eis radicem et germen
MAL|4|2|et orietur vobis timentibus nomen meum sol iustitiae et sanitas in pinnis eius et egrediemini et salietis sicut vituli de armento
MAL|4|3|et calcabitis impios cum fuerint cinis sub planta pedum vestrorum in die qua ego facio dicit Dominus exercituum
MAL|4|4|mementote legis Mosi servi mei quam mandavi ei in Choreb ad omnem Israhel praecepta et iudicia
MAL|4|5|ecce ego mittam vobis Heliam prophetam antequam veniat dies Domini magnus et horribilis
MAL|4|6|et convertet cor patrum ad filios et cor filiorum ad patres eorum ne forte veniam et percutiam terram anathemate
