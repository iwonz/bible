HEB|1|1|Бог, многократно и многообразно говоривший издревле отцам в пророках,
HEB|1|2|в последние дни сии говорил нам в Сыне, Которого поставил наследником всего, чрез Которого и веки сотворил.
HEB|1|3|Сей, будучи сияние славы и образ ипостаси Его и держа все словом силы Своей, совершив Собою очищение грехов наших, воссел одесную престола величия на высоте,
HEB|1|4|будучи столько превосходнее Ангелов, сколько славнейшее пред ними наследовал имя.
HEB|1|5|Ибо кому когда из Ангелов сказал [Бог]: Ты Сын Мой, Я ныне родил Тебя? И еще: Я буду Ему Отцем, и Он будет Мне Сыном?
HEB|1|6|Также, когда вводит Первородного во вселенную, говорит: и да поклонятся Ему все Ангелы Божии.
HEB|1|7|Об Ангелах сказано: Ты творишь Ангелами Своими духов и служителями Своими пламенеющий огонь.
HEB|1|8|А о Сыне: престол Твой, Боже, в век века; жезл царствия Твоего – жезл правоты.
HEB|1|9|Ты возлюбил правду и возненавидел беззаконие, посему помазал Тебя, Боже, Бог Твой елеем радости более соучастников Твоих.
HEB|1|10|И: в начале Ты, Господи, основал землю, и небеса – дело рук Твоих;
HEB|1|11|они погибнут, а Ты пребываешь; и все обветшают, как риза,
HEB|1|12|и как одежду свернешь их, и изменятся; но Ты тот же, и лета Твои не кончатся.
HEB|1|13|Кому когда из Ангелов сказал [Бог]: седи одесную Меня, доколе положу врагов Твоих в подножие ног Твоих?
HEB|1|14|Не все ли они суть служебные духи, посылаемые на служение для тех, которые имеют наследовать спасение?
HEB|2|1|Посему мы должны быть особенно внимательны к слышанному, чтобы не отпасть.
HEB|2|2|Ибо, если через Ангелов возвещенное слово было твердо, и всякое преступление и непослушание получало праведное воздаяние,
HEB|2|3|то как мы избежим, вознерадев о толиком спасении, которое, быв сначала проповедано Господом, в нас утвердилось слышавшими [от Него],
HEB|2|4|при засвидетельствовании от Бога знамениями и чудесами, и различными силами, и раздаянием Духа Святаго по Его воле?
HEB|2|5|Ибо не Ангелам Бог покорил будущую вселенную, о которой говорим;
HEB|2|6|напротив некто негде засвидетельствовал, говоря: что значит человек, что Ты помнишь его? или сын человеческий, что Ты посещаешь его?
HEB|2|7|Не много Ты унизил его пред Ангелами; славою и честью увенчал его, и поставил его над делами рук Твоих,
HEB|2|8|все покорил под ноги его. Когда же покорил ему все, то не оставил ничего непокоренным ему. Ныне же еще не видим, чтобы все было ему покорено;
HEB|2|9|но видим, что за претерпение смерти увенчан славою и честью Иисус, Который не много был унижен пред Ангелами, дабы Ему, по благодати Божией, вкусить смерть за всех.
HEB|2|10|Ибо надлежало, чтобы Тот, для Которого все и от Которого все, приводящего многих сынов в славу, вождя спасения их совершил через страдания.
HEB|2|11|Ибо и освящающий и освящаемые, все – от Единого; поэтому Он не стыдится называть их братиями, говоря:
HEB|2|12|возвещу имя Твое братиям Моим, посреди церкви воспою Тебя.
HEB|2|13|И еще: Я буду уповать на Него. И еще: вот Я и дети, которых дал Мне Бог.
HEB|2|14|А как дети причастны плоти и крови, то и Он также воспринял оные, дабы смертью лишить силы имеющего державу смерти, то есть диавола,
HEB|2|15|и избавить тех, которые от страха смерти через всю жизнь были подвержены рабству.
HEB|2|16|Ибо не Ангелов восприемлет Он, но восприемлет семя Авраамово.
HEB|2|17|Посему Он должен был во всем уподобиться братиям, чтобы быть милостивым и верным первосвященником пред Богом, для умилостивления за грехи народа.
HEB|2|18|Ибо, как Сам Он претерпел, быв искушен, то может и искушаемым помочь.
HEB|3|1|Итак, братия святые, участники в небесном звании, уразумейте Посланника и Первосвященника исповедания нашего, Иисуса Христа,
HEB|3|2|Который верен Поставившему Его, как и Моисей во всем доме Его.
HEB|3|3|Ибо Он достоин тем большей славы пред Моисеем, чем большую честь имеет в сравнении с домом тот, кто устроил его,
HEB|3|4|ибо всякий дом устрояется кем–либо; а устроивший все [есть] Бог.
HEB|3|5|И Моисей верен во всем доме Его, как служитель, для засвидетельствования того, что надлежало возвестить;
HEB|3|6|а Христос – как Сын в доме Его; дом же Его – мы, если только дерзновение и упование, которым хвалимся, твердо сохраним до конца.
HEB|3|7|Почему, как говорит Дух Святый, ныне, когда услышите глас Его,
HEB|3|8|не ожесточите сердец ваших, как во время ропота, в день искушения в пустыне,
HEB|3|9|где искушали Меня отцы ваши, испытывали Меня, и видели дела Мои сорок лет.
HEB|3|10|Посему Я вознегодовал на оный род и сказал: непрестанно заблуждаются сердцем, не познали они путей Моих;
HEB|3|11|посему Я поклялся во гневе Моем, что они не войдут в покой Мой.
HEB|3|12|Смотрите, братия, чтобы не было в ком из вас сердца лукавого и неверного, дабы вам не отступить от Бога живаго.
HEB|3|13|Но наставляйте друг друга каждый день, доколе можно говорить: "ныне", чтобы кто из вас не ожесточился, обольстившись грехом.
HEB|3|14|Ибо мы сделались причастниками Христу, если только начатую жизнь твердо сохраним до конца,
HEB|3|15|доколе говорится: "ныне, когда услышите глас Его, не ожесточите сердец ваших, как во время ропота".
HEB|3|16|Ибо некоторые из слышавших возроптали; но не все вышедшие из Египта с Моисеем.
HEB|3|17|На кого же негодовал Он сорок лет? Не на согрешивших ли, которых кости пали в пустыне?
HEB|3|18|Против кого же клялся, что не войдут в покой Его, как не против непокорных?
HEB|3|19|Итак видим, что они не могли войти за неверие.
HEB|4|1|Посему будем опасаться, чтобы, когда еще остается обетование войти в покой Его, не оказался кто из вас опоздавшим.
HEB|4|2|Ибо и нам оно возвещено, как и тем; но не принесло им пользы слово слышанное, не растворенное верою слышавших.
HEB|4|3|А входим в покой мы уверовавшие, так как Он сказал: "Я поклялся в гневе Моем, что они не войдут в покой Мой", хотя дела [Его] были совершены еще в начале мира.
HEB|4|4|Ибо негде сказано о седьмом [дне] так: и почил Бог в день седьмый от всех дел Своих.
HEB|4|5|И еще здесь: "не войдут в покой Мой".
HEB|4|6|Итак, как некоторым остается войти в него, а те, которым прежде возвещено, не вошли в него за непокорность,
HEB|4|7|[то] еще определяет некоторый день, "ныне", говоря через Давида, после столь долгого времени, как выше сказано: "ныне, когда услышите глас Его, не ожесточите сердец ваших".
HEB|4|8|Ибо если бы Иисус [Навин] доставил им покой, то не было бы сказано после того о другом дне.
HEB|4|9|Посему для народа Божия еще остается субботство.
HEB|4|10|Ибо, кто вошел в покой Его, тот и сам успокоился от дел своих, как и Бог от Своих.
HEB|4|11|Итак постараемся войти в покой оный, чтобы кто по тому же примеру не впал в непокорность.
HEB|4|12|Ибо слово Божие живо и действенно и острее всякого меча обоюдоострого: оно проникает до разделения души и духа, составов и мозгов, и судит помышления и намерения сердечные.
HEB|4|13|И нет твари, сокровенной от Него, но все обнажено и открыто перед очами Его: Ему дадим отчет.
HEB|4|14|Итак, имея Первосвященника великого, прошедшего небеса, Иисуса Сына Божия, будем твердо держаться исповедания [нашего].
HEB|4|15|Ибо мы имеем не такого первосвященника, который не может сострадать нам в немощах наших, но Который, подобно [нам], искушен во всем, кроме греха.
HEB|4|16|Посему да приступаем с дерзновением к престолу благодати, чтобы получить милость и обрести благодать для благовременной помощи.
HEB|5|1|Ибо всякий первосвященник, из человеков избираемый, для человеков поставляется на служение Богу, чтобы приносить дары и жертвы за грехи,
HEB|5|2|могущий снисходить невежествующим и заблуждающим, потому что и сам обложен немощью,
HEB|5|3|и посему он должен как за народ, так и за себя приносить [жертвы] о грехах.
HEB|5|4|И никто сам собою не приемлет этой чести, но призываемый Богом, как и Аарон.
HEB|5|5|Так и Христос не Сам Себе присвоил славу быть первосвященником, но Тот, Кто сказал Ему: Ты Сын Мой, Я ныне родил Тебя;
HEB|5|6|как и в другом [месте] говорит: Ты священник вовек по чину Мелхиседека.
HEB|5|7|Он, во дни плоти Своей, с сильным воплем и со слезами принес молитвы и моления Могущему спасти Его от смерти; и услышан был за [Свое] благоговение;
HEB|5|8|хотя Он и Сын, однако страданиями навык послушанию,
HEB|5|9|и, совершившись, сделался для всех послушных Ему виновником спасения вечного,
HEB|5|10|быв наречен от Бога Первосвященником по чину Мелхиседека.
HEB|5|11|О сем надлежало бы нам говорить много; но трудно истолковать, потому что вы сделались неспособны слушать.
HEB|5|12|Ибо, [судя] по времени, вам надлежало быть учителями; но вас снова нужно учить первым началам слова Божия, и для вас нужно молоко, а не твердая пища.
HEB|5|13|Всякий, питаемый молоком, несведущ в слове правды, потому что он младенец;
HEB|5|14|твердая же пища свойственна совершенным, у которых чувства навыком приучены к различению добра и зла.
HEB|6|1|Посему, оставив начатки учения Христова, поспешим к совершенству; и не станем снова полагать основание обращению от мертвых дел и вере в Бога,
HEB|6|2|учению о крещениях, о возложении рук, о воскресении мертвых и о суде вечном.
HEB|6|3|И это сделаем, если Бог позволит.
HEB|6|4|Ибо невозможно – однажды просвещенных, и вкусивших дара небесного, и соделавшихся причастниками Духа Святаго,
HEB|6|5|и вкусивших благого глагола Божия и сил будущего века,
HEB|6|6|и отпадших, опять обновлять покаянием, когда они снова распинают в себе Сына Божия и ругаются [Ему].
HEB|6|7|Земля, пившая многократно сходящий на нее дождь и произращающая злак, полезный тем, для которых и возделывается, получает благословение от Бога;
HEB|6|8|а производящая терния и волчцы негодна и близка к проклятию, которого конец – сожжение.
HEB|6|9|Впрочем о вас, возлюбленные, мы надеемся, что вы в лучшем [состоянии] и держитесь спасения, хотя и говорим так.
HEB|6|10|Ибо не неправеден Бог, чтобы забыл дело ваше и труд любви, которую вы оказали во имя Его, послужив и служа святым.
HEB|6|11|Желаем же, чтобы каждый из вас, для совершенной уверенности в надежде, оказывал такую же ревность до конца,
HEB|6|12|дабы вы не обленились, но подражали тем, которые верою и долготерпением наследуют обетования.
HEB|6|13|Бог, давая обетование Аврааму, как не мог никем высшим клясться, клялся Самим Собою,
HEB|6|14|говоря: истинно благословляя благословлю тебя и размножая размножу тебя.
HEB|6|15|И так Авраам, долготерпев, получил обещанное.
HEB|6|16|Люди клянутся высшим, и клятва во удостоверение оканчивает всякий спор их.
HEB|6|17|Посему и Бог, желая преимущественнее показать наследникам обетования непреложность Своей воли, употребил в посредство клятву,
HEB|6|18|дабы в двух непреложных вещах, в которых невозможно Богу солгать, твердое утешение имели мы, прибегшие взяться за предлежащую надежду,
HEB|6|19|которая для души есть как бы якорь безопасный и крепкий, и входит во внутреннейшее за завесу,
HEB|6|20|куда предтечею за нас вошел Иисус, сделавшись Первосвященником навек по чину Мелхиседека.
HEB|7|1|Ибо Мелхиседек, царь Салима, священник Бога Всевышнего, тот, который встретил Авраама и благословил его, возвращающегося после поражения царей,
HEB|7|2|которому и десятину отделил Авраам от всего, – во–первых, по знаменованию [имени] царь правды, а потом и царь Салима, то есть царь мира,
HEB|7|3|без отца, без матери, без родословия, не имеющий ни начала дней, ни конца жизни, уподобляясь Сыну Божию, пребывает священником навсегда.
HEB|7|4|Видите, как велик тот, которому и Авраам патриарх дал десятину из лучших добыч своих.
HEB|7|5|Получающие священство из сынов Левииных имеют заповедь – брать по закону десятину с народа, то есть со своих братьев, хотя и сии произошли от чресл Авраамовых.
HEB|7|6|Но сей, не происходящий от рода их, получил десятину от Авраама и благословил имевшего обетования.
HEB|7|7|Без всякого же прекословия меньший благословляется большим.
HEB|7|8|И здесь десятины берут человеки смертные, а там – имеющий о себе свидетельство, что он живет.
HEB|7|9|И, так сказать, сам Левий, принимающий десятины, в [лице] Авраама дал десятину:
HEB|7|10|ибо он был еще в чреслах отца, когда Мелхиседек встретил его.
HEB|7|11|Итак, если бы совершенство достигалось посредством левитского священства, – ибо с ним сопряжен закон народа, – то какая бы еще нужда была восставать иному священнику по чину Мелхиседека, а не по чину Аарона именоваться?
HEB|7|12|Потому что с переменою священства необходимо быть перемене и закона.
HEB|7|13|Ибо Тот, о Котором говорится сие, принадлежал к иному колену, из которого никто не приступал к жертвеннику.
HEB|7|14|Ибо известно, что Господь наш воссиял из колена Иудина, о котором Моисей ничего не сказал относительно священства.
HEB|7|15|И это еще яснее видно [из того], что по подобию Мелхиседека восстает Священник иной,
HEB|7|16|Который таков не по закону заповеди плотской, но по силе жизни непрестающей.
HEB|7|17|Ибо засвидетельствовано: Ты священник вовек по чину Мелхиседека.
HEB|7|18|Отменение же прежде бывшей заповеди бывает по причине ее немощи и бесполезности,
HEB|7|19|ибо закон ничего не довел до совершенства; но вводится лучшая надежда, посредством которой мы приближаемся к Богу.
HEB|7|20|И как [сие было] не без клятвы, –
HEB|7|21|ибо те были священниками без клятвы, а Сей с клятвою, потому что о Нем сказано: клялся Господь, и не раскается: Ты священник вовек по чину Мелхиседека, –
HEB|7|22|то лучшего завета поручителем соделался Иисус.
HEB|7|23|Притом тех священников было много, потому что смерть не допускала пребывать одному;
HEB|7|24|а Сей, как пребывающий вечно, имеет и священство непреходящее,
HEB|7|25|посему и может всегда спасать приходящих чрез Него к Богу, будучи всегда жив, чтобы ходатайствовать за них.
HEB|7|26|Таков и должен быть у нас Первосвященник: святой, непричастный злу, непорочный, отделенный от грешников и превознесенный выше небес,
HEB|7|27|Который не имеет нужды ежедневно, как те первосвященники, приносить жертвы сперва за свои грехи, потом за грехи народа, ибо Он совершил это однажды, принеся [в жертву] Себя Самого.
HEB|7|28|Ибо закон поставляет первосвященниками человеков, имеющих немощи; а слово клятвенное, после закона, [поставило] Сына, на веки совершенного.
HEB|8|1|Главное же в том, о чем говорим, есть то: мы имеем такого Первосвященника, Который воссел одесную престола величия на небесах
HEB|8|2|и [есть] священнодействователь святилища и скинии истинной, которую воздвиг Господь, а не человек.
HEB|8|3|Всякий первосвященник поставляется для приношения даров и жертв; а потому нужно было, чтобы и Сей также имел, что принести.
HEB|8|4|Если бы Он оставался на земле, то не был бы и священником, потому что [здесь] такие священники, которые по закону приносят дары,
HEB|8|5|которые служат образу и тени небесного, как сказано было Моисею, когда он приступал к совершению скинии: смотри, сказано, сделай все по образу, показанному тебе на горе.
HEB|8|6|Но Сей [Первосвященник] получил служение тем превосходнейшее, чем лучшего Он ходатай завета, который утвержден на лучших обетованиях.
HEB|8|7|Ибо, если бы первый [завет] был без недостатка, то не было бы нужды искать места другому.
HEB|8|8|Но [пророк], укоряя их, говорит: вот, наступают дни, говорит Господь, когда Я заключу с домом Израиля и с домом Иуды новый завет,
HEB|8|9|не такой завет, какой Я заключил с отцами их в то время, когда взял их за руку, чтобы вывести их из земли Египетской, потому что они не пребыли в том завете Моем, и Я пренебрег их, говорит Господь.
HEB|8|10|Вот завет, который завещаю дому Израилеву после тех дней, говорит Господь: вложу законы Мои в мысли их, и напишу их на сердцах их; и буду их Богом, а они будут Моим народом.
HEB|8|11|И не будет учить каждый ближнего своего и каждый брата своего, говоря: познай Господа; потому что все, от малого до большого, будут знать Меня,
HEB|8|12|потому что Я буду милостив к неправдам их, и грехов их и беззаконий их не воспомяну более.
HEB|8|13|Говоря "новый", показал ветхость первого; а ветшающее и стареющее близко к уничтожению.
HEB|9|1|И первый завет имел постановление о Богослужении и святилище земное:
HEB|9|2|ибо устроена была скиния первая, в которой был светильник, и трапеза, и предложение хлебов, и которая называется "святое".
HEB|9|3|За второю же завесою была скиния, называемая "Святое–святых",
HEB|9|4|имевшая золотую кадильницу и обложенный со всех сторон золотом ковчег завета, где были золотой сосуд с манною, жезл Ааронов расцветший и скрижали завета,
HEB|9|5|а над ним херувимы славы, осеняющие очистилище; о чем не нужно теперь говорить подробно.
HEB|9|6|При таком устройстве, в первую скинию всегда входят священники совершать Богослужение;
HEB|9|7|а во вторую – однажды в год один только первосвященник, не без крови, которую приносит за себя и за грехи неведения народа.
HEB|9|8|[Сим] Дух Святый показывает, что еще не открыт путь во святилище, доколе стоит прежняя скиния.
HEB|9|9|Она есть образ настоящего времени, в которое приносятся дары и жертвы, не могущие сделать в совести совершенным приносящего,
HEB|9|10|и которые с яствами и питиями, и различными омовениями и обрядами, [относящимися] до плоти, установлены были только до времени исправления.
HEB|9|11|Но Христос, Первосвященник будущих благ, придя с большею и совершеннейшею скиниею, нерукотворенною, то есть не такового устроения,
HEB|9|12|и не с кровью козлов и тельцов, но со Своею Кровию, однажды вошел во святилище и приобрел вечное искупление.
HEB|9|13|Ибо если кровь тельцов и козлов и пепел телицы, через окропление, освящает оскверненных, дабы чисто было тело,
HEB|9|14|то кольми паче Кровь Христа, Который Духом Святым принес Себя непорочного Богу, очистит совесть нашу от мертвых дел, для служения Богу живому и истинному!
HEB|9|15|И потому Он есть ходатай нового завета, дабы вследствие смерти [Его], бывшей для искупления от преступлений, сделанных в первом завете, призванные к вечному наследию получили обетованное.
HEB|9|16|Ибо, где завещание, там необходимо, чтобы последовала смерть завещателя,
HEB|9|17|потому что завещание действительно после умерших: оно не имеет силы, когда завещатель жив.
HEB|9|18|Почему и первый [завет] был утвержден не без крови.
HEB|9|19|Ибо Моисей, произнеся все заповеди по закону перед всем народом, взял кровь тельцов и козлов с водою и шерстью червленою и иссопом, и окропил как самую книгу, так и весь народ,
HEB|9|20|говоря: это кровь завета, который заповедал вам Бог.
HEB|9|21|Также окропил кровью и скинию и все сосуды Богослужебные.
HEB|9|22|Да и все почти по закону очищается кровью, и без пролития крови не бывает прощения.
HEB|9|23|Итак образы небесного должны были очищаться сими, самое же небесное лучшими сих жертвами.
HEB|9|24|Ибо Христос вошел не в рукотворенное святилище, по образу истинного [устроенное], но в самое небо, чтобы предстать ныне за нас пред лице Божие,
HEB|9|25|и не для того, чтобы многократно приносить Себя, как первосвященник входит во святилище каждогодно с чужою кровью;
HEB|9|26|иначе надлежало бы Ему многократно страдать от начала мира; Он же однажды, к концу веков, явился для уничтожения греха жертвою Своею.
HEB|9|27|И как человекам положено однажды умереть, а потом суд,
HEB|9|28|так и Христос, однажды принеся Себя в жертву, чтобы подъять грехи многих, во второй раз явится не [для очищения] греха, а для ожидающих Его во спасение.
HEB|10|1|Закон, имея тень будущих благ, а не самый образ вещей, одними и теми же жертвами, каждый год постоянно приносимыми, никогда не может сделать совершенными приходящих [с ними].
HEB|10|2|Иначе перестали бы приносить [их], потому что приносящие жертву, быв очищены однажды, не имели бы уже никакого сознания грехов.
HEB|10|3|Но жертвами каждогодно напоминается о грехах,
HEB|10|4|ибо невозможно, чтобы кровь тельцов и козлов уничтожала грехи.
HEB|10|5|Посему [Христос], входя в мир, говорит: жертвы и приношения Ты не восхотел, но тело уготовал Мне.
HEB|10|6|Всесожжения и [жертвы] за грех неугодны Тебе.
HEB|10|7|Тогда Я сказал: вот, иду, [как] в начале книги написано о Мне, исполнить волю Твою, Боже.
HEB|10|8|Сказав прежде, что "ни жертвы, ни приношения, ни всесожжений, ни [жертвы] за грех, – которые приносятся по закону, – Ты не восхотел и не благоизволил",
HEB|10|9|потом прибавил: "вот, иду исполнить волю Твою, Боже". Отменяет первое, чтобы постановить второе.
HEB|10|10|По сей–то воле освящены мы единократным принесением тела Иисуса Христа.
HEB|10|11|И всякий священник ежедневно стоит в служении, и многократно приносит одни и те же жертвы, которые никогда не могут истребить грехов.
HEB|10|12|Он же, принеся одну жертву за грехи, навсегда воссел одесную Бога,
HEB|10|13|ожидая затем, доколе враги Его будут положены в подножие ног Его.
HEB|10|14|Ибо Он одним приношением навсегда сделал совершенными освящаемых.
HEB|10|15|[О сем] свидетельствует нам и Дух Святый; ибо сказано:
HEB|10|16|Вот завет, который завещаю им после тех дней, говорит Господь: вложу законы Мои в сердца их, и в мыслях их напишу их,
HEB|10|17|и грехов их и беззаконий их не воспомяну более.
HEB|10|18|А где прощение грехов, там не нужно приношение за них.
HEB|10|19|Итак, братия, имея дерзновение входить во святилище посредством Крови Иисуса Христа, путем новым и живым,
HEB|10|20|который Он вновь открыл нам через завесу, то есть плоть Свою,
HEB|10|21|и [имея] великого Священника над домом Божиим,
HEB|10|22|да приступаем с искренним сердцем, с полною верою, кроплением очистив сердца от порочной совести, и омыв тело водою чистою,
HEB|10|23|будем держаться исповедания упования неуклонно, ибо верен Обещавший.
HEB|10|24|Будем внимательны друг ко другу, поощряя к любви и добрым делам.
HEB|10|25|Не будем оставлять собрания своего, как есть у некоторых обычай; но будем увещевать [друг друга], и тем более, чем более усматриваете приближение дня оного.
HEB|10|26|Ибо если мы, получив познание истины, произвольно грешим, то не остается более жертвы за грехи,
HEB|10|27|но некое страшное ожидание суда и ярость огня, готового пожрать противников.
HEB|10|28|[Если] отвергшийся закона Моисеева, при двух или трех свидетелях, без милосердия [наказывается] смертью,
HEB|10|29|то сколь тягчайшему, думаете, наказанию повинен будет тот, кто попирает Сына Божия и не почитает за святыню Кровь завета, которою освящен, и Духа благодати оскорбляет?
HEB|10|30|Мы знаем Того, Кто сказал: у Меня отмщение, Я воздам, говорит Господь. И еще: Господь будет судить народ Свой.
HEB|10|31|Страшно впасть в руки Бога живаго!
HEB|10|32|Вспомните прежние дни ваши, когда вы, быв просвещены, выдержали великий подвиг страданий,
HEB|10|33|то сами среди поношений и скорбей служа зрелищем [для других], то принимая участие в других, находившихся в таком же [состоянии];
HEB|10|34|ибо вы и моим узам сострадали и расхищение имения вашего приняли с радостью, зная, что есть у вас на небесах имущество лучшее и непреходящее.
HEB|10|35|Итак не оставляйте упования вашего, которому предстоит великое воздаяние.
HEB|10|36|Терпение нужно вам, чтобы, исполнив волю Божию, получить обещанное;
HEB|10|37|ибо еще немного, очень немного, и Грядущий придет и не умедлит.
HEB|10|38|Праведный верою жив будет; а если [кто] поколеблется, не благоволит к тому душа Моя.
HEB|10|39|Мы же не из колеблющихся на погибель, но [стоим] в вере к спасению души.
HEB|11|1|Вера же есть осуществление ожидаемого и уверенность в невидимом.
HEB|11|2|В ней свидетельствованы древние.
HEB|11|3|Верою познаем, что веки устроены словом Божиим, так что из невидимого произошло видимое.
HEB|11|4|Верою Авель принес Богу жертву лучшую, нежели Каин; ею получил свидетельство, что он праведен, как засвидетельствовал Бог о дарах его; ею он и по смерти говорит еще.
HEB|11|5|Верою Енох переселен был так, что не видел смерти; и не стало его, потому что Бог переселил его. Ибо прежде переселения своего получил он свидетельство, что угодил Богу.
HEB|11|6|А без веры угодить Богу невозможно; ибо надобно, чтобы приходящий к Богу веровал, что Он есть, и ищущим Его воздает.
HEB|11|7|Верою Ной, получив откровение о том, что еще не было видимо, благоговея приготовил ковчег для спасения дома своего; ею осудил он (весь) мир, и сделался наследником праведности по вере.
HEB|11|8|Верою Авраам повиновался призванию идти в страну, которую имел получить в наследие, и пошел, не зная, куда идет.
HEB|11|9|Верою обитал он на земле обетованной, как на чужой, и жил в шатрах с Исааком и Иаковом, сонаследниками того же обетования;
HEB|11|10|ибо он ожидал города, имеющего основание, которого художник и строитель Бог.
HEB|11|11|Верою и сама Сарра (будучи неплодна) получила силу к принятию семени, и не по времени возраста родила, ибо знала, что верен Обещавший.
HEB|11|12|И потому от одного, и притом омертвелого, родилось так много, как [много] звезд на небе и как бесчислен песок на берегу морском.
HEB|11|13|Все сии умерли в вере, не получив обетований, а только издали видели оные, и радовались, и говорили о себе, что они странники и пришельцы на земле;
HEB|11|14|ибо те, которые так говорят, показывают, что они ищут отечества.
HEB|11|15|И если бы они в мыслях имели то [отечество], из которого вышли, то имели бы время возвратиться;
HEB|11|16|но они стремились к лучшему, то есть к небесному; посему и Бог не стыдится их, называя Себя их Богом: ибо Он приготовил им город.
HEB|11|17|Верою Авраам, будучи искушаем, принес в жертву Исаака и, имея обетование, принес единородного,
HEB|11|18|о котором было сказано: в Исааке наречется тебе семя.
HEB|11|19|Ибо он думал, что Бог силен и из мертвых воскресить, почему и получил его в предзнаменование.
HEB|11|20|Верою в будущее Исаак благословил Иакова и Исава.
HEB|11|21|Верою Иаков, умирая, благословил каждого сына Иосифова и поклонился на верх жезла своего.
HEB|11|22|Верою Иосиф, при кончине, напоминал об исходе сынов Израилевых и завещал о костях своих.
HEB|11|23|Верою Моисей по рождении три месяца скрываем был родителями своими, ибо видели они, что дитя прекрасно, и не устрашились царского повеления.
HEB|11|24|Верою Моисей, придя в возраст, отказался называться сыном дочери фараоновой,
HEB|11|25|и лучше захотел страдать с народом Божиим, нежели иметь временное греховное наслаждение,
HEB|11|26|и поношение Христово почел большим для себя богатством, нежели Египетские сокровища; ибо он взирал на воздаяние.
HEB|11|27|Верою оставил он Египет, не убоявшись гнева царского, ибо он, как бы видя Невидимого, был тверд.
HEB|11|28|Верою совершил он Пасху и пролитие крови, дабы истребитель первенцев не коснулся их.
HEB|11|29|Верою перешли они Чермное море, как по суше, – на что покусившись, Египтяне потонули.
HEB|11|30|Верою пали стены Иерихонские, по семидневном обхождении.
HEB|11|31|Верою Раав блудница, с миром приняв соглядатаев (и проводив их другим путем), не погибла с неверными.
HEB|11|32|И что еще скажу? Недостанет мне времени, чтобы повествовать о Гедеоне, о Вараке, о Самсоне и Иеффае, о Давиде, Самуиле и (других) пророках,
HEB|11|33|которые верою побеждали царства, творили правду, получали обетования, заграждали уста львов,
HEB|11|34|угашали силу огня, избегали острия меча, укреплялись от немощи, были крепки на войне, прогоняли полки чужих;
HEB|11|35|жены получали умерших своих воскресшими; иные же замучены были, не приняв освобождения, дабы получить лучшее воскресение;
HEB|11|36|другие испытали поругания и побои, а также узы и темницу,
HEB|11|37|были побиваемы камнями, перепиливаемы, подвергаемы пытке, умирали от меча, скитались в милотях и козьих кожах, терпя недостатки, скорби, озлобления;
HEB|11|38|те, которых весь мир не был достоин, скитались по пустыням и горам, по пещерам и ущельям земли.
HEB|11|39|И все сии, свидетельствованные в вере, не получили обещанного,
HEB|11|40|потому что Бог предусмотрел о нас нечто лучшее, дабы они не без нас достигли совершенства.
HEB|12|1|Посему и мы, имея вокруг себя такое облако свидетелей, свергнем с себя всякое бремя и запинающий нас грех и с терпением будем проходить предлежащее нам поприще,
HEB|12|2|взирая на начальника и совершителя веры Иисуса, Который, вместо предлежавшей Ему радости, претерпел крест, пренебрегши посрамление, и воссел одесную престола Божия.
HEB|12|3|Помыслите о Претерпевшем такое над Собою поругание от грешников, чтобы вам не изнемочь и не ослабеть душами вашими.
HEB|12|4|Вы еще не до крови сражались, подвизаясь против греха,
HEB|12|5|и забыли утешение, которое предлагается вам, как сынам: сын мой! не пренебрегай наказания Господня, и не унывай, когда Он обличает тебя.
HEB|12|6|Ибо Господь, кого любит, того наказывает; бьет же всякого сына, которого принимает.
HEB|12|7|Если вы терпите наказание, то Бог поступает с вами, как с сынами. Ибо есть ли какой сын, которого бы не наказывал отец?
HEB|12|8|Если же остаетесь без наказания, которое всем обще, то вы незаконные дети, а не сыны.
HEB|12|9|Притом, [если] мы, будучи наказываемы плотскими родителями нашими, боялись их, то не гораздо ли более должны покориться Отцу духов, чтобы жить?
HEB|12|10|Те наказывали нас по своему произволу для немногих дней; а Сей – для пользы, чтобы нам иметь участие в святости Его.
HEB|12|11|Всякое наказание в настоящее время кажется не радостью, а печалью; но после наученным через него доставляет мирный плод праведности.
HEB|12|12|Итак укрепите опустившиеся руки и ослабевшие колени
HEB|12|13|и ходите прямо ногами вашими, дабы хромлющее не совратилось, а лучше исправилось.
HEB|12|14|Старайтесь иметь мир со всеми и святость, без которой никто не увидит Господа.
HEB|12|15|Наблюдайте, чтобы кто не лишился благодати Божией; чтобы какой горький корень, возникнув, не причинил вреда, и чтобы им не осквернились многие;
HEB|12|16|чтобы не было [между вами] какого блудника, или нечестивца, который бы, как Исав, за одну снедь отказался от своего первородства.
HEB|12|17|Ибо вы знаете, что после того он, желая наследовать благословение, был отвержен; не мог переменить мыслей [отца], хотя и просил о том со слезами.
HEB|12|18|Вы приступили не к горе, осязаемой и пылающей огнем, не ко тьме и мраку и буре,
HEB|12|19|не к трубному звуку и гласу глаголов, который слышавшие просили, чтобы к ним более не было продолжаемо слово,
HEB|12|20|ибо они не могли стерпеть того, что заповедуемо было: если и зверь прикоснется к горе, будет побит камнями (или поражен стрелою);
HEB|12|21|и столь ужасно было это видение, [что и] Моисей сказал: "я в страхе и трепете".
HEB|12|22|Но вы приступили к горе Сиону и ко граду Бога живаго, к небесному Иерусалиму и тьмам Ангелов,
HEB|12|23|к торжествующему собору и церкви первенцев, написанных на небесах, и к Судии всех Богу, и к духам праведников, достигших совершенства,
HEB|12|24|и к Ходатаю нового завета Иисусу, и к Крови кропления, говорящей лучше, нежели Авелева.
HEB|12|25|Смотрите, не отвратитесь и вы от говорящего. Если те, не послушав глаголавшего на земле, не избегли [наказания], то тем более [не] [избежим] мы, если отвратимся от [Глаголющего] с небес,
HEB|12|26|Которого глас тогда поколебал землю, и Который ныне дал такое обещание: еще раз поколеблю не только землю, но и небо.
HEB|12|27|Слова: "еще раз" означают изменение колеблемого, как сотворенного, чтобы пребыло непоколебимое.
HEB|12|28|Итак мы, приемля царство непоколебимое, будем хранить благодать, которою будем служить благоугодно Богу, с благоговением и страхом,
HEB|12|29|потому что Бог наш есть огнь поядающий.
HEB|13|1|Братолюбие [между вами] да пребывает.
HEB|13|2|Страннолюбия не забывайте, ибо через него некоторые, не зная, оказали гостеприимство Ангелам.
HEB|13|3|Помните узников, как бы и вы с ними были в узах, и страждущих, как и сами находитесь в теле.
HEB|13|4|Брак у всех [да будет] честен и ложе непорочно; блудников же и прелюбодеев судит Бог.
HEB|13|5|Имейте нрав несребролюбивый, довольствуясь тем, что есть. Ибо Сам сказал: не оставлю тебя и не покину тебя,
HEB|13|6|так что мы смело говорим: Господь мне помощник, и не убоюсь: что сделает мне человек?
HEB|13|7|Поминайте наставников ваших, которые проповедывали вам слово Божие, и, взирая на кончину их жизни, подражайте вере их.
HEB|13|8|Иисус Христос вчера и сегодня и во веки Тот же.
HEB|13|9|Учениями различными и чуждыми не увлекайтесь; ибо хорошо благодатью укреплять сердца, а не яствами, от которых не получили пользы занимающиеся ими.
HEB|13|10|Мы имеем жертвенник, от которого не имеют права питаться служащие скинии.
HEB|13|11|Так как тела животных, которых кровь для [очищения] греха вносится первосвященником во святилище, сжигаются вне стана, –
HEB|13|12|то и Иисус, дабы освятить людей Кровию Своею, пострадал вне врат.
HEB|13|13|Итак выйдем к Нему за стан, нося Его поругание;
HEB|13|14|ибо не имеем здесь постоянного града, но ищем будущего.
HEB|13|15|Итак будем через Него непрестанно приносить Богу жертву хвалы, то есть плод уст, прославляющих имя Его.
HEB|13|16|Не забывайте также благотворения и общительности, ибо таковые жертвы благоугодны Богу.
HEB|13|17|Повинуйтесь наставникам вашим и будьте покорны, ибо они неусыпно пекутся о душах ваших, как обязанные дать отчет; чтобы они делали это с радостью, а не воздыхая, ибо это для вас неполезно.
HEB|13|18|Молитесь о нас; ибо мы уверены, что имеем добрую совесть, потому что во всем желаем вести себя честно.
HEB|13|19|Особенно же прошу делать это, дабы я скорее возвращен был вам.
HEB|13|20|Бог же мира, воздвигший из мертвых Пастыря овец великого Кровию завета вечного, Господа нашего Иисуса (Христа),
HEB|13|21|да усовершит вас во всяком добром деле, к исполнению воли Его, производя в вас благоугодное Ему через Иисуса Христа. Ему слава во веки веков! Аминь.
HEB|13|22|Прошу вас, братия, примите сие слово увещания; я же не много и написал вам.
HEB|13|23|Знайте, что брат наш Тимофей освобожден, и я вместе с ним, если он скоро придет, увижу вас.
HEB|13|24|Приветствуйте всех наставников ваших и всех святых. Приветствуют вас Италийские.
HEB|13|25|Благодать со всеми вами. Аминь.
