COL|1|1|奉上帝旨意，作基督耶穌使徒的 保羅 ，和我們的弟兄 提摩太 ，
COL|1|2|寫信給 歌羅西 的聖徒，在基督裏忠心的弟兄。願恩惠、平安 從我們的父上帝歸給你們！
COL|1|3|我們為你們禱告的時候，常常感謝我們主耶穌基督的父上帝 ，
COL|1|4|因為聽見你們對基督耶穌的信心，並對眾聖徒有的愛心。
COL|1|5|這都是因著那給你們存在天上的盼望，它就是你們從前所聽見真理的道，就是福音；
COL|1|6|這福音傳到你們那裏，也傳到普天下，並且繼續增長，不斷結果，正如自從你們聽見福音，真正知道上帝恩惠的日子起，在你們中間也是這樣。
COL|1|7|這福音是你們從我們所親愛、一同作僕人的 以巴弗 學到的。他為我們 作了基督的忠心僕役，
COL|1|8|也把聖靈賜給你們的愛告訴我們。
COL|1|9|因此，我們自從聽見的日子就不住地為你們禱告和祈求，願你們滿有一切屬靈的智慧和悟性，真正知道上帝的旨意，
COL|1|10|好使你們行事為人對得起主，凡事蒙他喜悅，在一切善事上結果子，對上帝的認識更有長進。
COL|1|11|願你們從他榮耀的權能中，得以在一切事上力上加力，好使你們凡事歡歡喜喜地忍耐寬容，
COL|1|12|又感謝父，使你們配與眾聖徒在光明中分享基業。
COL|1|13|他救了我們脫離黑暗的權勢，遷移到他愛子的國度裏。
COL|1|14|藉著他的愛子，我們得蒙救贖，罪得赦免。
COL|1|15|愛子是那看不見的上帝之像， 是首生的 ，在一切被造的以先。
COL|1|16|因為萬有都是在他裏面 造的， 無論是天上的、地上的， 能看見的、不能看見的， 或是有權位的、統治的， 或是執政的、掌權的， 一概都是藉著他為著他造的。
COL|1|17|他在萬有之先； 萬有也靠他而存在。
COL|1|18|他是身體（教會）的頭； 他是元始， 是從死人中復活的首生者， 好讓他在萬有中居首位。
COL|1|19|因為上帝喜歡使一切的豐盛在他裏面居住，
COL|1|20|藉著他 ，上帝使萬有與自己和好， 無論是地上的、天上的， 都藉著他在十字架上所流的血促成了和平。
COL|1|21|從前你們與上帝隔絕，心思上與他為敵，行為邪惡；
COL|1|22|但如今，他藉著他兒子肉身的死，已經使你們與他自己和好了 ，把你們獻在他的面前，成為聖潔，沒有瑕疵，無可指責。
COL|1|23|只要你們持守信仰，根基穩固，堅定不移，不致動搖，離開了你們從前所聽見的福音的盼望；這福音也是傳給天下一切被造之物的，我— 保羅 作了這福音的僕役。
COL|1|24|現在我為你們受苦，倒很快樂；並且為基督的身體，就是為教會，我要在自己的肉身上補滿基督未盡的苦難。
COL|1|25|我照上帝為你們所賜我的職分作了教會的僕役，要把上帝的道傳得完滿；
COL|1|26|這道就是歷世歷代所隱藏的奧祕，但如今向他的聖徒顯明了。
COL|1|27|上帝要讓他們知道，這奧祕在外邦人中有何等豐盛的榮耀；就是基督在你們心裏 成了得榮耀的盼望。
COL|1|28|我們傳揚他，是用諸般的智慧，勸戒各人，教導各人，要把各人在基督裏完完全全地獻上 。
COL|1|29|我也為此勞苦，照著他在我裏面運用的大能盡心竭力。
COL|2|1|我要你們知道，我為你們和 老底嘉 人，和所有沒有與我見過面的人，是何等地勤奮；
COL|2|2|為要使他們的心得安慰，因愛心互相聯絡，以致有從確實了解所產生的豐盛，好深知上帝的奧祕，就是基督；
COL|2|3|在他裏面蘊藏著一切智慧和知識。
COL|2|4|我說這話，免得有人用花言巧語迷惑你們。
COL|2|5|雖然我身體不在你們那裏，心卻與你們同在，很高興見你們循規蹈矩，對基督的信心也堅固。
COL|2|6|既然你們接受了主基督耶穌，就要靠著他而生活，
COL|2|7|照著你們所領受的教導，在他裏面生根建造，信心堅固，充滿著感謝的心。
COL|2|8|你們要謹慎，免得有人用他的哲學和虛空的廢話，不照著基督，而是照人間的傳統和世上粗淺的學說 ，把你們擄去。
COL|2|9|因為上帝本性一切的豐盛都有形有體地居住在基督裏面；
COL|2|10|你們在他裏面也已經成為豐盛。他是所有執政掌權者的元首。
COL|2|11|你們也在他裏面受了不是人手所行的割禮，而是使你們脫去肉體情慾的基督的割禮。
COL|2|12|你們既受洗與他一同埋葬，也就在此禮上，因信那使他從死人中復活的上帝的作為跟他一同復活。
COL|2|13|你們從前在過犯和未受割禮的肉體中死了，上帝卻赦免了你們一切的過犯，使你們與基督一同活過來，
COL|2|14|塗去了在律例上所寫、敵對我們、束縛我們的字據，把它撤去，釘在十字架上。
COL|2|15|基督既將一切執政者、掌權者的權勢解除了，就在凱旋的行列中，將他們公開示眾，仗著十字架誇勝。
COL|2|16|所以，不要讓任何人在飲食上，或節期、初一、安息日等事上評斷你們。
COL|2|17|這些原是未來的事的影子，真體卻是屬基督的。
COL|2|18|不要讓人藉著故作謙虛和敬拜天使奪去你們的獎賞。這等人拘泥在所見過的幻象 ，隨著自己的慾望無故地自高自大，
COL|2|19|不緊隨元首；其實，由於他全身藉著關節筋絡才得到滋養，互相聯絡，靠上帝所賜的成長而成長。
COL|2|20|既然你們與基督同死而脫離了世上粗淺的學說，為甚麼仍像生活在世俗中一樣，去服從那「不可拿、不可嘗、不可摸」等類的規條呢？
COL|2|21|
COL|2|22|這些都是根據人的命令和教導，論到這一切都是一經使用就都敗壞了。
COL|2|23|這些規條使人徒有智慧之名，用私意崇拜，自表謙卑，苦待己身，其實在克制肉體的情慾上毫無功效。
COL|3|1|所以，既然你們已經與基督一同復活，就當求上面的事；那裏有基督，坐在上帝的右邊。
COL|3|2|你們要思考上面的事，不要思考地上的事。
COL|3|3|因為你們已經死了，你們的生命與基督一同藏在上帝裏面。
COL|3|4|基督是你們的生命，他顯現的時候，你們也要與他一同在榮耀裏顯現。
COL|3|5|所以，要治死你們在地上的肢體；就如淫亂、污穢、邪情、惡慾和貪婪—貪婪就是拜偶像。
COL|3|6|因這些事，上帝的憤怒必臨到那些悖逆的人 。
COL|3|7|當你們在這些事中活著的時候，你們的行為也曾是這樣的。
COL|3|8|但現在你們要棄絕這一切的事，就是惱恨、憤怒、惡毒、毀謗和口中污穢的言語。
COL|3|9|不要彼此說謊，因為你們已經脫去舊人和舊人的行為，
COL|3|10|穿上了新人，這新人照著造他的主的形像在知識上不斷地更新。
COL|3|11|在這事上並不分 希臘 人和 猶太 人，受割禮的和未受割禮的，未開化的人、 西古提 人、為奴的、自主的；惟獨基督是一切，又在一切之內。
COL|3|12|所以，你們既是上帝的選民，聖潔、蒙愛的人，要穿上憐憫、恩慈、謙虛、溫柔和忍耐。
COL|3|13|倘若這人與那人有嫌隙，總要彼此容忍，彼此饒恕；主 怎樣饒恕了你們，你們也要怎樣饒恕人。
COL|3|14|除此以外，還要穿上愛心，因為愛是貫通全德的。
COL|3|15|你們要讓基督所賜的和平在你們心裏作主，也為此蒙召，歸為一體。你們還要存感謝的心。
COL|3|16|當用各樣的智慧，把基督的道豐豐富富的存在心裏，用詩篇、讚美詩、靈歌，彼此教導，互相勸戒，以感恩的心歌頌上帝。
COL|3|17|你們無論做甚麼，或說話或行事，都要奉主耶穌的名，藉著他感謝父上帝。
COL|3|18|你們作妻子的，要順服自己的丈夫，這在主裏面是合宜的。
COL|3|19|你們作丈夫的，要愛你們的妻子，不可虐待她們。
COL|3|20|你們作兒女的，要凡事聽從父母，因為這是主所喜悅的。
COL|3|21|你們作父親的，不要惹兒女生氣，恐怕他們會灰心。
COL|3|22|你們作僕人的，要凡事聽從你們肉身的主人，不要只在眼前服事，像是討人喜歡的，總要心存誠實，因為你們敬畏主。
COL|3|23|你們無論做甚麼，都要從心裏做，像是為主做的，不是為人做的；
COL|3|24|因為你們知道，從主那裏必得著基業作為賞賜。你們要服侍的是主基督。
COL|3|25|行不義的人必受不義的報應；主並不偏待人。
COL|4|1|你們作主人的，待僕人要公正，因為知道，你們也有一位主在天上。
COL|4|2|你們要恆切禱告，在禱告中警醒感恩。
COL|4|3|同時，也要為我們禱告，求上帝給我們開傳道的門，能宣講基督的奧祕，
COL|4|4|使我能按著所該說的話將這奧祕顯明出來，我為此而被捆鎖。
COL|4|5|你們要把握時機，用智慧與外人來往。
COL|4|6|你們的言談要時常帶著溫和，好像用鹽調味，讓你們知道該怎樣應對每一個人。
COL|4|7|推基古 是我親愛的弟兄，忠心的僕役，和我一同作主的僕人；他要把我一切的事都告訴你們。
COL|4|8|我特意打發他到你們那裏去，好讓你們知道我們的情況，又讓他安慰你們的心。
COL|4|9|我又打發一位親愛忠心的弟兄 阿尼西謀 同去；他也是你們那裏的人。他們會把這裏一切的事都告訴你們。
COL|4|10|與我一同坐牢的 亞里達古 問候你們。 巴拿巴 的表弟 馬可 也問候你們。關於他，你們已經得到指示；他若到你們那裏，你們要接待他。
COL|4|11|稱為 猶士都 的 耶數 也問候你們。奉割禮的人中，只有這三個人是為上帝的國與我作同工的，也是使我心裏得安慰的。
COL|4|12|有一位你們那裏的人，作基督耶穌 僕人的 以巴弗 問候你們。他禱告的時候常為你們竭力祈求，願你們能站穩而成熟，充分確信上帝一切的旨意。
COL|4|13|他為你們、 老底嘉 和 希拉坡里 的弟兄多多勞苦，這是我可以為他作見證的。
COL|4|14|親愛的醫生 路加 和 底馬 問候你們。
COL|4|15|請問候 老底嘉 的弟兄以及 寧法 ，和她家裏 的教會。
COL|4|16|你們宣讀了這書信，也要交給 老底嘉 的教會宣讀；你們也要宣讀從 老底嘉 轉來的書信。
COL|4|17|你們要對 亞基布 說：「務要完成你從主所領受的職分。」
COL|4|18|我— 保羅 親筆問候你們。要記念我在捆鎖中。願恩惠與你們同在！
