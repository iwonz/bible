MATT|1|1|Родословие Иисуса Христа, Сына Давидова, Сына Авраамова.
MATT|1|2|Авраам родил Исаака; Исаак родил Иакова; Иаков родил Иуду и братьев его;
MATT|1|3|Иуда родил Фареса и Зару от Фамари; Фарес родил Есрома; Есром родил Арама;
MATT|1|4|Арам родил Аминадава; Аминадав родил Наассона; Наассон родил Салмона;
MATT|1|5|Салмон родил Вооза от Рахавы; Вооз родил Овида от Руфи; Овид родил Иессея;
MATT|1|6|Иессей родил Давида царя; Давид царь родил Соломона от бывшей за Уриею;
MATT|1|7|Соломон родил Ровоама; Ровоам родил Авию; Авия родил Асу;
MATT|1|8|Аса родил Иосафата; Иосафат родил Иорама; Иорам родил Озию;
MATT|1|9|Озия родил Иоафама; Иоафам родил Ахаза; Ахаз родил Езекию;
MATT|1|10|Езекия родил Манассию; Манассия родил Амона; Амон родил Иосию;
MATT|1|11|Иосия родил Иоакима; Иоаким родил Иехонию и братьев его, перед переселением в Вавилон.
MATT|1|12|По переселении же в Вавилон, Иехония родил Салафииля; Салафииль родил Зоровавеля;
MATT|1|13|Зоровавель родил Авиуда; Авиуд родил Елиакима; Елиаким родил Азора;
MATT|1|14|Азор родил Садока; Садок родил Ахима; Ахим родил Елиуда;
MATT|1|15|Елиуд родил Елеазара; Елеазар родил Матфана; Матфан родил Иакова;
MATT|1|16|Иаков родил Иосифа, мужа Марии, от Которой родился Иисус, называемый Христос.
MATT|1|17|Итак всех родов от Авраама до Давида четырнадцать родов; и от Давида до переселения в Вавилон четырнадцать родов; и от переселения в Вавилон до Христа четырнадцать родов.
MATT|1|18|Рождество Иисуса Христа было так: по обручении Матери Его Марии с Иосифом, прежде нежели сочетались они, оказалось, что Она имеет во чреве от Духа Святаго.
MATT|1|19|Иосиф же муж Ее, будучи праведен и не желая огласить Ее, хотел тайно отпустить Ее.
MATT|1|20|Но когда он помыслил это, – се, Ангел Господень явился ему во сне и сказал: Иосиф, сын Давидов! не бойся принять Марию, жену твою, ибо родившееся в Ней есть от Духа Святаго;
MATT|1|21|родит же Сына, и наречешь Ему имя Иисус, ибо Он спасет людей Своих от грехов их.
MATT|1|22|А все сие произошло, да сбудется реченное Господом через пророка, который говорит:
MATT|1|23|се, Дева во чреве приимет и родит Сына, и нарекут имя Ему Еммануил, что значит: с нами Бог.
MATT|1|24|Встав от сна, Иосиф поступил, как повелел ему Ангел Господень, и принял жену свою,
MATT|1|25|и не знал Ее. Как наконец Она родила Сына Своего первенца, и он нарек Ему имя: Иисус.
MATT|2|1|Когда же Иисус родился в Вифлееме Иудейском во дни царя Ирода, пришли в Иерусалим волхвы с востока и говорят:
MATT|2|2|где родившийся Царь Иудейский? ибо мы видели звезду Его на востоке и пришли поклониться Ему.
MATT|2|3|Услышав это, Ирод царь встревожился, и весь Иерусалим с ним.
MATT|2|4|И, собрав всех первосвященников и книжников народных, спрашивал у них: где должно родиться Христу?
MATT|2|5|Они же сказали ему: в Вифлееме Иудейском, ибо так написано через пророка:
MATT|2|6|и ты, Вифлеем, земля Иудина, ничем не меньше воеводств Иудиных, ибо из тебя произойдет Вождь, Который упасет народ Мой, Израиля.
MATT|2|7|Тогда Ирод, тайно призвав волхвов, выведал от них время появления звезды
MATT|2|8|и, послав их в Вифлеем, сказал: пойдите, тщательно разведайте о Младенце и, когда найдете, известите меня, чтобы и мне пойти поклониться Ему.
MATT|2|9|Они, выслушав царя, пошли. И се, звезда, которую видели они на востоке, шла перед ними, [как] наконец пришла и остановилась над [местом], где был Младенец.
MATT|2|10|Увидев же звезду, они возрадовались радостью весьма великою,
MATT|2|11|и, войдя в дом, увидели Младенца с Мариею, Матерью Его, и, пав, поклонились Ему; и, открыв сокровища свои, принесли Ему дары: золото, ладан и смирну.
MATT|2|12|И, получив во сне откровение не возвращаться к Ироду, иным путем отошли в страну свою.
MATT|2|13|Когда же они отошли, – се, Ангел Господень является во сне Иосифу и говорит: встань, возьми Младенца и Матерь Его и беги в Египет, и будь там, доколе не скажу тебе, ибо Ирод хочет искать Младенца, чтобы погубить Его.
MATT|2|14|Он встал, взял Младенца и Матерь Его ночью и пошел в Египет,
MATT|2|15|и там был до смерти Ирода, да сбудется реченное Господом через пророка, который говорит: из Египта воззвал Я Сына Моего.
MATT|2|16|Тогда Ирод, увидев себя осмеянным волхвами, весьма разгневался, и послал избить всех младенцев в Вифлееме и во всех пределах его, от двух лет и ниже, по времени, которое выведал от волхвов.
MATT|2|17|Тогда сбылось реченное через пророка Иеремию, который говорит:
MATT|2|18|глас в Раме слышен, плач и рыдание и вопль великий; Рахиль плачет о детях своих и не хочет утешиться, ибо их нет.
MATT|2|19|По смерти же Ирода, – се, Ангел Господень во сне является Иосифу в Египте
MATT|2|20|и говорит: встань, возьми Младенца и Матерь Его и иди в землю Израилеву, ибо умерли искавшие души Младенца.
MATT|2|21|Он встал, взял Младенца и Матерь Его и пришел в землю Израилеву.
MATT|2|22|Услышав же, что Архелай царствует в Иудее вместо Ирода, отца своего, убоялся туда идти; но, получив во сне откровение, пошел в пределы Галилейские
MATT|2|23|и, придя, поселился в городе, называемом Назарет, да сбудется реченное через пророков, что Он Назореем наречется.
MATT|3|1|В те дни приходит Иоанн Креститель и проповедует в пустыне Иудейской
MATT|3|2|и говорит: покайтесь, ибо приблизилось Царство Небесное.
MATT|3|3|Ибо он тот, о котором сказал пророк Исаия: глас вопиющего в пустыне: приготовьте путь Господу, прямыми сделайте стези Ему.
MATT|3|4|Сам же Иоанн имел одежду из верблюжьего волоса и пояс кожаный на чреслах своих, а пищею его были акриды и дикий мед.
MATT|3|5|Тогда Иерусалим и вся Иудея и вся окрестность Иорданская выходили к нему
MATT|3|6|и крестились от него в Иордане, исповедуя грехи свои.
MATT|3|7|Увидев же Иоанн многих фарисеев и саддукеев, идущих к нему креститься, сказал им: порождения ехиднины! кто внушил вам бежать от будущего гнева?
MATT|3|8|сотворите же достойный плод покаяния
MATT|3|9|и не думайте говорить в себе: "отец у нас Авраам", ибо говорю вам, что Бог может из камней сих воздвигнуть детей Аврааму.
MATT|3|10|Уже и секира при корне дерев лежит: всякое дерево, не приносящее доброго плода, срубают и бросают в огонь.
MATT|3|11|Я крещу вас в воде в покаяние, но Идущий за мною сильнее меня; я не достоин понести обувь Его; Он будет крестить вас Духом Святым и огнем;
MATT|3|12|лопата Его в руке Его, и Он очистит гумно Свое и соберет пшеницу Свою в житницу, а солому сожжет огнем неугасимым.
MATT|3|13|Тогда приходит Иисус из Галилеи на Иордан к Иоанну креститься от него.
MATT|3|14|Иоанн же удерживал Его и говорил: мне надобно креститься от Тебя, и Ты ли приходишь ко мне?
MATT|3|15|Но Иисус сказал ему в ответ: оставь теперь, ибо так надлежит нам исполнить всякую правду. Тогда [Иоанн] допускает Его.
MATT|3|16|И, крестившись, Иисус тотчас вышел из воды, – и се, отверзлись Ему небеса, и увидел [Иоанн] Духа Божия, Который сходил, как голубь, и ниспускался на Него.
MATT|3|17|И се, глас с небес глаголющий: Сей есть Сын Мой возлюбленный, в Котором Мое благоволение.
MATT|4|1|Тогда Иисус возведен был Духом в пустыню, для искушения от диавола,
MATT|4|2|и, постившись сорок дней и сорок ночей, напоследок взалкал.
MATT|4|3|И приступил к Нему искуситель и сказал: если Ты Сын Божий, скажи, чтобы камни сии сделались хлебами.
MATT|4|4|Он же сказал ему в ответ: написано: не хлебом одним будет жить человек, но всяким словом, исходящим из уст Божиих.
MATT|4|5|Потом берет Его диавол в святой город и поставляет Его на крыле храма,
MATT|4|6|и говорит Ему: если Ты Сын Божий, бросься вниз, ибо написано: Ангелам Своим заповедает о Тебе, и на руках понесут Тебя, да не преткнешься о камень ногою Твоею.
MATT|4|7|Иисус сказал ему: написано также: не искушай Господа Бога твоего.
MATT|4|8|Опять берет Его диавол на весьма высокую гору и показывает Ему все царства мира и славу их,
MATT|4|9|и говорит Ему: все это дам Тебе, если, пав, поклонишься мне.
MATT|4|10|Тогда Иисус говорит ему: отойди от Меня, сатана, ибо написано: Господу Богу твоему поклоняйся и Ему одному служи.
MATT|4|11|Тогда оставляет Его диавол, и се, Ангелы приступили и служили Ему.
MATT|4|12|Услышав же Иисус, что Иоанн отдан [под стражу], удалился в Галилею
MATT|4|13|и, оставив Назарет, пришел и поселился в Капернауме приморском, в пределах Завулоновых и Неффалимовых,
MATT|4|14|да сбудется реченное через пророка Исаию, который говорит:
MATT|4|15|земля Завулонова и земля Неффалимова, на пути приморском, за Иорданом, Галилея языческая,
MATT|4|16|народ, сидящий во тьме, увидел свет великий, и сидящим в стране и тени смертной воссиял свет.
MATT|4|17|С того времени Иисус начал проповедывать и говорить: покайтесь, ибо приблизилось Царство Небесное.
MATT|4|18|Проходя же близ моря Галилейского, Он увидел двух братьев: Симона, называемого Петром, и Андрея, брата его, закидывающих сети в море, ибо они были рыболовы,
MATT|4|19|и говорит им: идите за Мною, и Я сделаю вас ловцами человеков.
MATT|4|20|И они тотчас, оставив сети, последовали за Ним.
MATT|4|21|Оттуда, идя далее, увидел Он других двух братьев, Иакова Зеведеева и Иоанна, брата его, в лодке с Зеведеем, отцом их, починивающих сети свои, и призвал их.
MATT|4|22|И они тотчас, оставив лодку и отца своего, последовали за Ним.
MATT|4|23|И ходил Иисус по всей Галилее, уча в синагогах их и проповедуя Евангелие Царствия, и исцеляя всякую болезнь и всякую немощь в людях.
MATT|4|24|И прошел о Нем слух по всей Сирии; и приводили к Нему всех немощных, одержимых различными болезнями и припадками, и бесноватых, и лунатиков, и расслабленных, и Он исцелял их.
MATT|4|25|И следовало за Ним множество народа из Галилеи и Десятиградия, и Иерусалима, и Иудеи, и из–за Иордана.
MATT|5|1|Увидев народ, Он взошел на гору; и, когда сел, приступили к Нему ученики Его.
MATT|5|2|И Он, отверзши уста Свои, учил их, говоря:
MATT|5|3|Блаженны нищие духом, ибо их есть Царство Небесное.
MATT|5|4|Блаженны плачущие, ибо они утешатся.
MATT|5|5|Блаженны кроткие, ибо они наследуют землю.
MATT|5|6|Блаженны алчущие и жаждущие правды, ибо они насытятся.
MATT|5|7|Блаженны милостивые, ибо они помилованы будут.
MATT|5|8|Блаженны чистые сердцем, ибо они Бога узрят.
MATT|5|9|Блаженны миротворцы, ибо они будут наречены сынами Божиими.
MATT|5|10|Блаженны изгнанные за правду, ибо их есть Царство Небесное.
MATT|5|11|Блаженны вы, когда будут поносить вас и гнать и всячески неправедно злословить за Меня.
MATT|5|12|Радуйтесь и веселитесь, ибо велика ваша награда на небесах: так гнали [и] пророков, бывших прежде вас.
MATT|5|13|Вы – соль земли. Если же соль потеряет силу, то чем сделаешь ее соленою? Она уже ни к чему негодна, как разве выбросить ее вон на попрание людям.
MATT|5|14|Вы – свет мира. Не может укрыться город, стоящий на верху горы.
MATT|5|15|И, зажегши свечу, не ставят ее под сосудом, но на подсвечнике, и светит всем в доме.
MATT|5|16|Так да светит свет ваш пред людьми, чтобы они видели ваши добрые дела и прославляли Отца вашего Небесного.
MATT|5|17|Не думайте, что Я пришел нарушить закон или пророков: не нарушить пришел Я, но исполнить.
MATT|5|18|Ибо истинно говорю вам: доколе не прейдет небо и земля, ни одна иота или ни одна черта не прейдет из закона, пока не исполнится все.
MATT|5|19|Итак, кто нарушит одну из заповедей сих малейших и научит так людей, тот малейшим наречется в Царстве Небесном; а кто сотворит и научит, тот великим наречется в Царстве Небесном.
MATT|5|20|Ибо, говорю вам, если праведность ваша не превзойдет праведности книжников и фарисеев, то вы не войдете в Царство Небесное.
MATT|5|21|Вы слышали, что сказано древним: не убивай, кто же убьет, подлежит суду.
MATT|5|22|А Я говорю вам, что всякий, гневающийся на брата своего напрасно, подлежит суду; кто же скажет брату своему: "рака", подлежит синедриону; а кто скажет: "безумный", подлежит геенне огненной.
MATT|5|23|Итак, если ты принесешь дар твой к жертвеннику и там вспомнишь, что брат твой имеет что–нибудь против тебя,
MATT|5|24|оставь там дар твой пред жертвенником, и пойди прежде примирись с братом твоим, и тогда приди и принеси дар твой.
MATT|5|25|Мирись с соперником твоим скорее, пока ты еще на пути с ним, чтобы соперник не отдал тебя судье, а судья не отдал бы тебя слуге, и не ввергли бы тебя в темницу;
MATT|5|26|истинно говорю тебе: ты не выйдешь оттуда, пока не отдашь до последнего кодранта.
MATT|5|27|Вы слышали, что сказано древним: не прелюбодействуй.
MATT|5|28|А Я говорю вам, что всякий, кто смотрит на женщину с вожделением, уже прелюбодействовал с нею в сердце своем.
MATT|5|29|Если же правый глаз твой соблазняет тебя, вырви его и брось от себя, ибо лучше для тебя, чтобы погиб один из членов твоих, а не все тело твое было ввержено в геенну.
MATT|5|30|И если правая твоя рука соблазняет тебя, отсеки ее и брось от себя, ибо лучше для тебя, чтобы погиб один из членов твоих, а не все тело твое было ввержено в геенну.
MATT|5|31|Сказано также, что если кто разведется с женою своею, пусть даст ей разводную.
MATT|5|32|А Я говорю вам: кто разводится с женою своею, кроме вины прелюбодеяния, тот подает ей повод прелюбодействовать; и кто женится на разведенной, тот прелюбодействует.
MATT|5|33|Еще слышали вы, что сказано древним: не преступай клятвы, но исполняй пред Господом клятвы твои.
MATT|5|34|А Я говорю вам: не клянись вовсе: ни небом, потому что оно престол Божий;
MATT|5|35|ни землею, потому что она подножие ног Его; ни Иерусалимом, потому что он город великого Царя;
MATT|5|36|ни головою твоею не клянись, потому что не можешь ни одного волоса сделать белым или черным.
MATT|5|37|Но да будет слово ваше: да, да; нет, нет; а что сверх этого, то от лукавого.
MATT|5|38|Вы слышали, что сказано: око за око и зуб за зуб.
MATT|5|39|А Я говорю вам: не противься злому. Но кто ударит тебя в правую щеку твою, обрати к нему и другую;
MATT|5|40|и кто захочет судиться с тобою и взять у тебя рубашку, отдай ему и верхнюю одежду;
MATT|5|41|и кто принудит тебя идти с ним одно поприще, иди с ним два.
MATT|5|42|Просящему у тебя дай, и от хотящего занять у тебя не отвращайся.
MATT|5|43|Вы слышали, что сказано: люби ближнего твоего и ненавидь врага твоего.
MATT|5|44|А Я говорю вам: любите врагов ваших, благословляйте проклинающих вас, благотворите ненавидящим вас и молитесь за обижающих вас и гонящих вас,
MATT|5|45|да будете сынами Отца вашего Небесного, ибо Он повелевает солнцу Своему восходить над злыми и добрыми и посылает дождь на праведных и неправедных.
MATT|5|46|Ибо если вы будете любить любящих вас, какая вам награда? Не то же ли делают и мытари?
MATT|5|47|И если вы приветствуете только братьев ваших, что особенного делаете? Не так же ли поступают и язычники?
MATT|5|48|Итак будьте совершенны, как совершен Отец ваш Небесный.
MATT|6|1|Смотрите, не творите милостыни вашей пред людьми с тем, чтобы они видели вас: иначе не будет вам награды от Отца вашего Небесного.
MATT|6|2|Итак, когда творишь милостыню, не труби перед собою, как делают лицемеры в синагогах и на улицах, чтобы прославляли их люди. Истинно говорю вам: они уже получают награду свою.
MATT|6|3|У тебя же, когда творишь милостыню, пусть левая рука твоя не знает, что делает правая,
MATT|6|4|чтобы милостыня твоя была втайне; и Отец твой, видящий тайное, воздаст тебе явно.
MATT|6|5|И, когда молишься, не будь, как лицемеры, которые любят в синагогах и на углах улиц, останавливаясь, молиться, чтобы показаться перед людьми. Истинно говорю вам, что они уже получают награду свою.
MATT|6|6|Ты же, когда молишься, войди в комнату твою и, затворив дверь твою, помолись Отцу твоему, Который втайне; и Отец твой, видящий тайное, воздаст тебе явно.
MATT|6|7|А молясь, не говорите лишнего, как язычники, ибо они думают, что в многословии своем будут услышаны;
MATT|6|8|не уподобляйтесь им, ибо знает Отец ваш, в чем вы имеете нужду, прежде вашего прошения у Него.
MATT|6|9|Молитесь же так: Отче наш, сущий на небесах! да святится имя Твое;
MATT|6|10|да приидет Царствие Твое; да будет воля Твоя и на земле, как на небе;
MATT|6|11|хлеб наш насущный дай нам на сей день;
MATT|6|12|и прости нам долги наши, как и мы прощаем должникам нашим;
MATT|6|13|и не введи нас в искушение, но избавь нас от лукавого. Ибо Твое есть Царство и сила и слава во веки. Аминь.
MATT|6|14|Ибо если вы будете прощать людям согрешения их, то простит и вам Отец ваш Небесный,
MATT|6|15|а если не будете прощать людям согрешения их, то и Отец ваш не простит вам согрешений ваших.
MATT|6|16|Также, когда поститесь, не будьте унылы, как лицемеры, ибо они принимают на себя мрачные лица, чтобы показаться людям постящимися. Истинно говорю вам, что они уже получают награду свою.
MATT|6|17|А ты, когда постишься, помажь голову твою и умой лице твое,
MATT|6|18|чтобы явиться постящимся не пред людьми, но пред Отцом твоим, Который втайне; и Отец твой, видящий тайное, воздаст тебе явно.
MATT|6|19|Не собирайте себе сокровищ на земле, где моль и ржа истребляют и где воры подкапывают и крадут,
MATT|6|20|но собирайте себе сокровища на небе, где ни моль, ни ржа не истребляют и где воры не подкапывают и не крадут,
MATT|6|21|ибо где сокровище ваше, там будет и сердце ваше.
MATT|6|22|Светильник для тела есть око. Итак, если око твое будет чисто, то все тело твое будет светло;
MATT|6|23|если же око твое будет худо, то все тело твое будет темно. Итак, если свет, который в тебе, тьма, то какова же тьма?
MATT|6|24|Никто не может служить двум господам: ибо или одного будет ненавидеть, а другого любить; или одному станет усердствовать, а о другом нерадеть. Не можете служить Богу и маммоне.
MATT|6|25|Посему говорю вам: не заботьтесь для души вашей, что вам есть и что пить, ни для тела вашего, во что одеться. Душа не больше ли пищи, и тело одежды?
MATT|6|26|Взгляните на птиц небесных: они ни сеют, ни жнут, ни собирают в житницы; и Отец ваш Небесный питает их. Вы не гораздо ли лучше их?
MATT|6|27|Да и кто из вас, заботясь, может прибавить себе росту [хотя] на один локоть?
MATT|6|28|И об одежде что заботитесь? Посмотрите на полевые лилии, как они растут: ни трудятся, ни прядут;
MATT|6|29|но говорю вам, что и Соломон во всей славе своей не одевался так, как всякая из них;
MATT|6|30|если же траву полевую, которая сегодня есть, а завтра будет брошена в печь, Бог так одевает, кольми паче вас, маловеры!
MATT|6|31|Итак не заботьтесь и не говорите: что нам есть? или что пить? или во что одеться?
MATT|6|32|потому что всего этого ищут язычники, и потому что Отец ваш Небесный знает, что вы имеете нужду во всем этом.
MATT|6|33|Ищите же прежде Царства Божия и правды Его, и это все приложится вам.
MATT|6|34|Итак не заботьтесь о завтрашнем дне, ибо завтрашний [сам] будет заботиться о своем: довольно для [каждого] дня своей заботы.
MATT|7|1|Не судите, да не судимы будете,
MATT|7|2|ибо каким судом судите, [таким] будете судимы; и какою мерою мерите, [такою] и вам будут мерить.
MATT|7|3|И что ты смотришь на сучок в глазе брата твоего, а бревна в твоем глазе не чувствуешь?
MATT|7|4|Или как скажешь брату твоему: "дай, я выну сучок из глаза твоего", а вот, в твоем глазе бревно?
MATT|7|5|Лицемер! вынь прежде бревно из твоего глаза и тогда увидишь, [как] вынуть сучок из глаза брата твоего.
MATT|7|6|Не давайте святыни псам и не бросайте жемчуга вашего перед свиньями, чтобы они не попрали его ногами своими и, обратившись, не растерзали вас.
MATT|7|7|Просите, и дано будет вам; ищите, и найдете; стучите, и отворят вам;
MATT|7|8|ибо всякий просящий получает, и ищущий находит, и стучащему отворят.
MATT|7|9|Есть ли между вами такой человек, который, когда сын его попросит у него хлеба, подал бы ему камень?
MATT|7|10|и когда попросит рыбы, подал бы ему змею?
MATT|7|11|Итак если вы, будучи злы, умеете даяния благие давать детям вашим, тем более Отец ваш Небесный даст блага просящим у Него.
MATT|7|12|Итак во всем, как хотите, чтобы с вами поступали люди, так поступайте и вы с ними, ибо в этом закон и пророки.
MATT|7|13|Входите тесными вратами, потому что широки врата и пространен путь, ведущие в погибель, и многие идут ими;
MATT|7|14|потому что тесны врата и узок путь, ведущие в жизнь, и немногие находят их.
MATT|7|15|Берегитесь лжепророков, которые приходят к вам в овечьей одежде, а внутри суть волки хищные.
MATT|7|16|По плодам их узнаете их. Собирают ли с терновника виноград, или с репейника смоквы?
MATT|7|17|Так всякое дерево доброе приносит и плоды добрые, а худое дерево приносит и плоды худые.
MATT|7|18|Не может дерево доброе приносить плоды худые, ни дерево худое приносить плоды добрые.
MATT|7|19|Всякое дерево, не приносящее плода доброго, срубают и бросают в огонь.
MATT|7|20|Итак по плодам их узнаете их.
MATT|7|21|Не всякий, говорящий Мне: "Господи! Господи!", войдет в Царство Небесное, но исполняющий волю Отца Моего Небесного.
MATT|7|22|Многие скажут Мне в тот день: Господи! Господи! не от Твоего ли имени мы пророчествовали? и не Твоим ли именем бесов изгоняли? и не Твоим ли именем многие чудеса творили?
MATT|7|23|И тогда объявлю им: Я никогда не знал вас; отойдите от Меня, делающие беззаконие.
MATT|7|24|Итак всякого, кто слушает слова Мои сии и исполняет их, уподоблю мужу благоразумному, который построил дом свой на камне;
MATT|7|25|и пошел дождь, и разлились реки, и подули ветры, и устремились на дом тот, и он не упал, потому что основан был на камне.
MATT|7|26|А всякий, кто слушает сии слова Мои и не исполняет их, уподобится человеку безрассудному, который построил дом свой на песке;
MATT|7|27|и пошел дождь, и разлились реки, и подули ветры, и налегли на дом тот; и он упал, и было падение его великое.
MATT|7|28|И когда Иисус окончил слова сии, народ дивился учению Его,
MATT|7|29|ибо Он учил их, как власть имеющий, а не как книжники и фарисеи.
MATT|8|1|Когда же сошел Он с горы, за Ним последовало множество народа.
MATT|8|2|И вот подошел прокаженный и, кланяясь Ему, сказал: Господи! если хочешь, можешь меня очистить.
MATT|8|3|Иисус, простерши руку, коснулся его и сказал: хочу, очистись. И он тотчас очистился от проказы.
MATT|8|4|И говорит ему Иисус: смотри, никому не сказывай, но пойди, покажи себя священнику и принеси дар, какой повелел Моисей, во свидетельство им.
MATT|8|5|Когда же вошел Иисус в Капернаум, к Нему подошел сотник и просил Его:
MATT|8|6|Господи! слуга мой лежит дома в расслаблении и жестоко страдает.
MATT|8|7|Иисус говорит ему: Я приду и исцелю его.
MATT|8|8|Сотник же, отвечая, сказал: Господи! я недостоин, чтобы Ты вошел под кров мой, но скажи только слово, и выздоровеет слуга мой;
MATT|8|9|ибо я и подвластный человек, но, имея у себя в подчинении воинов, говорю одному: пойди, и идет; и другому: приди, и приходит; и слуге моему: сделай то, и делает.
MATT|8|10|Услышав сие, Иисус удивился и сказал идущим за Ним: истинно говорю вам, и в Израиле не нашел Я такой веры.
MATT|8|11|Говорю же вам, что многие придут с востока и запада и возлягут с Авраамом, Исааком и Иаковом в Царстве Небесном;
MATT|8|12|а сыны царства извержены будут во тьму внешнюю: там будет плач и скрежет зубов.
MATT|8|13|И сказал Иисус сотнику: иди, и, как ты веровал, да будет тебе. И выздоровел слуга его в тот час.
MATT|8|14|Придя в дом Петров, Иисус увидел тещу его, лежащую в горячке,
MATT|8|15|и коснулся руки ее, и горячка оставила ее; и она встала и служила им.
MATT|8|16|Когда же настал вечер, к Нему привели многих бесноватых, и Он изгнал духов словом и исцелил всех больных,
MATT|8|17|да сбудется реченное через пророка Исаию, который говорит: Он взял на Себя наши немощи и понес болезни.
MATT|8|18|Увидев же Иисус вокруг Себя множество народа, велел ученикам отплыть на другую сторону.
MATT|8|19|Тогда один книжник, подойдя, сказал Ему: Учитель! я пойду за Тобою, куда бы Ты ни пошел.
MATT|8|20|И говорит ему Иисус: лисицы имеют норы и птицы небесные – гнезда, а Сын Человеческий не имеет, где приклонить голову.
MATT|8|21|Другой же из учеников Его сказал Ему: Господи! позволь мне прежде пойти и похоронить отца моего.
MATT|8|22|Но Иисус сказал ему: иди за Мною, и предоставь мертвым погребать своих мертвецов.
MATT|8|23|И когда вошел Он в лодку, за Ним последовали ученики Его.
MATT|8|24|И вот, сделалось великое волнение на море, так что лодка покрывалась волнами; а Он спал.
MATT|8|25|Тогда ученики Его, подойдя к Нему, разбудили Его и сказали: Господи! спаси нас, погибаем.
MATT|8|26|И говорит им: что вы [так] боязливы, маловерные? Потом, встав, запретил ветрам и морю, и сделалась великая тишина.
MATT|8|27|Люди же, удивляясь, говорили: кто это, что и ветры и море повинуются Ему?
MATT|8|28|И когда Он прибыл на другой берег в страну Гергесинскую, Его встретили два бесноватые, вышедшие из гробов, весьма свирепые, так что никто не смел проходить тем путем.
MATT|8|29|И вот, они закричали: что Тебе до нас, Иисус, Сын Божий? пришел Ты сюда прежде времени мучить нас.
MATT|8|30|Вдали же от них паслось большое стадо свиней.
MATT|8|31|И бесы просили Его: если выгонишь нас, то пошли нас в стадо свиней.
MATT|8|32|И Он сказал им: идите. И они, выйдя, пошли в стадо свиное. И вот, все стадо свиней бросилось с крутизны в море и погибло в воде.
MATT|8|33|Пастухи же побежали и, придя в город, рассказали обо всем, и о том, что было с бесноватыми.
MATT|8|34|И вот, весь город вышел навстречу Иисусу; и, увидев Его, просили, чтобы Он отошел от пределов их.
MATT|9|1|Тогда Он, войдя в лодку, переправился [обратно] и прибыл в Свой город.
MATT|9|2|И вот, принесли к Нему расслабленного, положенного на постели. И, видя Иисус веру их, сказал расслабленному: дерзай, чадо! прощаются тебе грехи твои.
MATT|9|3|При сем некоторые из книжников сказали сами в себе: Он богохульствует.
MATT|9|4|Иисус же, видя помышления их, сказал: для чего вы мыслите худое в сердцах ваших?
MATT|9|5|ибо что легче сказать: прощаются тебе грехи, или сказать: встань и ходи?
MATT|9|6|Но чтобы вы знали, что Сын Человеческий имеет власть на земле прощать грехи, – тогда говорит расслабленному: встань, возьми постель твою, и иди в дом твой.
MATT|9|7|И он встал, [взял постель свою] и пошел в дом свой.
MATT|9|8|Народ же, видев это, удивился и прославил Бога, давшего такую власть человекам.
MATT|9|9|Проходя оттуда, Иисус увидел человека, сидящего у сбора пошлин, по имени Матфея, и говорит ему: следуй за Мною. И он встал и последовал за Ним.
MATT|9|10|И когда Иисус возлежал в доме, многие мытари и грешники пришли и возлегли с Ним и учениками Его.
MATT|9|11|Увидев то, фарисеи сказали ученикам Его: для чего Учитель ваш ест и пьет с мытарями и грешниками?
MATT|9|12|Иисус же, услышав это, сказал им: не здоровые имеют нужду во враче, но больные,
MATT|9|13|пойдите, научитесь, что значит: милости хочу, а не жертвы? Ибо Я пришел призвать не праведников, но грешников к покаянию.
MATT|9|14|Тогда приходят к Нему ученики Иоанновы и говорят: почему мы и фарисеи постимся много, а Твои ученики не постятся?
MATT|9|15|И сказал им Иисус: могут ли печалиться сыны чертога брачного, пока с ними жених? Но придут дни, когда отнимется у них жених, и тогда будут поститься.
MATT|9|16|И никто к ветхой одежде не приставляет заплаты из небеленой ткани, ибо вновь пришитое отдерет от старого, и дыра будет еще хуже.
MATT|9|17|Не вливают также вина молодого в мехи ветхие; а иначе прорываются мехи, и вино вытекает, и мехи пропадают, но вино молодое вливают в новые мехи, и сберегается то и другое.
MATT|9|18|Когда Он говорил им сие, подошел к Нему некоторый начальник и, кланяясь Ему, говорил: дочь моя теперь умирает; но приди, возложи на нее руку Твою, и она будет жива.
MATT|9|19|И встав, Иисус пошел за ним, и ученики Его.
MATT|9|20|И вот, женщина, двенадцать лет страдавшая кровотечением, подойдя сзади, прикоснулась к краю одежды Его,
MATT|9|21|ибо она говорила сама в себе: если только прикоснусь к одежде Его, выздоровею.
MATT|9|22|Иисус же, обратившись и увидев ее, сказал: дерзай, дщерь! вера твоя спасла тебя. Женщина с того часа стала здорова.
MATT|9|23|И когда пришел Иисус в дом начальника и увидел свирельщиков и народ в смятении,
MATT|9|24|сказал им: выйдите вон, ибо не умерла девица, но спит. И смеялись над Ним.
MATT|9|25|Когда же народ был выслан, Он, войдя, взял ее за руку, и девица встала.
MATT|9|26|И разнесся слух о сем по всей земле той.
MATT|9|27|Когда Иисус шел оттуда, за Ним следовали двое слепых и кричали: помилуй нас, Иисус, сын Давидов!
MATT|9|28|Когда же Он пришел в дом, слепые приступили к Нему. И говорит им Иисус: веруете ли, что Я могу это сделать? Они говорят Ему: ей, Господи!
MATT|9|29|Тогда Он коснулся глаз их и сказал: по вере вашей да будет вам.
MATT|9|30|И открылись глаза их; и Иисус строго сказал им: смотрите, чтобы никто не узнал.
MATT|9|31|А они, выйдя, разгласили о Нем по всей земле той.
MATT|9|32|Когда же те выходили, то привели к Нему человека немого бесноватого.
MATT|9|33|И когда бес был изгнан, немой стал говорить. И народ, удивляясь, говорил: никогда не бывало такого явления в Израиле.
MATT|9|34|А фарисеи говорили: Он изгоняет бесов силою князя бесовского.
MATT|9|35|И ходил Иисус по всем городам и селениям, уча в синагогах их, проповедуя Евангелие Царствия и исцеляя всякую болезнь и всякую немощь в людях.
MATT|9|36|Видя толпы народа, Он сжалился над ними, что они были изнурены и рассеяны, как овцы, не имеющие пастыря.
MATT|9|37|Тогда говорит ученикам Своим: жатвы много, а делателей мало;
MATT|9|38|итак молите Господина жатвы, чтобы выслал делателей на жатву Свою.
MATT|10|1|И призвав двенадцать учеников Своих, Он дал им власть над нечистыми духами, чтобы изгонять их и врачевать всякую болезнь и всякую немощь.
MATT|10|2|Двенадцати же Апостолов имена суть сии: первый Симон, называемый Петром, и Андрей, брат его, Иаков Зеведеев и Иоанн, брат его,
MATT|10|3|Филипп и Варфоломей, Фома и Матфей мытарь, Иаков Алфеев и Леввей, прозванный Фаддеем,
MATT|10|4|Симон Кананит и Иуда Искариот, который и предал Его.
MATT|10|5|Сих двенадцать послал Иисус, и заповедал им, говоря: на путь к язычникам не ходите, и в город Самарянский не входите;
MATT|10|6|а идите наипаче к погибшим овцам дома Израилева;
MATT|10|7|ходя же, проповедуйте, что приблизилось Царство Небесное;
MATT|10|8|больных исцеляйте, прокаженных очищайте, мертвых воскрешайте, бесов изгоняйте; даром получили, даром давайте.
MATT|10|9|Не берите с собою ни золота, ни серебра, ни меди в поясы свои,
MATT|10|10|ни сумы на дорогу, ни двух одежд, ни обуви, ни посоха, ибо трудящийся достоин пропитания.
MATT|10|11|В какой бы город или селение ни вошли вы, наведывайтесь, кто в нем достоин, и там оставайтесь, пока не выйдете;
MATT|10|12|а входя в дом, приветствуйте его, говоря: мир дому сему;
MATT|10|13|и если дом будет достоин, то мир ваш придет на него; если же не будет достоин, то мир ваш к вам возвратится.
MATT|10|14|А если кто не примет вас и не послушает слов ваших, то, выходя из дома или из города того, отрясите прах от ног ваших;
MATT|10|15|истинно говорю вам: отраднее будет земле Содомской и Гоморрской в день суда, нежели городу тому.
MATT|10|16|Вот, Я посылаю вас, как овец среди волков: итак будьте мудры, как змии, и просты, как голуби.
MATT|10|17|Остерегайтесь же людей: ибо они будут отдавать вас в судилища и в синагогах своих будут бить вас,
MATT|10|18|и поведут вас к правителям и царям за Меня, для свидетельства перед ними и язычниками.
MATT|10|19|Когда же будут предавать вас, не заботьтесь, как или что сказать; ибо в тот час дано будет вам, что сказать,
MATT|10|20|ибо не вы будете говорить, но Дух Отца вашего будет говорить в вас.
MATT|10|21|Предаст же брат брата на смерть, и отец – сына; и восстанут дети на родителей, и умертвят их;
MATT|10|22|и будете ненавидимы всеми за имя Мое; претерпевший же до конца спасется.
MATT|10|23|Когда же будут гнать вас в одном городе, бегите в другой. Ибо истинно говорю вам: не успеете обойти городов Израилевых, как приидет Сын Человеческий.
MATT|10|24|Ученик не выше учителя, и слуга не выше господина своего:
MATT|10|25|довольно для ученика, чтобы он был, как учитель его, и для слуги, чтобы он был, как господин его. Если хозяина дома назвали веельзевулом, не тем ли более домашних его?
MATT|10|26|Итак не бойтесь их, ибо нет ничего сокровенного, что не открылось бы, и тайного, что не было бы узнано.
MATT|10|27|Что говорю вам в темноте, говорите при свете; и что на ухо слышите, проповедуйте на кровлях.
MATT|10|28|И не бойтесь убивающих тело, души же не могущих убить; а бойтесь более Того, Кто может и душу и тело погубить в геенне.
MATT|10|29|Не две ли малые птицы продаются за ассарий? И ни одна из них не упадет на землю без [воли] Отца вашего;
MATT|10|30|у вас же и волосы на голове все сочтены;
MATT|10|31|не бойтесь же: вы лучше многих малых птиц.
MATT|10|32|Итак всякого, кто исповедает Меня пред людьми, того исповедаю и Я пред Отцем Моим Небесным;
MATT|10|33|а кто отречется от Меня пред людьми, отрекусь от того и Я пред Отцем Моим Небесным.
MATT|10|34|Не думайте, что Я пришел принести мир на землю; не мир пришел Я принести, но меч,
MATT|10|35|ибо Я пришел разделить человека с отцом его, и дочь с матерью ее, и невестку со свекровью ее.
MATT|10|36|И враги человеку – домашние его.
MATT|10|37|Кто любит отца или мать более, нежели Меня, не достоин Меня; и кто любит сына или дочь более, нежели Меня, не достоин Меня;
MATT|10|38|и кто не берет креста своего и следует за Мною, тот не достоин Меня.
MATT|10|39|Сберегший душу свою потеряет ее; а потерявший душу свою ради Меня сбережет ее.
MATT|10|40|Кто принимает вас, принимает Меня, а кто принимает Меня, принимает Пославшего Меня;
MATT|10|41|кто принимает пророка, во имя пророка, получит награду пророка; и кто принимает праведника, во имя праведника, получит награду праведника.
MATT|10|42|И кто напоит одного из малых сих только чашею холодной воды, во имя ученика, истинно говорю вам, не потеряет награды своей.
MATT|11|1|И когда окончил Иисус наставления двенадцати ученикам Своим, перешел оттуда учить и проповедывать в городах их.
MATT|11|2|Иоанн же, услышав в темнице о делах Христовых, послал двоих из учеников своих
MATT|11|3|сказать Ему: Ты ли Тот, Который должен придти, или ожидать нам другого?
MATT|11|4|И сказал им Иисус в ответ: пойдите, скажите Иоанну, что слышите и видите:
MATT|11|5|слепые прозревают и хромые ходят, прокаженные очищаются и глухие слышат, мертвые воскресают и нищие благовествуют;
MATT|11|6|и блажен, кто не соблазнится о Мне.
MATT|11|7|Когда же они пошли, Иисус начал говорить народу об Иоанне: что смотреть ходили вы в пустыню? трость ли, ветром колеблемую?
MATT|11|8|Что же смотреть ходили вы? человека ли, одетого в мягкие одежды? Носящие мягкие одежды находятся в чертогах царских.
MATT|11|9|Что же смотреть ходили вы? пророка? Да, говорю вам, и больше пророка.
MATT|11|10|Ибо он тот, о котором написано: се, Я посылаю Ангела Моего пред лицем Твоим, который приготовит путь Твой пред Тобою.
MATT|11|11|Истинно говорю вам: из рожденных женами не восставал больший Иоанна Крестителя; но меньший в Царстве Небесном больше его.
MATT|11|12|От дней же Иоанна Крестителя доныне Царство Небесное силою берется, и употребляющие усилие восхищают его,
MATT|11|13|ибо все пророки и закон прорекли до Иоанна.
MATT|11|14|И если хотите принять, он есть Илия, которому должно придти.
MATT|11|15|Кто имеет уши слышать, да слышит!
MATT|11|16|Но кому уподоблю род сей? Он подобен детям, которые сидят на улице и, обращаясь к своим товарищам,
MATT|11|17|говорят: мы играли вам на свирели, и вы не плясали; мы пели вам печальные песни, и вы не рыдали.
MATT|11|18|Ибо пришел Иоанн, ни ест, ни пьет; и говорят: в нем бес.
MATT|11|19|Пришел Сын Человеческий, ест и пьет; и говорят: вот человек, который любит есть и пить вино, друг мытарям и грешникам. И оправдана премудрость чадами ее.
MATT|11|20|Тогда начал Он укорять города, в которых наиболее явлено было сил Его, за то, что они не покаялись:
MATT|11|21|горе тебе, Хоразин! горе тебе, Вифсаида! ибо если бы в Тире и Сидоне явлены были силы, явленные в вас, то давно бы они во вретище и пепле покаялись,
MATT|11|22|но говорю вам: Тиру и Сидону отраднее будет в день суда, нежели вам.
MATT|11|23|И ты, Капернаум, до неба вознесшийся, до ада низвергнешься, ибо если бы в Содоме явлены были силы, явленные в тебе, то он оставался бы до сего дня;
MATT|11|24|но говорю вам, что земле Содомской отраднее будет в день суда, нежели тебе.
MATT|11|25|В то время, продолжая речь, Иисус сказал: славлю Тебя, Отче, Господи неба и земли, что Ты утаил сие от мудрых и разумных и открыл то младенцам;
MATT|11|26|ей, Отче! ибо таково было Твое благоволение.
MATT|11|27|Все предано Мне Отцем Моим, и никто не знает Сына, кроме Отца; и Отца не знает никто, кроме Сына, и кому Сын хочет открыть.
MATT|11|28|Придите ко Мне все труждающиеся и обремененные, и Я успокою вас;
MATT|11|29|возьмите иго Мое на себя и научитесь от Меня, ибо Я кроток и смирен сердцем, и найдете покой душам вашим;
MATT|11|30|ибо иго Мое благо, и бремя Мое легко.
MATT|12|1|В то время проходил Иисус в субботу засеянными полями; ученики же Его взалкали и начали срывать колосья и есть.
MATT|12|2|Фарисеи, увидев это, сказали Ему: вот, ученики Твои делают, чего не должно делать в субботу.
MATT|12|3|Он же сказал им: разве вы не читали, что сделал Давид, когда взалкал сам и бывшие с ним?
MATT|12|4|как он вошел в дом Божий и ел хлебы предложения, которых не должно было есть ни ему, ни бывшим с ним, а только одним священникам?
MATT|12|5|Или не читали ли вы в законе, что в субботы священники в храме нарушают субботу, однако невиновны?
MATT|12|6|Но говорю вам, что здесь Тот, Кто больше храма;
MATT|12|7|если бы вы знали, что значит: милости хочу, а не жертвы, то не осудили бы невиновных,
MATT|12|8|ибо Сын Человеческий есть господин и субботы.
MATT|12|9|И, отойдя оттуда, вошел Он в синагогу их.
MATT|12|10|И вот, там был человек, имеющий сухую руку. И спросили Иисуса, чтобы обвинить Его: можно ли исцелять в субботы?
MATT|12|11|Он же сказал им: кто из вас, имея одну овцу, если она в субботу упадет в яму, не возьмет ее и не вытащит?
MATT|12|12|Сколько же лучше человек овцы! Итак можно в субботы делать добро.
MATT|12|13|Тогда говорит человеку тому: протяни руку твою. И он протянул, и стала она здорова, как другая.
MATT|12|14|Фарисеи же, выйдя, имели совещание против Него, как бы погубить Его. Но Иисус, узнав, удалился оттуда.
MATT|12|15|И последовало за Ним множество народа, и Он исцелил их всех
MATT|12|16|и запретил им объявлять о Нем,
MATT|12|17|да сбудется реченное через пророка Исаию, который говорит:
MATT|12|18|Се, Отрок Мой, Которого Я избрал, Возлюбленный Мой, Которому благоволит душа Моя. Положу дух Мой на Него, и возвестит народам суд;
MATT|12|19|не воспрекословит, не возопиет, и никто не услышит на улицах голоса Его;
MATT|12|20|трости надломленной не переломит, и льна курящегося не угасит, доколе не доставит суду победы;
MATT|12|21|и на имя Его будут уповать народы.
MATT|12|22|Тогда привели к Нему бесноватого слепого и немого; и исцелил его, так что слепой и немой стал и говорить и видеть.
MATT|12|23|И дивился весь народ и говорил: не это ли Христос, сын Давидов?
MATT|12|24|Фарисеи же, услышав [сие], сказали: Он изгоняет бесов не иначе, как [силою] веельзевула, князя бесовского.
MATT|12|25|Но Иисус, зная помышления их, сказал им: всякое царство, разделившееся само в себе, опустеет; и всякий город или дом, разделившийся сам в себе, не устоит.
MATT|12|26|И если сатана сатану изгоняет, то он разделился сам с собою: как же устоит царство его?
MATT|12|27|И если Я [силою] веельзевула изгоняю бесов, то сыновья ваши чьею [силою] изгоняют? Посему они будут вам судьями.
MATT|12|28|Если же Я Духом Божиим изгоняю бесов, то конечно достигло до вас Царствие Божие.
MATT|12|29|Или, как может кто войти в дом сильного и расхитить вещи его, если прежде не свяжет сильного? и тогда расхитит дом его.
MATT|12|30|Кто не со Мною, тот против Меня; и кто не собирает со Мною, тот расточает.
MATT|12|31|Посему говорю вам: всякий грех и хула простятся человекам, а хула на Духа не простится человекам;
MATT|12|32|если кто скажет слово на Сына Человеческого, простится ему; если же кто скажет на Духа Святаго, не простится ему ни в сем веке, ни в будущем.
MATT|12|33|Или признайте дерево хорошим и плод его хорошим; или признайте дерево худым и плод его худым, ибо дерево познается по плоду.
MATT|12|34|Порождения ехиднины! как вы можете говорить доброе, будучи злы? Ибо от избытка сердца говорят уста.
MATT|12|35|Добрый человек из доброго сокровища выносит доброе, а злой человек из злого сокровища выносит злое.
MATT|12|36|Говорю же вам, что за всякое праздное слово, какое скажут люди, дадут они ответ в день суда:
MATT|12|37|ибо от слов своих оправдаешься, и от слов своих осудишься.
MATT|12|38|Тогда некоторые из книжников и фарисеев сказали: Учитель! хотелось бы нам видеть от Тебя знамение.
MATT|12|39|Но Он сказал им в ответ: род лукавый и прелюбодейный ищет знамения; и знамение не дастся ему, кроме знамения Ионы пророка;
MATT|12|40|ибо как Иона был во чреве кита три дня и три ночи, так и Сын Человеческий будет в сердце земли три дня и три ночи.
MATT|12|41|Ниневитяне восстанут на суд с родом сим и осудят его, ибо они покаялись от проповеди Иониной; и вот, здесь больше Ионы.
MATT|12|42|Царица южная восстанет на суд с родом сим и осудит его, ибо она приходила от пределов земли послушать мудрости Соломоновой; и вот, здесь больше Соломона.
MATT|12|43|Когда нечистый дух выйдет из человека, то ходит по безводным местам, ища покоя, и не находит;
MATT|12|44|тогда говорит: возвращусь в дом мой, откуда я вышел. И, придя, находит [его] незанятым, выметенным и убранным;
MATT|12|45|тогда идет и берет с собою семь других духов, злейших себя, и, войдя, живут там; и бывает для человека того последнее хуже первого. Так будет и с этим злым родом.
MATT|12|46|Когда же Он еще говорил к народу, Матерь и братья Его стояли вне [дома], желая говорить с Ним.
MATT|12|47|И некто сказал Ему: вот Матерь Твоя и братья Твои стоят вне, желая говорить с Тобою.
MATT|12|48|Он же сказал в ответ говорившему: кто Матерь Моя? и кто братья Мои?
MATT|12|49|И, указав рукою Своею на учеников Своих, сказал: вот матерь Моя и братья Мои;
MATT|12|50|ибо, кто будет исполнять волю Отца Моего Небесного, тот Мне брат, и сестра, и матерь.
MATT|13|1|Выйдя же в день тот из дома, Иисус сел у моря.
MATT|13|2|И собралось к Нему множество народа, так что Он вошел в лодку и сел; а весь народ стоял на берегу.
MATT|13|3|И поучал их много притчами, говоря: вот, вышел сеятель сеять;
MATT|13|4|и когда он сеял, иное упало при дороге, и налетели птицы и поклевали то;
MATT|13|5|иное упало на места каменистые, где немного было земли, и скоро взошло, потому что земля была неглубока.
MATT|13|6|Когда же взошло солнце, увяло, и, как не имело корня, засохло;
MATT|13|7|иное упало в терние, и выросло терние и заглушило его;
MATT|13|8|иное упало на добрую землю и принесло плод: одно во сто крат, а другое в шестьдесят, иное же в тридцать.
MATT|13|9|Кто имеет уши слышать, да слышит!
MATT|13|10|И, приступив, ученики сказали Ему: для чего притчами говоришь им?
MATT|13|11|Он сказал им в ответ: для того, что вам дано знать тайны Царствия Небесного, а им не дано,
MATT|13|12|ибо кто имеет, тому дано будет и приумножится, а кто не имеет, у того отнимется и то, что имеет;
MATT|13|13|потому говорю им притчами, что они видя не видят, и слыша не слышат, и не разумеют;
MATT|13|14|и сбывается над ними пророчество Исаии, которое говорит: слухом услышите – и не уразумеете, и глазами смотреть будете – и не увидите,
MATT|13|15|ибо огрубело сердце людей сих и ушами с трудом слышат, и глаза свои сомкнули, да не увидят глазами и не услышат ушами, и не уразумеют сердцем, и да не обратятся, чтобы Я исцелил их.
MATT|13|16|Ваши же блаженны очи, что видят, и уши ваши, что слышат,
MATT|13|17|ибо истинно говорю вам, что многие пророки и праведники желали видеть, что вы видите, и не видели, и слышать, что вы слышите, и не слышали.
MATT|13|18|Вы же выслушайте [значение] притчи о сеятеле:
MATT|13|19|ко всякому, слушающему слово о Царствии и не разумеющему, приходит лукавый и похищает посеянное в сердце его – вот кого означает посеянное при дороге.
MATT|13|20|А посеянное на каменистых местах означает того, кто слышит слово и тотчас с радостью принимает его;
MATT|13|21|но не имеет в себе корня и непостоянен: когда настанет скорбь или гонение за слово, тотчас соблазняется.
MATT|13|22|А посеянное в тернии означает того, кто слышит слово, но забота века сего и обольщение богатства заглушает слово, и оно бывает бесплодно.
MATT|13|23|Посеянное же на доброй земле означает слышащего слово и разумеющего, который и бывает плодоносен, так что иной приносит плод во сто крат, иной в шестьдесят, а иной в тридцать.
MATT|13|24|Другую притчу предложил Он им, говоря: Царство Небесное подобно человеку, посеявшему доброе семя на поле своем;
MATT|13|25|когда же люди спали, пришел враг его и посеял между пшеницею плевелы и ушел;
MATT|13|26|когда взошла зелень и показался плод, тогда явились и плевелы.
MATT|13|27|Придя же, рабы домовладыки сказали ему: господин! не доброе ли семя сеял ты на поле твоем? откуда же на нем плевелы?
MATT|13|28|Он же сказал им: враг человека сделал это. А рабы сказали ему: хочешь ли, мы пойдем, выберем их?
MATT|13|29|Но он сказал: нет, – чтобы, выбирая плевелы, вы не выдергали вместе с ними пшеницы,
MATT|13|30|оставьте расти вместе то и другое до жатвы; и во время жатвы я скажу жнецам: соберите прежде плевелы и свяжите их в связки, чтобы сжечь их, а пшеницу уберите в житницу мою.
MATT|13|31|Иную притчу предложил Он им, говоря: Царство Небесное подобно зерну горчичному, которое человек взял и посеял на поле своем,
MATT|13|32|которое, хотя меньше всех семян, но, когда вырастет, бывает больше всех злаков и становится деревом, так что прилетают птицы небесные и укрываются в ветвях его.
MATT|13|33|Иную притчу сказал Он им: Царство Небесное подобно закваске, которую женщина, взяв, положила в три меры муки, доколе не вскисло все.
MATT|13|34|Все сие Иисус говорил народу притчами, и без притчи не говорил им,
MATT|13|35|да сбудется реченное через пророка, который говорит: отверзу в притчах уста Мои; изреку сокровенное от создания мира.
MATT|13|36|Тогда Иисус, отпустив народ, вошел в дом. И, приступив к Нему, ученики Его сказали: изъясни нам притчу о плевелах на поле.
MATT|13|37|Он же сказал им в ответ: сеющий доброе семя есть Сын Человеческий;
MATT|13|38|поле есть мир; доброе семя, это сыны Царствия, а плевелы – сыны лукавого;
MATT|13|39|враг, посеявший их, есть диавол; жатва есть кончина века, а жнецы суть Ангелы.
MATT|13|40|Посему как собирают плевелы и огнем сжигают, так будет при кончине века сего:
MATT|13|41|пошлет Сын Человеческий Ангелов Своих, и соберут из Царства Его все соблазны и делающих беззаконие,
MATT|13|42|и ввергнут их в печь огненную; там будет плач и скрежет зубов;
MATT|13|43|тогда праведники воссияют, как солнце, в Царстве Отца их. Кто имеет уши слышать, да слышит!
MATT|13|44|Еще подобно Царство Небесное сокровищу, скрытому на поле, которое, найдя, человек утаил, и от радости о нем идет и продает все, что имеет, и покупает поле то.
MATT|13|45|Еще подобно Царство Небесное купцу, ищущему хороших жемчужин,
MATT|13|46|который, найдя одну драгоценную жемчужину, пошел и продал все, что имел, и купил ее.
MATT|13|47|Еще подобно Царство Небесное неводу, закинутому в море и захватившему рыб всякого рода,
MATT|13|48|который, когда наполнился, вытащили на берег и, сев, хорошее собрали в сосуды, а худое выбросили вон.
MATT|13|49|Так будет при кончине века: изыдут Ангелы, и отделят злых из среды праведных,
MATT|13|50|и ввергнут их в печь огненную: там будет плач и скрежет зубов.
MATT|13|51|И спросил их Иисус: поняли ли вы все это? Они говорят Ему: так, Господи!
MATT|13|52|Он же сказал им: поэтому всякий книжник, наученный Царству Небесному, подобен хозяину, который выносит из сокровищницы своей новое и старое.
MATT|13|53|И, когда окончил Иисус притчи сии, пошел оттуда.
MATT|13|54|И, придя в отечество Свое, учил их в синагоге их, так что они изумлялись и говорили: откуда у Него такая премудрость и силы?
MATT|13|55|не плотников ли Он сын? не Его ли Мать называется Мария, и братья Его Иаков и Иосий, и Симон, и Иуда?
MATT|13|56|и сестры Его не все ли между нами? откуда же у Него все это?
MATT|13|57|И соблазнялись о Нем. Иисус же сказал им: не бывает пророк без чести, разве только в отечестве своем и в доме своем.
MATT|13|58|И не совершил там многих чудес по неверию их.
MATT|14|1|В то время Ирод четвертовластник услышал молву об Иисусе
MATT|14|2|и сказал служащим при нем: это Иоанн Креститель; он воскрес из мертвых, и потому чудеса делаются им.
MATT|14|3|Ибо Ирод, взяв Иоанна, связал его и посадил в темницу за Иродиаду, жену Филиппа, брата своего,
MATT|14|4|потому что Иоанн говорил ему: не должно тебе иметь ее.
MATT|14|5|И хотел убить его, но боялся народа, потому что его почитали за пророка.
MATT|14|6|Во время же [празднования] дня рождения Ирода дочь Иродиады плясала перед собранием и угодила Ироду,
MATT|14|7|посему он с клятвою обещал ей дать, чего она ни попросит.
MATT|14|8|Она же, по наущению матери своей, сказала: дай мне здесь на блюде голову Иоанна Крестителя.
MATT|14|9|И опечалился царь, но, ради клятвы и возлежащих с ним, повелел дать ей,
MATT|14|10|и послал отсечь Иоанну голову в темнице.
MATT|14|11|И принесли голову его на блюде и дали девице, а она отнесла матери своей.
MATT|14|12|Ученики же его, придя, взяли тело его и погребли его; и пошли, возвестили Иисусу.
MATT|14|13|И, услышав, Иисус удалился оттуда на лодке в пустынное место один; а народ, услышав о том, пошел за Ним из городов пешком.
MATT|14|14|И, выйдя, Иисус увидел множество людей и сжалился над ними, и исцелил больных их.
MATT|14|15|Когда же настал вечер, приступили к Нему ученики Его и сказали: место здесь пустынное и время уже позднее; отпусти народ, чтобы они пошли в селения и купили себе пищи.
MATT|14|16|Но Иисус сказал им: не нужно им идти, вы дайте им есть.
MATT|14|17|Они же говорят Ему: у нас здесь только пять хлебов и две рыбы.
MATT|14|18|Он сказал: принесите их Мне сюда.
MATT|14|19|И велел народу возлечь на траву и, взяв пять хлебов и две рыбы, воззрел на небо, благословил и, преломив, дал хлебы ученикам, а ученики народу.
MATT|14|20|И ели все и насытились; и набрали оставшихся кусков двенадцать коробов полных;
MATT|14|21|а евших было около пяти тысяч человек, кроме женщин и детей.
MATT|14|22|И тотчас понудил Иисус учеников Своих войти в лодку и отправиться прежде Его на другую сторону, пока Он отпустит народ.
MATT|14|23|И, отпустив народ, Он взошел на гору помолиться наедине; и вечером оставался там один.
MATT|14|24|А лодка была уже на средине моря, и ее било волнами, потому что ветер был противный.
MATT|14|25|В четвертую же стражу ночи пошел к ним Иисус, идя по морю.
MATT|14|26|И ученики, увидев Его идущего по морю, встревожились и говорили: это призрак; и от страха вскричали.
MATT|14|27|Но Иисус тотчас заговорил с ними и сказал: ободритесь; это Я, не бойтесь.
MATT|14|28|Петр сказал Ему в ответ: Господи! если это Ты, повели мне придти к Тебе по воде.
MATT|14|29|Он же сказал: иди. И, выйдя из лодки, Петр пошел по воде, чтобы подойти к Иисусу,
MATT|14|30|но, видя сильный ветер, испугался и, начав утопать, закричал: Господи! спаси меня.
MATT|14|31|Иисус тотчас простер руку, поддержал его и говорит ему: маловерный! зачем ты усомнился?
MATT|14|32|И, когда вошли они в лодку, ветер утих.
MATT|14|33|Бывшие же в лодке подошли, поклонились Ему и сказали: истинно Ты Сын Божий.
MATT|14|34|И, переправившись, прибыли в землю Геннисаретскую.
MATT|14|35|Жители того места, узнав Его, послали во всю окрестность ту и принесли к Нему всех больных,
MATT|14|36|и просили Его, чтобы только прикоснуться к краю одежды Его; и которые прикасались, исцелялись.
MATT|15|1|Тогда приходят к Иисусу Иерусалимские книжники и фарисеи и говорят:
MATT|15|2|зачем ученики Твои преступают предание старцев? ибо не умывают рук своих, когда едят хлеб.
MATT|15|3|Он же сказал им в ответ: зачем и вы преступаете заповедь Божию ради предания вашего?
MATT|15|4|Ибо Бог заповедал: почитай отца и мать; и: злословящий отца или мать смертью да умрет.
MATT|15|5|А вы говорите: если кто скажет отцу или матери: дар [Богу] то, чем бы ты от меня пользовался,
MATT|15|6|тот может и не почтить отца своего или мать свою; таким образом вы устранили заповедь Божию преданием вашим.
MATT|15|7|Лицемеры! хорошо пророчествовал о вас Исаия, говоря:
MATT|15|8|приближаются ко Мне люди сии устами своими, и чтут Меня языком, сердце же их далеко отстоит от Меня;
MATT|15|9|но тщетно чтут Меня, уча учениям, заповедям человеческим.
MATT|15|10|И, призвав народ, сказал им: слушайте и разумейте!
MATT|15|11|не то, что входит в уста, оскверняет человека, но то, что выходит из уст, оскверняет человека.
MATT|15|12|Тогда ученики Его, приступив, сказали Ему: знаешь ли, что фарисеи, услышав слово сие, соблазнились?
MATT|15|13|Он же сказал в ответ: всякое растение, которое не Отец Мой Небесный насадил, искоренится;
MATT|15|14|оставьте их: они – слепые вожди слепых; а если слепой ведет слепого, то оба упадут в яму.
MATT|15|15|Петр же, отвечая, сказал Ему: изъясни нам притчу сию.
MATT|15|16|Иисус сказал: неужели и вы еще не разумеете?
MATT|15|17|еще ли не понимаете, что все, входящее в уста, проходит в чрево и извергается вон?
MATT|15|18|а исходящее из уст – из сердца исходит – сие оскверняет человека,
MATT|15|19|ибо из сердца исходят злые помыслы, убийства, прелюбодеяния, любодеяния, кражи, лжесвидетельства, хуления –
MATT|15|20|это оскверняет человека; а есть неумытыми руками – не оскверняет человека.
MATT|15|21|И, выйдя оттуда, Иисус удалился в страны Тирские и Сидонские.
MATT|15|22|И вот, женщина Хананеянка, выйдя из тех мест, кричала Ему: помилуй меня, Господи, сын Давидов, дочь моя жестоко беснуется.
MATT|15|23|Но Он не отвечал ей ни слова. И ученики Его, приступив, просили Его: отпусти ее, потому что кричит за нами.
MATT|15|24|Он же сказал в ответ: Я послан только к погибшим овцам дома Израилева.
MATT|15|25|А она, подойдя, кланялась Ему и говорила: Господи! помоги мне.
MATT|15|26|Он же сказал в ответ: нехорошо взять хлеб у детей и бросить псам.
MATT|15|27|Она сказала: так, Господи! но и псы едят крохи, которые падают со стола господ их.
MATT|15|28|Тогда Иисус сказал ей в ответ: о, женщина! велика вера твоя; да будет тебе по желанию твоему. И исцелилась дочь ее в тот час.
MATT|15|29|Перейдя оттуда, пришел Иисус к морю Галилейскому и, взойдя на гору, сел там.
MATT|15|30|И приступило к Нему множество народа, имея с собою хромых, слепых, немых, увечных и иных многих, и повергли их к ногам Иисусовым; и Он исцелил их;
MATT|15|31|так что народ дивился, видя немых говорящими, увечных здоровыми, хромых ходящими и слепых видящими; и прославлял Бога Израилева.
MATT|15|32|Иисус же, призвав учеников Своих, сказал им: жаль Мне народа, что уже три дня находятся при Мне, и нечего им есть; отпустить же их неевшими не хочу, чтобы не ослабели в дороге.
MATT|15|33|И говорят Ему ученики Его: откуда нам взять в пустыне столько хлебов, чтобы накормить столько народа?
MATT|15|34|Говорит им Иисус: сколько у вас хлебов? Они же сказали: семь, и немного рыбок.
MATT|15|35|Тогда велел народу возлечь на землю.
MATT|15|36|И, взяв семь хлебов и рыбы, воздал благодарение, преломил и дал ученикам Своим, а ученики народу.
MATT|15|37|И ели все и насытились; и набрали оставшихся кусков семь корзин полных,
MATT|15|38|а евших было четыре тысячи человек, кроме женщин и детей.
MATT|15|39|И, отпустив народ, Он вошел в лодку и прибыл в пределы Магдалинские.
MATT|16|1|И приступили фарисеи и саддукеи и, искушая Его, просили показать им знамение с неба.
MATT|16|2|Он же сказал им в ответ: вечером вы говорите: будет ведро, потому что небо красно;
MATT|16|3|и поутру: сегодня ненастье, потому что небо багрово. Лицемеры! различать лице неба вы умеете, а знамений времен не можете.
MATT|16|4|Род лукавый и прелюбодейный знамения ищет, и знамение не дастся ему, кроме знамения Ионы пророка. И, оставив их, отошел.
MATT|16|5|Переправившись на другую сторону, ученики Его забыли взять хлебов.
MATT|16|6|Иисус сказал им: смотрите, берегитесь закваски фарисейской и саддукейской.
MATT|16|7|Они же помышляли в себе и говорили: [это значит], что хлебов мы не взяли.
MATT|16|8|Уразумев то, Иисус сказал им: что помышляете в себе, маловерные, что хлебов не взяли?
MATT|16|9|Еще ли не понимаете и не помните о пяти хлебах на пять тысяч [человек], и сколько коробов вы набрали?
MATT|16|10|ни о семи хлебах на четыре тысячи, и сколько корзин вы набрали?
MATT|16|11|как не разумеете, что не о хлебе сказал Я вам: берегитесь закваски фарисейской и саддукейской?
MATT|16|12|Тогда они поняли, что Он говорил им беречься не закваски хлебной, но учения фарисейского и саддукейского.
MATT|16|13|Придя же в страны Кесарии Филипповой, Иисус спрашивал учеников Своих: за кого люди почитают Меня, Сына Человеческого?
MATT|16|14|Они сказали: одни за Иоанна Крестителя, другие за Илию, а иные за Иеремию, или за одного из пророков.
MATT|16|15|Он говорит им: а вы за кого почитаете Меня?
MATT|16|16|Симон же Петр, отвечая, сказал: Ты – Христос, Сын Бога Живаго.
MATT|16|17|Тогда Иисус сказал ему в ответ: блажен ты, Симон, сын Ионин, потому что не плоть и кровь открыли тебе это, но Отец Мой, Сущий на небесах;
MATT|16|18|и Я говорю тебе: ты – Петр, и на сем камне Я создам Церковь Мою, и врата ада не одолеют ее;
MATT|16|19|и дам тебе ключи Царства Небесного: и что свяжешь на земле, то будет связано на небесах, и что разрешишь на земле, то будет разрешено на небесах.
MATT|16|20|Тогда Иисус запретил ученикам Своим, чтобы никому не сказывали, что Он есть Иисус Христос.
MATT|16|21|С того времени Иисус начал открывать ученикам Своим, что Ему должно идти в Иерусалим и много пострадать от старейшин и первосвященников и книжников, и быть убиту, и в третий день воскреснуть.
MATT|16|22|И, отозвав Его, Петр начал прекословить Ему: будь милостив к Себе, Господи! да не будет этого с Тобою!
MATT|16|23|Он же, обратившись, сказал Петру: отойди от Меня, сатана! ты Мне соблазн! потому что думаешь не о том, что Божие, но что человеческое.
MATT|16|24|Тогда Иисус сказал ученикам Своим: если кто хочет идти за Мною, отвергнись себя, и возьми крест свой, и следуй за Мною,
MATT|16|25|ибо кто хочет душу свою сберечь, тот потеряет ее, а кто потеряет душу свою ради Меня, тот обретет ее;
MATT|16|26|какая польза человеку, если он приобретет весь мир, а душе своей повредит? или какой выкуп даст человек за душу свою?
MATT|16|27|ибо приидет Сын Человеческий во славе Отца Своего с Ангелами Своими и тогда воздаст каждому по делам его.
MATT|16|28|Истинно говорю вам: есть некоторые из стоящих здесь, которые не вкусят смерти, как уже увидят Сына Человеческого, грядущего в Царствии Своем.
MATT|17|1|По прошествии дней шести, взял Иисус Петра, Иакова и Иоанна, брата его, и возвел их на гору высокую одних,
MATT|17|2|и преобразился пред ними: и просияло лице Его, как солнце, одежды же Его сделались белыми, как свет.
MATT|17|3|И вот, явились им Моисей и Илия, с Ним беседующие.
MATT|17|4|При сем Петр сказал Иисусу: Господи! хорошо нам здесь быть; если хочешь, сделаем здесь три кущи: Тебе одну, и Моисею одну, и одну Илии.
MATT|17|5|Когда он еще говорил, се, облако светлое осенило их; и се, глас из облака глаголющий: Сей есть Сын Мой Возлюбленный, в Котором Мое благоволение; Его слушайте.
MATT|17|6|И, услышав, ученики пали на лица свои и очень испугались.
MATT|17|7|Но Иисус, приступив, коснулся их и сказал: встаньте и не бойтесь.
MATT|17|8|Возведя же очи свои, они никого не увидели, кроме одного Иисуса.
MATT|17|9|И когда сходили они с горы, Иисус запретил им, говоря: никому не сказывайте о сем видении, доколе Сын Человеческий не воскреснет из мертвых.
MATT|17|10|И спросили Его ученики Его: как же книжники говорят, что Илии надлежит придти прежде?
MATT|17|11|Иисус сказал им в ответ: правда, Илия должен придти прежде и устроить все;
MATT|17|12|но говорю вам, что Илия уже пришел, и не узнали его, а поступили с ним, как хотели; так и Сын Человеческий пострадает от них.
MATT|17|13|Тогда ученики поняли, что Он говорил им об Иоанне Крестителе.
MATT|17|14|Когда они пришли к народу, то подошел к Нему человек и, преклоняя пред Ним колени,
MATT|17|15|сказал: Господи! помилуй сына моего; он в новолуния [беснуется] и тяжко страдает, ибо часто бросается в огонь и часто в воду,
MATT|17|16|я приводил его к ученикам Твоим, и они не могли исцелить его.
MATT|17|17|Иисус же, отвечая, сказал: о, род неверный и развращенный! доколе буду с вами? доколе буду терпеть вас? приведите его ко Мне сюда.
MATT|17|18|И запретил ему Иисус, и бес вышел из него; и отрок исцелился в тот час.
MATT|17|19|Тогда ученики, приступив к Иисусу наедине, сказали: почему мы не могли изгнать его?
MATT|17|20|Иисус же сказал им: по неверию вашему; ибо истинно говорю вам: если вы будете иметь веру с горчичное зерно и скажете горе сей: "перейди отсюда туда", и она перейдет; и ничего не будет невозможного для вас;
MATT|17|21|сей же род изгоняется только молитвою и постом.
MATT|17|22|Во время пребывания их в Галилее, Иисус сказал им: Сын Человеческий предан будет в руки человеческие,
MATT|17|23|и убьют Его, и в третий день воскреснет. И они весьма опечалились.
MATT|17|24|Когда же пришли они в Капернаум, то подошли к Петру собиратели дидрахм и сказали: Учитель ваш не даст ли дидрахмы?
MATT|17|25|Он говорит: да. И когда вошел он в дом, то Иисус, предупредив его, сказал: как тебе кажется, Симон? цари земные с кого берут пошлины или подати? с сынов ли своих, или с посторонних?
MATT|17|26|Петр говорит Ему: с посторонних. Иисус сказал ему: итак сыны свободны;
MATT|17|27|но, чтобы нам не соблазнить их, пойди на море, брось уду, и первую рыбу, которая попадется, возьми, и, открыв у ней рот, найдешь статир; возьми его и отдай им за Меня и за себя.
MATT|18|1|В то время ученики приступили к Иисусу и сказали: кто больше в Царстве Небесном?
MATT|18|2|Иисус, призвав дитя, поставил его посреди них
MATT|18|3|и сказал: истинно говорю вам, если не обратитесь и не будете как дети, не войдете в Царство Небесное;
MATT|18|4|итак, кто умалится, как это дитя, тот и больше в Царстве Небесном;
MATT|18|5|и кто примет одно такое дитя во имя Мое, тот Меня принимает;
MATT|18|6|а кто соблазнит одного из малых сих, верующих в Меня, тому лучше было бы, если бы повесили ему мельничный жернов на шею и потопили его во глубине морской.
MATT|18|7|Горе миру от соблазнов, ибо надобно придти соблазнам; но горе тому человеку, через которого соблазн приходит.
MATT|18|8|Если же рука твоя или нога твоя соблазняет тебя, отсеки их и брось от себя: лучше тебе войти в жизнь без руки или без ноги, нежели с двумя руками и с двумя ногами быть ввержену в огонь вечный;
MATT|18|9|и если глаз твой соблазняет тебя, вырви его и брось от себя: лучше тебе с одним глазом войти в жизнь, нежели с двумя глазами быть ввержену в геенну огненную.
MATT|18|10|Смотрите, не презирайте ни одного из малых сих; ибо говорю вам, что Ангелы их на небесах всегда видят лице Отца Моего Небесного.
MATT|18|11|Ибо Сын Человеческий пришел взыскать и спасти погибшее.
MATT|18|12|Как вам кажется? Если бы у кого было сто овец, и одна из них заблудилась, то не оставит ли он девяносто девять в горах и не пойдет ли искать заблудившуюся?
MATT|18|13|и если случится найти ее, то, истинно говорю вам, он радуется о ней более, нежели о девяноста девяти незаблудившихся.
MATT|18|14|Так, нет воли Отца вашего Небесного, чтобы погиб один из малых сих.
MATT|18|15|Если же согрешит против тебя брат твой, пойди и обличи его между тобою и им одним; если послушает тебя, то приобрел ты брата твоего;
MATT|18|16|если же не послушает, возьми с собою еще одного или двух, дабы устами двух или трех свидетелей подтвердилось всякое слово;
MATT|18|17|если же не послушает их, скажи церкви; а если и церкви не послушает, то да будет он тебе, как язычник и мытарь.
MATT|18|18|Истинно говорю вам: что вы свяжете на земле, то будет связано на небе; и что разрешите на земле, то будет разрешено на небе.
MATT|18|19|Истинно также говорю вам, что если двое из вас согласятся на земле просить о всяком деле, то, чего бы ни попросили, будет им от Отца Моего Небесного,
MATT|18|20|ибо, где двое или трое собраны во имя Мое, там Я посреди них.
MATT|18|21|Тогда Петр приступил к Нему и сказал: Господи! сколько раз прощать брату моему, согрешающему против меня? до семи ли раз?
MATT|18|22|Иисус говорит ему: не говорю тебе: до семи раз, но до седмижды семидесяти раз.
MATT|18|23|Посему Царство Небесное подобно царю, который захотел сосчитаться с рабами своими;
MATT|18|24|когда начал он считаться, приведен был к нему некто, который должен был ему десять тысяч талантов;
MATT|18|25|а как он не имел, чем заплатить, то государь его приказал продать его, и жену его, и детей, и все, что он имел, и заплатить;
MATT|18|26|тогда раб тот пал, и, кланяясь ему, говорил: государь! потерпи на мне, и все тебе заплачу.
MATT|18|27|Государь, умилосердившись над рабом тем, отпустил его и долг простил ему.
MATT|18|28|Раб же тот, выйдя, нашел одного из товарищей своих, который должен был ему сто динариев, и, схватив его, душил, говоря: отдай мне, что должен.
MATT|18|29|Тогда товарищ его пал к ногам его, умолял его и говорил: потерпи на мне, и все отдам тебе.
MATT|18|30|Но тот не захотел, а пошел и посадил его в темницу, пока не отдаст долга.
MATT|18|31|Товарищи его, видев происшедшее, очень огорчились и, придя, рассказали государю своему все бывшее.
MATT|18|32|Тогда государь его призывает его и говорит: злой раб! весь долг тот я простил тебе, потому что ты упросил меня;
MATT|18|33|не надлежало ли и тебе помиловать товарища твоего, как и я помиловал тебя?
MATT|18|34|И, разгневавшись, государь его отдал его истязателям, пока не отдаст ему всего долга.
MATT|18|35|Так и Отец Мой Небесный поступит с вами, если не простит каждый из вас от сердца своего брату своему согрешений его.
MATT|19|1|Когда Иисус окончил слова сии, то вышел из Галилеи и пришел в пределы Иудейские, за Иорданскою стороною.
MATT|19|2|За Ним последовало много людей, и Он исцелил их там.
MATT|19|3|И приступили к Нему фарисеи и, искушая Его, говорили Ему: по всякой ли причине позволительно человеку разводиться с женою своею?
MATT|19|4|Он сказал им в ответ: не читали ли вы, что Сотворивший вначале мужчину и женщину сотворил их?
MATT|19|5|И сказал: посему оставит человек отца и мать и прилепится к жене своей, и будут два одною плотью,
MATT|19|6|так что они уже не двое, но одна плоть. Итак, что Бог сочетал, того человек да не разлучает.
MATT|19|7|Они говорят Ему: как же Моисей заповедал давать разводное письмо и разводиться с нею?
MATT|19|8|Он говорит им: Моисей по жестокосердию вашему позволил вам разводиться с женами вашими, а сначала не было так;
MATT|19|9|но Я говорю вам: кто разведется с женою своею не за прелюбодеяние и женится на другой, [тот] прелюбодействует; и женившийся на разведенной прелюбодействует.
MATT|19|10|Говорят Ему ученики Его: если такова обязанность человека к жене, то лучше не жениться.
MATT|19|11|Он же сказал им: не все вмещают слово сие, но кому дано,
MATT|19|12|ибо есть скопцы, которые из чрева матернего родились так; и есть скопцы, которые оскоплены от людей; и есть скопцы, которые сделали сами себя скопцами для Царства Небесного. Кто может вместить, да вместит.
MATT|19|13|Тогда приведены были к Нему дети, чтобы Он возложил на них руки и помолился; ученики же возбраняли им.
MATT|19|14|Но Иисус сказал: пустите детей и не препятствуйте им приходить ко Мне, ибо таковых есть Царство Небесное.
MATT|19|15|И, возложив на них руки, пошел оттуда.
MATT|19|16|И вот, некто, подойдя, сказал Ему: Учитель благий! что сделать мне доброго, чтобы иметь жизнь вечную?
MATT|19|17|Он же сказал ему: что ты называешь Меня благим? Никто не благ, как только один Бог. Если же хочешь войти в жизнь [вечную], соблюди заповеди.
MATT|19|18|Говорит Ему: какие? Иисус же сказал: не убивай; не прелюбодействуй; не кради; не лжесвидетельствуй;
MATT|19|19|почитай отца и мать; и: люби ближнего твоего, как самого себя.
MATT|19|20|Юноша говорит Ему: все это сохранил я от юности моей; чего еще недостает мне?
MATT|19|21|Иисус сказал ему: если хочешь быть совершенным, пойди, продай имение твое и раздай нищим; и будешь иметь сокровище на небесах; и приходи и следуй за Мною.
MATT|19|22|Услышав слово сие, юноша отошел с печалью, потому что у него было большое имение.
MATT|19|23|Иисус же сказал ученикам Своим: истинно говорю вам, что трудно богатому войти в Царство Небесное;
MATT|19|24|и еще говорю вам: удобнее верблюду пройти сквозь игольные уши, нежели богатому войти в Царство Божие.
MATT|19|25|Услышав это, ученики Его весьма изумились и сказали: так кто же может спастись?
MATT|19|26|А Иисус, воззрев, сказал им: человекам это невозможно, Богу же все возможно.
MATT|19|27|Тогда Петр, отвечая, сказал Ему: вот, мы оставили все и последовали за Тобою; что же будет нам?
MATT|19|28|Иисус же сказал им: истинно говорю вам, что вы, последовавшие за Мною, – в пакибытии, когда сядет Сын Человеческий на престоле славы Своей, сядете и вы на двенадцати престолах судить двенадцать колен Израилевых.
MATT|19|29|И всякий, кто оставит домы, или братьев, или сестер, или отца, или мать, или жену, или детей, или земли, ради имени Моего, получит во сто крат и наследует жизнь вечную.
MATT|19|30|Многие же будут первые последними, и последние первыми.
MATT|20|1|Ибо Царство Небесное подобно хозяину дома, который вышел рано поутру нанять работников в виноградник свой
MATT|20|2|и, договорившись с работниками по динарию на день, послал их в виноградник свой;
MATT|20|3|выйдя около третьего часа, он увидел других, стоящих на торжище праздно,
MATT|20|4|и им сказал: идите и вы в виноградник мой, и что следовать будет, дам вам. Они пошли.
MATT|20|5|Опять выйдя около шестого и девятого часа, сделал то же.
MATT|20|6|Наконец, выйдя около одиннадцатого часа, он нашел других, стоящих праздно, и говорит им: что вы стоите здесь целый день праздно?
MATT|20|7|Они говорят ему: никто нас не нанял. Он говорит им: идите и вы в виноградник мой, и что следовать будет, получите.
MATT|20|8|Когда же наступил вечер, говорит господин виноградника управителю своему: позови работников и отдай им плату, начав с последних до первых.
MATT|20|9|И пришедшие около одиннадцатого часа получили по динарию.
MATT|20|10|Пришедшие же первыми думали, что они получат больше, но получили и они по динарию;
MATT|20|11|и, получив, стали роптать на хозяина дома
MATT|20|12|и говорили: эти последние работали один час, и ты сравнял их с нами, перенесшими тягость дня и зной.
MATT|20|13|Он же в ответ сказал одному из них: друг! я не обижаю тебя; не за динарий ли ты договорился со мною?
MATT|20|14|возьми свое и пойди; я же хочу дать этому последнему [то же], что и тебе;
MATT|20|15|разве я не властен в своем делать, что хочу? или глаз твой завистлив от того, что я добр?
MATT|20|16|Так будут последние первыми, и первые последними, ибо много званых, а мало избранных.
MATT|20|17|И, восходя в Иерусалим, Иисус дорогою отозвал двенадцать учеников одних, и сказал им:
MATT|20|18|вот, мы восходим в Иерусалим, и Сын Человеческий предан будет первосвященникам и книжникам, и осудят Его на смерть;
MATT|20|19|и предадут Его язычникам на поругание и биение и распятие; и в третий день воскреснет.
MATT|20|20|Тогда приступила к Нему мать сыновей Зеведеевых с сыновьями своими, кланяясь и чего–то прося у Него.
MATT|20|21|Он сказал ей: чего ты хочешь? Она говорит Ему: скажи, чтобы сии два сына мои сели у Тебя один по правую сторону, а другой по левую в Царстве Твоем.
MATT|20|22|Иисус сказал в ответ: не знаете, чего просите. Можете ли пить чашу, которую Я буду пить, или креститься крещением, которым Я крещусь? Они говорят Ему: можем.
MATT|20|23|И говорит им: чашу Мою будете пить, и крещением, которым Я крещусь, будете креститься, но дать сесть у Меня по правую сторону и по левую – не от Меня [зависит], но кому уготовано Отцем Моим.
MATT|20|24|Услышав [сие, прочие] десять [учеников] вознегодовали на двух братьев.
MATT|20|25|Иисус же, подозвав их, сказал: вы знаете, что князья народов господствуют над ними, и вельможи властвуют ими;
MATT|20|26|но между вами да не будет так: а кто хочет между вами быть большим, да будет вам слугою;
MATT|20|27|и кто хочет между вами быть первым, да будет вам рабом;
MATT|20|28|так как Сын Человеческий не [для того] пришел, чтобы Ему служили, но чтобы послужить и отдать душу Свою для искупления многих.
MATT|20|29|И когда выходили они из Иерихона, за Ним следовало множество народа.
MATT|20|30|И вот, двое слепых, сидевшие у дороги, услышав, что Иисус идет мимо, начали кричать: помилуй нас, Господи, Сын Давидов!
MATT|20|31|Народ же заставлял их молчать; но они еще громче стали кричать: помилуй нас, Господи, Сын Давидов!
MATT|20|32|Иисус, остановившись, подозвал их и сказал: чего вы хотите от Меня?
MATT|20|33|Они говорят Ему: Господи! чтобы открылись глаза наши.
MATT|20|34|Иисус же, умилосердившись, прикоснулся к глазам их; и тотчас прозрели глаза их, и они пошли за Ним.
MATT|21|1|И когда приблизились к Иерусалиму и пришли в Виффагию к горе Елеонской, тогда Иисус послал двух учеников,
MATT|21|2|сказав им: пойдите в селение, которое прямо перед вами; и тотчас найдете ослицу привязанную и молодого осла с нею; отвязав, приведите ко Мне;
MATT|21|3|и если кто скажет вам что–нибудь, отвечайте, что они надобны Господу; и тотчас пошлет их.
MATT|21|4|Все же сие было, да сбудется реченное через пророка, который говорит:
MATT|21|5|Скажите дщери Сионовой: се, Царь твой грядет к тебе кроткий, сидя на ослице и молодом осле, сыне подъяремной.
MATT|21|6|Ученики пошли и поступили так, как повелел им Иисус:
MATT|21|7|привели ослицу и молодого осла и положили на них одежды свои, и Он сел поверх их.
MATT|21|8|Множество же народа постилали свои одежды по дороге, а другие резали ветви с дерев и постилали по дороге;
MATT|21|9|народ же, предшествовавший и сопровождавший, восклицал: осанна Сыну Давидову! благословен Грядущий во имя Господне! осанна в вышних!
MATT|21|10|И когда вошел Он в Иерусалим, весь город пришел в движение и говорил: кто Сей?
MATT|21|11|Народ же говорил: Сей есть Иисус, Пророк из Назарета Галилейского.
MATT|21|12|И вошел Иисус в храм Божий и выгнал всех продающих и покупающих в храме, и опрокинул столы меновщиков и скамьи продающих голубей,
MATT|21|13|и говорил им: написано, – дом Мой домом молитвы наречется; а вы сделали его вертепом разбойников.
MATT|21|14|И приступили к Нему в храме слепые и хромые, и Он исцелил их.
MATT|21|15|Видев же первосвященники и книжники чудеса, которые Он сотворил, и детей, восклицающих в храме и говорящих: осанна Сыну Давидову! – вознегодовали
MATT|21|16|и сказали Ему: слышишь ли, что они говорят? Иисус же говорит им: да! разве вы никогда не читали: из уст младенцев и грудных детей Ты устроил хвалу?
MATT|21|17|И, оставив их, вышел вон из города в Вифанию и провел там ночь.
MATT|21|18|Поутру же, возвращаясь в город, взалкал;
MATT|21|19|и увидев при дороге одну смоковницу, подошел к ней и, ничего не найдя на ней, кроме одних листьев, говорит ей: да не будет же впредь от тебя плода вовек. И смоковница тотчас засохла.
MATT|21|20|Увидев это, ученики удивились и говорили: как это тотчас засохла смоковница?
MATT|21|21|Иисус же сказал им в ответ: истинно говорю вам, если будете иметь веру и не усомнитесь, не только сделаете то, что [сделано] со смоковницею, но если и горе сей скажете: поднимись и ввергнись в море, – будет;
MATT|21|22|и все, чего ни попросите в молитве с верою, получите.
MATT|21|23|И когда пришел Он в храм и учил, приступили к Нему первосвященники и старейшины народа и сказали: какой властью Ты это делаешь? и кто Тебе дал такую власть?
MATT|21|24|Иисус сказал им в ответ: спрошу и Я вас об одном; если о том скажете Мне, то и Я вам скажу, какою властью это делаю;
MATT|21|25|крещение Иоанново откуда было: с небес, или от человеков? Они же рассуждали между собою: если скажем: с небес, то Он скажет нам: почему же вы не поверили ему?
MATT|21|26|а если сказать: от человеков, – боимся народа, ибо все почитают Иоанна за пророка.
MATT|21|27|И сказали в ответ Иисусу: не знаем. Сказал им и Он: и Я вам не скажу, какою властью это делаю.
MATT|21|28|А как вам кажется? У одного человека было два сына; и он, подойдя к первому, сказал: сын! пойди сегодня работай в винограднике моем.
MATT|21|29|Но он сказал в ответ: не хочу; а после, раскаявшись, пошел.
MATT|21|30|И подойдя к другому, он сказал то же. Этот сказал в ответ: иду, государь, и не пошел.
MATT|21|31|Который из двух исполнил волю отца? Говорят Ему: первый. Иисус говорит им: истинно говорю вам, что мытари и блудницы вперед вас идут в Царство Божие,
MATT|21|32|ибо пришел к вам Иоанн путем праведности, и вы не поверили ему, а мытари и блудницы поверили ему; вы же, и видев это, не раскаялись после, чтобы поверить ему.
MATT|21|33|Выслушайте другую притчу: был некоторый хозяин дома, который насадил виноградник, обнес его оградою, выкопал в нем точило, построил башню и, отдав его виноградарям, отлучился.
MATT|21|34|Когда же приблизилось время плодов, он послал своих слуг к виноградарям взять свои плоды;
MATT|21|35|виноградари, схватив слуг его, иного прибили, иного убили, а иного побили камнями.
MATT|21|36|Опять послал он других слуг, больше прежнего; и с ними поступили так же.
MATT|21|37|Наконец, послал он к ним своего сына, говоря: постыдятся сына моего.
MATT|21|38|Но виноградари, увидев сына, сказали друг другу: это наследник; пойдем, убьем его и завладеем наследством его.
MATT|21|39|И, схватив его, вывели вон из виноградника и убили.
MATT|21|40|Итак, когда придет хозяин виноградника, что сделает он с этими виноградарями?
MATT|21|41|Говорят Ему: злодеев сих предаст злой смерти, а виноградник отдаст другим виноградарям, которые будут отдавать ему плоды во времена свои.
MATT|21|42|Иисус говорит им: неужели вы никогда не читали в Писании: камень, который отвергли строители, тот самый сделался главою угла? Это от Господа, и есть дивно в очах наших?
MATT|21|43|Потому сказываю вам, что отнимется от вас Царство Божие и дано будет народу, приносящему плоды его;
MATT|21|44|и тот, кто упадет на этот камень, разобьется, а на кого он упадет, того раздавит.
MATT|21|45|И слышав притчи Его, первосвященники и фарисеи поняли, что Он о них говорит,
MATT|21|46|и старались схватить Его, но побоялись народа, потому что Его почитали за Пророка.
MATT|22|1|Иисус, продолжая говорить им притчами, сказал:
MATT|22|2|Царство Небесное подобно человеку царю, который сделал брачный пир для сына своего
MATT|22|3|и послал рабов своих звать званых на брачный пир; и не хотели придти.
MATT|22|4|Опять послал других рабов, сказав: скажите званым: вот, я приготовил обед мой, тельцы мои и что откормлено, заколото, и все готово; приходите на брачный пир.
MATT|22|5|Но они, пренебрегши то, пошли, кто на поле свое, а кто на торговлю свою;
MATT|22|6|прочие же, схватив рабов его, оскорбили и убили [их].
MATT|22|7|Услышав о сем, царь разгневался, и, послав войска свои, истребил убийц оных и сжег город их.
MATT|22|8|Тогда говорит он рабам своим: брачный пир готов, а званые не были достойны;
MATT|22|9|итак пойдите на распутия и всех, кого найдете, зовите на брачный пир.
MATT|22|10|И рабы те, выйдя на дороги, собрали всех, кого только нашли, и злых и добрых; и брачный пир наполнился возлежащими.
MATT|22|11|Царь, войдя посмотреть возлежащих, увидел там человека, одетого не в брачную одежду,
MATT|22|12|и говорит ему: друг! как ты вошел сюда не в брачной одежде? Он же молчал.
MATT|22|13|Тогда сказал царь слугам: связав ему руки и ноги, возьмите его и бросьте во тьму внешнюю; там будет плач и скрежет зубов;
MATT|22|14|ибо много званых, а мало избранных.
MATT|22|15|Тогда фарисеи пошли и совещались, как бы уловить Его в словах.
MATT|22|16|И посылают к Нему учеников своих с иродианами, говоря: Учитель! мы знаем, что Ты справедлив, и истинно пути Божию учишь, и не заботишься об угождении кому–либо, ибо не смотришь ни на какое лице;
MATT|22|17|итак скажи нам: как Тебе кажется? позволительно ли давать подать кесарю, или нет?
MATT|22|18|Но Иисус, видя лукавство их, сказал: что искушаете Меня, лицемеры?
MATT|22|19|покажите Мне монету, которою платится подать. Они принесли Ему динарий.
MATT|22|20|И говорит им: чье это изображение и надпись?
MATT|22|21|Говорят Ему: кесаревы. Тогда говорит им: итак отдавайте кесарево кесарю, а Божие Богу.
MATT|22|22|Услышав это, они удивились и, оставив Его, ушли.
MATT|22|23|В тот день приступили к Нему саддукеи, которые говорят, что нет воскресения, и спросили Его:
MATT|22|24|Учитель! Моисей сказал: если кто умрет, не имея детей, то брат его пусть возьмет за себя жену его и восстановит семя брату своему;
MATT|22|25|было у нас семь братьев; первый, женившись, умер и, не имея детей, оставил жену свою брату своему;
MATT|22|26|подобно и второй, и третий, даже до седьмого;
MATT|22|27|после же всех умерла и жена;
MATT|22|28|итак, в воскресении, которого из семи будет она женою? ибо все имели ее.
MATT|22|29|Иисус сказал им в ответ: заблуждаетесь, не зная Писаний, ни силы Божией,
MATT|22|30|ибо в воскресении ни женятся, ни выходят замуж, но пребывают, как Ангелы Божии на небесах.
MATT|22|31|А о воскресении мертвых не читали ли вы реченного вам Богом:
MATT|22|32|Я Бог Авраама, и Бог Исаака, и Бог Иакова? Бог не есть Бог мертвых, но живых.
MATT|22|33|И, слыша, народ дивился учению Его.
MATT|22|34|А фарисеи, услышав, что Он привел саддукеев в молчание, собрались вместе.
MATT|22|35|И один из них, законник, искушая Его, спросил, говоря:
MATT|22|36|Учитель! какая наибольшая заповедь в законе?
MATT|22|37|Иисус сказал ему: возлюби Господа Бога твоего всем сердцем твоим и всею душею твоею и всем разумением твоим:
MATT|22|38|сия есть первая и наибольшая заповедь;
MATT|22|39|вторая же подобная ей: возлюби ближнего твоего, как самого себя;
MATT|22|40|на сих двух заповедях утверждается весь закон и пророки.
MATT|22|41|Когда же собрались фарисеи, Иисус спросил их:
MATT|22|42|что вы думаете о Христе? чей Он сын? Говорят Ему: Давидов.
MATT|22|43|Говорит им: как же Давид, по вдохновению, называет Его Господом, когда говорит:
MATT|22|44|сказал Господь Господу моему: седи одесную Меня, доколе положу врагов Твоих в подножие ног Твоих?
MATT|22|45|Итак, если Давид называет Его Господом, как же Он сын ему?
MATT|22|46|И никто не мог отвечать Ему ни слова; и с того дня никто уже не смел спрашивать Его.
MATT|23|1|Тогда Иисус начал говорить народу и ученикам Своим
MATT|23|2|и сказал: на Моисеевом седалище сели книжники и фарисеи;
MATT|23|3|итак все, что они велят вам соблюдать, соблюдайте и делайте; по делам же их не поступайте, ибо они говорят, и не делают:
MATT|23|4|связывают бремена тяжелые и неудобоносимые и возлагают на плечи людям, а сами не хотят и перстом двинуть их;
MATT|23|5|все же дела свои делают с тем, чтобы видели их люди: расширяют хранилища свои и увеличивают воскрилия одежд своих;
MATT|23|6|также любят предвозлежания на пиршествах и председания в синагогах
MATT|23|7|и приветствия в народных собраниях, и чтобы люди звали их: учитель! учитель!
MATT|23|8|А вы не называйтесь учителями, ибо один у вас Учитель – Христос, все же вы – братья;
MATT|23|9|и отцом себе не называйте никого на земле, ибо один у вас Отец, Который на небесах;
MATT|23|10|и не называйтесь наставниками, ибо один у вас Наставник – Христос.
MATT|23|11|Больший из вас да будет вам слуга:
MATT|23|12|ибо, кто возвышает себя, тот унижен будет, а кто унижает себя, тот возвысится.
MATT|23|13|Горе вам, книжники и фарисеи, лицемеры, что затворяете Царство Небесное человекам, ибо сами не входите и хотящих войти не допускаете.
MATT|23|14|Горе вам, книжники и фарисеи, лицемеры, что поедаете домы вдов и лицемерно долго молитесь: за то примете тем большее осуждение.
MATT|23|15|Горе вам, книжники и фарисеи, лицемеры, что обходите море и сушу, дабы обратить хотя одного; и когда это случится, делаете его сыном геенны, вдвое худшим вас.
MATT|23|16|Горе вам, вожди слепые, которые говорите: если кто поклянется храмом, то ничего, а если кто поклянется золотом храма, то повинен.
MATT|23|17|Безумные и слепые! что больше: золото, или храм, освящающий золото?
MATT|23|18|Также: если кто поклянется жертвенником, то ничего, если же кто поклянется даром, который на нем, то повинен.
MATT|23|19|Безумные и слепые! что больше: дар, или жертвенник, освящающий дар?
MATT|23|20|Итак клянущийся жертвенником клянется им и всем, что на нем;
MATT|23|21|и клянущийся храмом клянется им и Живущим в нем;
MATT|23|22|и клянущийся небом клянется Престолом Божиим и Сидящим на нем.
MATT|23|23|Горе вам, книжники и фарисеи, лицемеры, что даете десятину с мяты, аниса и тмина, и оставили важнейшее в законе: суд, милость и веру; сие надлежало делать, и того не оставлять.
MATT|23|24|Вожди слепые, оцеживающие комара, а верблюда поглощающие!
MATT|23|25|Горе вам, книжники и фарисеи, лицемеры, что очищаете внешность чаши и блюда, между тем как внутри они полны хищения и неправды.
MATT|23|26|Фарисей слепой! очисти прежде внутренность чаши и блюда, чтобы чиста была и внешность их.
MATT|23|27|Горе вам, книжники и фарисеи, лицемеры, что уподобляетесь окрашенным гробам, которые снаружи кажутся красивыми, а внутри полны костей мертвых и всякой нечистоты;
MATT|23|28|так и вы по наружности кажетесь людям праведными, а внутри исполнены лицемерия и беззакония.
MATT|23|29|Горе вам, книжники и фарисеи, лицемеры, что строите гробницы пророкам и украшаете памятники праведников,
MATT|23|30|и говорите: если бы мы были во дни отцов наших, то не были бы сообщниками их в [пролитии] крови пророков;
MATT|23|31|таким образом вы сами против себя свидетельствуете, что вы сыновья тех, которые избили пророков;
MATT|23|32|дополняйте же меру отцов ваших.
MATT|23|33|Змии, порождения ехиднины! как убежите вы от осуждения в геенну?
MATT|23|34|Посему, вот, Я посылаю к вам пророков, и мудрых, и книжников; и вы иных убьете и распнете, а иных будете бить в синагогах ваших и гнать из города в город;
MATT|23|35|да придет на вас вся кровь праведная, пролитая на земле, от крови Авеля праведного до крови Захарии, сына Варахиина, которого вы убили между храмом и жертвенником.
MATT|23|36|Истинно говорю вам, что все сие придет на род сей.
MATT|23|37|Иерусалим, Иерусалим, избивающий пророков и камнями побивающий посланных к тебе! сколько раз хотел Я собрать детей твоих, как птица собирает птенцов своих под крылья, и вы не захотели!
MATT|23|38|Се, оставляется вам дом ваш пуст.
MATT|23|39|Ибо сказываю вам: не увидите Меня отныне, доколе не воскликнете: благословен Грядый во имя Господне!
MATT|24|1|И выйдя, Иисус шел от храма; и приступили ученики Его, чтобы показать Ему здания храма.
MATT|24|2|Иисус же сказал им: видите ли все это? Истинно говорю вам: не останется здесь камня на камне; все будет разрушено.
MATT|24|3|Когда же сидел Он на горе Елеонской, то приступили к Нему ученики наедине и спросили: скажи нам, когда это будет? и какой признак Твоего пришествия и кончины века?
MATT|24|4|Иисус сказал им в ответ: берегитесь, чтобы кто не прельстил вас,
MATT|24|5|ибо многие придут под именем Моим, и будут говорить: "Я Христос", и многих прельстят.
MATT|24|6|Также услышите о войнах и о военных слухах. Смотрите, не ужасайтесь, ибо надлежит всему тому быть, но это еще не конец:
MATT|24|7|ибо восстанет народ на народ, и царство на царство; и будут глады, моры и землетрясения по местам;
MATT|24|8|все же это – начало болезней.
MATT|24|9|Тогда будут предавать вас на мучения и убивать вас; и вы будете ненавидимы всеми народами за имя Мое;
MATT|24|10|и тогда соблазнятся многие, и друг друга будут предавать, и возненавидят друг друга;
MATT|24|11|и многие лжепророки восстанут, и прельстят многих;
MATT|24|12|и, по причине умножения беззакония, во многих охладеет любовь;
MATT|24|13|претерпевший же до конца спасется.
MATT|24|14|И проповедано будет сие Евангелие Царствия по всей вселенной, во свидетельство всем народам; и тогда придет конец.
MATT|24|15|Итак, когда увидите мерзость запустения, реченную через пророка Даниила, стоящую на святом месте, – читающий да разумеет, –
MATT|24|16|тогда находящиеся в Иудее да бегут в горы;
MATT|24|17|и кто на кровле, тот да не сходит взять что–нибудь из дома своего;
MATT|24|18|и кто на поле, тот да не обращается назад взять одежды свои.
MATT|24|19|Горе же беременным и питающим сосцами в те дни!
MATT|24|20|Молитесь, чтобы не случилось бегство ваше зимою или в субботу,
MATT|24|21|ибо тогда будет великая скорбь, какой не было от начала мира доныне, и не будет.
MATT|24|22|И если бы не сократились те дни, то не спаслась бы никакая плоть; но ради избранных сократятся те дни.
MATT|24|23|Тогда, если кто скажет вам: вот, здесь Христос, или там, – не верьте.
MATT|24|24|Ибо восстанут лжехристы и лжепророки, и дадут великие знамения и чудеса, чтобы прельстить, если возможно, и избранных.
MATT|24|25|Вот, Я наперед сказал вам.
MATT|24|26|Итак, если скажут вам: "вот, [Он] в пустыне", – не выходите; "вот, [Он] в потаенных комнатах", – не верьте;
MATT|24|27|ибо, как молния исходит от востока и видна бывает даже до запада, так будет пришествие Сына Человеческого;
MATT|24|28|ибо, где будет труп, там соберутся орлы.
MATT|24|29|И вдруг, после скорби дней тех, солнце померкнет, и луна не даст света своего, и звезды спадут с неба, и силы небесные поколеблются;
MATT|24|30|тогда явится знамение Сына Человеческого на небе; и тогда восплачутся все племена земные и увидят Сына Человеческого, грядущего на облаках небесных с силою и славою великою;
MATT|24|31|и пошлет Ангелов Своих с трубою громогласною, и соберут избранных Его от четырех ветров, от края небес до края их.
MATT|24|32|От смоковницы возьмите подобие: когда ветви ее становятся уже мягки и пускают листья, то знаете, что близко лето;
MATT|24|33|так, когда вы увидите все сие, знайте, что близко, при дверях.
MATT|24|34|Истинно говорю вам: не прейдет род сей, как все сие будет;
MATT|24|35|небо и земля прейдут, но слова Мои не прейдут.
MATT|24|36|О дне же том и часе никто не знает, ни Ангелы небесные, а только Отец Мой один;
MATT|24|37|но, как было во дни Ноя, так будет и в пришествие Сына Человеческого:
MATT|24|38|ибо, как во дни перед потопом ели, пили, женились и выходили замуж, до того дня, как вошел Ной в ковчег,
MATT|24|39|и не думали, пока не пришел потоп и не истребил всех, – так будет и пришествие Сына Человеческого;
MATT|24|40|тогда будут двое на поле: один берется, а другой оставляется;
MATT|24|41|две мелющие в жерновах: одна берется, а другая оставляется.
MATT|24|42|Итак бодрствуйте, потому что не знаете, в который час Господь ваш приидет.
MATT|24|43|Но это вы знаете, что, если бы ведал хозяин дома, в какую стражу придет вор, то бодрствовал бы и не дал бы подкопать дома своего.
MATT|24|44|Потому и вы будьте готовы, ибо в который час не думаете, приидет Сын Человеческий.
MATT|24|45|Кто же верный и благоразумный раб, которого господин его поставил над слугами своими, чтобы давать им пищу во время?
MATT|24|46|Блажен тот раб, которого господин его, придя, найдет поступающим так;
MATT|24|47|истинно говорю вам, что над всем имением своим поставит его.
MATT|24|48|Если же раб тот, будучи зол, скажет в сердце своем: не скоро придет господин мой,
MATT|24|49|и начнет бить товарищей своих и есть и пить с пьяницами, –
MATT|24|50|то придет господин раба того в день, в который он не ожидает, и в час, в который не думает,
MATT|24|51|и рассечет его, и подвергнет его одной участи с лицемерами; там будет плач и скрежет зубов.
MATT|25|1|Тогда подобно будет Царство Небесное десяти девам, которые, взяв светильники свои, вышли навстречу жениху.
MATT|25|2|Из них пять было мудрых и пять неразумных.
MATT|25|3|Неразумные, взяв светильники свои, не взяли с собою масла.
MATT|25|4|Мудрые же, вместе со светильниками своими, взяли масла в сосудах своих.
MATT|25|5|И как жених замедлил, то задремали все и уснули.
MATT|25|6|Но в полночь раздался крик: вот, жених идет, выходите навстречу ему.
MATT|25|7|Тогда встали все девы те и поправили светильники свои.
MATT|25|8|Неразумные же сказали мудрым: дайте нам вашего масла, потому что светильники наши гаснут.
MATT|25|9|А мудрые отвечали: чтобы не случилось недостатка и у нас и у вас, пойдите лучше к продающим и купите себе.
MATT|25|10|Когда же пошли они покупать, пришел жених, и готовые вошли с ним на брачный пир, и двери затворились;
MATT|25|11|после приходят и прочие девы, и говорят: Господи! Господи! отвори нам.
MATT|25|12|Он же сказал им в ответ: истинно говорю вам: не знаю вас.
MATT|25|13|Итак, бодрствуйте, потому что не знаете ни дня, ни часа, в который приидет Сын Человеческий.
MATT|25|14|Ибо [Он поступит], как человек, который, отправляясь в чужую страну, призвал рабов своих и поручил им имение свое:
MATT|25|15|и одному дал он пять талантов, другому два, иному один, каждому по его силе; и тотчас отправился.
MATT|25|16|Получивший пять талантов пошел, употребил их в дело и приобрел другие пять талантов;
MATT|25|17|точно так же и получивший два таланта приобрел другие два;
MATT|25|18|получивший же один талант пошел и закопал [его] в землю и скрыл серебро господина своего.
MATT|25|19|По долгом времени, приходит господин рабов тех и требует у них отчета.
MATT|25|20|И, подойдя, получивший пять талантов принес другие пять талантов и говорит: господин! пять талантов ты дал мне; вот, другие пять талантов я приобрел на них.
MATT|25|21|Господин его сказал ему: хорошо, добрый и верный раб! в малом ты был верен, над многим тебя поставлю; войди в радость господина твоего.
MATT|25|22|Подошел также и получивший два таланта и сказал: господин! два таланта ты дал мне; вот, другие два таланта я приобрел на них.
MATT|25|23|Господин его сказал ему: хорошо, добрый и верный раб! в малом ты был верен, над многим тебя поставлю; войди в радость господина твоего.
MATT|25|24|Подошел и получивший один талант и сказал: господин! я знал тебя, что ты человек жестокий, жнешь, где не сеял, и собираешь, где не рассыпал,
MATT|25|25|и, убоявшись, пошел и скрыл талант твой в земле; вот тебе твое.
MATT|25|26|Господин же его сказал ему в ответ: лукавый раб и ленивый! ты знал, что я жну, где не сеял, и собираю, где не рассыпал;
MATT|25|27|посему надлежало тебе отдать серебро мое торгующим, и я, придя, получил бы мое с прибылью;
MATT|25|28|итак, возьмите у него талант и дайте имеющему десять талантов,
MATT|25|29|ибо всякому имеющему дастся и приумножится, а у неимеющего отнимется и то, что имеет;
MATT|25|30|а негодного раба выбросьте во тьму внешнюю: там будет плач и скрежет зубов. Сказав сие, возгласил: кто имеет уши слышать, да слышит!
MATT|25|31|Когда же приидет Сын Человеческий во славе Своей и все святые Ангелы с Ним, тогда сядет на престоле славы Своей,
MATT|25|32|и соберутся пред Ним все народы; и отделит одних от других, как пастырь отделяет овец от козлов;
MATT|25|33|и поставит овец по правую Свою сторону, а козлов – по левую.
MATT|25|34|Тогда скажет Царь тем, которые по правую сторону Его: приидите, благословенные Отца Моего, наследуйте Царство, уготованное вам от создания мира:
MATT|25|35|ибо алкал Я, и вы дали Мне есть; жаждал, и вы напоили Меня; был странником, и вы приняли Меня;
MATT|25|36|был наг, и вы одели Меня; был болен, и вы посетили Меня; в темнице был, и вы пришли ко Мне.
MATT|25|37|Тогда праведники скажут Ему в ответ: Господи! когда мы видели Тебя алчущим, и накормили? или жаждущим, и напоили?
MATT|25|38|когда мы видели Тебя странником, и приняли? или нагим, и одели?
MATT|25|39|когда мы видели Тебя больным, или в темнице, и пришли к Тебе?
MATT|25|40|И Царь скажет им в ответ: истинно говорю вам: так как вы сделали это одному из сих братьев Моих меньших, то сделали Мне.
MATT|25|41|Тогда скажет и тем, которые по левую сторону: идите от Меня, проклятые, в огонь вечный, уготованный диаволу и ангелам его:
MATT|25|42|ибо алкал Я, и вы не дали Мне есть; жаждал, и вы не напоили Меня;
MATT|25|43|был странником, и не приняли Меня; был наг, и не одели Меня; болен и в темнице, и не посетили Меня.
MATT|25|44|Тогда и они скажут Ему в ответ: Господи! когда мы видели Тебя алчущим, или жаждущим, или странником, или нагим, или больным, или в темнице, и не послужили Тебе?
MATT|25|45|Тогда скажет им в ответ: истинно говорю вам: так как вы не сделали этого одному из сих меньших, то не сделали Мне.
MATT|25|46|И пойдут сии в муку вечную, а праведники в жизнь вечную.
MATT|26|1|Когда Иисус окончил все слова сии, то сказал ученикам Своим:
MATT|26|2|вы знаете, что через два дня будет Пасха, и Сын Человеческий предан будет на распятие.
MATT|26|3|Тогда собрались первосвященники и книжники и старейшины народа во двор первосвященника, по имени Каиафы,
MATT|26|4|и положили в совете взять Иисуса хитростью и убить;
MATT|26|5|но говорили: только не в праздник, чтобы не сделалось возмущения в народе.
MATT|26|6|Когда же Иисус был в Вифании, в доме Симона прокаженного,
MATT|26|7|приступила к Нему женщина с алавастровым сосудом мира драгоценного и возливала Ему возлежащему на голову.
MATT|26|8|Увидев это, ученики Его вознегодовали и говорили: к чему такая трата?
MATT|26|9|Ибо можно было бы продать это миро за большую цену и дать нищим.
MATT|26|10|Но Иисус, уразумев сие, сказал им: что смущаете женщину? она доброе дело сделала для Меня:
MATT|26|11|ибо нищих всегда имеете с собою, а Меня не всегда имеете;
MATT|26|12|возлив миро сие на тело Мое, она приготовила Меня к погребению;
MATT|26|13|истинно говорю вам: где ни будет проповедано Евангелие сие в целом мире, сказано будет в память ее и о том, что она сделала.
MATT|26|14|Тогда один из двенадцати, называемый Иуда Искариот, пошел к первосвященникам
MATT|26|15|и сказал: что вы дадите мне, и я вам предам Его? Они предложили ему тридцать сребренников;
MATT|26|16|и с того времени он искал удобного случая предать Его.
MATT|26|17|В первый же день опресночный приступили ученики к Иисусу и сказали Ему: где велишь нам приготовить Тебе пасху?
MATT|26|18|Он сказал: пойдите в город к такому–то и скажите ему: Учитель говорит: время Мое близко; у тебя совершу пасху с учениками Моими.
MATT|26|19|Ученики сделали, как повелел им Иисус, и приготовили пасху.
MATT|26|20|Когда же настал вечер, Он возлег с двенадцатью учениками;
MATT|26|21|и когда они ели, сказал: истинно говорю вам, что один из вас предаст Меня.
MATT|26|22|Они весьма опечалились, и начали говорить Ему, каждый из них: не я ли, Господи?
MATT|26|23|Он же сказал в ответ: опустивший со Мною руку в блюдо, этот предаст Меня;
MATT|26|24|впрочем Сын Человеческий идет, как писано о Нем, но горе тому человеку, которым Сын Человеческий предается: лучше было бы этому человеку не родиться.
MATT|26|25|При сем и Иуда, предающий Его, сказал: не я ли, Равви? [Иисус] говорит ему: ты сказал.
MATT|26|26|И когда они ели, Иисус взял хлеб и, благословив, преломил и, раздавая ученикам, сказал: приимите, ядите: сие есть Тело Мое.
MATT|26|27|И, взяв чашу и благодарив, подал им и сказал: пейте из нее все,
MATT|26|28|ибо сие есть Кровь Моя Нового Завета, за многих изливаемая во оставление грехов.
MATT|26|29|Сказываю же вам, что отныне не буду пить от плода сего виноградного до того дня, когда буду пить с вами новое [вино] в Царстве Отца Моего.
MATT|26|30|И, воспев, пошли на гору Елеонскую.
MATT|26|31|Тогда говорит им Иисус: все вы соблазнитесь о Мне в эту ночь, ибо написано: поражу пастыря, и рассеются овцы стада;
MATT|26|32|по воскресении же Моем предварю вас в Галилее.
MATT|26|33|Петр сказал Ему в ответ: если и все соблазнятся о Тебе, я никогда не соблазнюсь.
MATT|26|34|Иисус сказал ему: истинно говорю тебе, что в эту ночь, прежде нежели пропоет петух, трижды отречешься от Меня.
MATT|26|35|Говорит Ему Петр: хотя бы надлежало мне и умереть с Тобою, не отрекусь от Тебя. Подобное говорили и все ученики.
MATT|26|36|Потом приходит с ними Иисус на место, называемое Гефсимания, и говорит ученикам: посидите тут, пока Я пойду, помолюсь там.
MATT|26|37|И, взяв с Собою Петра и обоих сыновей Зеведеевых, начал скорбеть и тосковать.
MATT|26|38|Тогда говорит им Иисус: душа Моя скорбит смертельно; побудьте здесь и бодрствуйте со Мною.
MATT|26|39|И, отойдя немного, пал на лице Свое, молился и говорил: Отче Мой! если возможно, да минует Меня чаша сия; впрочем не как Я хочу, но как Ты.
MATT|26|40|И приходит к ученикам и находит их спящими, и говорит Петру: так ли не могли вы один час бодрствовать со Мною?
MATT|26|41|бодрствуйте и молитесь, чтобы не впасть в искушение: дух бодр, плоть же немощна.
MATT|26|42|Еще, отойдя в другой раз, молился, говоря: Отче Мой! если не может чаша сия миновать Меня, чтобы Мне не пить ее, да будет воля Твоя.
MATT|26|43|И, придя, находит их опять спящими, ибо у них глаза отяжелели.
MATT|26|44|И, оставив их, отошел опять и помолился в третий раз, сказав то же слово.
MATT|26|45|Тогда приходит к ученикам Своим и говорит им: вы все еще спите и почиваете? вот, приблизился час, и Сын Человеческий предается в руки грешников;
MATT|26|46|встаньте, пойдем: вот, приблизился предающий Меня.
MATT|26|47|И, когда еще говорил Он, вот Иуда, один из двенадцати, пришел, и с ним множество народа с мечами и кольями, от первосвященников и старейшин народных.
MATT|26|48|Предающий же Его дал им знак, сказав: Кого я поцелую, Тот и есть, возьмите Его.
MATT|26|49|И, тотчас подойдя к Иисусу, сказал: радуйся, Равви! И поцеловал Его.
MATT|26|50|Иисус же сказал ему: друг, для чего ты пришел? Тогда подошли и возложили руки на Иисуса, и взяли Его.
MATT|26|51|И вот, один из бывших с Иисусом, простерши руку, извлек меч свой и, ударив раба первосвященникова, отсек ему ухо.
MATT|26|52|Тогда говорит ему Иисус: возврати меч твой в его место, ибо все, взявшие меч, мечом погибнут;
MATT|26|53|или думаешь, что Я не могу теперь умолить Отца Моего, и Он представит Мне более, нежели двенадцать легионов Ангелов?
MATT|26|54|как же сбудутся Писания, что так должно быть?
MATT|26|55|В тот час сказал Иисус народу: как будто на разбойника вышли вы с мечами и кольями взять Меня; каждый день с вами сидел Я, уча в храме, и вы не брали Меня.
MATT|26|56|Сие же все было, да сбудутся писания пророков. Тогда все ученики, оставив Его, бежали.
MATT|26|57|А взявшие Иисуса отвели Его к Каиафе первосвященнику, куда собрались книжники и старейшины.
MATT|26|58|Петр же следовал за Ним издали, до двора первосвященникова; и, войдя внутрь, сел со служителями, чтобы видеть конец.
MATT|26|59|Первосвященники и старейшины и весь синедрион искали лжесвидетельства против Иисуса, чтобы предать Его смерти,
MATT|26|60|и не находили; и, хотя много лжесвидетелей приходило, не нашли. Но наконец пришли два лжесвидетеля
MATT|26|61|и сказали: Он говорил: могу разрушить храм Божий и в три дня создать его.
MATT|26|62|И, встав, первосвященник сказал Ему: [что же] ничего не отвечаешь? что они против Тебя свидетельствуют?
MATT|26|63|Иисус молчал. И первосвященник сказал Ему: заклинаю Тебя Богом живым, скажи нам, Ты ли Христос, Сын Божий?
MATT|26|64|Иисус говорит ему: ты сказал; даже сказываю вам: отныне узрите Сына Человеческого, сидящего одесную силы и грядущего на облаках небесных.
MATT|26|65|Тогда первосвященник разодрал одежды свои и сказал: Он богохульствует! на что еще нам свидетелей? вот, теперь вы слышали богохульство Его!
MATT|26|66|как вам кажется? Они же сказали в ответ: повинен смерти.
MATT|26|67|Тогда плевали Ему в лице и заушали Его; другие же ударяли Его по ланитам
MATT|26|68|и говорили: прореки нам, Христос, кто ударил Тебя?
MATT|26|69|Петр же сидел вне на дворе. И подошла к нему одна служанка и сказала: и ты был с Иисусом Галилеянином.
MATT|26|70|Но он отрекся перед всеми, сказав: не знаю, что ты говоришь.
MATT|26|71|Когда же он выходил за ворота, увидела его другая, и говорит бывшим там: и этот был с Иисусом Назореем.
MATT|26|72|И он опять отрекся с клятвою, что не знает Сего Человека.
MATT|26|73|Немного спустя подошли стоявшие там и сказали Петру: точно и ты из них, ибо и речь твоя обличает тебя.
MATT|26|74|Тогда он начал клясться и божиться, что не знает Сего Человека. И вдруг запел петух.
MATT|26|75|И вспомнил Петр слово, сказанное ему Иисусом: прежде нежели пропоет петух, трижды отречешься от Меня. И выйдя вон, плакал горько.
MATT|27|1|Когда же настало утро, все первосвященники и старейшины народа имели совещание об Иисусе, чтобы предать Его смерти;
MATT|27|2|и, связав Его, отвели и предали Его Понтию Пилату, правителю.
MATT|27|3|Тогда Иуда, предавший Его, увидев, что Он осужден, и, раскаявшись, возвратил тридцать сребренников первосвященникам и старейшинам,
MATT|27|4|говоря: согрешил я, предав кровь невинную. Они же сказали ему: что нам до того? смотри сам.
MATT|27|5|И, бросив сребренники в храме, он вышел, пошел и удавился.
MATT|27|6|Первосвященники, взяв сребренники, сказали: непозволительно положить их в сокровищницу церковную, потому что это цена крови.
MATT|27|7|Сделав же совещание, купили на них землю горшечника, для погребения странников;
MATT|27|8|посему и называется земля та "землею крови" до сего дня.
MATT|27|9|Тогда сбылось реченное через пророка Иеремию, который говорит: и взяли тридцать сребренников, цену Оцененного, Которого оценили сыны Израиля,
MATT|27|10|и дали их за землю горшечника, как сказал мне Господь.
MATT|27|11|Иисус же стал пред правителем. И спросил Его правитель: Ты Царь Иудейский? Иисус сказал ему: ты говоришь.
MATT|27|12|И когда обвиняли Его первосвященники и старейшины, Он ничего не отвечал.
MATT|27|13|Тогда говорит Ему Пилат: не слышишь, сколько свидетельствуют против Тебя?
MATT|27|14|И не отвечал ему ни на одно слово, так что правитель весьма дивился.
MATT|27|15|На праздник же [Пасхи] правитель имел обычай отпускать народу одного узника, которого хотели.
MATT|27|16|Был тогда у них известный узник, называемый Варавва;
MATT|27|17|итак, когда собрались они, сказал им Пилат: кого хотите, чтобы я отпустил вам: Варавву, или Иисуса, называемого Христом?
MATT|27|18|ибо знал, что предали Его из зависти.
MATT|27|19|Между тем, как сидел он на судейском месте, жена его послала ему сказать: не делай ничего Праведнику Тому, потому что я ныне во сне много пострадала за Него.
MATT|27|20|Но первосвященники и старейшины возбудили народ просить Варавву, а Иисуса погубить.
MATT|27|21|Тогда правитель спросил их: кого из двух хотите, чтобы я отпустил вам? Они сказали: Варавву.
MATT|27|22|Пилат говорит им: что же я сделаю Иисусу, называемому Христом? Говорят ему все: да будет распят.
MATT|27|23|Правитель сказал: какое же зло сделал Он? Но они еще сильнее кричали: да будет распят.
MATT|27|24|Пилат, видя, что ничто не помогает, но смятение увеличивается, взял воды и умыл руки перед народом, и сказал: невиновен я в крови Праведника Сего; смотрите вы.
MATT|27|25|И, отвечая, весь народ сказал: кровь Его на нас и на детях наших.
MATT|27|26|Тогда отпустил им Варавву, а Иисуса, бив, предал на распятие.
MATT|27|27|Тогда воины правителя, взяв Иисуса в преторию, собрали на Него весь полк
MATT|27|28|и, раздев Его, надели на Него багряницу;
MATT|27|29|и, сплетши венец из терна, возложили Ему на голову и дали Ему в правую руку трость; и, становясь пред Ним на колени, насмехались над Ним, говоря: радуйся, Царь Иудейский!
MATT|27|30|и плевали на Него и, взяв трость, били Его по голове.
MATT|27|31|И когда насмеялись над Ним, сняли с Него багряницу, и одели Его в одежды Его, и повели Его на распятие.
MATT|27|32|Выходя, они встретили одного Киринеянина, по имени Симона; сего заставили нести крест Его.
MATT|27|33|И, придя на место, называемое Голгофа, что значит: Лобное место,
MATT|27|34|дали Ему пить уксуса, смешанного с желчью; и, отведав, не хотел пить.
MATT|27|35|Распявшие же Его делили одежды Его, бросая жребий;
MATT|27|36|и, сидя, стерегли Его там;
MATT|27|37|и поставили над головою Его надпись, означающую вину Его: Сей есть Иисус, Царь Иудейский.
MATT|27|38|Тогда распяты с Ним два разбойника: один по правую сторону, а другой по левую.
MATT|27|39|Проходящие же злословили Его, кивая головами своими
MATT|27|40|и говоря: Разрушающий храм и в три дня Созидающий! спаси Себя Самого; если Ты Сын Божий, сойди с креста.
MATT|27|41|Подобно и первосвященники с книжниками и старейшинами и фарисеями, насмехаясь, говорили:
MATT|27|42|других спасал, а Себя Самого не может спасти; если Он Царь Израилев, пусть теперь сойдет с креста, и уверуем в Него;
MATT|27|43|уповал на Бога; пусть теперь избавит Его, если Он угоден Ему. Ибо Он сказал: Я Божий Сын.
MATT|27|44|Также и разбойники, распятые с Ним, поносили Его.
MATT|27|45|От шестого же часа тьма была по всей земле до часа девятого;
MATT|27|46|а около девятого часа возопил Иисус громким голосом: Или, Или! лама савахфани? то есть: Боже Мой, Боже Мой! для чего Ты Меня оставил?
MATT|27|47|Некоторые из стоявших там, слыша это, говорили: Илию зовет Он.
MATT|27|48|И тотчас побежал один из них, взял губку, наполнил уксусом и, наложив на трость, давал Ему пить;
MATT|27|49|а другие говорили: постой, посмотрим, придет ли Илия спасти Его.
MATT|27|50|Иисус же, опять возопив громким голосом, испустил дух.
MATT|27|51|И вот, завеса в храме раздралась надвое, сверху донизу; и земля потряслась; и камни расселись;
MATT|27|52|и гробы отверзлись; и многие тела усопших святых воскресли
MATT|27|53|и, выйдя из гробов по воскресении Его, вошли во святый град и явились многим.
MATT|27|54|Сотник же и те, которые с ним стерегли Иисуса, видя землетрясение и все бывшее, устрашились весьма и говорили: воистину Он был Сын Божий.
MATT|27|55|Там были также и смотрели издали многие женщины, которые следовали за Иисусом из Галилеи, служа Ему;
MATT|27|56|между ними были Мария Магдалина и Мария, мать Иакова и Иосии, и мать сыновей Зеведеевых.
MATT|27|57|Когда же настал вечер, пришел богатый человек из Аримафеи, именем Иосиф, который также учился у Иисуса;
MATT|27|58|он, придя к Пилату, просил тела Иисусова. Тогда Пилат приказал отдать тело;
MATT|27|59|и, взяв тело, Иосиф обвил его чистою плащаницею
MATT|27|60|и положил его в новом своем гробе, который высек он в скале; и, привалив большой камень к двери гроба, удалился.
MATT|27|61|Была же там Мария Магдалина и другая Мария, которые сидели против гроба.
MATT|27|62|На другой день, который следует за пятницею, собрались первосвященники и фарисеи к Пилату
MATT|27|63|и говорили: господин! Мы вспомнили, что обманщик тот, еще будучи в живых, сказал: после трех дней воскресну;
MATT|27|64|итак прикажи охранять гроб до третьего дня, чтобы ученики Его, придя ночью, не украли Его и не сказали народу: воскрес из мертвых; и будет последний обман хуже первого.
MATT|27|65|Пилат сказал им: имеете стражу; пойдите, охраняйте, как знаете.
MATT|27|66|Они пошли и поставили у гроба стражу, и приложили к камню печать.
MATT|28|1|По прошествии же субботы, на рассвете первого дня недели, пришла Мария Магдалина и другая Мария посмотреть гроб.
MATT|28|2|И вот, сделалось великое землетрясение, ибо Ангел Господень, сошедший с небес, приступив, отвалил камень от двери гроба и сидел на нем;
MATT|28|3|вид его был, как молния, и одежда его бела, как снег;
MATT|28|4|устрашившись его, стерегущие пришли в трепет и стали, как мертвые;
MATT|28|5|Ангел же, обратив речь к женщинам, сказал: не бойтесь, ибо знаю, что вы ищете Иисуса распятого;
MATT|28|6|Его нет здесь – Он воскрес, как сказал. Подойдите, посмотрите место, где лежал Господь,
MATT|28|7|и пойдите скорее, скажите ученикам Его, что Он воскрес из мертвых и предваряет вас в Галилее; там Его увидите. Вот, я сказал вам.
MATT|28|8|И, выйдя поспешно из гроба, они со страхом и радостью великою побежали возвестить ученикам Его.
MATT|28|9|Когда же шли они возвестить ученикам Его, и се Иисус встретил их и сказал: радуйтесь! И они, приступив, ухватились за ноги Его и поклонились Ему.
MATT|28|10|Тогда говорит им Иисус: не бойтесь; пойдите, возвестите братьям Моим, чтобы шли в Галилею, и там они увидят Меня.
MATT|28|11|Когда же они шли, то некоторые из стражи, войдя в город, объявили первосвященникам о всем бывшем.
MATT|28|12|И сии, собравшись со старейшинами и сделав совещание, довольно денег дали воинам,
MATT|28|13|и сказали: скажите, что ученики Его, придя ночью, украли Его, когда мы спали;
MATT|28|14|и, если слух об этом дойдет до правителя, мы убедим его, и вас от неприятности избавим.
MATT|28|15|Они, взяв деньги, поступили, как научены были; и пронеслось слово сие между иудеями до сего дня.
MATT|28|16|Одиннадцать же учеников пошли в Галилею, на гору, куда повелел им Иисус,
MATT|28|17|и, увидев Его, поклонились Ему, а иные усомнились.
MATT|28|18|И приблизившись Иисус сказал им: дана Мне всякая власть на небе и на земле.
MATT|28|19|Итак идите, научите все народы, крестя их во имя Отца и Сына и Святаго Духа,
MATT|28|20|уча их соблюдать все, что Я повелел вам; и се, Я с вами во все дни до скончания века. Аминь.
