MARK|1|1|Начало Евангелия Иисуса Христа, Сына Божия,
MARK|1|2|как написано у пророков: вот, Я посылаю Ангела Моего пред лицем Твоим, который приготовит путь Твой пред Тобою.
MARK|1|3|Глас вопиющего в пустыне: приготовьте путь Господу, прямыми сделайте стези Ему.
MARK|1|4|Явился Иоанн, крестя в пустыне и проповедуя крещение покаяния для прощения грехов.
MARK|1|5|И выходили к нему вся страна Иудейская и Иерусалимляне, и крестились от него все в реке Иордане, исповедуя грехи свои.
MARK|1|6|Иоанн же носил одежду из верблюжьего волоса и пояс кожаный на чреслах своих, и ел акриды и дикий мед.
MARK|1|7|И проповедывал, говоря: идет за мною Сильнейший меня, у Которого я недостоин, наклонившись, развязать ремень обуви Его;
MARK|1|8|я крестил вас водою, а Он будет крестить вас Духом Святым.
MARK|1|9|И было в те дни, пришел Иисус из Назарета Галилейского и крестился от Иоанна в Иордане.
MARK|1|10|И когда выходил из воды, тотчас увидел [Иоанн] разверзающиеся небеса и Духа, как голубя, сходящего на Него.
MARK|1|11|И глас был с небес: Ты Сын Мой возлюбленный, в Котором Мое благоволение.
MARK|1|12|Немедленно после того Дух ведет Его в пустыню.
MARK|1|13|И был Он там в пустыне сорок дней, искушаемый сатаною, и был со зверями; и Ангелы служили Ему.
MARK|1|14|После же того, как предан был Иоанн, пришел Иисус в Галилею, проповедуя Евангелие Царствия Божия
MARK|1|15|и говоря, что исполнилось время и приблизилось Царствие Божие: покайтесь и веруйте в Евангелие.
MARK|1|16|Проходя же близ моря Галилейского, увидел Симона и Андрея, брата его, закидывающих сети в море, ибо они были рыболовы.
MARK|1|17|И сказал им Иисус: идите за Мною, и Я сделаю, что вы будете ловцами человеков.
MARK|1|18|И они тотчас, оставив свои сети, последовали за Ним.
MARK|1|19|И, пройдя оттуда немного, Он увидел Иакова Зеведеева и Иоанна, брата его, также в лодке починивающих сети;
MARK|1|20|и тотчас призвал их. И они, оставив отца своего Зеведея в лодке с работниками, последовали за Ним.
MARK|1|21|И приходят в Капернаум; и вскоре в субботу вошел Он в синагогу и учил.
MARK|1|22|И дивились Его учению, ибо Он учил их, как власть имеющий, а не как книжники.
MARK|1|23|В синагоге их был человек, [одержимый] духом нечистым, и вскричал:
MARK|1|24|оставь! что Тебе до нас, Иисус Назарянин? Ты пришел погубить нас! знаю Тебя, кто Ты, Святый Божий.
MARK|1|25|Но Иисус запретил ему, говоря: замолчи и выйди из него.
MARK|1|26|Тогда дух нечистый, сотрясши его и вскричав громким голосом, вышел из него.
MARK|1|27|И все ужаснулись, так что друг друга спрашивали: что это? что это за новое учение, что Он и духам нечистым повелевает со властью, и они повинуются Ему?
MARK|1|28|И скоро разошлась о Нем молва по всей окрестности в Галилее.
MARK|1|29|Выйдя вскоре из синагоги, пришли в дом Симона и Андрея, с Иаковом и Иоанном.
MARK|1|30|Теща же Симонова лежала в горячке; и тотчас говорят Ему о ней.
MARK|1|31|Подойдя, Он поднял ее, взяв ее за руку; и горячка тотчас оставила ее, и она стала служить им.
MARK|1|32|При наступлении же вечера, когда заходило солнце, приносили к Нему всех больных и бесноватых.
MARK|1|33|И весь город собрался к дверям.
MARK|1|34|И Он исцелил многих, страдавших различными болезнями; изгнал многих бесов, и не позволял бесам говорить, что они знают, что Он Христос.
MARK|1|35|А утром, встав весьма рано, вышел и удалился в пустынное место, и там молился.
MARK|1|36|Симон и бывшие с ним пошли за Ним
MARK|1|37|и, найдя Его, говорят Ему: все ищут Тебя.
MARK|1|38|Он говорит им: пойдем в ближние селения и города, чтобы Мне и там проповедывать, ибо Я для того пришел.
MARK|1|39|И Он проповедывал в синагогах их по всей Галилее и изгонял бесов.
MARK|1|40|Приходит к Нему прокаженный и, умоляя Его и падая пред Ним на колени, говорит Ему: если хочешь, можешь меня очистить.
MARK|1|41|Иисус, умилосердившись над ним, простер руку, коснулся его и сказал ему: хочу, очистись.
MARK|1|42|После сего слова проказа тотчас сошла с него, и он стал чист.
MARK|1|43|И, посмотрев на него строго, тотчас отослал его
MARK|1|44|и сказал ему: смотри, никому ничего не говори, но пойди, покажись священнику и принеси за очищение твое, что повелел Моисей, во свидетельство им.
MARK|1|45|А он, выйдя, начал провозглашать и рассказывать о происшедшем, так что [Иисус] не мог уже явно войти в город, но находился вне, в местах пустынных. И приходили к Нему отовсюду.
MARK|2|1|Через [несколько] дней опять пришел Он в Капернаум; и слышно стало, что Он в доме.
MARK|2|2|Тотчас собрались многие, так что уже и у дверей не было места; и Он говорил им слово.
MARK|2|3|И пришли к Нему с расслабленным, которого несли четверо;
MARK|2|4|и, не имея возможности приблизиться к Нему за многолюдством, раскрыли кровлю [дома], где Он находился, и, прокопав ее, спустили постель, на которой лежал расслабленный.
MARK|2|5|Иисус, видя веру их, говорит расслабленному: чадо! прощаются тебе грехи твои.
MARK|2|6|Тут сидели некоторые из книжников и помышляли в сердцах своих:
MARK|2|7|что Он так богохульствует? кто может прощать грехи, кроме одного Бога?
MARK|2|8|Иисус, тотчас узнав духом Своим, что они так помышляют в себе, сказал им: для чего так помышляете в сердцах ваших?
MARK|2|9|Что легче? сказать ли расслабленному: прощаются тебе грехи? или сказать: встань, возьми свою постель и ходи?
MARK|2|10|Но чтобы вы знали, что Сын Человеческий имеет власть на земле прощать грехи, – говорит расслабленному:
MARK|2|11|тебе говорю: встань, возьми постель твою и иди в дом твой.
MARK|2|12|Он тотчас встал и, взяв постель, вышел перед всеми, так что все изумлялись и прославляли Бога, говоря: никогда ничего такого мы не видали.
MARK|2|13|И вышел [Иисус] опять к морю; и весь народ пошел к Нему, и Он учил их.
MARK|2|14|Проходя, увидел Он Левия Алфеева, сидящего у сбора пошлин, и говорит ему: следуй за Мною. И [он], встав, последовал за Ним.
MARK|2|15|И когда Иисус возлежал в доме его, возлежали с Ним и ученики Его и многие мытари и грешники: ибо много их было, и они следовали за Ним.
MARK|2|16|Книжники и фарисеи, увидев, что Он ест с мытарями и грешниками, говорили ученикам Его: как это Он ест и пьет с мытарями и грешниками.
MARK|2|17|Услышав [сие], Иисус говорит им: не здоровые имеют нужду во враче, но больные; Я пришел призвать не праведников, но грешников к покаянию.
MARK|2|18|Ученики Иоанновы и фарисейские постились. Приходят к Нему и говорят: почему ученики Иоанновы и фарисейские постятся, а Твои ученики не постятся?
MARK|2|19|И сказал им Иисус: могут ли поститься сыны чертога брачного, когда с ними жених? Доколе с ними жених, не могут поститься,
MARK|2|20|но придут дни, когда отнимется у них жених, и тогда будут поститься в те дни.
MARK|2|21|Никто к ветхой одежде не приставляет заплаты из небеленой ткани: иначе вновь пришитое отдерет от старого, и дыра будет еще хуже.
MARK|2|22|Никто не вливает вина молодого в мехи ветхие: иначе молодое вино прорвет мехи, и вино вытечет, и мехи пропадут; но вино молодое надобно вливать в мехи новые.
MARK|2|23|И случилось Ему в субботу проходить засеянными [полями], и ученики Его дорогою начали срывать колосья.
MARK|2|24|И фарисеи сказали Ему: смотри, что они делают в субботу, чего не должно [делать]?
MARK|2|25|Он сказал им: неужели вы не читали никогда, что сделал Давид, когда имел нужду и взалкал сам и бывшие с ним?
MARK|2|26|как вошел он в дом Божий при первосвященнике Авиафаре и ел хлебы предложения, которых не должно было есть никому, кроме священников, и дал и бывшим с ним?
MARK|2|27|И сказал им: суббота для человека, а не человек для субботы;
MARK|2|28|посему Сын Человеческий есть господин и субботы.
MARK|3|1|И пришел опять в синагогу; там был человек, имевший иссохшую руку.
MARK|3|2|И наблюдали за Ним, не исцелит ли его в субботу, чтобы обвинить Его.
MARK|3|3|Он же говорит человеку, имевшему иссохшую руку: стань на средину.
MARK|3|4|А им говорит: должно ли в субботу добро делать, или зло делать? душу спасти, или погубить? Но они молчали.
MARK|3|5|И, воззрев на них с гневом, скорбя об ожесточении сердец их, говорит тому человеку: протяни руку твою. Он протянул, и стала рука его здорова, как другая.
MARK|3|6|Фарисеи, выйдя, немедленно составили с иродианами совещание против Него, как бы погубить Его.
MARK|3|7|Но Иисус с учениками Своими удалился к морю; и за Ним последовало множество народа из Галилеи, Иудеи,
MARK|3|8|Иерусалима, Идумеи и из–за Иордана. И [живущие] в окрестностях Тира и Сидона, услышав, что Он делал, шли к Нему в великом множестве.
MARK|3|9|И сказал ученикам Своим, чтобы готова была для Него лодка по причине многолюдства, дабы не теснили Его.
MARK|3|10|Ибо многих Он исцелил, так что имевшие язвы бросались к Нему, чтобы коснуться Его.
MARK|3|11|И духи нечистые, когда видели Его, падали пред Ним и кричали: Ты Сын Божий.
MARK|3|12|Но Он строго запрещал им, чтобы не делали Его известным.
MARK|3|13|Потом взошел на гору и позвал к Себе, кого Сам хотел; и пришли к Нему.
MARK|3|14|И поставил [из них] двенадцать, чтобы с Ним были и чтобы посылать их на проповедь,
MARK|3|15|и чтобы они имели власть исцелять от болезней и изгонять бесов;
MARK|3|16|[поставил] Симона, нарекши ему имя Петр,
MARK|3|17|Иакова Зеведеева и Иоанна, брата Иакова, нарекши им имена Воанергес, то есть "сыны громовы",
MARK|3|18|Андрея, Филиппа, Варфоломея, Матфея, Фому, Иакова Алфеева, Фаддея, Симона Кананита
MARK|3|19|и Иуду Искариотского, который и предал Его.
MARK|3|20|Приходят в дом; и опять сходится народ, так что им невозможно было и хлеба есть.
MARK|3|21|И, услышав, ближние Его пошли взять Его, ибо говорили, что Он вышел из себя.
MARK|3|22|А книжники, пришедшие из Иерусалима, говорили, что Он имеет [в] [Себе] веельзевула и что изгоняет бесов силою бесовского князя.
MARK|3|23|И, призвав их, говорил им притчами: как может сатана изгонять сатану?
MARK|3|24|Если царство разделится само в себе, не может устоять царство то;
MARK|3|25|и если дом разделится сам в себе, не может устоять дом тот;
MARK|3|26|и если сатана восстал на самого себя и разделился, не может устоять, но пришел конец его.
MARK|3|27|Никто, войдя в дом сильного, не может расхитить вещей его, если прежде не свяжет сильного, и тогда расхитит дом его.
MARK|3|28|Истинно говорю вам: будут прощены сынам человеческим все грехи и хуления, какими бы ни хулили;
MARK|3|29|но кто будет хулить Духа Святаго, тому не будет прощения вовек, но подлежит он вечному осуждению.
MARK|3|30|[Сие сказал Он], потому что говорили: в Нем нечистый дух.
MARK|3|31|И пришли Матерь и братья Его и, стоя [вне] дома, послали к Нему звать Его.
MARK|3|32|Около Него сидел народ. И сказали Ему: вот, Матерь Твоя и братья Твои и сестры Твои, [вне] дома, спрашивают Тебя.
MARK|3|33|И отвечал им: кто матерь Моя и братья Мои?
MARK|3|34|И обозрев сидящих вокруг Себя, говорит: вот матерь Моя и братья Мои;
MARK|3|35|ибо кто будет исполнять волю Божию, тот Мне брат, и сестра, и матерь.
MARK|4|1|И опять начал учить при море; и собралось к Нему множество народа, так что Он вошел в лодку и сидел на море, а весь народ был на земле, у моря.
MARK|4|2|И учил их притчами много, и в учении Своем говорил им:
MARK|4|3|слушайте: вот, вышел сеятель сеять;
MARK|4|4|и, когда сеял, случилось, что иное упало при дороге, и налетели птицы и поклевали то.
MARK|4|5|Иное упало на каменистое [место], где немного было земли, и скоро взошло, потому что земля была неглубока;
MARK|4|6|когда же взошло солнце, увяло и, как не имело корня, засохло.
MARK|4|7|Иное упало в терние, и терние выросло, и заглушило [семя], и оно не дало плода.
MARK|4|8|И иное упало на добрую землю и дало плод, который взошел и вырос, и принесло иное тридцать, иное шестьдесят, и иное сто.
MARK|4|9|И сказал им: кто имеет уши слышать, да слышит!
MARK|4|10|Когда же остался без народа, окружающие Его, вместе с двенадцатью, спросили Его о притче.
MARK|4|11|И сказал им: вам дано знать тайны Царствия Божия, а тем внешним все бывает в притчах;
MARK|4|12|так что они своими глазами смотрят, и не видят; своими ушами слышат, и не разумеют, да не обратятся, и прощены будут им грехи.
MARK|4|13|И говорит им: не понимаете этой притчи? Как же вам уразуметь все притчи?
MARK|4|14|Сеятель слово сеет.
MARK|4|15|[Посеянное] при дороге означает тех, в которых сеется слово, но [к которым], когда услышат, тотчас приходит сатана и похищает слово, посеянное в сердцах их.
MARK|4|16|Подобным образом и посеянное на каменистом [месте] означает тех, которые, когда услышат слово, тотчас с радостью принимают его,
MARK|4|17|но не имеют в себе корня и непостоянны; потом, когда настанет скорбь или гонение за слово, тотчас соблазняются.
MARK|4|18|Посеянное в тернии означает слышащих слово,
MARK|4|19|но в которых заботы века сего, обольщение богатством и другие пожелания, входя в них, заглушают слово, и оно бывает без плода.
MARK|4|20|А посеянное на доброй земле означает тех, которые слушают слово и принимают, и приносят плод, один в тридцать, другой в шестьдесят, иной во сто крат.
MARK|4|21|И сказал им: для того ли приносится свеча, чтобы поставить ее под сосуд или под кровать? не для того ли, чтобы поставить ее на подсвечнике?
MARK|4|22|Нет ничего тайного, что не сделалось бы явным, и ничего не бывает потаенного, что не вышло бы наружу.
MARK|4|23|Если кто имеет уши слышать, да слышит!
MARK|4|24|И сказал им: замечайте, что слышите: какою мерою мерите, такою отмерено будет вам и прибавлено будет вам, слушающим.
MARK|4|25|Ибо кто имеет, тому дано будет, а кто не имеет, у того отнимется и то, что имеет.
MARK|4|26|И сказал: Царствие Божие подобно тому, как если человек бросит семя в землю,
MARK|4|27|и спит, и встает ночью и днем; и как семя всходит и растет, не знает он,
MARK|4|28|ибо земля сама собою производит сперва зелень, потом колос, потом полное зерно в колосе.
MARK|4|29|Когда же созреет плод, немедленно посылает серп, потому что настала жатва.
MARK|4|30|И сказал: чему уподобим Царствие Божие? или какою притчею изобразим его?
MARK|4|31|Оно – как зерно горчичное, которое, когда сеется в землю, есть меньше всех семян на земле;
MARK|4|32|а когда посеяно, всходит и становится больше всех злаков, и пускает большие ветви, так что под тенью его могут укрываться птицы небесные.
MARK|4|33|И таковыми многими притчами проповедывал им слово, сколько они могли слышать.
MARK|4|34|Без притчи же не говорил им, а ученикам наедине изъяснял все.
MARK|4|35|Вечером того дня сказал им: переправимся на ту сторону.
MARK|4|36|И они, отпустив народ, взяли Его с собою, как Он был в лодке; с Ним были и другие лодки.
MARK|4|37|И поднялась великая буря; волны били в лодку, так что она уже наполнялась [водою].
MARK|4|38|А Он спал на корме на возглавии. Его будят и говорят Ему: Учитель! неужели Тебе нужды нет, что мы погибаем?
MARK|4|39|И, встав, Он запретил ветру и сказал морю: умолкни, перестань. И ветер утих, и сделалась великая тишина.
MARK|4|40|И сказал им: что вы так боязливы? как у вас нет веры?
MARK|4|41|И убоялись страхом великим и говорили между собою: кто же Сей, что и ветер и море повинуются Ему?
MARK|5|1|И пришли на другой берег моря, в страну Гадаринскую.
MARK|5|2|И когда вышел Он из лодки, тотчас встретил Его вышедший из гробов человек, [одержимый] нечистым духом,
MARK|5|3|он имел жилище в гробах, и никто не мог его связать даже цепями,
MARK|5|4|потому что многократно был он скован оковами и цепями, но разрывал цепи и разбивал оковы, и никто не в силах был укротить его;
MARK|5|5|всегда, ночью и днем, в горах и гробах, кричал он и бился о камни;
MARK|5|6|увидев же Иисуса издалека, прибежал и поклонился Ему,
MARK|5|7|и, вскричав громким голосом, сказал: что Тебе до меня, Иисус, Сын Бога Всевышнего? заклинаю Тебя Богом, не мучь меня!
MARK|5|8|Ибо [Иисус] сказал ему: выйди, дух нечистый, из сего человека.
MARK|5|9|И спросил его: как тебе имя? И он сказал в ответ: легион имя мне, потому что нас много.
MARK|5|10|И много просили Его, чтобы не высылал их вон из страны той.
MARK|5|11|Паслось же там при горе большое стадо свиней.
MARK|5|12|И просили Его все бесы, говоря: пошли нас в свиней, чтобы нам войти в них.
MARK|5|13|Иисус тотчас позволил им. И нечистые духи, выйдя, вошли в свиней; и устремилось стадо с крутизны в море, а их было около двух тысяч; и потонули в море.
MARK|5|14|Пасущие же свиней побежали и рассказали в городе и в деревнях. И [жители] вышли посмотреть, что случилось.
MARK|5|15|Приходят к Иисусу и видят, что бесновавшийся, в котором был легион, сидит и одет, и в здравом уме; и устрашились.
MARK|5|16|Видевшие рассказали им о том, как это произошло с бесноватым, и о свиньях.
MARK|5|17|И начали просить Его, чтобы отошел от пределов их.
MARK|5|18|И когда Он вошел в лодку, бесновавшийся просил Его, чтобы быть с Ним.
MARK|5|19|Но Иисус не дозволил ему, а сказал: иди домой к своим и расскажи им, что сотворил с тобою Господь и [как] помиловал тебя.
MARK|5|20|И пошел и начал проповедывать в Десятиградии, что сотворил с ним Иисус; и все дивились.
MARK|5|21|Когда Иисус опять переправился в лодке на другой берег, собралось к Нему множество народа. Он был у моря.
MARK|5|22|И вот, приходит один из начальников синагоги, по имени Иаир, и, увидев Его, падает к ногам Его
MARK|5|23|и усильно просит Его, говоря: дочь моя при смерти; приди и возложи на нее руки, чтобы она выздоровела и осталась жива.
MARK|5|24|[Иисус] пошел с ним. За Ним следовало множество народа, и теснили Его.
MARK|5|25|Одна женщина, которая страдала кровотечением двенадцать лет,
MARK|5|26|много потерпела от многих врачей, истощила все, что было у ней, и не получила никакой пользы, но пришла еще в худшее состояние, –
MARK|5|27|услышав об Иисусе, подошла сзади в народе и прикоснулась к одежде Его,
MARK|5|28|ибо говорила: если хотя к одежде Его прикоснусь, то выздоровею.
MARK|5|29|И тотчас иссяк у ней источник крови, и она ощутила в теле, что исцелена от болезни.
MARK|5|30|В то же время Иисус, почувствовав Сам в Себе, что вышла из Него сила, обратился в народе и сказал: кто прикоснулся к Моей одежде?
MARK|5|31|Ученики сказали Ему: Ты видишь, что народ теснит Тебя, и говоришь: кто прикоснулся ко Мне?
MARK|5|32|Но Он смотрел вокруг, чтобы видеть ту, которая сделала это.
MARK|5|33|Женщина в страхе и трепете, зная, что с нею произошло, подошла, пала пред Ним и сказала Ему всю истину.
MARK|5|34|Он же сказал ей: дщерь! вера твоя спасла тебя; иди в мире и будь здорова от болезни твоей.
MARK|5|35|Когда Он еще говорил сие, приходят от начальника синагоги и говорят: дочь твоя умерла; что еще утруждаешь Учителя?
MARK|5|36|Но Иисус, услышав сии слова, тотчас говорит начальнику синагоги: не бойся, только веруй.
MARK|5|37|И не позволил никому следовать за Собою, кроме Петра, Иакова и Иоанна, брата Иакова.
MARK|5|38|Приходит в дом начальника синагоги и видит смятение и плачущих и вопиющих громко.
MARK|5|39|И, войдя, говорит им: что смущаетесь и плачете? девица не умерла, но спит.
MARK|5|40|И смеялись над Ним. Но Он, выслав всех, берет с Собою отца и мать девицы и бывших с Ним и входит туда, где девица лежала.
MARK|5|41|И, взяв девицу за руку, говорит ей: "талифа куми", что значит: девица, тебе говорю, встань.
MARK|5|42|И девица тотчас встала и начала ходить, ибо была лет двенадцати. [Видевшие] пришли в великое изумление.
MARK|5|43|И Он строго приказал им, чтобы никто об этом не знал, и сказал, чтобы дали ей есть.
MARK|6|1|Оттуда вышел Он и пришел в Свое отечество; за Ним следовали ученики Его.
MARK|6|2|Когда наступила суббота, Он начал учить в синагоге; и многие слышавшие с изумлением говорили: откуда у Него это? что за премудрость дана Ему, и как такие чудеса совершаются руками Его?
MARK|6|3|Не плотник ли Он, сын Марии, брат Иакова, Иосии, Иуды и Симона? Не здесь ли, между нами, Его сестры? И соблазнялись о Нем.
MARK|6|4|Иисус же сказал им: не бывает пророк без чести, разве только в отечестве своем и у сродников и в доме своем.
MARK|6|5|И не мог совершить там никакого чуда, только на немногих больных возложив руки, исцелил [их].
MARK|6|6|И дивился неверию их; потом ходил по окрестным селениям и учил.
MARK|6|7|И, призвав двенадцать, начал посылать их по два, и дал им власть над нечистыми духами.
MARK|6|8|И заповедал им ничего не брать в дорогу, кроме одного посоха: ни сумы, ни хлеба, ни меди в поясе,
MARK|6|9|но обуваться в простую обувь и не носить двух одежд.
MARK|6|10|И сказал им: если где войдете в дом, оставайтесь в нем, доколе не выйдете из того места.
MARK|6|11|И если кто не примет вас и не будет слушать вас, то, выходя оттуда, отрясите прах от ног ваших, во свидетельство на них. Истинно говорю вам: отраднее будет Содому и Гоморре в день суда, нежели тому городу.
MARK|6|12|Они пошли и проповедывали покаяние;
MARK|6|13|изгоняли многих бесов и многих больных мазали маслом и исцеляли.
MARK|6|14|Царь Ирод, услышав [об Иисусе], – ибо имя Его стало гласно, – говорил: это Иоанн Креститель воскрес из мертвых, и потому чудеса делаются им.
MARK|6|15|Другие говорили: это Илия, а иные говорили: это пророк, или как один из пророков.
MARK|6|16|Ирод же, услышав, сказал: это Иоанн, которого я обезглавил; он воскрес из мертвых.
MARK|6|17|Ибо сей Ирод, послав, взял Иоанна и заключил его в темницу за Иродиаду, жену Филиппа, брата своего, потому что женился на ней.
MARK|6|18|Ибо Иоанн говорил Ироду: не должно тебе иметь жену брата твоего.
MARK|6|19|Иродиада же, злобясь на него, желала убить его; но не могла.
MARK|6|20|Ибо Ирод боялся Иоанна, зная, что он муж праведный и святой, и берег его; многое делал, слушаясь его, и с удовольствием слушал его.
MARK|6|21|Настал удобный день, когда Ирод, по случаю [дня] рождения своего, делал пир вельможам своим, тысяченачальникам и старейшинам Галилейским, –
MARK|6|22|дочь Иродиады вошла, плясала и угодила Ироду и возлежавшим с ним; царь сказал девице: проси у меня, чего хочешь, и дам тебе;
MARK|6|23|и клялся ей: чего ни попросишь у меня, дам тебе, даже до половины моего царства.
MARK|6|24|Она вышла и спросила у матери своей: чего просить? Та отвечала: головы Иоанна Крестителя.
MARK|6|25|И она тотчас пошла с поспешностью к царю и просила, говоря: хочу, чтобы ты дал мне теперь же на блюде голову Иоанна Крестителя.
MARK|6|26|Царь опечалился, но ради клятвы и возлежавших с ним не захотел отказать ей.
MARK|6|27|И тотчас, послав оруженосца, царь повелел принести голову его.
MARK|6|28|Он пошел, отсек ему голову в темнице, и принес голову его на блюде, и отдал ее девице, а девица отдала ее матери своей.
MARK|6|29|Ученики его, услышав, пришли и взяли тело его, и положили его во гробе.
MARK|6|30|И собрались Апостолы к Иисусу и рассказали Ему все, и что сделали, и чему научили.
MARK|6|31|Он сказал им: пойдите вы одни в пустынное место и отдохните немного, – ибо много было приходящих и отходящих, так что и есть им было некогда.
MARK|6|32|И отправились в пустынное место в лодке одни.
MARK|6|33|Народ увидел, [как] они отправлялись, и многие узнали их; и бежали туда пешие из всех городов, и предупредили их, и собрались к Нему.
MARK|6|34|Иисус, выйдя, увидел множество народа и сжалился над ними, потому что они были, как овцы, не имеющие пастыря; и начал учить их много.
MARK|6|35|И как времени прошло много, ученики Его, приступив к Нему, говорят: место [здесь] пустынное, а времени уже много, –
MARK|6|36|отпусти их, чтобы они пошли в окрестные деревни и селения и купили себе хлеба, ибо им нечего есть.
MARK|6|37|Он сказал им в ответ: вы дайте им есть. И сказали Ему: разве нам пойти купить хлеба динариев на двести и дать им есть?
MARK|6|38|Но Он спросил их: сколько у вас хлебов? пойдите, посмотрите. Они, узнав, сказали: пять хлебов и две рыбы.
MARK|6|39|Тогда повелел им рассадить всех отделениями на зеленой траве.
MARK|6|40|И сели рядами, по сто и по пятидесяти.
MARK|6|41|Он взял пять хлебов и две рыбы, воззрев на небо, благословил и преломил хлебы и дал ученикам Своим, чтобы они раздали им; и две рыбы разделил на всех.
MARK|6|42|И ели все, и насытились.
MARK|6|43|И набрали кусков хлеба и [остатков] от рыб двенадцать полных коробов.
MARK|6|44|Было же евших хлебы около пяти тысяч мужей.
MARK|6|45|И тотчас понудил учеников Своих войти в лодку и отправиться вперед на другую сторону к Вифсаиде, пока Он отпустит народ.
MARK|6|46|И, отпустив их, пошел на гору помолиться.
MARK|6|47|Вечером лодка была посреди моря, а Он один на земле.
MARK|6|48|И увидел их бедствующих в плавании, потому что ветер им был противный; около же четвертой стражи ночи подошел к ним, идя по морю, и хотел миновать их.
MARK|6|49|Они, увидев Его идущего по морю, подумали, что это призрак, и вскричали.
MARK|6|50|Ибо все видели Его и испугались. И тотчас заговорил с ними и сказал им: ободритесь; это Я, не бойтесь.
MARK|6|51|И вошел к ним в лодку, и ветер утих. И они чрезвычайно изумлялись в себе и дивились,
MARK|6|52|ибо не вразумились [чудом] над хлебами, потому что сердце их было окаменено.
MARK|6|53|И, переправившись, прибыли в землю Геннисаретскую и пристали [к] [берегу].
MARK|6|54|Когда вышли они из лодки, тотчас [жители], узнав Его,
MARK|6|55|обежали всю окрестность ту и начали на постелях приносить больных туда, где Он, как слышно было, находился.
MARK|6|56|И куда ни приходил Он, в селения ли, в города ли, в деревни ли, клали больных на открытых местах и просили Его, чтобы им прикоснуться хотя к краю одежды Его; и которые прикасались к Нему, исцелялись.
MARK|7|1|Собрались к Нему фарисеи и некоторые из книжников, пришедшие из Иерусалима,
MARK|7|2|и, увидев некоторых из учеников Его, евших хлеб нечистыми, то есть неумытыми, руками, укоряли.
MARK|7|3|Ибо фарисеи и все Иудеи, держась предания старцев, не едят, не умыв тщательно рук;
MARK|7|4|и, [придя] с торга, не едят не омывшись. Есть и многое другое, чего они приняли держаться: наблюдать омовение чаш, кружек, котлов и скамей.
MARK|7|5|Потом спрашивают Его фарисеи и книжники: зачем ученики Твои не поступают по преданию старцев, но неумытыми руками едят хлеб?
MARK|7|6|Он сказал им в ответ: хорошо пророчествовал о вас, лицемерах, Исаия, как написано: люди сии чтут Меня устами, сердце же их далеко отстоит от Меня,
MARK|7|7|но тщетно чтут Меня, уча учениям, заповедям человеческим.
MARK|7|8|Ибо вы, оставив заповедь Божию, держитесь предания человеческого, омовения кружек и чаш, и делаете многое другое, сему подобное.
MARK|7|9|И сказал им: хорошо ли, [что] вы отменяете заповедь Божию, чтобы соблюсти свое предание?
MARK|7|10|Ибо Моисей сказал: почитай отца своего и мать свою; и: злословящий отца или мать смертью да умрет.
MARK|7|11|А вы говорите: кто скажет отцу или матери: корван, то есть дар [Богу] то, чем бы ты от меня пользовался,
MARK|7|12|тому вы уже попускаете ничего не делать для отца своего или матери своей,
MARK|7|13|устраняя слово Божие преданием вашим, которое вы установили; и делаете многое сему подобное.
MARK|7|14|И, призвав весь народ, говорил им: слушайте Меня все и разумейте:
MARK|7|15|ничто, входящее в человека извне, не может осквернить его; но что исходит из него, то оскверняет человека.
MARK|7|16|Если кто имеет уши слышать, да слышит!
MARK|7|17|И когда Он от народа вошел в дом, ученики Его спросили Его о притче.
MARK|7|18|Он сказал им: неужели и вы так непонятливы? Неужели не разумеете, что ничто, извне входящее в человека, не может осквернить его?
MARK|7|19|Потому что не в сердце его входит, а в чрево, и выходит вон, [чем] очищается всякая пища.
MARK|7|20|Далее сказал: исходящее из человека оскверняет человека.
MARK|7|21|Ибо извнутрь, из сердца человеческого, исходят злые помыслы, прелюбодеяния, любодеяния, убийства,
MARK|7|22|кражи, лихоимство, злоба, коварство, непотребство, завистливое око, богохульство, гордость, безумство, –
MARK|7|23|все это зло извнутрь исходит и оскверняет человека.
MARK|7|24|И, отправившись оттуда, пришел в пределы Тирские и Сидонские; и, войдя в дом, не хотел, чтобы кто узнал; но не мог утаиться.
MARK|7|25|Ибо услышала о Нем женщина, у которой дочь одержима была нечистым духом, и, придя, припала к ногам Его;
MARK|7|26|а женщина та была язычница, родом сирофиникиянка; и просила Его, чтобы изгнал беса из ее дочери.
MARK|7|27|Но Иисус сказал ей: дай прежде насытиться детям, ибо нехорошо взять хлеб у детей и бросить псам.
MARK|7|28|Она же сказала Ему в ответ: так, Господи; но и псы под столом едят крохи у детей.
MARK|7|29|И сказал ей: за это слово, пойди; бес вышел из твоей дочери.
MARK|7|30|И, придя в свой дом, она нашла, что бес вышел и дочь лежит на постели.
MARK|7|31|Выйдя из пределов Тирских и Сидонских, [Иисус] опять пошел к морю Галилейскому через пределы Десятиградия.
MARK|7|32|Привели к Нему глухого косноязычного и просили Его возложить на него руку.
MARK|7|33|[Иисус], отведя его в сторону от народа, вложил персты Свои в уши ему и, плюнув, коснулся языка его;
MARK|7|34|и, воззрев на небо, вздохнул и сказал ему: "еффафа", то есть: отверзись.
MARK|7|35|И тотчас отверзся у него слух и разрешились узы его языка, и стал говорить чисто.
MARK|7|36|И повелел им не сказывать никому. Но сколько Он ни запрещал им, они еще более разглашали.
MARK|7|37|И чрезвычайно дивились, и говорили: все хорошо делает, – и глухих делает слышащими, и немых – говорящими.
MARK|8|1|В те дни, когда собралось весьма много народа и нечего было им есть, Иисус, призвав учеников Своих, сказал им:
MARK|8|2|жаль Мне народа, что уже три дня находятся при Мне, и нечего им есть.
MARK|8|3|Если неевшими отпущу их в домы их, ослабеют в дороге, ибо некоторые из них пришли издалека.
MARK|8|4|Ученики Его отвечали Ему: откуда мог бы кто [взять] здесь в пустыне хлебов, чтобы накормить их?
MARK|8|5|И спросил их: сколько у вас хлебов? Они сказали: семь.
MARK|8|6|Тогда велел народу возлечь на землю; и, взяв семь хлебов и воздав благодарение, преломил и дал ученикам Своим, чтобы они раздали; и они раздали народу.
MARK|8|7|Было у них и немного рыбок: благословив, Он велел раздать и их.
MARK|8|8|И ели, и насытились; и набрали оставшихся кусков семь корзин.
MARK|8|9|Евших же было около четырех тысяч. И отпустил их.
MARK|8|10|И тотчас войдя в лодку с учениками Своими, прибыл в пределы Далмануфские.
MARK|8|11|Вышли фарисеи, начали с Ним спорить и требовали от Него знамения с неба, искушая Его.
MARK|8|12|И Он, глубоко вздохнув, сказал: для чего род сей требует знамения? Истинно говорю вам, не дастся роду сему знамение.
MARK|8|13|И, оставив их, опять вошел в лодку и отправился на ту сторону.
MARK|8|14|При сем ученики Его забыли взять хлебов и кроме одного хлеба не имели с собою в лодке.
MARK|8|15|А Он заповедал им, говоря: смотрите, берегитесь закваски фарисейской и закваски Иродовой.
MARK|8|16|И, рассуждая между собою, говорили: [это значит], что хлебов нет у нас.
MARK|8|17|Иисус, уразумев, говорит им: что рассуждаете о том, что нет у вас хлебов? Еще ли не понимаете и не разумеете? Еще ли окаменено у вас сердце?
MARK|8|18|Имея очи, не видите? имея уши, не слышите? и не помните?
MARK|8|19|Когда Я пять хлебов преломил для пяти тысяч [человек], сколько полных коробов набрали вы кусков? Говорят Ему: двенадцать.
MARK|8|20|А когда семь для четырех тысяч, сколько корзин набрали вы оставшихся кусков. Сказали: семь.
MARK|8|21|И сказал им: как же не разумеете?
MARK|8|22|Приходит в Вифсаиду; и приводят к Нему слепого и просят, чтобы прикоснулся к нему.
MARK|8|23|Он, взяв слепого за руку, вывел его вон из селения и, плюнув ему на глаза, возложил на него руки и спросил его: видит ли что?
MARK|8|24|Он, взглянув, сказал: вижу проходящих людей, как деревья.
MARK|8|25|Потом опять возложил руки на глаза ему и велел ему взглянуть. И он исцелел и стал видеть все ясно.
MARK|8|26|И послал его домой, сказав: не заходи в селение и не рассказывай никому в селении.
MARK|8|27|И пошел Иисус с учениками Своими в селения Кесарии Филипповой. Дорогою Он спрашивал учеников Своих: за кого почитают Меня люди?
MARK|8|28|Они отвечали: за Иоанна Крестителя; другие же – за Илию; а иные – за одного из пророков.
MARK|8|29|Он говорит им: а вы за кого почитаете Меня? Петр сказал Ему в ответ: Ты Христос.
MARK|8|30|И запретил им, чтобы никому не говорили о Нем.
MARK|8|31|И начал учить их, что Сыну Человеческому много должно пострадать, быть отвержену старейшинами, первосвященниками и книжниками, и быть убиту, и в третий день воскреснуть.
MARK|8|32|И говорил о сем открыто. Но Петр, отозвав Его, начал прекословить Ему.
MARK|8|33|Он же, обратившись и взглянув на учеников Своих, воспретил Петру, сказав: отойди от Меня, сатана, потому что ты думаешь не о том, что Божие, но что человеческое.
MARK|8|34|И, подозвав народ с учениками Своими, сказал им: кто хочет идти за Мною, отвергнись себя, и возьми крест свой, и следуй за Мною.
MARK|8|35|Ибо кто хочет душу свою сберечь, тот потеряет ее, а кто потеряет душу свою ради Меня и Евангелия, тот сбережет ее.
MARK|8|36|Ибо какая польза человеку, если он приобретет весь мир, а душе своей повредит?
MARK|8|37|Или какой выкуп даст человек за душу свою?
MARK|8|38|Ибо кто постыдится Меня и Моих слов в роде сем прелюбодейном и грешном, того постыдится и Сын Человеческий, когда приидет в славе Отца Своего со святыми Ангелами.
MARK|9|1|И сказал им: истинно говорю вам: есть некоторые из стоящих здесь, которые не вкусят смерти, как уже увидят Царствие Божие, пришедшее в силе.
MARK|9|2|И, по прошествии дней шести, взял Иисус Петра, Иакова и Иоанна, и возвел на гору высокую особо их одних, и преобразился перед ними.
MARK|9|3|Одежды Его сделались блистающими, весьма белыми, как снег, как на земле белильщик не может выбелить.
MARK|9|4|И явился им Илия с Моисеем; и беседовали с Иисусом.
MARK|9|5|При сем Петр сказал Иисусу: Равви! хорошо нам здесь быть; сделаем три кущи: Тебе одну, Моисею одну, и одну Илии.
MARK|9|6|Ибо не знал, что сказать; потому что они были в страхе.
MARK|9|7|И явилось облако, осеняющее их, и из облака исшел глас, глаголющий: Сей есть Сын Мой возлюбленный; Его слушайте.
MARK|9|8|И, внезапно посмотрев вокруг, никого более с собою не видели, кроме одного Иисуса.
MARK|9|9|Когда же сходили они с горы, Он не велел никому рассказывать о том, что видели, доколе Сын Человеческий не воскреснет из мертвых.
MARK|9|10|И они удержали это слово, спрашивая друг друга, что значит: воскреснуть из мертвых.
MARK|9|11|И спросили Его: как же книжники говорят, что Илии надлежит придти прежде?
MARK|9|12|Он сказал им в ответ: правда, Илия должен придти прежде и устроить все; и Сыну Человеческому, как написано о Нем, [надлежит] много пострадать и быть уничижену.
MARK|9|13|Но говорю вам, что и Илия пришел, и поступили с ним, как хотели, как написано о нем.
MARK|9|14|Придя к ученикам, увидел много народа около них и книжников, спорящих с ними.
MARK|9|15|Тотчас, увидев Его, весь народ изумился, и, подбегая, приветствовали Его.
MARK|9|16|Он спросил книжников: о чем спорите с ними?
MARK|9|17|Один из народа сказал в ответ: Учитель! я привел к Тебе сына моего, одержимого духом немым:
MARK|9|18|где ни схватывает его, повергает его на землю, и он испускает пену, и скрежещет зубами своими, и цепенеет. Говорил я ученикам Твоим, чтобы изгнали его, и они не могли.
MARK|9|19|Отвечая ему, Иисус сказал: о, род неверный! доколе буду с вами? доколе буду терпеть вас? Приведите его ко Мне.
MARK|9|20|И привели его к Нему. Как скоро [бесноватый] увидел Его, дух сотряс его; он упал на землю и валялся, испуская пену.
MARK|9|21|И спросил [Иисус] отца его: как давно это сделалось с ним? Он сказал: с детства;
MARK|9|22|и многократно [дух] бросал его и в огонь и в воду, чтобы погубить его; но, если что можешь, сжалься над нами и помоги нам.
MARK|9|23|Иисус сказал ему: если сколько–нибудь можешь веровать, все возможно верующему.
MARK|9|24|И тотчас отец отрока воскликнул со слезами: верую, Господи! помоги моему неверию.
MARK|9|25|Иисус, видя, что сбегается народ, запретил духу нечистому, сказав ему: дух немой и глухой! Я повелеваю тебе, выйди из него и впредь не входи в него.
MARK|9|26|И, вскрикнув и сильно сотрясши его, вышел; и он сделался, как мертвый, так что многие говорили, что он умер.
MARK|9|27|Но Иисус, взяв его за руку, поднял его; и он встал.
MARK|9|28|И как вошел [Иисус] в дом, ученики Его спрашивали Его наедине: почему мы не могли изгнать его?
MARK|9|29|И сказал им: сей род не может выйти иначе, как от молитвы и поста.
MARK|9|30|Выйдя оттуда, проходили через Галилею; и Он не хотел, чтобы кто узнал.
MARK|9|31|Ибо учил Своих учеников и говорил им, что Сын Человеческий предан будет в руки человеческие и убьют Его, и, по убиении, в третий день воскреснет.
MARK|9|32|Но они не разумели сих слов, а спросить Его боялись.
MARK|9|33|Пришел в Капернаум; и когда был в доме, спросил их: о чем дорогою вы рассуждали между собою?
MARK|9|34|Они молчали; потому что дорогою рассуждали между собою, кто больше.
MARK|9|35|И, сев, призвал двенадцать и сказал им: кто хочет быть первым, будь из всех последним и всем слугою.
MARK|9|36|И, взяв дитя, поставил его посреди них и, обняв его, сказал им:
MARK|9|37|кто примет одно из таких детей во имя Мое, тот принимает Меня; а кто Меня примет, тот не Меня принимает, но Пославшего Меня.
MARK|9|38|При сем Иоанн сказал: Учитель! мы видели человека, который именем Твоим изгоняет бесов, а не ходит за нами; и запретили ему, потому что не ходит за нами.
MARK|9|39|Иисус сказал: не запрещайте ему, ибо никто, сотворивший чудо именем Моим, не может вскоре злословить Меня.
MARK|9|40|Ибо кто не против вас, тот за вас.
MARK|9|41|И кто напоит вас чашею воды во имя Мое, потому что вы Христовы, истинно говорю вам, не потеряет награды своей.
MARK|9|42|А кто соблазнит одного из малых сих, верующих в Меня, тому лучше было бы, если бы повесили ему жерновный камень на шею и бросили его в море.
MARK|9|43|И если соблазняет тебя рука твоя, отсеки ее: лучше тебе увечному войти в жизнь, нежели с двумя руками идти в геенну, в огонь неугасимый,
MARK|9|44|где червь их не умирает и огонь не угасает.
MARK|9|45|И если нога твоя соблазняет тебя, отсеки ее: лучше тебе войти в жизнь хромому, нежели с двумя ногами быть ввержену в геенну, в огонь неугасимый,
MARK|9|46|где червь их не умирает и огонь не угасает.
MARK|9|47|И если глаз твой соблазняет тебя, вырви его: лучше тебе с одним глазом войти в Царствие Божие, нежели с двумя глазами быть ввержену в геенну огненную,
MARK|9|48|где червь их не умирает и огонь не угасает.
MARK|9|49|Ибо всякий огнем осолится, и всякая жертва солью осолится.
MARK|9|50|Соль – добрая [вещь]; но ежели соль не солона будет, чем вы ее поправите? Имейте в себе соль, и мир имейте между собою.
MARK|10|1|Отправившись оттуда, приходит в пределы Иудейские за Иорданскою стороною. Опять собирается к Нему народ, и, по обычаю Своему, Он опять учил их.
MARK|10|2|Подошли фарисеи и спросили, искушая Его: позволительно ли разводиться мужу с женою?
MARK|10|3|Он сказал им в ответ: что заповедал вам Моисей?
MARK|10|4|Они сказали: Моисей позволил писать разводное письмо и разводиться.
MARK|10|5|Иисус сказал им в ответ: по жестокосердию вашему он написал вам сию заповедь.
MARK|10|6|В начале же создания, Бог мужчину и женщину сотворил их.
MARK|10|7|Посему оставит человек отца своего и мать
MARK|10|8|и прилепится к жене своей, и будут два одною плотью; так что они уже не двое, но одна плоть.
MARK|10|9|Итак, что Бог сочетал, того человек да не разлучает.
MARK|10|10|В доме ученики Его опять спросили Его о том же.
MARK|10|11|Он сказал им: кто разведется с женою своею и женится на другой, тот прелюбодействует от нее;
MARK|10|12|и если жена разведется с мужем своим и выйдет за другого, прелюбодействует.
MARK|10|13|Приносили к Нему детей, чтобы Он прикоснулся к ним; ученики же не допускали приносящих.
MARK|10|14|Увидев [то], Иисус вознегодовал и сказал им: пустите детей приходить ко Мне и не препятствуйте им, ибо таковых есть Царствие Божие.
MARK|10|15|Истинно говорю вам: кто не примет Царствия Божия, как дитя, тот не войдет в него.
MARK|10|16|И, обняв их, возложил руки на них и благословил их.
MARK|10|17|Когда выходил Он в путь, подбежал некто, пал пред Ним на колени и спросил Его: Учитель благий! что мне делать, чтобы наследовать жизнь вечную?
MARK|10|18|Иисус сказал ему: что ты называешь Меня благим? Никто не благ, как только один Бог.
MARK|10|19|Знаешь заповеди: не прелюбодействуй, не убивай, не кради, не лжесвидетельствуй, не обижай, почитай отца твоего и мать.
MARK|10|20|Он же сказал Ему в ответ: Учитель! все это сохранил я от юности моей.
MARK|10|21|Иисус, взглянув на него, полюбил его и сказал ему: одного тебе недостает: пойди, все, что имеешь, продай и раздай нищим, и будешь иметь сокровище на небесах; и приходи, последуй за Мною, взяв крест.
MARK|10|22|Он же, смутившись от сего слова, отошел с печалью, потому что у него было большое имение.
MARK|10|23|И, посмотрев вокруг, Иисус говорит ученикам Своим: как трудно имеющим богатство войти в Царствие Божие!
MARK|10|24|Ученики ужаснулись от слов Его. Но Иисус опять говорит им в ответ: дети! как трудно надеющимся на богатство войти в Царствие Божие!
MARK|10|25|Удобнее верблюду пройти сквозь игольные уши, нежели богатому войти в Царствие Божие.
MARK|10|26|Они же чрезвычайно изумлялись и говорили между собою: кто же может спастись?
MARK|10|27|Иисус, воззрев на них, говорит: человекам это невозможно, но не Богу, ибо все возможно Богу.
MARK|10|28|И начал Петр говорить Ему: вот, мы оставили все и последовали за Тобою.
MARK|10|29|Иисус сказал в ответ: истинно говорю вам: нет никого, кто оставил бы дом, или братьев, или сестер, или отца, или мать, или жену, или детей, или земли, ради Меня и Евангелия,
MARK|10|30|и не получил бы ныне, во время сие, среди гонений, во сто крат более домов, и братьев и сестер, и отцов, и матерей, и детей, и земель, а в веке грядущем жизни вечной.
MARK|10|31|Многие же будут первые последними, и последние первыми.
MARK|10|32|Когда были они на пути, восходя в Иерусалим, Иисус шел впереди их, а они ужасались и, следуя за Ним, были в страхе. Подозвав двенадцать, Он опять начал им говорить о том, что будет с Ним:
MARK|10|33|вот, мы восходим в Иерусалим, и Сын Человеческий предан будет первосвященникам и книжникам, и осудят Его на смерть, и предадут Его язычникам,
MARK|10|34|и поругаются над Ним, и будут бить Его, и оплюют Его, и убьют Его; и в третий день воскреснет.
MARK|10|35|[Тогда] подошли к Нему сыновья Зеведеевы Иаков и Иоанн и сказали: Учитель! мы желаем, чтобы Ты сделал нам, о чем попросим.
MARK|10|36|Он сказал им: что хотите, чтобы Я сделал вам?
MARK|10|37|Они сказали Ему: дай нам сесть у Тебя, одному по правую сторону, а другому по левую в славе Твоей.
MARK|10|38|Но Иисус сказал им: не знаете, чего просите. Можете ли пить чашу, которую Я пью, и креститься крещением, которым Я крещусь?
MARK|10|39|Они отвечали: можем. Иисус же сказал им: чашу, которую Я пью, будете пить, и крещением, которым Я крещусь, будете креститься;
MARK|10|40|а дать сесть у Меня по правую сторону и по левую – не от Меня [зависит], но кому уготовано.
MARK|10|41|И, услышав, десять начали негодовать на Иакова и Иоанна.
MARK|10|42|Иисус же, подозвав их, сказал им: вы знаете, что почитающиеся князьями народов господствуют над ними, и вельможи их властвуют ими.
MARK|10|43|Но между вами да не будет так: а кто хочет быть большим между вами, да будем вам слугою;
MARK|10|44|и кто хочет быть первым между вами, да будет всем рабом.
MARK|10|45|Ибо и Сын Человеческий не для того пришел, чтобы Ему служили, но чтобы послужить и отдать душу Свою для искупления многих.
MARK|10|46|Приходят в Иерихон. И когда выходил Он из Иерихона с учениками Своими и множеством народа, Вартимей, сын Тимеев, слепой сидел у дороги, прося [милостыни].
MARK|10|47|Услышав, что это Иисус Назорей, он начал кричать и говорить: Иисус, Сын Давидов! помилуй меня.
MARK|10|48|Многие заставляли его молчать; но он еще более стал кричать: Сын Давидов! помилуй меня.
MARK|10|49|Иисус остановился и велел его позвать. Зовут слепого и говорят ему: не бойся, вставай, зовет тебя.
MARK|10|50|Он сбросил с себя верхнюю одежду, встал и пришел к Иисусу.
MARK|10|51|Отвечая ему, Иисус спросил: чего ты хочешь от Меня? Слепой сказал Ему: Учитель! чтобы мне прозреть.
MARK|10|52|Иисус сказал ему: иди, вера твоя спасла тебя. И он тотчас прозрел и пошел за Иисусом по дороге.
MARK|11|1|Когда приблизились к Иерусалиму, к Виффагии и Вифании, к горе Елеонской, [Иисус] посылает двух из учеников Своих
MARK|11|2|и говорит им: пойдите в селение, которое прямо перед вами; входя в него, тотчас найдете привязанного молодого осла, на которого никто из людей не садился; отвязав его, приведите.
MARK|11|3|И если кто скажет вам: что вы это делаете? – отвечайте, что он надобен Господу; и тотчас пошлет его сюда.
MARK|11|4|Они пошли, и нашли молодого осла, привязанного у ворот на улице, и отвязали его.
MARK|11|5|И некоторые из стоявших там говорили им: что делаете? [зачем] отвязываете осленка?
MARK|11|6|Они отвечали им, как повелел Иисус; и те отпустили их.
MARK|11|7|И привели осленка к Иисусу, и возложили на него одежды свои; [Иисус] сел на него.
MARK|11|8|Многие же постилали одежды свои по дороге; а другие резали ветви с дерев и постилали по дороге.
MARK|11|9|И предшествовавшие и сопровождавшие восклицали: осанна! благословен Грядущий во имя Господне!
MARK|11|10|благословенно грядущее во имя Господа царство отца нашего Давида! осанна в вышних!
MARK|11|11|И вошел Иисус в Иерусалим и в храм; и, осмотрев все, как время уже было позднее, вышел в Вифанию с двенадцатью.
MARK|11|12|На другой день, когда они вышли из Вифании, Он взалкал;
MARK|11|13|и, увидев издалека смоковницу, покрытую листьями, пошел, не найдет ли чего на ней; но, придя к ней, ничего не нашел, кроме листьев, ибо еще не время было [собирания] смокв.
MARK|11|14|И сказал ей Иисус: отныне да не вкушает никто от тебя плода вовек! И слышали то ученики Его.
MARK|11|15|Пришли в Иерусалим. Иисус, войдя в храм, начал выгонять продающих и покупающих в храме; и столы меновщиков и скамьи продающих голубей опрокинул;
MARK|11|16|и не позволял, чтобы кто пронес через храм какую–либо вещь.
MARK|11|17|И учил их, говоря: не написано ли: дом Мой домом молитвы наречется для всех народов? а вы сделали его вертепом разбойников.
MARK|11|18|Услышали [это] книжники и первосвященники, и искали, как бы погубить Его, ибо боялись Его, потому что весь народ удивлялся учению Его.
MARK|11|19|Когда же стало поздно, Он вышел вон из города.
MARK|11|20|Поутру, проходя мимо, увидели, что смоковница засохла до корня.
MARK|11|21|И, вспомнив, Петр говорит Ему: Равви! посмотри, смоковница, которую Ты проклял, засохла.
MARK|11|22|Иисус, отвечая, говорит им:
MARK|11|23|имейте веру Божию, ибо истинно говорю вам, если кто скажет горе сей: поднимись и ввергнись в море, и не усомнится в сердце своем, но поверит, что сбудется по словам его, – будет ему, что ни скажет.
MARK|11|24|Потому говорю вам: все, чего ни будете просить в молитве, верьте, что получите, – и будет вам.
MARK|11|25|И когда стоите на молитве, прощайте, если что имеете на кого, дабы и Отец ваш Небесный простил вам согрешения ваши.
MARK|11|26|Если же не прощаете, то и Отец ваш Небесный не простит вам согрешений ваших.
MARK|11|27|Пришли опять в Иерусалим. И когда Он ходил в храме, подошли к Нему первосвященники и книжники, и старейшины
MARK|11|28|и говорили Ему: какою властью Ты это делаешь? и кто Тебе дал власть делать это?
MARK|11|29|Иисус сказал им в ответ: спрошу и Я вас об одном, отвечайте Мне; [тогда] и Я скажу вам, какою властью это делаю.
MARK|11|30|Крещение Иоанново с небес было, или от человеков? отвечайте Мне.
MARK|11|31|Они рассуждали между собою: если скажем: с небес, – то Он скажет: почему же вы не поверили ему?
MARK|11|32|а сказать: от человеков – боялись народа, потому что все полагали, что Иоанн точно был пророк.
MARK|11|33|И сказали в ответ Иисусу: не знаем. Тогда Иисус сказал им в ответ: и Я не скажу вам, какою властью это делаю.
MARK|12|1|И начал говорить им притчами: некоторый человек насадил виноградник и обнес оградою, и выкопал точило, и построил башню, и, отдав его виноградарям, отлучился.
MARK|12|2|И послал в свое время к виноградарям слугу – принять от виноградарей плодов из виноградника.
MARK|12|3|Они же, схватив его, били, и отослали ни с чем.
MARK|12|4|Опять послал к ним другого слугу; и тому камнями разбили голову и отпустили его с бесчестьем.
MARK|12|5|И опять иного послал: и того убили; и многих других то били, то убивали.
MARK|12|6|Имея же еще одного сына, любезного ему, напоследок послал и его к ним, говоря: постыдятся сына моего.
MARK|12|7|Но виноградари сказали друг другу: это наследник; пойдем, убьем его, и наследство будет наше.
MARK|12|8|И, схватив его, убили и выбросили вон из виноградника.
MARK|12|9|Что же сделает хозяин виноградника? – Придет и предаст смерти виноградарей, и отдаст виноградник другим.
MARK|12|10|Неужели вы не читали сего в Писании: камень, который отвергли строители, тот самый сделался главою угла;
MARK|12|11|это от Господа, и есть дивно в очах наших.
MARK|12|12|И старались схватить Его, но побоялись народа, ибо поняли, что о них сказал притчу; и, оставив Его, отошли.
MARK|12|13|И посылают к Нему некоторых из фарисеев и иродиан, чтобы уловить Его в слове.
MARK|12|14|Они же, придя, говорят Ему: Учитель! мы знаем, что Ты справедлив и не заботишься об угождении кому–либо, ибо не смотришь ни на какое лице, но истинно пути Божию учишь. Позволительно ли давать подать кесарю или нет? давать ли нам или не давать?
MARK|12|15|Но Он, зная их лицемерие, сказал им: что искушаете Меня? принесите Мне динарий, чтобы Мне видеть его.
MARK|12|16|Они принесли. Тогда говорит им: чье это изображение и надпись? Они сказали Ему: кесаревы.
MARK|12|17|Иисус сказал им в ответ: отдавайте кесарево кесарю, а Божие Богу. И дивились Ему.
MARK|12|18|Потом пришли к Нему саддукеи, которые говорят, что нет воскресения, и спросили Его, говоря:
MARK|12|19|Учитель! Моисей написал нам: если у кого умрет брат и оставит жену, а детей не оставит, то брат его пусть возьмет жену его и восстановит семя брату своему.
MARK|12|20|Было семь братьев: первый взял жену и, умирая, не оставил детей.
MARK|12|21|Взял ее второй и умер, и он не оставил детей; также и третий.
MARK|12|22|Брали ее [за себя] семеро и не оставили детей. После всех умерла и жена.
MARK|12|23|Итак, в воскресении, когда воскреснут, которого из них будет она женою? Ибо семеро имели ее женою?
MARK|12|24|Иисус сказал им в ответ: этим ли приводитесь вы в заблуждение, не зная Писаний, ни силы Божией?
MARK|12|25|Ибо, когда из мертвых воскреснут, [тогда] не будут ни жениться, ни замуж выходить, но будут, как Ангелы на небесах.
MARK|12|26|А о мертвых, что они воскреснут, разве не читали вы в книге Моисея, как Бог при купине сказал ему: Я Бог Авраама, и Бог Исаака, и Бог Иакова?
MARK|12|27|[Бог] не есть Бог мертвых, но Бог живых. Итак, вы весьма заблуждаетесь.
MARK|12|28|Один из книжников, слыша их прения и видя, что [Иисус] хорошо им отвечал, подошел и спросил Его: какая первая из всех заповедей?
MARK|12|29|Иисус отвечал ему: первая из всех заповедей: слушай, Израиль! Господь Бог наш есть Господь единый;
MARK|12|30|и возлюби Господа Бога твоего всем сердцем твоим, и всею душею твоею, и всем разумением твоим, и всею крепостию твоею, – вот первая заповедь!
MARK|12|31|Вторая подобная ей: возлюби ближнего твоего, как самого себя. Иной большей сих заповеди нет.
MARK|12|32|Книжник сказал Ему: хорошо, Учитель! истину сказал Ты, что один есть Бог и нет иного, кроме Его;
MARK|12|33|и любить Его всем сердцем и всем умом, и всею душею, и всею крепостью, и любить ближнего, как самого себя, есть больше всех всесожжений и жертв.
MARK|12|34|Иисус, видя, что он разумно отвечал, сказал ему: недалеко ты от Царствия Божия. После того никто уже не смел спрашивать Его.
MARK|12|35|Продолжая учить в храме, Иисус говорил: как говорят книжники, что Христос есть Сын Давидов?
MARK|12|36|Ибо сам Давид сказал Духом Святым: сказал Господь Господу моему: седи одесную Меня, доколе положу врагов Твоих в подножие ног Твоих.
MARK|12|37|Итак, сам Давид называет Его Господом: как же Он Сын ему? И множество народа слушало Его с услаждением.
MARK|12|38|И говорил им в учении Своем: остерегайтесь книжников, любящих ходить в длинных одеждах и [принимать] приветствия в народных собраниях,
MARK|12|39|сидеть впереди в синагогах и возлежать на первом [месте] на пиршествах, –
MARK|12|40|сии, поядающие домы вдов и напоказ долго молящиеся, примут тягчайшее осуждение.
MARK|12|41|И сел Иисус против сокровищницы и смотрел, как народ кладет деньги в сокровищницу. Многие богатые клали много.
MARK|12|42|Придя же, одна бедная вдова положила две лепты, что составляет кодрант.
MARK|12|43|Подозвав учеников Своих, [Иисус] сказал им: истинно говорю вам, что эта бедная вдова положила больше всех, клавших в сокровищницу,
MARK|12|44|ибо все клали от избытка своего, а она от скудости своей положила все, что имела, все пропитание свое.
MARK|13|1|И когда выходил Он из храма, говорит Ему один из учеников его: Учитель! посмотри, какие камни и какие здания!
MARK|13|2|Иисус сказал ему в ответ: видишь сии великие здания? все это будет разрушено, так что не останется здесь камня на камне.
MARK|13|3|И когда Он сидел на горе Елеонской против храма, спрашивали Его наедине Петр, и Иаков, и Иоанн, и Андрей:
MARK|13|4|скажи нам, когда это будет, и какой признак, когда все сие должно совершиться?
MARK|13|5|Отвечая им, Иисус начал говорить: берегитесь, чтобы кто не прельстил вас,
MARK|13|6|ибо многие придут под именем Моим и будут говорить, что это Я; и многих прельстят.
MARK|13|7|Когда же услышите о войнах и о военных слухах, не ужасайтесь: ибо надлежит [сему] быть, – но [это] еще не конец.
MARK|13|8|Ибо восстанет народ на народ и царство на царство; и будут землетрясения по местам, и будут глады и смятения. Это – начало болезней.
MARK|13|9|Но вы смотрите за собою, ибо вас будут предавать в судилища и бить в синагогах, и перед правителями и царями поставят вас за Меня, для свидетельства перед ними.
MARK|13|10|И во всех народах прежде должно быть проповедано Евангелие.
MARK|13|11|Когда же поведут предавать вас, не заботьтесь наперед, что вам говорить, и не обдумывайте; но что дано будет вам в тот час, то и говорите, ибо не вы будете говорить, но Дух Святый.
MARK|13|12|Предаст же брат брата на смерть, и отец – детей; и восстанут дети на родителей и умертвят их.
MARK|13|13|И будете ненавидимы всеми за имя Мое; претерпевший же до конца спасется.
MARK|13|14|Когда же увидите мерзость запустения, реченную пророком Даниилом, стоящую, где не должно, – читающий да разумеет, – тогда находящиеся в Иудее да бегут в горы;
MARK|13|15|а кто на кровле, тот не сходи в дом и не входи взять что–нибудь из дома своего;
MARK|13|16|и кто на поле, не обращайся назад взять одежду свою.
MARK|13|17|Горе беременным и питающим сосцами в те дни.
MARK|13|18|Молитесь, чтобы не случилось бегство ваше зимою.
MARK|13|19|Ибо в те дни будет такая скорбь, какой не было от начала творения, которое сотворил Бог, даже доныне, и не будет.
MARK|13|20|И если бы Господь не сократил тех дней, то не спаслась бы никакая плоть; но ради избранных, которых Он избрал, сократил те дни.
MARK|13|21|Тогда, если кто вам скажет: вот, здесь Христос, или: вот, там, – не верьте.
MARK|13|22|Ибо восстанут лжехристы и лжепророки и дадут знамения и чудеса, чтобы прельстить, если возможно, и избранных.
MARK|13|23|Вы же берегитесь. Вот, Я наперед сказал вам все.
MARK|13|24|Но в те дни, после скорби той, солнце померкнет, и луна не даст света своего,
MARK|13|25|и звезды спадут с неба, и силы небесные поколеблются.
MARK|13|26|Тогда увидят Сына Человеческого, грядущего на облаках с силою многою и славою.
MARK|13|27|И тогда Он пошлет Ангелов Своих и соберет избранных Своих от четырех ветров, от края земли до края неба.
MARK|13|28|От смоковницы возьмите подобие: когда ветви ее становятся уже мягки и пускают листья, то знаете, что близко лето.
MARK|13|29|Так и когда вы увидите то сбывающимся, знайте, что близко, при дверях.
MARK|13|30|Истинно говорю вам: не прейдет род сей, как все это будет.
MARK|13|31|Небо и земля прейдут, но слова Мои не прейдут.
MARK|13|32|О дне же том, или часе, никто не знает, ни Ангелы небесные, ни Сын, но только Отец.
MARK|13|33|Смотрите, бодрствуйте, молитесь, ибо не знаете, когда наступит это время.
MARK|13|34|Подобно как бы кто, отходя в путь и оставляя дом свой, дал слугам своим власть и каждому свое дело, и приказал привратнику бодрствовать.
MARK|13|35|Итак бодрствуйте, ибо не знаете, когда придет хозяин дома: вечером, или в полночь, или в пение петухов, или поутру;
MARK|13|36|чтобы, придя внезапно, не нашел вас спящими.
MARK|13|37|А что вам говорю, говорю всем: бодрствуйте.
MARK|14|1|Через два дня [надлежало] быть [празднику] Пасхи и опресноков. И искали первосвященники и книжники, как бы взять Его хитростью и убить;
MARK|14|2|но говорили: [только] не в праздник, чтобы не произошло возмущения в народе.
MARK|14|3|И когда был Он в Вифании, в доме Симона прокаженного, и возлежал, – пришла женщина с алавастровым сосудом мира из нарда чистого, драгоценного и, разбив сосуд, возлила Ему на голову.
MARK|14|4|Некоторые же вознегодовали и говорили между собою: к чему сия трата мира?
MARK|14|5|Ибо можно было бы продать его более нежели за триста динариев и раздать нищим. И роптали на нее.
MARK|14|6|Но Иисус сказал: оставьте ее; что ее смущаете? Она доброе дело сделала для Меня.
MARK|14|7|Ибо нищих всегда имеете с собою и, когда захотите, можете им благотворить; а Меня не всегда имеете.
MARK|14|8|Она сделала, что могла: предварила помазать тело Мое к погребению.
MARK|14|9|Истинно говорю вам: где ни будет проповедано Евангелие сие в целом мире, сказано будет, в память ее, и о том, что она сделала.
MARK|14|10|И пошел Иуда Искариот, один из двенадцати, к первосвященникам, чтобы предать Его им.
MARK|14|11|Они же, услышав, обрадовались, и обещали дать ему сребренники. И он искал, как бы в удобное время предать Его.
MARK|14|12|В первый день опресноков, когда заколали пасхального [агнца], говорят Ему ученики Его: где хочешь есть пасху? мы пойдем и приготовим.
MARK|14|13|И посылает двух из учеников Своих и говорит им: пойдите в город; и встретится вам человек, несущий кувшин воды; последуйте за ним
MARK|14|14|и куда он войдет, скажите хозяину дома того: Учитель говорит: где комната, в которой бы Мне есть пасху с учениками Моими?
MARK|14|15|И он покажет вам горницу большую, устланную, готовую: там приготовьте нам.
MARK|14|16|И пошли ученики Его, и пришли в город, и нашли, как сказал им; и приготовили пасху.
MARK|14|17|Когда настал вечер, Он приходит с двенадцатью.
MARK|14|18|И, когда они возлежали и ели, Иисус сказал: истинно говорю вам, один из вас, ядущий со Мною, предаст Меня.
MARK|14|19|Они опечалились и стали говорить Ему, один за другим: не я ли? и другой: не я ли?
MARK|14|20|Он же сказал им в ответ: один из двенадцати, обмакивающий со Мною в блюдо.
MARK|14|21|Впрочем Сын Человеческий идет, как писано о Нем; но горе тому человеку, которым Сын Человеческий предается: лучше было бы тому человеку не родиться.
MARK|14|22|И когда они ели, Иисус, взяв хлеб, благословил, преломил, дал им и сказал: приимите, ядите; сие есть Тело Мое.
MARK|14|23|И, взяв чашу, благодарив, подал им: и пили из нее все.
MARK|14|24|И сказал им: сие есть Кровь Моя Нового Завета, за многих изливаемая.
MARK|14|25|Истинно говорю вам: Я уже не буду пить от плода виноградного до того дня, когда буду пить новое вино в Царствии Божием.
MARK|14|26|И, воспев, пошли на гору Елеонскую.
MARK|14|27|И говорит им Иисус: все вы соблазнитесь о Мне в эту ночь; ибо написано: поражу пастыря, и рассеются овцы.
MARK|14|28|По воскресении же Моем, Я предваряю вас в Галилее.
MARK|14|29|Петр сказал Ему: если и все соблазнятся, но не я.
MARK|14|30|И говорит ему Иисус: истинно говорю тебе, что ты ныне, в эту ночь, прежде нежели дважды пропоет петух, трижды отречешься от Меня.
MARK|14|31|Но он еще с большим усилием говорил: хотя бы мне надлежало и умереть с Тобою, не отрекусь от Тебя. То же и все говорили.
MARK|14|32|Пришли в селение, называемое Гефсимания; и Он сказал ученикам Своим: посидите здесь, пока Я помолюсь.
MARK|14|33|И взял с Собою Петра, Иакова и Иоанна; и начал ужасаться и тосковать.
MARK|14|34|И сказал им: душа Моя скорбит смертельно; побудьте здесь и бодрствуйте.
MARK|14|35|И, отойдя немного, пал на землю и молился, чтобы, если возможно, миновал Его час сей;
MARK|14|36|и говорил: Авва Отче! все возможно Тебе; пронеси чашу сию мимо Меня; но не чего Я хочу, а чего Ты.
MARK|14|37|Возвращается и находит их спящими, и говорит Петру: Симон! ты спишь? не мог ты бодрствовать один час?
MARK|14|38|Бодрствуйте и молитесь, чтобы не впасть в искушение: дух бодр, плоть же немощна.
MARK|14|39|И, опять отойдя, молился, сказав то же слово.
MARK|14|40|И, возвратившись, опять нашел их спящими, ибо глаза у них отяжелели, и они не знали, что Ему отвечать.
MARK|14|41|И приходит в третий раз и говорит им: вы все еще спите и почиваете? Кончено, пришел час: вот, предается Сын Человеческий в руки грешников.
MARK|14|42|Встаньте, пойдем; вот, приблизился предающий Меня.
MARK|14|43|И тотчас, как Он еще говорил, приходит Иуда, один из двенадцати, и с ним множество народа с мечами и кольями, от первосвященников и книжников и старейшин.
MARK|14|44|Предающий же Его дал им знак, сказав: Кого я поцелую, Тот и есть, возьмите Его и ведите осторожно.
MARK|14|45|И, придя, тотчас подошел к Нему и говорит: Равви! Равви! и поцеловал Его.
MARK|14|46|А они возложили на Него руки свои и взяли Его.
MARK|14|47|Один же из стоявших тут извлек меч, ударил раба первосвященникова и отсек ему ухо.
MARK|14|48|Тогда Иисус сказал им: как будто на разбойника вышли вы с мечами и кольями, чтобы взять Меня.
MARK|14|49|Каждый день бывал Я с вами в храме и учил, и вы не брали Меня. Но да сбудутся Писания.
MARK|14|50|Тогда, оставив Его, все бежали.
MARK|14|51|Один юноша, завернувшись по нагому телу в покрывало, следовал за Ним; и воины схватили его.
MARK|14|52|Но он, оставив покрывало, нагой убежал от них.
MARK|14|53|И привели Иисуса к первосвященнику; и собрались к нему все первосвященники и старейшины и книжники.
MARK|14|54|Петр издали следовал за Ним, даже внутрь двора первосвященникова; и сидел со служителями, и грелся у огня.
MARK|14|55|Первосвященники же и весь синедрион искали свидетельства на Иисуса, чтобы предать Его смерти; и не находили.
MARK|14|56|Ибо многие лжесвидетельствовали на Него, но свидетельства сии не были достаточны.
MARK|14|57|И некоторые, встав, лжесвидетельствовали против Него и говорили:
MARK|14|58|мы слышали, как Он говорил: Я разрушу храм сей рукотворенный, и через три дня воздвигну другой, нерукотворенный.
MARK|14|59|Но и такое свидетельство их не было достаточно.
MARK|14|60|Тогда первосвященник стал посреди и спросил Иисуса: что Ты ничего не отвечаешь? что они против Тебя свидетельствуют?
MARK|14|61|Но Он молчал и не отвечал ничего. Опять первосвященник спросил Его и сказал Ему: Ты ли Христос, Сын Благословенного?
MARK|14|62|Иисус сказал: Я; и вы узрите Сына Человеческого, сидящего одесную силы и грядущего на облаках небесных.
MARK|14|63|Тогда первосвященник, разодрав одежды свои, сказал: на что еще нам свидетелей?
MARK|14|64|Вы слышали богохульство; как вам кажется? Они же все признали Его повинным смерти.
MARK|14|65|И некоторые начали плевать на Него и, закрывая Ему лице, ударять Его и говорить Ему: прореки. И слуги били Его по ланитам.
MARK|14|66|Когда Петр был на дворе внизу, пришла одна из служанок первосвященника
MARK|14|67|и, увидев Петра греющегося и всмотревшись в него, сказала: и ты был с Иисусом Назарянином.
MARK|14|68|Но он отрекся, сказав: не знаю и не понимаю, что ты говоришь. И вышел вон на передний двор; и запел петух.
MARK|14|69|Служанка, увидев его опять, начала говорить стоявшим тут: этот из них.
MARK|14|70|Он опять отрекся. Спустя немного, стоявшие тут опять стали говорить Петру: точно ты из них; ибо ты Галилеянин, и наречие твое сходно.
MARK|14|71|Он же начал клясться и божиться: не знаю Человека Сего, о Котором говорите.
MARK|14|72|Тогда петух запел во второй раз. И вспомнил Петр слово, сказанное ему Иисусом: прежде нежели петух пропоет дважды, трижды отречешься от Меня; и начал плакать.
MARK|15|1|Немедленно поутру первосвященники со старейшинами и книжниками и весь синедрион составили совещание и, связав Иисуса, отвели и предали Пилату.
MARK|15|2|Пилат спросил Его: Ты Царь Иудейский? Он же сказал ему в ответ: ты говоришь.
MARK|15|3|И первосвященники обвиняли Его во многом.
MARK|15|4|Пилат же опять спросил Его: Ты ничего не отвечаешь? видишь, как много против Тебя обвинений.
MARK|15|5|Но Иисус и на это ничего не отвечал, так что Пилат дивился.
MARK|15|6|На всякий же праздник отпускал он им одного узника, о котором просили.
MARK|15|7|Тогда был в узах [некто], по имени Варавва, со своими сообщниками, которые во время мятежа сделали убийство.
MARK|15|8|И народ начал кричать и просить [Пилата] о том, что он всегда делал для них.
MARK|15|9|Он сказал им в ответ: хотите ли, отпущу вам Царя Иудейского?
MARK|15|10|Ибо знал, что первосвященники предали Его из зависти.
MARK|15|11|Но первосвященники возбудили народ [просить], чтобы отпустил им лучше Варавву.
MARK|15|12|Пилат, отвечая, опять сказал им: что же хотите, чтобы я сделал с Тем, Которого вы называете Царем Иудейским?
MARK|15|13|Они опять закричали: распни Его.
MARK|15|14|Пилат сказал им: какое же зло сделал Он? Но они еще сильнее закричали: распни Его.
MARK|15|15|Тогда Пилат, желая сделать угодное народу, отпустил им Варавву, а Иисуса, бив, предал на распятие.
MARK|15|16|А воины отвели Его внутрь двора, то есть в преторию, и собрали весь полк,
MARK|15|17|и одели Его в багряницу, и, сплетши терновый венец, возложили на Него;
MARK|15|18|и начали приветствовать Его: радуйся, Царь Иудейский!
MARK|15|19|И били Его по голове тростью, и плевали на Него, и, становясь на колени, кланялись Ему.
MARK|15|20|Когда же насмеялись над Ним, сняли с Него багряницу, одели Его в собственные одежды Его и повели Его, чтобы распять Его.
MARK|15|21|И заставили проходящего некоего Киринеянина Симона, отца Александрова и Руфова, идущего с поля, нести крест Его.
MARK|15|22|И привели Его на место Голгофу, что значит: Лобное место.
MARK|15|23|И давали Ему пить вино со смирною; но Он не принял.
MARK|15|24|Распявшие Его делили одежды Его, бросая жребий, кому что взять.
MARK|15|25|Был час третий, и распяли Его.
MARK|15|26|И была надпись вины Его: Царь Иудейский.
MARK|15|27|С Ним распяли двух разбойников, одного по правую, а другого по левую [сторону] Его.
MARK|15|28|И сбылось слово Писания: и к злодеям причтен.
MARK|15|29|Проходящие злословили Его, кивая головами своими и говоря: э! разрушающий храм, и в три дня созидающий!
MARK|15|30|спаси Себя Самого и сойди со креста.
MARK|15|31|Подобно и первосвященники с книжниками, насмехаясь, говорили друг другу: других спасал, а Себя не может спасти.
MARK|15|32|Христос, Царь Израилев, пусть сойдет теперь с креста, чтобы мы видели, и уверуем. И распятые с Ним поносили Его.
MARK|15|33|В шестом же часу настала тьма по всей земле и [продолжалась] до часа девятого.
MARK|15|34|В девятом часу возопил Иисус громким голосом: Элои! Элои! ламма савахфани? – что значит: Боже Мой! Боже Мой! для чего Ты Меня оставил?
MARK|15|35|Некоторые из стоявших тут, услышав, говорили: вот, Илию зовет.
MARK|15|36|А один побежал, наполнил губку уксусом и, наложив на трость, давал Ему пить, говоря: постойте, посмотрим, придет ли Илия снять Его.
MARK|15|37|Иисус же, возгласив громко, испустил дух.
MARK|15|38|И завеса в храме раздралась надвое, сверху донизу.
MARK|15|39|Сотник, стоявший напротив Его, увидев, что Он, так возгласив, испустил дух, сказал: истинно Человек Сей был Сын Божий.
MARK|15|40|Были [тут] и женщины, которые смотрели издали: между ними была и Мария Магдалина, и Мария, мать Иакова меньшего и Иосии, и Саломия,
MARK|15|41|которые и тогда, как Он был в Галилее, следовали за Ним и служили Ему, и другие многие, вместе с Ним пришедшие в Иерусалим.
MARK|15|42|И как уже настал вечер, – потому что была пятница, то есть [день] перед субботою, –
MARK|15|43|пришел Иосиф из Аримафеи, знаменитый член совета, который и сам ожидал Царствия Божия, осмелился войти к Пилату, и просил тела Иисусова.
MARK|15|44|Пилат удивился, что Он уже умер, и, призвав сотника, спросил его, давно ли умер?
MARK|15|45|И, узнав от сотника, отдал тело Иосифу.
MARK|15|46|Он, купив плащаницу и сняв Его, обвил плащаницею, и положил Его во гробе, который был высечен в скале, и привалил камень к двери гроба.
MARK|15|47|Мария же Магдалина и Мария Иосиева смотрели, где Его полагали.
MARK|16|1|По прошествии субботы Мария Магдалина и Мария Иаковлева и Саломия купили ароматы, чтобы идти помазать Его.
MARK|16|2|И весьма рано, в первый [день] недели, приходят ко гробу, при восходе солнца,
MARK|16|3|и говорят между собою: кто отвалит нам камень от двери гроба?
MARK|16|4|И, взглянув, видят, что камень отвален; а он был весьма велик.
MARK|16|5|И, войдя во гроб, увидели юношу, сидящего на правой стороне, облеченного в белую одежду; и ужаснулись.
MARK|16|6|Он же говорит им: не ужасайтесь. Иисуса ищете Назарянина, распятого; Он воскрес, Его нет здесь. Вот место, где Он был положен.
MARK|16|7|Но идите, скажите ученикам Его и Петру, что Он предваряет вас в Галилее; там Его увидите, как Он сказал вам.
MARK|16|8|И, выйдя, побежали от гроба; их объял трепет и ужас, и никому ничего не сказали, потому что боялись.
MARK|16|9|Воскреснув рано в первый [день] недели, [Иисус] явился сперва Марии Магдалине, из которой изгнал семь бесов.
MARK|16|10|Она пошла и возвестила бывшим с Ним, плачущим и рыдающим;
MARK|16|11|но они, услышав, что Он жив и она видела Его, – не поверили.
MARK|16|12|После сего явился в ином образе двум из них на дороге, когда они шли в селение.
MARK|16|13|И те, возвратившись, возвестили прочим; но и им не поверили.
MARK|16|14|Наконец, явился самим одиннадцати, возлежавшим [на вечери], и упрекал их за неверие и жестокосердие, что видевшим Его воскресшего не поверили.
MARK|16|15|И сказал им: идите по всему миру и проповедуйте Евангелие всей твари.
MARK|16|16|Кто будет веровать и креститься, спасен будет; а кто не будет веровать, осужден будет.
MARK|16|17|Уверовавших же будут сопровождать сии знамения: именем Моим будут изгонять бесов; будут говорить новыми языками;
MARK|16|18|будут брать змей; и если что смертоносное выпьют, не повредит им; возложат руки на больных, и они будут здоровы.
MARK|16|19|И так Господь, после беседования с ними, вознесся на небо и воссел одесную Бога.
MARK|16|20|А они пошли и проповедывали везде, при Господнем содействии и подкреплении слова последующими знамениями. Аминь.
