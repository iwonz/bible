1SAM|1|1|以法蓮 山區有一個 拉瑪 的 瑣非 人 ，名叫 以利加拿 ，他是 蘇弗 的玄孫， 託戶 的曾孫， 以利戶 的孫子， 耶羅罕 的兒子，是 以法蓮 人。
1SAM|1|2|他有兩個妻子：一個名叫 哈拿 ，另一個名叫 毗尼拿 。 毗尼拿 有孩子， 哈拿 卻沒有孩子。
1SAM|1|3|這人每年從本城上到 示羅 ，敬拜萬軍之耶和華，向他獻祭。在那裏有 以利 的兩個兒子 何弗尼 和 非尼哈 當耶和華的祭司。
1SAM|1|4|每逢獻祭的日子， 以利加拿 把祭肉分給他的妻子 毗尼拿 和 毗尼拿 所生的兒女。
1SAM|1|5|他給 哈拿 的卻是雙分，因為他愛 哈拿 。耶和華卻不使 哈拿 生育。
1SAM|1|6|她的對頭 毗尼拿 因耶和華不使 哈拿 生育，就常常惹她發怒，要使她生氣。
1SAM|1|7|年年都是如此。每當她上到耶和華殿的時候， 毗尼拿 就這樣惹她發怒，以致她哭泣不吃飯。
1SAM|1|8|她丈夫 以利加拿 對她說：「 哈拿 ，你為何哭泣？為何不吃飯？為何傷心難過呢？有我不比有十個兒子更好嗎？」
1SAM|1|9|他們在 示羅 吃喝完了， 哈拿 就站起來。祭司 以利 坐在耶和華殿門框旁邊的位子上。
1SAM|1|10|哈拿 心裏愁苦，就痛痛哭泣，向耶和華祈禱。
1SAM|1|11|她許願說：「萬軍之耶和華啊，你若垂顧你使女的苦情，眷念不忘你的使女，賜你的使女一個子嗣，我必使他終生歸給耶和華，不用剃刀剃他的頭。」
1SAM|1|12|哈拿 在耶和華面前不住地祈禱， 以利 注意她的嘴。
1SAM|1|13|哈拿 心中默禱，只動嘴唇，聽不到她的聲音，因此 以利 以為她喝醉了。
1SAM|1|14|以利 對她說：「你要醉到幾時呢？不要再喝酒了！」
1SAM|1|15|哈拿 回答說：「我主啊，不是這樣。我是心裏愁苦的婦人，清酒烈酒都沒有喝，只在耶和華面前傾心吐意。
1SAM|1|16|不要將你的使女看作不正經的女子。我因極其難過和生氣，所以一直禱告到如今。」
1SAM|1|17|以利 回答說：「平平安安地回去吧。願 以色列 的上帝允准你向他所求的！」
1SAM|1|18|哈拿 說：「願你的婢女在你眼前蒙恩。」於是婦人上路，去吃飯，臉上不再帶愁容了。
1SAM|1|19|他們清早起來，在耶和華面前敬拜，就回去，往 拉瑪 自己的家裏。 以利加拿 和妻子 哈拿 同房，耶和華顧念 哈拿 。
1SAM|1|20|時候到了， 哈拿 懷孕生了一個兒子， 哈拿 給他起名叫 撒母耳 ，說：「這是我從耶和華那裏求來的。」
1SAM|1|21|以利加拿 和他全家都上去，要向耶和華獻年祭和還願祭。
1SAM|1|22|哈拿 卻沒有上去，因為她對丈夫說：「等孩子斷了奶，我就帶他上去朝見耶和華，讓他永遠住在那裏。」
1SAM|1|23|她丈夫 以利加拿 對她說：「就照你看為好的去做吧！可以留到兒子斷了奶，願耶和華應驗他的話。」於是婦人留在家裏乳養兒子，直到斷了奶。
1SAM|1|24|斷奶之後，她就帶著孩子，連同一頭三歲的公牛 ，一伊法細麵 ，一皮袋酒，上 示羅 耶和華的殿去。那時，孩子還小。
1SAM|1|25|他們宰了公牛，就領孩子到 以利 面前。
1SAM|1|26|婦人說：「我主啊，請容許我說，我向你，我的主起誓，從前在你這裏站著祈求耶和華的那婦人就是我。
1SAM|1|27|我祈求為要得這孩子，耶和華已將我向他所求的賜給我了。
1SAM|1|28|所以，我將這孩子獻給耶和華，使他終生歸給耶和華。」 他就在那裏敬拜耶和華。
1SAM|2|1|哈拿 禱告說： 「我的心因耶和華快樂， 我的角因耶和華高舉。 我的口向仇敵張開； 我因你的救恩歡欣。
1SAM|2|2|「沒有一位聖者像耶和華， 除你以外沒有別的了， 也沒有磐石像我們的上帝。
1SAM|2|3|不要誇口說驕傲的話， 也不要口出狂妄的言語， 因耶和華是有知識的上帝， 人的行為被他衡量。
1SAM|2|4|勇士的弓折斷， 跌倒的人以力量束腰。
1SAM|2|5|飽足的人作雇工求食； 飢餓的人也不再飢餓。 不生育的生了七個； 兒女多的反倒孤獨。
1SAM|2|6|耶和華使人死，也使人活， 使人下陰間，也使人往上升。
1SAM|2|7|耶和華使人貧窮，也使人富足； 使人降卑，也使人升高。
1SAM|2|8|他從灰塵裏抬舉貧寒人， 從糞堆中提拔貧窮人， 使他們與貴族同坐， 繼承榮耀的座位。 地的柱子屬耶和華， 他將世界立在其上。
1SAM|2|9|「他必保護他聖民的腳步， 但惡人卻在黑暗中毀滅， 因為人不是靠力量得勝。
1SAM|2|10|與耶和華相爭的，必被打碎； 他必從天上打雷攻擊他們。 耶和華審判地極的人， 將力量賜給所立的王， 高舉受膏者的角。」
1SAM|2|11|以利加拿 往 拉瑪 回自己的家去了。那孩子在 以利 祭司面前事奉耶和華。
1SAM|2|12|以利 的兩個兒子是無賴，不認識耶和華。
1SAM|2|13|這二祭司對待百姓的規矩是這樣：凡有人獻祭，正煮肉的時候，祭司的僕人就手拿三齒的叉子來，
1SAM|2|14|將叉子往盆裏，或鍋裏，或釜裏，或壺裏一插，插上來的肉，祭司都拿了去。他們對所有上到 示羅 的 以色列 人都這樣做。
1SAM|2|15|甚至在未燒脂肪之前，祭司的僕人就來對獻祭的人說：「把肉給祭司，讓他烤吧。他不要拿你煮過的肉，要生的。」
1SAM|2|16|獻祭的人若說：「他們必須先燒脂肪，然後你才可以隨意拿。」僕人就說：「不，你立刻給我，不然我就要搶了。」
1SAM|2|17|這些年輕人的罪在耶和華面前非常嚴重，因為這些人藐視耶和華的祭物。
1SAM|2|18|那時， 撒母耳 還是孩子，穿著細麻布的以弗得，侍立在耶和華面前。
1SAM|2|19|他母親每年為他做一件小外袍，同丈夫上來獻年祭的時候帶來給他。
1SAM|2|20|以利 為 以利加拿 和他妻子祝福，說：「願耶和華由這婦人再賜你後裔，代替從耶和華求來的孩子。」他們就回自己的地方去了。
1SAM|2|21|耶和華眷顧 哈拿 ，她就懷孕生了三個兒子，兩個女兒。那孩子 撒母耳 在耶和華面前漸漸長大。
1SAM|2|22|以利 年紀老邁，聽見他兩個兒子對 以色列 眾人所做一切的事，又聽見他們與會幕門前伺候的婦人同寢，
1SAM|2|23|就對他們說：「你們為何做這樣的事呢？我從這眾百姓聽見了你們的惡行。
1SAM|2|24|我兒啊，不可這樣！我聽到耶和華的百姓傳出你們不好的名聲 。
1SAM|2|25|人若得罪人，有上帝 可以裁決；人若得罪耶和華，誰能為他代求呢？」然而他們還是不聽父親的話，因為耶和華想要他們死。
1SAM|2|26|撒母耳 這孩子漸漸長大，耶和華與人越發喜愛他。
1SAM|2|27|有神人來見 以利 ，對他說：「耶和華如此說：『你祖宗的家在 埃及 法老家 的時候，我不是向他們顯現嗎？
1SAM|2|28|在 以色列 眾支派中，我不是揀選他作我的祭司，上我的祭壇，燒香，在我面前穿以弗得嗎？我不是將 以色列 人所獻的火祭都賜給你祖宗的家嗎？
1SAM|2|29|你們為何踐踏我所吩咐獻在我居所的祭物和供物呢 ？你為何尊重你的兒子過於尊重我，將我百姓 以色列 所獻美好的祭物都拿去養肥你們自己呢？』
1SAM|2|30|因此，耶和華－ 以色列 的上帝說：『我確實說過，你和你祖宗的家必永遠行在我面前，但現在耶和華卻說，我絕不會這樣做。因為尊重我的，我必尊重他；藐視我的，他必被輕視。
1SAM|2|31|看哪，日子將到，我要折斷你的膀臂和你祖宗家的膀臂，使你家中沒有一個老年人。
1SAM|2|32|你在 以色列 人享福的時候必看見我居所的衰敗 ，你家中必永遠沒有一個老年人。
1SAM|2|33|你家中的人，我沒有從我壇前剪除的，必使你眼睛失明，心中憂傷。你家中所添的人口都必夭折。
1SAM|2|34|你的兩個兒子 何弗尼 、 非尼哈 所遭遇的事是給你的預兆：他們二人必在同一日死亡。
1SAM|2|35|我要為自己立一個忠心的祭司，他行事必照我的心、如我的意。我要為他建立堅固的家，他必天天行走在我受膏者的面前。
1SAM|2|36|你家所剩下的人都必來叩拜他，求一塊銀子，一個餅，說：求你給我一個祭司的職分，好使我得點餅吃。』」
1SAM|3|1|那孩子 撒母耳 在 以利 面前事奉耶和華。在那些日子，耶和華的言語稀少，不常有異象。
1SAM|3|2|那時， 以利 在自己的地方睡覺；他眼目開始昏花，不能看見。
1SAM|3|3|上帝的燈還沒有熄滅， 撒母耳 睡在耶和華的殿內，上帝的約櫃就在那裏。
1SAM|3|4|耶和華呼喚 撒母耳 ， 撒母耳 說：「我在這裏！」
1SAM|3|5|他跑到 以利 那裏，說：「你叫我嗎？我在這裏。」 以利 說：「我沒有叫你，回去睡吧。」他就回去睡了。
1SAM|3|6|耶和華又呼喚 撒母耳 。 撒母耳 起來，到 以利 那裏，說：「你叫我嗎？我在這裏。」 以利 說：「我兒，我沒有叫你，回去睡吧。」
1SAM|3|7|那時 撒母耳 還未認識耶和華，耶和華的話也未曾向他啟示。
1SAM|3|8|耶和華第三次再呼喚 撒母耳 。 撒母耳 起來，到 以利 那裏，說：「你叫我嗎？我在這裏。」 以利 才明白是耶和華呼喚這小孩。
1SAM|3|9|以利 對 撒母耳 說：「你回去睡吧。他若再叫你，你就說：『耶和華啊，請說，僕人敬聽！』」 撒母耳 就回去，仍睡在原處。
1SAM|3|10|耶和華來站著，像前幾次呼喚：「 撒母耳 ！ 撒母耳 ！」 撒母耳 說：「請說，僕人敬聽！」
1SAM|3|11|耶和華對 撒母耳 說：「看哪，我在 以色列 中必行一件事，凡聽見的人都必雙耳齊鳴。
1SAM|3|12|我指著 以利 家所說的話，到了時候，必從頭到尾應驗在 以利 身上。
1SAM|3|13|我曾告訴他，我必永遠懲罰他的家，因為他知道自己的兒子作惡，褻瀆上帝 ，卻不禁止他們。
1SAM|3|14|所以我向 以利 家起誓：『 以利 家的罪孽，就是獻祭物和供物，也永不得贖。』」
1SAM|3|15|撒母耳 睡到天亮，就開了耶和華殿的門。 撒母耳 害怕，不敢將異象告訴 以利 。
1SAM|3|16|以利 呼喚 撒母耳 說：「我兒 撒母耳 ！」 撒母耳 說：「我在這裏！」
1SAM|3|17|以利 說：「他對你說了甚麼話，你不要向我隱瞞。你若將他對你所說的話向我隱瞞一句，願上帝重重懲罰你。」
1SAM|3|18|撒母耳 就把一切話都告訴 以利 ，並沒有隱瞞。 以利 說：「他是耶和華，願他照他看為好的去做。」
1SAM|3|19|撒母耳 長大了，耶和華與他同在，使他所說的話一句都不落空。
1SAM|3|20|從 但 到 別是巴 ，所有的 以色列 人都知道耶和華立 撒母耳 為先知。
1SAM|3|21|耶和華又在 示羅 顯現，因為耶和華在 示羅 藉他的話向 撒母耳 啟示他自己。
1SAM|4|1|撒母耳 的話傳遍了全 以色列 。 以色列 人出去與 非利士 人打仗，安營在 以便‧以謝 ， 非利士 人安營在 亞弗 。
1SAM|4|2|非利士 人向 以色列 人擺陣。兩軍交戰的時候， 以色列 人敗在 非利士 人面前； 非利士 人在戰場上殺了他們約四千人。
1SAM|4|3|百姓回到營裏， 以色列 的長老說：「耶和華今日為何使我們敗在 非利士 人面前呢？我們要將耶和華的約櫃從 示羅 抬到我們這裏來，好讓他來到我們中間，救我們脫離敵人的手掌。」
1SAM|4|4|於是百姓派人到 示羅 ，從那裏將坐在二基路伯上萬軍之耶和華的約櫃抬來。 以利 的兩個兒子 何弗尼 、 非尼哈 也與上帝的約櫃同來。
1SAM|4|5|耶和華的約櫃到了營中，全 以色列 就大聲歡呼，連地都震動。
1SAM|4|6|非利士 人聽見歡呼的聲音，就說：「為何 希伯來 人在營裏這麼大聲歡呼呢？」他們知道耶和華的約櫃到了營中。
1SAM|4|7|非利士 人就懼怕，說：「有神明到了他們營中。」又說：「我們有禍了！從來不曾有這樣的事。
1SAM|4|8|我們有禍了！誰能救我們脫離這些大能之神明的手呢？從前在曠野用各樣災禍擊打 埃及 人的，就是這些神明。
1SAM|4|9|非利士 人哪，要剛強，要作大丈夫，免得作 希伯來 人的奴僕，如同他們作你們的奴僕一樣。你們要作大丈夫，與他們爭戰。」
1SAM|4|10|非利士 人進攻， 以色列 人敗了，各往自己的家逃跑。被殺的人很多， 以色列 倒下的步兵有三萬。
1SAM|4|11|上帝的約櫃被擄去， 以利 的兩個兒子 何弗尼 、 非尼哈 也都被殺了。
1SAM|4|12|有一個 便雅憫 人從戰場上逃跑，衣服撕裂，頭蒙灰塵，當日來到 示羅 。
1SAM|4|13|他到了的時候，看哪， 以利 正坐在路旁的位子上觀望，為上帝的約櫃心裏擔憂。那人進城報信，全城的人就都呼喊起來。
1SAM|4|14|以利 聽見呼喊的聲音就說：「這喧嚷的聲音是甚麼呢？」那人急忙來報信給 以利 。
1SAM|4|15|那時 以利 九十八歲了，兩眼發直，不能看見。
1SAM|4|16|那人對 以利 說：「我是從戰場上來的，今日剛從戰場上逃回來。」 以利 說：「我兒，事情怎樣了？」
1SAM|4|17|報信的回答說：「 以色列 人在 非利士 人面前逃跑，百姓中被殺的很多！你的兩個兒子 何弗尼 和 非尼哈 也都死了，並且上帝的約櫃已經被擄去了。」
1SAM|4|18|他一提到上帝的約櫃， 以利 就從城門旁自己的位子上往後跌倒，折斷頸項而死，因為他年紀老邁，身體沉重。 以利 作 以色列 的士師四十年。
1SAM|4|19|以利 的媳婦， 非尼哈 的妻子懷孕將到產期，她聽見上帝的約櫃被擄，公公和丈夫都死了，就曲身生產，極其疼痛。
1SAM|4|20|她將要死的時候，旁邊站著的婦人們對她說：「不要怕！你生了男孩了。」她不回答，也不放在心上。
1SAM|4|21|她給孩子起名叫 以迦博 ，說：「榮耀離開 以色列 了！」這是因為上帝的約櫃被擄去，又因為她公公和丈夫都死了。
1SAM|4|22|她又說：「榮耀離開 以色列 ，因為上帝的約櫃被擄去了。」
1SAM|5|1|非利士 人擄去上帝的約櫃，從 以便‧以謝 帶到 亞實突 。
1SAM|5|2|非利士 人擄了上帝的約櫃，帶進 大袞 廟，放在 大袞 的旁邊。
1SAM|5|3|次日， 亞實突 人清早起來，看哪， 大袞 仆倒在耶和華的約櫃前，臉伏於地，他們就扶起 大袞 ，把它放回原處。
1SAM|5|4|又次日，他們清早起來，看哪， 大袞 仆倒在耶和華的約櫃前，臉伏於地，並且 大袞 的頭和兩手都在門檻上折斷，只剩下 大袞 的軀幹。
1SAM|5|5|因此， 大袞 的祭司和所有進 大袞 廟的人，都不踏 亞實突 的 大袞 廟的門檻，直到今日。
1SAM|5|6|耶和華的手重重擊打 亞實突 人，使他們恐懼，使 亞實突 和 亞實突 周圍的人都生痔瘡。
1SAM|5|7|亞實突 人見這情況，就說：「 以色列 上帝的約櫃不可留在我們這裏，因為他的手重重擊打我們和我們的神明 大袞 」。
1SAM|5|8|他們就派人去請 非利士 的眾領袖來聚集，對他們說：「我們向 以色列 上帝的約櫃應當怎樣做呢？」他們說：「可以把 以色列 上帝的約櫃運到 迦特 去。」於是他們把 以色列 上帝的約櫃運到那裏。
1SAM|5|9|運到之後，耶和華的手擊打那城，使那城的人非常驚慌，無論大小都生痔瘡。
1SAM|5|10|他們就把上帝的約櫃送到 以革倫 。上帝的約櫃到了 以革倫 ， 以革倫 人就呼喊說：「他們把 以色列 上帝的約櫃運到我這裏，要害我和我的百姓！」
1SAM|5|11|於是他們派人去請 非利士 的眾領袖來，說：「請你們把 以色列 上帝的約櫃送回原處，免得害死我和我的百姓！」原來上帝的手重重攻擊那城，死亡的恐懼瀰漫全城，
1SAM|5|12|沒有死的人都受痔瘡的折磨。城裏的哀聲上達於天。
1SAM|6|1|耶和華的約櫃在 非利士 人之地七個月。
1SAM|6|2|非利士 人召了祭司和占卜的來，說：「我們向耶和華的約櫃應當怎樣做呢？請指示我們要用甚麼方法把約櫃送回原處。」
1SAM|6|3|他們說：「若要將 以色列 上帝的約櫃送回去，不可空手送回，一定要給他獻賠罪的禮物，然後你們才可以得痊癒，並且知道他的手為何不離開你們。」
1SAM|6|4|非利士 人說：「應當用甚麼獻為賠罪的禮物呢？」他們說：「當按照 非利士 領袖的數目，獻五個金痔瘡和五個金老鼠，因為你們眾人和領袖所遭遇的都是一樣的災禍。
1SAM|6|5|當製造你們痔瘡的像和毀壞田地老鼠的像，並要將榮耀歸給 以色列 的上帝，或者他向你們和你們的神明，以及你們的田地，把手放輕些。
1SAM|6|6|你們為何硬著心，像 埃及 人和法老硬著心一樣呢？上帝豈不是嚴厲對付 埃及 ，使 埃及 人釋放 以色列 人，他們就走了嗎？
1SAM|6|7|現在你們應當造一輛新車，把兩頭未曾負軛，還在哺乳的母牛套在車上，趕牛犢離開母牛，回家去。
1SAM|6|8|你們要把耶和華的約櫃放在車上，把所獻賠罪的金器裝在匣子裏，放在櫃旁，送走櫃子，讓它去。
1SAM|6|9|你們要觀察：車若直行過 以色列 的邊界，上到 伯‧示麥 去，這大災禍就是耶和華降在我們身上的；若不然，我們就知道，這不是他的手擊打我們，而是我們偶然遭遇的。」
1SAM|6|10|非利士 人就照樣做了。他們取了兩頭哺乳的母牛套在車上，把牛犢關在家裏，
1SAM|6|11|把耶和華的約櫃和裝金老鼠以及金痔瘡像的匣子都放在車上。
1SAM|6|12|牛直行大路，在往 伯‧示麥 的一條大道上，一面走一面叫，不偏左右。 非利士 的領袖跟在後面，直到 伯‧示麥 的地界。
1SAM|6|13|那時， 伯‧示麥 人正在平原收割麥子，舉目看見約櫃，就歡歡喜喜地迎見它。
1SAM|6|14|車到了 伯‧示麥 人 約書亞 的田間，就在那裏停了。在那裏有一塊大磐石，他們把車的木頭劈了，把兩頭母牛獻給耶和華為燔祭。
1SAM|6|15|利未 人將耶和華的約櫃和櫃子旁邊裝金器的匣子拿下來，放在大磐石上。當日 伯‧示麥 人獻上燔祭，又獻其他祭物給耶和華。
1SAM|6|16|非利士 人的五個領袖看見了，當日就回 以革倫 去。
1SAM|6|17|非利士 人獻給耶和華作賠罪的金痔瘡像如下：一個為 亞實突 ，一個為 迦薩 ，一個為 亞實基倫 ，一個為 迦特 ，一個為 以革倫 。
1SAM|6|18|金老鼠的數目是按照 非利士 五個領袖的城鎮，就是堅固的城鎮和鄉村，以及大磐石。這磐石是安放耶和華約櫃的，到今日還在 伯‧示麥 人 約書亞 的田間。
1SAM|6|19|耶和華擊殺 伯‧示麥 人，因為他們觀看他的約櫃。他擊殺了百姓七十人 。百姓因耶和華大大擊殺他們，就哀哭了。
1SAM|6|20|伯‧示麥 人說：「誰能在耶和華這位聖潔的上帝面前侍立呢？這約櫃可以從我們這裏上到誰那裏去呢？」
1SAM|6|21|於是他們派使者到 基列‧耶琳 的居民那裏，說：「 非利士 人將耶和華的約櫃送回來了，你們下來將約櫃接了，上到你們那裏去吧！」
1SAM|7|1|基列‧耶琳 人就來了，將耶和華的約櫃接上去，抬到山上 亞比拿達 的家中，將他兒子 以利亞撒 分別為聖，看守耶和華的約櫃。
1SAM|7|2|從約櫃留在 基列‧耶琳 的那天起，經過了許多日子，有二十年； 以色列 全家都哀哭歸向耶和華。
1SAM|7|3|撒母耳 對 以色列 全家說：「你們若全心回轉歸向耶和華，就要從你們中間除掉外邦的神明和 亞斯她錄 ，預備你們的心歸向耶和華，單單事奉他，他必救你們脫離 非利士 人的手。」
1SAM|7|4|以色列 人就除掉諸 巴力 和 亞斯她錄 ，單單事奉耶和華。
1SAM|7|5|撒母耳 說：「要召集 以色列 眾人到 米斯巴 去，我好為你們向耶和華禱告。」
1SAM|7|6|他們就聚集在 米斯巴 ，打水澆在耶和華面前。當日他們禁食，說：「我們得罪了耶和華。」 撒母耳 在 米斯巴 作 以色列 人的士師。
1SAM|7|7|非利士 人聽見 以色列 人聚集在 米斯巴 ， 非利士 的領袖就上來要攻擊 以色列 。 以色列 人聽見，就懼怕 非利士 人。
1SAM|7|8|以色列 人對 撒母耳 說：「願你不住為我們呼求耶和華－我們的上帝，救我們脫離 非利士 人的手。」
1SAM|7|9|撒母耳 就把一隻吃奶的羔羊獻給耶和華作全牲的燔祭，為 以色列 人呼求耶和華，耶和華就應允他。
1SAM|7|10|撒母耳 正獻燔祭的時候， 非利士 人前來要與 以色列 爭戰。當日，耶和華打雷，發出極大的聲音，使 非利士 人潰亂，他們就敗在 以色列 面前。
1SAM|7|11|以色列 人從 米斯巴 出來，追趕 非利士 人，擊殺他們，直到 伯‧甲 的下邊。
1SAM|7|12|撒母耳 拿一塊石頭立在 米斯巴 和 善 的中間，給石頭起名叫 以便‧以謝 ，說：「到如今耶和華都幫助我們。」
1SAM|7|13|因此， 非利士 人被制伏了，不再入侵 以色列 境內。 撒母耳 有生之年，耶和華的手攻擊 非利士 人。
1SAM|7|14|非利士 人所奪取 以色列 的城鎮，從 以革倫 直到 迦特 ，都歸回 以色列 了。 以色列 也從 非利士 人手中收回這些城所屬的地界。那時 以色列 與 亞摩利 人和平相處。
1SAM|7|15|撒母耳 一生作 以色列 的士師。
1SAM|7|16|他每年巡行到 伯特利 、 吉甲 、 米斯巴 ，在這些地方審判 以色列 人。
1SAM|7|17|隨後他回到 拉瑪 ，因為他的家在那裏；他在那裏審判 以色列 人，並且在那裏為耶和華築了一座壇。
1SAM|8|1|撒母耳 年紀老邁，就立他的兒子作 以色列 的士師。
1SAM|8|2|他的長子名叫 約珥 ，次子名叫 亞比亞 ；他們在 別是巴 作士師。
1SAM|8|3|他的兒子不行他的道，貪圖財利，收取賄賂，屈枉正直。
1SAM|8|4|以色列 的長老都聚集在 拉瑪 ，來到 撒母耳 那裏，
1SAM|8|5|對他說：「看哪，你年紀老了，你的兒子又不行你的道。現在請你為我們立一個王治理我們，像列國一樣。」
1SAM|8|6|撒母耳 不喜悅他們說「立一個王治理我們」，他就向耶和華禱告。
1SAM|8|7|耶和華對 撒母耳 說：「你只管聽從百姓向你說的一切話，因為他們不是厭棄你，而是厭棄我，不要我作他們的王。
1SAM|8|8|自從我領他們出 埃及 的日子到如今，他們離棄我，事奉別神；正像他們從前所做的一切事，現在他們也照樣向你做了。
1SAM|8|9|現在你只管聽從他們的話，不過要嚴厲警告他們，告訴他們將來王會用甚麼方式管轄他們。」
1SAM|8|10|撒母耳 將耶和華一切的話轉告求他立王的百姓。
1SAM|8|11|他說：「管轄你們的王必用這樣的方式：他必派你們的兒子為他駕車，趕馬，在他的戰車前奔跑。
1SAM|8|12|他要為自己立千夫長、五十夫長；耕種他的田地，收割他的莊稼；打造他的兵器和車上的器械。
1SAM|8|13|他必叫你們的女兒為他製造香膏，作廚師與烤餅的，
1SAM|8|14|也必取你們最好的田地、葡萄園、橄欖園，賜給他的臣僕。
1SAM|8|15|你們的糧食和葡萄園所出產的，他必徵收十分之一給他的官員和臣僕，
1SAM|8|16|又必叫你們的僕人婢女，健壯的青年和你們的驢為他做工。
1SAM|8|17|你們的羊群，他必徵收十分之一，你們自己也必作他的僕人。
1SAM|8|18|那日，你們必因自己所選的王哀求耶和華，但那日耶和華卻不應允你們。」
1SAM|8|19|百姓卻不肯聽 撒母耳 的話，說：「不！我們一定要一個王治理我們，
1SAM|8|20|使我們像列國一樣，有王治理我們，率領我們，為我們爭戰。」
1SAM|8|21|撒母耳 聽見百姓這一切話，就稟告給耶和華聽。
1SAM|8|22|耶和華對 撒母耳 說：「你只管聽從他們的話，為他們立一個王。」 撒母耳 對 以色列 人說：「去，你們各歸各城吧！」
1SAM|9|1|有一個 便雅憫 人名叫 基士 ，是 便雅憫 人 亞斐亞 的玄孫， 比歌拉 的曾孫， 洗羅 的孫子， 亞別 的兒子，是個大能的勇士 。
1SAM|9|2|他有一個兒子名叫 掃羅 ，又健壯、又英俊，在 以色列 人中沒有一個可以與他相比；他比眾百姓高出一個頭 。
1SAM|9|3|掃羅 的父親 基士 丟失了幾匹母驢，他就吩咐兒子 掃羅 說：「起來，帶一個僕人去尋找驢子。」
1SAM|9|4|掃羅 走過 以法蓮 山區，又過 沙利沙 地，都沒有找著。他們走過 沙琳 地，驢不在那裏，又走過 便雅憫 地，也沒有找到。
1SAM|9|5|到了 蘇弗 地， 掃羅 對跟隨他的僕人說：「我們不如回去，免得我父親不為驢掛慮，反為我們擔憂。」
1SAM|9|6|僕人對他說：「看哪，這城裏有一位神人，受人敬重，凡他所說的全都應驗。現在讓我們到他那裏去，或者他能指示我們當走的路。」
1SAM|9|7|掃羅 對僕人說：「看哪，我們若去，送甚麼給那人呢？我們袋子裏的食物都吃完了，也沒有禮物可以送給神人，我們還有些甚麼呢？」
1SAM|9|8|僕人又回答 掃羅 說：「看哪，我手裏還有四分之一舍客勒的銀子，可以送給神人，請他指示我們當走的路。」
1SAM|9|9|從前 以色列 中，若有人去求問上帝，就這麼說：「來，我們到先見那裏去吧！」因現在的先知，從前稱為先見。
1SAM|9|10|掃羅 對僕人說：「好主意！來，我們去吧。」於是他們往神人所住的城裏去了。
1SAM|9|11|他們上坡要進城，遇見幾個少女出來打水，就問她們說：「先見有沒有在這裏呢？」
1SAM|9|12|她們回答說：「有的，看哪，他就在你們前面。快！他今日正來到城裏，因為今日百姓要在丘壇獻祭。
1SAM|9|13|你們一進城，他還沒有上丘壇吃祭物之前，就會遇見他。因為他沒有到，百姓不能吃，必須等他先為祭物祝謝，然後受邀的人才可以吃。現在就上去吧，因為這時候你們會遇見他。」
1SAM|9|14|他們就上到那城，進入城中的時候，看哪， 撒母耳 正迎著他們來，要上丘壇去。
1SAM|9|15|掃羅 還沒有到的前一日，耶和華已經對 撒母耳 啟示說：
1SAM|9|16|「明日這時候，我必使一個人從 便雅憫 地到你這裏來，你要膏他作我百姓 以色列 的君王。他必救我的百姓脫離 非利士 人的手，因為我眷顧我的百姓 ，他們的哀聲已上達於我。」
1SAM|9|17|撒母耳 看見 掃羅 的時候，耶和華對他說：「看哪，這就是我對你所說的人，他必治理我的百姓。」
1SAM|9|18|掃羅 在城門中走到 撒母耳 跟前，說：「請告訴我，先見的家在哪裏？」
1SAM|9|19|撒母耳 回答掃羅說：「我就是先見。你在我前面先上丘壇去，因為你們今日必跟我同席。明日早晨我送你走，會把你心裏一切的事都告訴你。
1SAM|9|20|至於你前三日所丟失的幾匹母驢，你心裏不必掛慮，都已經找到了。 以色列 眾人所仰慕的是誰呢？不是仰慕你和你父的全家嗎？」
1SAM|9|21|掃羅 回答說：「我不是 以色列 支派中最小的 便雅憫 人嗎？我的家族不是 便雅憫 支派中最小的家族嗎？你為何對我說這樣的話呢？」
1SAM|9|22|撒母耳 領 掃羅 和他的僕人進了大廳，使他們在受邀的人中坐首位；受邀者約有三十個。
1SAM|9|23|撒母耳 對廚師說：「我交給你的那一份祭肉，吩咐你收存的，現在可以拿來。」
1SAM|9|24|廚師就舉起祭肉的腿和腿上的部分 ，擺在 掃羅 面前。 撒母耳 說：「看哪，所存留的擺在你面前了。吃吧！因為這是為你保留到這特定的時候的，好讓你說，是我請了這百姓來，」 當日， 掃羅 就與 撒母耳 同席。
1SAM|9|25|他們從丘壇下來進城， 撒母耳 和 掃羅 在房頂上說話。
1SAM|9|26|次日他們清早起來。黎明的時候， 撒母耳 呼叫在房頂上的 掃羅 ，說：「起來，我好送你回去。」 掃羅 就起來，和 撒母耳 二人一同到外面去。
1SAM|9|27|二人下到城邊， 撒母耳 對 掃羅 說：「你要吩咐僕人先走，僕人走了以後， 你要留在這裏，這時候我要將上帝的話傳給你聽。」
1SAM|10|1|撒母耳 拿一瓶膏油倒在 掃羅 的頭上，親吻他，說：「耶和華豈不是膏你作他產業的君王嗎？
1SAM|10|2|你今日離開我之後，會在 便雅憫 境內的 謝撒 ，靠近 拉結 的墳墓，遇見兩個人。他們會對你說：『你要找的幾匹母驢已經找到了。看哪，你父親不為驢子的事掛慮，反為你擔憂，說：我為兒子該做些甚麼呢？』
1SAM|10|3|你從那裏往前走，到了 他泊 的橡樹那裏，會遇見三個往 伯特利 去敬拜上帝的人：一個帶著三隻小山羊，一個帶著三個餅，一個帶著一皮袋酒。
1SAM|10|4|他們會向你問安，給你兩個餅，你就從他們手中接過來。
1SAM|10|5|然後你要到上帝的山去，在那裏有 非利士 的駐軍。你到了城裏的時候，會遇見一隊先知從丘壇下來，前面有鼓瑟的、擊鼓的、吹笛的、彈琴的，他們都受感說話。
1SAM|10|6|耶和華的靈必大大感動你，你就與他們一同受感說話，轉變成另一個人。
1SAM|10|7|這徵兆臨到你，你就要趁機做該做的事，因為上帝與你同在。
1SAM|10|8|你要在我以先下到 吉甲 。看哪，我必下到你那裏獻燔祭和平安祭。你要等候七日，等我到你那裏指示你當做的事。」
1SAM|10|9|掃羅 轉身離開 撒母耳 ，上帝就改變他，賜給他另一顆心。當日這一切徵兆都應驗了。
1SAM|10|10|他們來到那座山，看哪，有一隊先知遇見 掃羅 。上帝的靈大大感動他，他就在先知中受感說話。
1SAM|10|11|所有先前認識 掃羅 的人看見了，看哪，他和先知一同受感說話，百姓就彼此說：「 基士 的兒子遇見了甚麼呢？ 掃羅 也在先知中嗎？」
1SAM|10|12|那地方有一個人說：「這些人的父親是誰呢？」因此就有一句俗語說：「 掃羅 也在先知中嗎？」
1SAM|10|13|掃羅 受感說完了話，就上丘壇去了。
1SAM|10|14|掃羅 的叔叔問 掃羅 和他的僕人說：「你們到哪裏去了？」他說：「我們找驢子去了。但我們找不到，就去了 撒母耳 那裏。」
1SAM|10|15|掃羅 的叔叔說：「告訴我 撒母耳 對你們說了些甚麼。」
1SAM|10|16|掃羅 對他的叔叔說：「他明明告訴我們，驢子已經找到了。」至於 撒母耳 所說君王的事， 掃羅 沒有告訴叔叔。
1SAM|10|17|撒母耳 召集百姓到 米斯巴 耶和華那裏。
1SAM|10|18|他對 以色列 眾人說：「耶和華－ 以色列 的上帝如此說：『我領 以色列 出 埃及 ，救你們脫離 埃及 人的手，以及脫離欺壓你們各國之人的手。』
1SAM|10|19|你們今日卻厭棄救你們脫離一切災禍和患難的上帝，對他說：『求你立一個王治理我們。』現在你們應當按支派和宗族站在耶和華面前。」
1SAM|10|20|於是， 撒母耳 叫 以色列 眾支派近前來抽籤，抽到了 便雅憫 支派。
1SAM|10|21|然後，他叫 便雅憫 支派按宗族近前來，抽到了 瑪特利 族，接著又抽到了 基士 的兒子 掃羅 。眾人尋找他卻找不到，
1SAM|10|22|就再問耶和華說：「那人來到這裏了沒有？」耶和華說：「看哪，他藏在物品堆中。」
1SAM|10|23|眾人就跑去從那裏領他出來。他站在百姓中間，比眾百姓高出一個頭。
1SAM|10|24|撒母耳 對眾百姓說：「你們看到了耶和華所揀選的人嗎？眾百姓中沒有人可以與他相比。」眾百姓就歡呼說：「願王萬歲！」
1SAM|10|25|撒母耳 將君王的典章對百姓說明，又記在書上，放在耶和華面前，然後 撒母耳 遣散眾百姓，各回自己的家去了。
1SAM|10|26|掃羅 也往 基比亞 自己的家去，有一群心中被上帝感動的勇士跟隨他。
1SAM|10|27|但有些無賴之輩說：「這人怎麼能救我們呢？」他們就藐視他，不送禮物給他。 掃羅 卻保持沉默。
1SAM|11|1|亞捫 人 拿轄 上來，對著 基列 的 雅比 安營。 雅比 眾人對 拿轄 說：「你與我們立約，我們就服事你。」
1SAM|11|2|亞捫 人 拿轄 對他們說：「你們若由我挖出你們各人的右眼，以此凌辱 以色列 眾人，我就與你們立約。」
1SAM|11|3|雅比 的長老對他說：「求你寬容我們七日，等我們派人到 以色列 的全境去。若沒有人來救我們，我們就出來歸順你。」
1SAM|11|4|使者到了 掃羅 住的 基比亞 ，把這事說給百姓聽，眾百姓就都放聲大哭。
1SAM|11|5|看哪， 掃羅 正從田間趕牛回來，說：「百姓為甚麼哭呢？」眾人把 雅比 人的話告訴他。
1SAM|11|6|掃羅 聽見這些話，就被上帝的靈催逼，大發怒氣。
1SAM|11|7|他把一對牛切成小塊，吩咐使者傳送到 以色列 全境，說：「凡不出來跟隨 掃羅 和 撒母耳 的，就必這樣待他的牛。」耶和華使百姓懼怕，他們就都出來如同一人。
1SAM|11|8|掃羅 在 比色 數點他們： 以色列 人有三十萬， 猶大 人有三萬。
1SAM|11|9|他們對那些來的使者說：「你們要對 基列 的 雅比 人這樣說，明天太陽快到中午的時候，你們必得解救。」使者回去告訴 雅比 人，他們就歡喜了。
1SAM|11|10|於是 雅比 人對 亞捫 人說：「明日我們出來歸順你們，可以照你們看為好的待我們。」
1SAM|11|11|第二日， 掃羅 把百姓分為三隊，在清晨換崗哨的時候入侵 亞捫 人的軍營，擊殺他們直到中午的時候。逃脫的人都分散了，甚至沒有兩個人同在一起。
1SAM|11|12|百姓對 撒母耳 說：「那說『 掃羅 豈能作我們的王』的是誰呢？把他們交出來，我們好處死他們。」
1SAM|11|13|掃羅 說：「今日耶和華在 以色列 中施行拯救，所以今日不可處死人。」
1SAM|11|14|撒母耳 對百姓說：「來，我們到 吉甲 去，在那裏開始新的王國。」
1SAM|11|15|眾百姓到了 吉甲 那裏，在耶和華面前擁立 掃羅 為王，又在耶和華面前獻平安祭。 掃羅 和 以色列 眾人在那裏都非常歡喜。
1SAM|12|1|撒母耳 對 以色列 眾人說：「看哪，我已聽了你們對我所說一切的話，為你們立了一個王。
1SAM|12|2|現在，看哪，有這王行走在你們前面。我已年老髮白，看哪，我的兒子都在你們這裏。我從幼年直到今日都行走在你們前面。
1SAM|12|3|我在這裏，你們要在耶和華和他的受膏者面前為我作證，我奪過誰的牛，搶過誰的驢，欺負過誰，虐待過誰，從誰手裏收過賄賂而蒙蔽自己的眼目呢？若有，我必償還。」
1SAM|12|4|眾人說：「你未曾欺負我們，虐待我們，也未曾從任何人手裏收過任何東西。」
1SAM|12|5|撒母耳 對他們說：「你們在我手裏沒有找著甚麼，有耶和華在你們中間作證，也有他的受膏者今日作證。」他們說 ：「願耶和華作證。」
1SAM|12|6|撒母耳 對百姓說：「從前立 摩西 和 亞倫 ，又領你們祖先出 埃及 地的是耶和華。
1SAM|12|7|現在你們要站住，讓我在耶和華面前，以耶和華向你們和你們祖先所行一切公義的事來和你們爭辯。
1SAM|12|8|從前 雅各 到了 埃及 ，後來你們的祖先呼求耶和華，耶和華就差遣 摩西 和 亞倫 領你們的祖先出 埃及 ，來到這地方居住。
1SAM|12|9|他們卻忘記耶和華－他們的上帝，他就把他們交給 夏瑣 將軍 西西拉 的手中，以及 非利士 人和 摩押 王的手中 。於是這些人常來攻擊他們。
1SAM|12|10|他們呼求耶和華說：『我們離棄了耶和華去事奉諸 巴力 和 亞斯她錄 ，我們有罪了。現在求你救我們脫離仇敵的手，我們必事奉你。』
1SAM|12|11|耶和華就差遣 耶路巴力 、 比但 、 耶弗他 、 撒母耳 救你們脫離四圍仇敵的手，你們才安然居住。
1SAM|12|12|你們見 亞捫 人的王 拿轄 來攻擊你們，就對我說：『不，要有一個王治理我們。』其實耶和華－你們的上帝是你們的王。
1SAM|12|13|現在，看哪，這就是你們所選的、你們所求的王。看哪，耶和華已經為你們立王了。
1SAM|12|14|你們若敬畏耶和華，事奉他，聽從他的話，不違背耶和華的命令，你們和治理你們的王也都跟從耶和華－你們的上帝就好了。
1SAM|12|15|倘若不聽從耶和華的話，違背他的命令，耶和華的手必攻擊你們，像從前攻擊你們祖先一樣。
1SAM|12|16|現在你們要站住，看耶和華在你們眼前要行的一件大事。
1SAM|12|17|這不是割麥子的時候嗎？我求告耶和華，他必打雷降雨，讓你們知道並且看出，你們為自己求立王的事在耶和華眼前是犯大罪了。」
1SAM|12|18|於是 撒母耳 求告耶和華，耶和華就在這日打雷降雨，眾百姓就非常懼怕耶和華和 撒母耳 。
1SAM|12|19|眾百姓對 撒母耳 說：「請你為僕人向耶和華－你的上帝禱告，免得我們死亡，因為我們求立王的事，正是罪上加罪了。」
1SAM|12|20|撒母耳 對百姓說：「不要懼怕！你們雖然行了這惡，卻不要偏離耶和華，只要盡心事奉他。
1SAM|12|21|不可偏離去隨從那沒有益處、不能救人的虛無的神明 ，因為它們是虛無的。
1SAM|12|22|耶和華必因他大名的緣故不撇棄他的子民，因為耶和華喜悅你們作他的子民。
1SAM|12|23|至於我，我如果停止為你們禱告，就得罪耶和華了，我絕不會這樣做。我必以善道正路指教你們。
1SAM|12|24|但你們要敬畏耶和華，誠誠實實地盡心事奉他，因你們要留意，他向你們所行的事何等大。
1SAM|12|25|你們若不斷作惡，你們和你們的王必一同滅亡。」
1SAM|13|1|掃羅 登基的時候年三十 歲，作 以色列 王二年 。
1SAM|13|2|掃羅 從 以色列 中選出三千人：二千跟隨 掃羅 在 密抹 和 伯特利 山區，一千跟隨 約拿單 在 便雅憫 的 基比亞 。其餘的百姓， 掃羅 打發他們各自回自己的帳棚去了。
1SAM|13|3|約拿單 攻擊 非利士 人在 迦巴 的駐軍， 非利士 人聽見了這事。 掃羅 就在遍地吹角，說：「讓 希伯來 人都聽見。」
1SAM|13|4|以色列 眾人聽見 掃羅 攻擊 非利士 的駐軍，又聽見 以色列 為 非利士 人所憎惡，百姓就跟隨 掃羅 ，在 吉甲 集合。
1SAM|13|5|非利士 人集合，要與 以色列 人作戰。他們有戰車三萬輛，騎兵六千，士兵像海邊的沙那樣多。他們上來，在 伯‧亞文 東邊的 密抹 安營。
1SAM|13|6|以色列 人見自己危急，軍隊被圍攻，百姓就藏在山洞、叢林、巖隙、地窖和深坑中。
1SAM|13|7|有些 希伯來 人過了 約旦河 ，逃到 迦得 和 基列 地。 掃羅 還在 吉甲 ，所有的人都戰戰兢兢地跟隨他。
1SAM|13|8|掃羅 照著 撒母耳 所定的日期等了七日。但是， 撒母耳 還沒有來到 吉甲 ，百姓就離開 掃羅 散去了。
1SAM|13|9|於是 掃羅 說：「把燔祭和平安祭帶到我這裏來。」 掃羅 就獻上燔祭。
1SAM|13|10|他剛獻完燔祭，看哪， 撒母耳 就到了。 掃羅 出去迎接他，向他問安。
1SAM|13|11|撒母耳 說：「你做了甚麼事啊？」 掃羅 說：「因為我見百姓離開我散去，你又不照所定的日期來到，而且 非利士 人已在 密抹 集合；
1SAM|13|12|我說：『現在 非利士 人已經下到 吉甲 來攻擊我，可是我還沒有向耶和華禱告。』所以我就勉強獻上燔祭。」
1SAM|13|13|撒母耳 對 掃羅 說：「你做了糊塗事了，沒有遵守耶和華－你上帝吩咐你的命令。不然，耶和華會在 以色列 中堅立你的國度，直到永遠。
1SAM|13|14|現在你的國度必不長久。耶和華已經尋著一個合他心意的人，立他作百姓的君王，因為你沒有遵守耶和華所吩咐你的。」
1SAM|13|15|撒母耳 就起來，從 吉甲 上到 便雅憫 的 基比亞 。 掃羅 數點跟隨他的百姓，約有六百人。
1SAM|13|16|掃羅 和他兒子 約拿單 ，以及跟隨他們的百姓，都住在 便雅憫 的 迦巴 ， 非利士 人卻在 密抹 安營。
1SAM|13|17|有突擊隊從 非利士 營中出來，分成三隊：一隊往 俄弗拉 到 書亞 地去，
1SAM|13|18|一隊往 伯‧和崙 去，一隊往邊界，下望朝著曠野的 洗波音谷 。
1SAM|13|19|那時， 以色列 全地找不到一個鐵匠，因為 非利士 人說：「恐怕 希伯來 人製造刀槍。」
1SAM|13|20|以色列 眾人要磨鋤、犁、斧、鏟，就各自下到 非利士 人那裏去磨。
1SAM|13|21|磨鋤或犁的價錢是三分之二舍客勒，磨斧或修整刺棒的價錢是三分之一舍客勒。
1SAM|13|22|所以到了戰爭的日子，所有跟隨 掃羅 和 約拿單 的百姓找不到一個手裏有刀有槍的，惟 掃羅 和他兒子 約拿單 有。
1SAM|13|23|非利士 人的一隊駐軍出來，到 密抹 的隘口。
1SAM|14|1|有一日， 掃羅 的兒子 約拿單 對拿他兵器的青年說：「來，我們過去到 非利士 的駐軍那裏。」但他沒有告訴父親。
1SAM|14|2|掃羅 在 基比亞 的郊外，坐在 米磯崙 的石榴樹下，跟隨他的百姓約有六百人。
1SAM|14|3|在那裏有 亞希突 的兒子 亞希亞 ，穿著以弗得。 亞希突 是 以迦博 的哥哥， 非尼哈 的兒子， 以利 的孫子。 以利 從前在 示羅 作耶和華的祭司。 約拿單 去了，百姓卻不知道。
1SAM|14|4|約拿單 要從隘口過到 非利士 駐軍那裏去。這隘口兩邊各有一座齒狀峭壁：一座名叫 播薛 ，另一座名叫 西尼 ；
1SAM|14|5|一座向北，對著 密抹 ，一座向南，對著 迦巴 。
1SAM|14|6|約拿單 對拿兵器的青年說：「來，我們過去到那些未受割禮之人的駐軍那裏，或者耶和華為我們施展能力，因為耶和華使人得勝，不在乎人多人少 。」
1SAM|14|7|拿兵器的對他說：「隨你的心意做吧。你上去，看哪，我一定跟隨你，與你同心。」
1SAM|14|8|約拿單 說：「看哪，我們要過去到那些人那裏，在他們那裏展現我們自己。
1SAM|14|9|他們若對我們這麼說：『站住，等我們到你們那裏去』，我們就站在原地，不上他們那裏去；
1SAM|14|10|但他們若這麼說：『上到我們這裏來吧』，我們就上去，因為耶和華把他們交在我們手裏了。這就是我們的憑據。」
1SAM|14|11|二人就讓 非利士 的駐軍看見。 非利士 人說：「看哪， 希伯來 人從躲藏的洞穴裏出來了！」
1SAM|14|12|站崗的士兵對 約拿單 和拿兵器的人說：「上到這裏來，我們有一件事要告訴你們。」 約拿單 就對拿兵器的人說：「跟我上去，因為耶和華把他們交在 以色列 人手裏了。」
1SAM|14|13|約拿單 手腳並用爬上去，拿兵器的人跟隨他。 非利士 人仆倒在 約拿單 面前，拿兵器的人跟著他，殺死他們。
1SAM|14|14|約拿單 和拿兵器的人第一次擊殺的約有二十人，都在一畝 地的半犁溝之內。
1SAM|14|15|於是在軍營、在田野、在眾百姓中，人心惶惶，駐軍和突擊隊都戰兢；地也震動，這是從上帝那裏來的驚恐 。
1SAM|14|16|在 便雅憫 的 基比亞 ， 掃羅 的哨兵觀看，看哪， 非利士 全軍潰亂，四處亂竄。
1SAM|14|17|掃羅 就對跟隨他的百姓說：「你們去數點人數，看是誰從我們這裏出去。」他們一數點，看哪， 約拿單 和拿兵器的人不在其中。
1SAM|14|18|那時上帝的約櫃 在 以色列 人那裏。 掃羅 對 亞希亞 說：「你把上帝的約櫃請到這裏來。」
1SAM|14|19|掃羅 正與祭司說話的時候， 非利士 營中的騷亂越來越劇烈； 掃羅 就對祭司說：「停手吧！」
1SAM|14|20|掃羅 和所有跟隨他的百姓都集合，來到戰場，看哪， 非利士 人用刀互相擊殺，大大混亂。
1SAM|14|21|那先前由四方來跟隨 非利士 人、在他們營中的 希伯來 人，現在也轉過來幫助跟隨 掃羅 和 約拿單 的 以色列 人了。
1SAM|14|22|那藏在 以法蓮 山區的 以色列 眾人聽說 非利士 人逃跑，就出來緊緊地追擊他們。
1SAM|14|23|那日，耶和華使 以色列 人得勝，戰爭一直打到 伯‧亞文 。
1SAM|14|24|那日， 以色列 人非常困憊，因為 掃羅 叫百姓起誓說：「凡不等到晚上我向敵人報完了仇就吃東西的，必受詛咒。」因此所有的百姓都沒有嘗食物。
1SAM|14|25|所有的百姓 進入樹林，見地面上有蜜。
1SAM|14|26|百姓進了樹林，看哪，有蜜流出來，卻沒有人敢用手取蜜入口，因為百姓怕那誓言。
1SAM|14|27|約拿單 沒有聽見他父親叫百姓起誓，所以他伸出手中的杖，以杖頭蘸在蜂房裏，用手取回送入口內，他的眼睛就明亮了。
1SAM|14|28|百姓中有一人對他說：「你父親曾叫百姓嚴嚴地起誓說，今日吃東西的人必受詛咒；因此百姓就疲乏了。」
1SAM|14|29|約拿單 說：「我父親給這地添麻煩了。你們看，我嘗了這一點蜜，眼睛就明亮了。
1SAM|14|30|今日百姓若隨意吃了從仇敵奪來的東西，現在擊殺的 非利士 人豈不更多嗎？」
1SAM|14|31|這日， 以色列 人擊殺 非利士 人，從 密抹 直到 亞雅崙 。但百姓非常疲乏，
1SAM|14|32|就急著撲向掠物，奪取牛羊和牛犢，宰於地上，連肉帶血吃了。
1SAM|14|33|有人告訴 掃羅 說：「看哪，百姓吃帶血的肉，得罪耶和華了。」 掃羅 說：「你們行了詭詐，今日把一塊大石頭滾到我這裏來吧。」
1SAM|14|34|掃羅 又說：「你們分散到百姓中，對他們說，你們各人把牛羊牽到我這裏來宰了吃，不可吃帶血的肉得罪耶和華。」那夜，所有的百姓把自己手中的牛 牽到那裏宰了。
1SAM|14|35|掃羅 為耶和華築了一座壇，這是他開始為耶和華築的壇。
1SAM|14|36|掃羅 說：「我們要在夜裏下去追趕 非利士 人，搶掠他們，直到天亮，不給他們留下一人。」眾百姓說：「你看怎樣好就做吧！」祭司說：「我們要先在這裏親近上帝。」
1SAM|14|37|掃羅 求問上帝說：「我可以下去追趕 非利士 人嗎？你把他們交在 以色列 人手裏嗎？」這日上帝沒有回答他。
1SAM|14|38|掃羅 說：「百姓中的眾領袖，你們都要近前來到這裏，查明今日這罪是怎樣發生的。
1SAM|14|39|我指著拯救 以色列 的永生的耶和華起誓，就是我兒子 約拿單 犯了罪，他也必被處死。」但眾百姓中無人回答他。
1SAM|14|40|掃羅 對 以色列 眾人說：「你們站在一邊，我與我兒子 約拿單 也站在一邊。」百姓對 掃羅 說：「你看怎樣好就做吧！」
1SAM|14|41|掃羅 向耶和華－ 以色列 的上帝禱告說：「求你指示正確的答案。」抽中的是 掃羅 和 約拿單 ，百姓盡都無事。
1SAM|14|42|掃羅 說：「你們再抽籤，看是我，還是我兒子 約拿單 。」抽中的是 約拿單 。
1SAM|14|43|掃羅 對 約拿單 說：「你告訴我，你做了甚麼事？」 約拿單 說：「我只是用手中的杖，以杖頭蘸了一點蜜嘗嘗，看哪，我就要死嗎？」
1SAM|14|44|掃羅 說：「 約拿單 哪，你一定要死！若不然，願上帝重重懲罰我。」
1SAM|14|45|百姓對 掃羅 說：「 約拿單 在 以色列 中大行拯救，豈可死呢？絕對不可！我們指著永生的耶和華起誓，連他的一根頭髮也不可落地，因為他今日與上帝一同做事。」於是百姓救 約拿單 免了死亡。
1SAM|14|46|掃羅 上去，不追趕 非利士 人， 非利士 人也回本地去了。
1SAM|14|47|掃羅 執掌 以色列 的國權，攻打他四圍所有的仇敵，就是 摩押 人、 亞捫 人、 以東 人和 瑣巴 諸王，以及 非利士 人。他無論往何處去，都打敗他們。
1SAM|14|48|掃羅 奮勇作戰，擊敗 亞瑪力 人，救了 以色列 脫離搶掠他們之人的手。
1SAM|14|49|掃羅 的兒子是 約拿單 、 亦施韋 、 麥基‧舒亞 。他的兩個女兒：長女名叫 米拉 ，次女名叫 米甲 。
1SAM|14|50|掃羅 的妻子名叫 亞希暖 ，是 亞希瑪斯 的女兒。 掃羅 軍隊的元帥名叫 押尼珥 ，是 掃羅 的叔叔 尼珥 的兒子。
1SAM|14|51|掃羅 的父親 基士 ， 押尼珥 的父親 尼珥 ，都是 亞別 的兒子。
1SAM|14|52|掃羅 有生之年常與 非利士 人激烈爭戰，他看到任何有能力的人或勇士，都招募來跟隨他。
1SAM|15|1|撒母耳 對 掃羅 說：「耶和華差遣我膏你為王，治理他的百姓 以色列 ，現在你要聽從耶和華的話。
1SAM|15|2|萬軍之耶和華如此說：『 以色列 人從 埃及 上來的時候，在路上 亞瑪力 人怎樣待他們，怎樣抵擋他們，我都要懲罰。
1SAM|15|3|現在你要去攻打 亞瑪力 人，滅盡他們所有的，不可憐惜他們，將男女、孩童、吃奶的，以及牛、羊、駱駝和驢全都殺死。』」
1SAM|15|4|於是 掃羅 在 提拉因 召集百姓，數點他們，共有二十萬步兵和一萬 猶大 人。
1SAM|15|5|掃羅 到了 亞瑪力 的京城，在谷中設下埋伏。
1SAM|15|6|掃羅 對 基尼 人說：「你們離開 亞瑪力 人下去吧，免得我把你們和 亞瑪力 人一同殺滅，因為 以色列 眾人從 埃及 上來的時候，你們曾恩待他們。」於是 基尼 人離開了 亞瑪力 人。
1SAM|15|7|掃羅 攻打 亞瑪力 人，從 哈腓拉 直到 埃及 東邊的 書珥 ，
1SAM|15|8|生擒了 亞瑪力 王 亞甲 ，用刀殺盡 亞瑪力 的眾百姓。
1SAM|15|9|掃羅 和百姓卻憐惜 亞甲 ，愛惜上好的牛、羊、牛犢、羔羊，以及一切美物，不肯滅絕。但是凡看不上眼和沒有價值的，他們盡都殺了。
1SAM|15|10|耶和華的話臨到 撒母耳 說：
1SAM|15|11|「我立 掃羅 為王，我感到遺憾，因為他轉去不跟從我，不遵守我的命令。」 撒母耳 就很生氣，終夜哀求耶和華。
1SAM|15|12|撒母耳 清早起來，去見 掃羅 。有人告訴 撒母耳 說：「 掃羅 到了 迦密 ，看哪，他在那裏為自己立了紀念碑，又轉身下到 吉甲 。」
1SAM|15|13|撒母耳 到了 掃羅 那裏， 掃羅 對他說：「願耶和華賜福給你，耶和華的命令我已遵守了。」
1SAM|15|14|撒母耳 說：「我耳中聽見有羊叫、牛鳴的聲音，又是甚麼呢？」
1SAM|15|15|掃羅 說：「這是百姓從 亞瑪力 人那裏帶來的，因為他們愛惜上好的牛羊，要獻給耶和華－你的上帝。其餘的，我們都滅盡了。」
1SAM|15|16|撒母耳 對 掃羅 說：「住口吧！等我把耶和華昨夜向我所說的話告訴你。」 掃羅 說：「請說。」
1SAM|15|17|撒母耳 說：「你雖然看自己為小，你豈不是作了 以色列 諸支派的元首嗎？耶和華膏你作了 以色列 的王。
1SAM|15|18|耶和華差遣你，吩咐你說：『你去除滅那些犯罪的 亞瑪力 人，攻打他們，直到把他們完全滅盡。』
1SAM|15|19|你為何沒有聽從耶和華的話呢？你為何急著撲向掠物，行耶和華眼中看為惡的事呢？」
1SAM|15|20|掃羅 對 撒母耳 說：「我聽從了耶和華的話，行了耶和華派我行的路，擒了 亞瑪力 王 亞甲 來，滅盡了 亞瑪力 人。
1SAM|15|21|百姓卻從掠物中取了牛羊，是當滅之物中最好的，要在 吉甲 獻給耶和華－你的上帝。」
1SAM|15|22|撒母耳 說： 「耶和華喜愛燔祭和祭物， 豈如喜愛人聽從他的話呢？ 看哪，聽命勝於獻祭， 順從勝於公羊的脂肪。
1SAM|15|23|悖逆與占卜的罪相等， 頑梗與拜偶像的罪孽相同。 因為你厭棄耶和華的命令， 耶和華也厭棄你作王。」
1SAM|15|24|掃羅 對 撒母耳 說：「我有罪了！我違背了耶和華的指示和你的命令；因為我懼怕百姓，聽從了他們的話。
1SAM|15|25|現在求你赦免我的罪，同我回去，我好敬拜耶和華。」
1SAM|15|26|撒母耳 對 掃羅 說：「我不同你回去，因為你厭棄耶和華的命令，耶和華也厭棄你作 以色列 的王。」
1SAM|15|27|撒母耳 轉身要走， 掃羅 抓住他外袍的衣角，外袍就斷裂了。
1SAM|15|28|撒母耳 對他說：「今日耶和華使 以色列 國與你斷絕，把這國賜給另一個比你更好的人。
1SAM|15|29|以色列 的大能者必不說謊，也不後悔，因為他不是世人，絕不後悔。」
1SAM|15|30|掃羅 說：「我有罪了。現在求你在我百姓的長老和 以色列 人面前尊重我，同我回去，我好敬拜耶和華－你的上帝。」
1SAM|15|31|於是 撒母耳 轉身跟隨 掃羅 回去， 掃羅 就敬拜耶和華。
1SAM|15|32|撒母耳 說：「把 亞瑪力 王 亞甲 帶到我這裏來。」 亞甲 就歡歡喜喜地來到他面前，說：「死亡的苦難必定過去了。」
1SAM|15|33|撒母耳 說：「你既用刀使婦人喪子，你母親在婦人中也必照樣喪子。」於是， 撒母耳 在 吉甲 耶和華面前把 亞甲 砍碎了。
1SAM|15|34|撒母耳 回了 拉瑪 。 掃羅 上他所住的 基比亞 ，回自己的家去了。
1SAM|15|35|撒母耳 直到死的日子，再沒有見 掃羅 。但 撒母耳 為 掃羅 悲傷，因為耶和華遺憾立 掃羅 為 以色列 的王。
1SAM|16|1|耶和華對 撒母耳 說：「我既厭棄 掃羅 作 以色列 的王，你為他悲傷要到幾時呢？你將膏油盛滿了角；來，我差遣你到 伯利恆 人 耶西 那裏去，因為我在他兒子中已看中了一個為我作王的。」
1SAM|16|2|撒母耳 說：「我怎麼能去呢？ 掃羅 一聽見，就會殺我。」耶和華說：「你可以手裏牽一頭小母牛去，說：『我來是要向耶和華獻祭。』
1SAM|16|3|你要請 耶西 來一同獻祭，我會指示你當做的事。我對你說的那個人，你要為我膏他。」
1SAM|16|4|撒母耳 遵照耶和華的話去做，來到 伯利恆 ，城裏的長老都戰戰兢兢出來迎接他，有人問他說：「你是為平安來的嗎？」
1SAM|16|5|他說：「為平安來的，我來是要向耶和華獻祭。你們要使自己分別為聖，來跟我一同獻祭。」 撒母耳 把 耶西 和他眾兒子分別為聖，請他們來一同獻祭。
1SAM|16|6|他們來的時候， 撒母耳 看見 以利押 ，就心裏說，耶和華的受膏者一定在耶和華面前了。
1SAM|16|7|耶和華卻對 撒母耳 說：「不要只看他的外貌和他身材高大，我不揀選他。因為耶和華不像人看人，人是看外貌 ，耶和華是看內心。」
1SAM|16|8|耶西 叫 亞比拿達 從 撒母耳 面前經過， 撒母耳 說：「耶和華也不揀選他。」
1SAM|16|9|耶西 又叫 沙瑪 經過， 撒母耳 說：「耶和華也不揀選他。」
1SAM|16|10|耶西 叫他七個兒子都從 撒母耳 面前經過， 撒母耳 對 耶西 說：「這些都不是耶和華所揀選的。」
1SAM|16|11|撒母耳 對 耶西 說：「你的兒子都在這裏了嗎？」他說：「還有一個最小的，看哪，他正在放羊。」 撒母耳 對 耶西 說：「你派人去叫他來；他若不來這裏，我們必不坐席。」
1SAM|16|12|耶西 就派人去叫他來。他面色紅潤，雙目清秀，容貌俊美。耶和華說：「起來，膏他，因為這就是他了。」
1SAM|16|13|撒母耳 就用角裏的膏油，在他的兄長中膏了他。從這日起，耶和華的靈就大大感動 大衛 。 撒母耳 起身回 拉瑪 去了。
1SAM|16|14|耶和華的靈離開 掃羅 ，有邪靈從耶和華那裏來擾亂他。
1SAM|16|15|掃羅 的臣僕對他說：「看哪，有邪靈從上帝那裏來擾亂你。
1SAM|16|16|我們的主可以吩咐你面前的臣僕，去找一個善於彈琴的來。上帝那裏來的邪靈臨到你身上的時候，他用手彈琴，你就會感覺爽快。」
1SAM|16|17|掃羅 對臣僕說：「你們給我找一個善於彈琴的，帶到我這裏來。」
1SAM|16|18|僕人中有一個回答說：「看哪，我曾見 伯利恆 人 耶西 的一個兒子善於彈琴，是大能的勇士，說話合宜，容貌俊美，耶和華也與他同在。」
1SAM|16|19|於是 掃羅 差遣使者到 耶西 那裏，說：「叫你放羊的兒子 大衛 到我這裏來。」
1SAM|16|20|耶西 把幾個餅和一皮袋酒，以及一隻小山羊，馱在驢上，由兒子 大衛 的手送給 掃羅 。
1SAM|16|21|大衛 到了 掃羅 那裏，就侍立在 掃羅 面前。 掃羅 很喜歡他，他就作了 掃羅 拿兵器的人。
1SAM|16|22|掃羅 派人到 耶西 那裏，說：「讓 大衛 侍立在我面前，因為他在我眼前蒙了恩寵。」
1SAM|16|23|從上帝那裏來的邪靈臨到 掃羅 身上的時候， 大衛 就拿琴，用手彈奏，使 掃羅 舒暢，感覺爽快，那邪靈就離開他了。
1SAM|17|1|非利士 人召集他們的軍隊來爭戰。他們聚集在 猶大 的 梭哥 ，在 梭哥 和 亞西加 中間的 以弗‧大憫 安營。
1SAM|17|2|掃羅 和 以色列 人也聚集，在 以拉谷 安營，擺陣迎戰，要與 非利士 人打仗。
1SAM|17|3|非利士 人站在這邊的山上， 以色列 人站在那邊的山上，當中有谷。
1SAM|17|4|從 非利士 營中出來一個挑戰的人，名叫 歌利亞 ，是 迦特 人，身高六肘一虎口。
1SAM|17|5|他頭戴銅盔，身穿鎧甲，甲重五千舍客勒銅。
1SAM|17|6|他腿上有銅護膝，兩肩之中背負銅矛。
1SAM|17|7|他的槍桿粗如織布機的軸，槍頭的鐵重六百舍客勒。有一個拿盾牌的人走在他前面。
1SAM|17|8|歌利亞 站著，對 以色列 的軍隊喊叫，對他們說：「你們出來擺陣作戰是為了甚麼呢？我不是 非利士 人嗎？你們不是 掃羅 的僕人嗎？你們選一個人出來，叫他下來到我這裏吧。
1SAM|17|9|他若能與我決鬥，把我殺死，我們就作你們的奴隸；我若勝了他，把他殺死，你們就作我們的奴隸，服事我們。」
1SAM|17|10|那 非利士 人又說：「我今日向 以色列 的軍隊罵陣。你們叫一個人出來，跟我決鬥吧。」
1SAM|17|11|掃羅 和 以色列 眾人聽見 非利士 人這些話就驚惶，非常害怕。
1SAM|17|12|大衛 是 猶大 伯利恆 的 以法他 人 耶西 的兒子， 耶西 有八個兒子。在 掃羅 的時候，這人年老，在眾人中受敬重 。
1SAM|17|13|耶西 最大的三個兒子跟隨 掃羅 出征。出征的三個兒子名字是：長子 以利押 ，次子 亞比拿達 ，三子 沙瑪 。
1SAM|17|14|大衛 是最小的，最大的三個兒子跟隨 掃羅 。
1SAM|17|15|大衛 有時離開 掃羅 ，回 伯利恆 為他父親放羊。
1SAM|17|16|那 非利士 人早晚都出來站著，共四十日。
1SAM|17|17|耶西 對他兒子 大衛 說：「你拿一伊法烘了的穗子和十個餅，跑到營裏去，交給你的哥哥，
1SAM|17|18|再拿這十塊奶餅，送給他們的千夫長，並要問你哥哥好，向他們要個憑據回來。」
1SAM|17|19|掃羅 和 大衛 的三個哥哥，以及 以色列 眾人，都在 以拉谷 與 非利士 人打仗。
1SAM|17|20|大衛 早晨起來，把羊交託一個看守的人，照 耶西 所吩咐的帶著食物去了。到了軍營，軍隊剛出到戰場，吶喊叫陣。
1SAM|17|21|以色列 人和 非利士 人都擺列陣勢，彼此相對。
1SAM|17|22|大衛 把東西留在看守物件的人手中，跑到戰場，問他哥哥好。
1SAM|17|23|他與他們說話的時候，看哪，那挑戰的人，就是 迦特 的 非利士 人 歌利亞 ，從 非利士 隊伍中上來，說了同樣的話， 大衛 聽見了。
1SAM|17|24|以色列 眾人看見那人就非常害怕，從他面前逃跑。
1SAM|17|25|以色列 人說：「這上來的人你看見了嗎？他上來是要向 以色列 人罵陣。若有人能殺他，王必賞賜他大財，將自己的女兒嫁給他，並在 以色列 人中免除他父家納糧服役。」
1SAM|17|26|大衛 對站在旁邊的人說：「若有人殺這 非利士 人，除掉 以色列 人的羞辱，他會怎樣呢？這未受割禮的 非利士 人是誰，竟敢向永生上帝的軍隊罵陣！」
1SAM|17|27|百姓照同樣的話對他說：「若有人殺了那人，必這樣待他。」
1SAM|17|28|大衛 的長兄 以利押 聽見 大衛 與他們所說的話，就向他發怒，說：「你下來做甚麼呢？在曠野的那幾隻羊，你交託誰了呢？我知道你的驕傲和你心裏的惡意，你下來只是為了看戰爭！」
1SAM|17|29|大衛 說：「我現在做了甚麼呢？只是問一句話也不可以嗎？」
1SAM|17|30|大衛 離開他轉向別人，問了同樣的事，百姓也照先前的話回答他。
1SAM|17|31|有人聽見 大衛 所說的話，就在 掃羅 面前報告； 掃羅 就派人叫他來。
1SAM|17|32|大衛 對 掃羅 說：「人不必因那 非利士 人灰心。你的僕人要去與他決鬥。」
1SAM|17|33|掃羅 對 大衛 說：「你不能去與那 非利士 人決鬥，因為你年紀太輕，他從小就是戰士。」
1SAM|17|34|大衛 對 掃羅 說：「你僕人為父親放羊，有時獅子來了，有時熊來了，從群中抓走一隻羔羊。
1SAM|17|35|我就追趕牠，擊打牠，把羔羊從牠口中救出來。牠起來攻擊我，我就揪牠的鬍子，打死牠。
1SAM|17|36|你僕人曾打死獅子和熊，這未受割禮的 非利士 人必像獅子和熊一樣，因為他向永生上帝的軍隊罵陣。」
1SAM|17|37|大衛 又說：「耶和華救我脫離獅子和熊的爪，他必救我脫離這 非利士 人的手。」 掃羅 對 大衛 說：「你去吧！耶和華必與你同在。」
1SAM|17|38|掃羅 把自己的戰衣給 大衛 穿上，將銅盔戴在他頭上，又給他穿上鎧甲。
1SAM|17|39|大衛 佩刀在戰衣上，試著走走看。因 大衛 沒有試過，就對 掃羅 說：「我穿戴這些不能走路，因為我沒有試過。」於是他脫下身上的這些軍裝。
1SAM|17|40|他手中拿杖，又在溪中挑選了五塊光滑的石子，放在袋裏，就是牧人帶的囊裏，手裏拿著甩石的機弦，迎向那 非利士 人。
1SAM|17|41|那 非利士 人漸漸走近 大衛 ，拿盾牌的人在他前面。
1SAM|17|42|非利士 人觀看，見了 大衛 ，就藐視他，因為他年輕，面色紅潤，容貌俊美。
1SAM|17|43|非利士 人對 大衛 說：「你拿著杖到我這裏來，我豈是狗嗎？」 非利士 人就指著自己的神明詛咒 大衛 。
1SAM|17|44|非利士 人又對 大衛 說：「來吧！我要把你的肉給空中的飛鳥和田野的走獸。」
1SAM|17|45|大衛 對 非利士 人說：「你來攻擊我，是靠著刀槍和銅矛，但我來攻擊你，是靠著萬軍之耶和華的名，就是你所辱罵、帶領 以色列 軍隊的上帝。
1SAM|17|46|今日耶和華必將你交在我手裏。我必殺你，砍下你的頭，今日我要把 非利士 軍兵的屍體給空中的飛鳥和地上的野獸，使全地的人都知道以色列中有上帝，
1SAM|17|47|又使這裏的全會眾知道，耶和華使人得勝，不是用刀用槍，因為戰爭全在乎耶和華。他必將你們交在我們手裏。」
1SAM|17|48|那 非利士 人起來，迎向 大衛 ，走近前來。 大衛 急忙往戰場，迎向 非利士 人跑去。
1SAM|17|49|大衛 伸手入囊中，從裏面掏出一塊石子來，用機弦甩去，擊中 非利士 人的前額，石子進入額內，他就仆倒，面伏於地。
1SAM|17|50|這樣， 大衛 用機弦和石子勝了那 非利士 人，擊中了他，把他殺死； 大衛 手中沒有刀。
1SAM|17|51|大衛 跑去，站在那 非利士 人身旁，把他的刀從鞘中拔出來，殺死他，用刀割下他的頭。 非利士 眾人看見他們的勇士死了，就都逃跑。
1SAM|17|52|以色列 人和 猶大 人就起來吶喊，追趕 非利士 人，直到 該 和 以革倫 的城門。被殺的 非利士 人倒在路上，從 沙拉音 直到 迦特 和 以革倫 。
1SAM|17|53|以色列 人追趕 非利士 人回來，搶奪了他們的軍營。
1SAM|17|54|大衛 拿著那 非利士 人的頭帶到 耶路撒冷 ，卻把那 非利士 人的軍裝放在自己的帳棚裏。
1SAM|17|55|掃羅 看見 大衛 去迎戰 非利士 人，就問 押尼珥 元帥說：「 押尼珥 ，那年輕人是誰的兒子？」 押尼珥 說：「王啊，我在你面前起誓，我不知道。」
1SAM|17|56|王說：「你可以問問那孩子是誰的兒子。」
1SAM|17|57|大衛 打死那 非利士 人回來， 押尼珥 領他到 掃羅 面前， 大衛 手中拿著 非利士 人的頭。
1SAM|17|58|掃羅 問他說：「年輕人，你是誰的兒子？」 大衛 說：「我是你僕人 伯利恆 人 耶西 的兒子。」
1SAM|18|1|大衛 對 掃羅 說完了話， 約拿單 的心與 大衛 的心深相契合。 約拿單 愛 大衛 ，如同愛自己的性命。
1SAM|18|2|那日 掃羅 留住 大衛 ，不讓他回父家。
1SAM|18|3|約拿單 愛 大衛 如同愛自己的性命，就與他立約。
1SAM|18|4|約拿單 從身上脫下外袍，給了 大衛 ，又把戰衣、刀、弓、腰帶都給了他。
1SAM|18|5|掃羅 無論差遣 大衛 往何處去，他都做事精明。 掃羅 立他作軍隊的指揮官，眾百姓和 掃羅 的臣僕都看為美。
1SAM|18|6|大衛 打死了那 非利士 人，同眾人回來的時候，婦女們從 以色列 各城裏出來，歡歡喜喜，打鼓奏樂，唱歌跳舞，迎接 掃羅 王。
1SAM|18|7|眾婦女歡樂唱和，說： 「 掃羅 殺死千千， 大衛 殺死萬萬。」
1SAM|18|8|掃羅 非常憤怒，不喜歡這話。他說：「將萬萬歸給 大衛 ，千千歸給我，只剩下王國沒有給他！」
1SAM|18|9|從這日起， 掃羅 就敵視 大衛 。
1SAM|18|10|次日，從上帝來的邪靈緊抓住 掃羅 ，他就在家中胡言亂語。 大衛 照常彈琴， 掃羅 手裏拿著槍。
1SAM|18|11|掃羅 把槍一擲，心裏說：「我要將 大衛 刺透，釘在牆上。」 大衛 閃避了他兩次。
1SAM|18|12|掃羅 懼怕 大衛 ，因為耶和華離開自己，與 大衛 同在。
1SAM|18|13|所以 掃羅 叫 大衛 離開自己，立他為千夫長，他就領兵出入。
1SAM|18|14|大衛 所做的每一件事都精明，耶和華也與他同在。
1SAM|18|15|掃羅 見 大衛 做事精明，就更怕他。
1SAM|18|16|但 以色列 和 猶大 眾人都愛 大衛 ，因為他領他們出入。
1SAM|18|17|掃羅 對 大衛 說：「看哪，我將大女兒 米拉 嫁給你，只要你作我的勇士，為耶和華爭戰。」 掃羅 心裏說：「我不好親手害他，要藉 非利士 人的手害他。」
1SAM|18|18|大衛 對 掃羅 說：「我是誰，我是甚麼出身，我父家在 以色列 中算甚麼，豈敢作王的女婿呢？」
1SAM|18|19|掃羅 的女兒 米拉 到了當嫁給 大衛 的時候， 掃羅 卻將她嫁給了 米何拉 人 亞得列 。
1SAM|18|20|掃羅 的女兒 米甲 愛 大衛 。有人告訴 掃羅 ，這件事在 掃羅 眼中看為合宜。
1SAM|18|21|掃羅 心裏說：「我把這女兒嫁給 大衛 ，作他的圈套，好藉 非利士 人的手害他。」所以 掃羅 第二次對 大衛 說：「你今日可以作我的女婿。」
1SAM|18|22|掃羅 吩咐臣僕：「你們暗中對 大衛 說：『看哪，王喜歡你，王的臣僕也都愛戴你，現在你就作王的女婿吧。』」
1SAM|18|23|掃羅 的臣僕照這話說給 大衛 聽。 大衛 說：「你們把作王的女婿看為小事嗎？我是貧窮卑微的人。」
1SAM|18|24|掃羅 的臣僕回奏說， 大衛 說了這樣的話。
1SAM|18|25|掃羅 說：「你們要對 大衛 這樣說：『王不要甚麼聘禮，只要一百 非利士 人的包皮，好在王的仇敵身上報仇。』」 掃羅 的意圖是要 大衛 落在 非利士 人的手中。
1SAM|18|26|掃羅 的臣僕把這話告訴 大衛 ， 大衛 就歡喜作王的女婿。日期還沒有到，
1SAM|18|27|大衛 和跟隨他的人起來前往，殺了二百 非利士 人，將包皮足數交給王，為要作王的女婿。於是 掃羅 將女兒 米甲 嫁給 大衛 。
1SAM|18|28|掃羅 見耶和華與 大衛 同在，女兒 米甲 又愛 大衛 ，
1SAM|18|29|就更怕 大衛 ，常常與 大衛 為敵。
1SAM|18|30|每逢 非利士 的軍官出來打仗， 大衛 做事比 掃羅 任何臣僕更精明，因此他的名極受尊重。
1SAM|19|1|掃羅 吩咐他兒子 約拿單 和眾臣僕要殺 大衛 ，但 掃羅 的兒子 約拿單 卻很喜愛 大衛 。
1SAM|19|2|約拿單 告訴 大衛 說：「我父 掃羅 想要殺你，現在你要小心，明日早晨留在一個僻靜的地方藏起來。
1SAM|19|3|我會出去，到你所藏的田裏，站在我父親旁邊，與父親談論到你。我看情形怎樣，會告訴你。」
1SAM|19|4|約拿單 向他父親 掃羅 說 大衛 的好話，對他說：「王不可得罪王的僕人 大衛 ，因為他未曾得罪你，他所行的對你都很有益處。
1SAM|19|5|他拚了命殺那 非利士 人，並且耶和華為全 以色列 大施拯救。那時你看見，也很歡喜，現在為何要犯罪，流無辜人的血，無緣無故殺 大衛 呢？」
1SAM|19|6|掃羅 聽了 約拿單 的話，就指著永生的耶和華起誓：「我絕不殺他。」
1SAM|19|7|約拿單 叫 大衛 來，把這一切事告訴他。 約拿單 帶他去見 掃羅 ，他就像以前一樣侍立在 掃羅 面前。
1SAM|19|8|此後又有戰爭， 大衛 出去與 非利士 人打仗。他大大擊敗他們，他們就在他面前逃跑。
1SAM|19|9|從耶和華來的邪靈又降在 掃羅 身上， 掃羅 手裏拿槍坐在屋裏， 大衛 正用手彈琴。
1SAM|19|10|掃羅 想要用槍刺透 大衛 ，把他釘在牆上，他卻躲開 掃羅 ， 掃羅 的槍刺入牆內。當夜 大衛 逃走，躲起來了。
1SAM|19|11|掃羅 派一些使者到 大衛 的房屋那裏守著他，等到天亮要殺他。 大衛 的妻子 米甲 對 大衛 說：「你今夜若不逃命，明日就要被殺。」
1SAM|19|12|於是 米甲 將 大衛 從窗戶縋下去，讓他走； 大衛 就逃走，躲起來了。
1SAM|19|13|米甲 把家中的神像放在床上，頭枕在山羊毛的枕頭上，用衣服蓋起來。
1SAM|19|14|掃羅 派一些使者去捉拿 大衛 ， 米甲 說：「他病了。」
1SAM|19|15|掃羅 又派一些使者去看 大衛 ，說：「把他連床一起抬到我這裏，我好殺他。」
1SAM|19|16|使者進去，看哪，神像在床上，頭枕在山羊毛的枕頭上。
1SAM|19|17|掃羅 對 米甲 說：「你為甚麼這樣欺騙我，放我仇敵逃走呢？」 米甲 對 掃羅 說：「他對我說：『你放我走吧，我何必要殺你呢？』」
1SAM|19|18|大衛 逃跑躲避，來到 拉瑪 的 撒母耳 那裏，把 掃羅 向他所行的事全告訴他。他和 撒母耳 就去，住在 拿約 。
1SAM|19|19|有人告訴 掃羅 說：「看哪， 大衛 在 拉瑪 的 拿約 」。
1SAM|19|20|掃羅 派一些使者去捉拿 大衛 。去的人見一隊先知受感說話， 撒母耳 站在當中領導他們， 掃羅 派去的使者也受上帝的靈感動說話。
1SAM|19|21|有人把這事告訴 掃羅 ，他又派另一些使者去，他們也受感說話。 掃羅 第三次派使者去，他們也受感說話。
1SAM|19|22|然後 掃羅 親自往 拉瑪 去，到了 西沽 的大井，問人說：「 撒母耳 和 大衛 在哪裏？」有人說：「看哪，在 拉瑪 的 拿約 。」
1SAM|19|23|他就往那裏去，到了 拉瑪 的 拿約 。上帝的靈也臨到他，他一面走一面受感說話，直到 拉瑪 的 拿約 。
1SAM|19|24|他也脫了衣服，也在 撒母耳 面前受感說話，一日一夜赤身躺臥。因此有人說：「 掃羅 也在先知中嗎？」
1SAM|20|1|大衛 從 拉瑪 的 拿約 逃跑，來到 約拿單 面前，對他說：「我做了甚麼，有甚麼罪孽，在你父親面前犯了甚麼罪，他竟要尋索我的性命呢？」
1SAM|20|2|約拿單 對他說：「絕無此事！你必不至於死。看哪，我父做事，無論大小，沒有不告訴我的。我父親為甚麼要隱瞞我這件事呢？不會這樣的！」
1SAM|20|3|大衛 又起誓說：「你父親確實知道我在你眼前蒙恩。所以他說，『這事不要讓 約拿單 知道，免得他愁煩。』我指著永生的耶和華起誓，又指著你的性命起誓，我離死只差一步而已。」
1SAM|20|4|約拿單 對 大衛 說：「你心裏所求的，我必為你成就。」
1SAM|20|5|大衛 對 約拿單 說：「看哪，明日是初一，我必須與王同席用餐，求你讓我去藏在田野，直到第三日傍晚。
1SAM|20|6|你父親若見我不在席上，你就說：『 大衛 懇求我允許他趕回本城 伯利恆 去，因為他全家在那裏獻年祭。』
1SAM|20|7|你父親若說好，你的僕人就平安了；他若大怒，你就知道他決意行惡。
1SAM|20|8|求你施恩於僕人，因你在耶和華面前曾與僕人立約。我若有罪孽，你就親自殺死我，何必把我交給你父親呢？」
1SAM|20|9|約拿單 說：「絕無此事！我若確實知道我父親決意害你，怎麼會不告訴你呢？」
1SAM|20|10|大衛 對 約拿單 說：「你父親若嚴厲回答你，誰來告訴我呢？」
1SAM|20|11|約拿單 對 大衛 說：「來，讓我們到田野去。」二人就往田野去了。
1SAM|20|12|約拿單 對 大衛 說：「願耶和華－ 以色列 的上帝作證。明日約在這時候，或第三日，我一探出我父親的心意，看哪，若對 大衛 是好意，我怎麼會不派人來告訴你呢？
1SAM|20|13|我父親若有意害你，而我不告訴你，送你平安地離開，願耶和華重重懲罰 約拿單 。願耶和華與你同在，如同從前與我父親同在一樣。
1SAM|20|14|你要照耶和華的慈愛恩待我，不但我活著的時候免我死亡，
1SAM|20|15|就是耶和華從地面逐一剪除 大衛 仇敵的時候，你也永不可向我家斷絕恩惠。」
1SAM|20|16|於是 約拿單 與 大衛 家立約：「願耶和華從 大衛 仇敵 的手來追討。」
1SAM|20|17|約拿單 因愛 大衛 如同愛自己的性命，就叫他再起誓。
1SAM|20|18|約拿單 對他說：「明日是初一，你的座位空著，人必察覺你不在。
1SAM|20|19|到第三日，就要走一段長路下去 ，去到你遇事那天所藏的地方，在 以色 磐石 的旁邊等候。
1SAM|20|20|我會向磐石旁邊射三箭，如同射箭靶一樣。
1SAM|20|21|看哪，我會派僮僕，說：『去把箭找來。』我若對僮僕喊說：『看哪，箭在你的這邊，把箭拿來』，你就可以平安回來；我指著永生的耶和華起誓，你一定沒有事。
1SAM|20|22|我若對孩子說：『看哪，箭在你的前方』，你就要離開，因為是耶和華差你去的。
1SAM|20|23|至於你和我，我們所說的話，看哪，耶和華在你我中間作證，直到永遠。」
1SAM|20|24|大衛 就去藏在田野。到了初一，王要坐席用餐。
1SAM|20|25|王照常坐在靠牆的位子上， 約拿單 在對面 ， 押尼珥 坐在 掃羅 旁邊， 大衛 的座位卻是空的。
1SAM|20|26|這日 掃羅 沒有說甚麼，因為他說：「 大衛 或許有事，偶染不潔，還未得潔淨。」
1SAM|20|27|初二， 大衛 的座位還空著。 掃羅 對他兒子 約拿單 說：「 耶西 的兒子為何昨日、今日都沒有來用餐呢？」
1SAM|20|28|約拿單 回答 掃羅 說：「 大衛 懇求我允許他回 伯利恆 去，
1SAM|20|29|說：『求你讓我去，因為我家在城裏有獻祭的事，我哥哥吩咐我去。如今我若在你眼前蒙恩，求你讓我去見我的兄弟。』所以 大衛 沒有來赴王的筵席。」
1SAM|20|30|掃羅 向 約拿單 怒氣大發，對他說：「你這頑梗悖逆之婦人所生的，我怎麼會不知道你選擇 耶西 的兒子 ，自取羞辱，也使你母親露體蒙羞呢？
1SAM|20|31|只要 耶西 的兒子還活在世上一天，你和你的國必保不住。現在你要派人去，把他帶到我這裏來，因為他是該死的。」
1SAM|20|32|約拿單 回答父親 掃羅 說：「他為甚麼該死呢？他做了甚麼呢？」
1SAM|20|33|掃羅 向 約拿單 擲槍要刺他， 約拿單 就知道他父親決意要殺死 大衛 。
1SAM|20|34|於是 約拿單 氣憤憤地從席上起來。他在初二這天沒有吃飯，因為他為 大衛 愁煩，又因為他父親羞辱了他。
1SAM|20|35|次日早晨， 約拿單 按著與 大衛 約定的時候到田野去，有一個小僮僕跟隨他。
1SAM|20|36|約拿單 對僮僕說：「你跑去把我所射的箭找來。」僮僕跑去， 約拿單 就把箭射在僮僕的前方。
1SAM|20|37|僮僕到了 約拿單 落箭之地， 約拿單 呼叫僮僕說：「箭不是在你的前方嗎？」
1SAM|20|38|約拿單 又呼叫僮僕說：「快去，不要站在那裏！」僮僕就撿起箭來，回到主人那裏。
1SAM|20|39|僮僕不知道這是甚麼意思，只有 約拿單 和 大衛 知道這事。
1SAM|20|40|約拿單 把他的弓箭交給僮僕，吩咐他說：「你拿到城裏去。」
1SAM|20|41|僮僕一去， 大衛 就從南邊 出來，俯伏在地，拜了三拜。他們彼此親吻，一起哭泣， 大衛 哭得更悲哀。
1SAM|20|42|約拿單 對 大衛 說：「你平平安安地去吧！因為我們二人曾指著耶和華的名起誓說：『願耶和華在你我中間，以及你我後裔中間作證，直到永遠。』」 大衛 就起身走了， 約拿單 也回城裏去了。
1SAM|21|1|大衛 到了 挪伯 的 亞希米勒 祭司那裏， 亞希米勒 戰戰兢兢地出來迎接他，對他說：「你為甚麼獨自一人，沒有人跟隨你呢？」
1SAM|21|2|大衛 對 亞希米勒 祭司說：「王吩咐我一件事，對我說：『我差遣你，吩咐你的這件事，不可讓任何人知道。』因此我已告訴一些僕人到某處去 。
1SAM|21|3|現在你手中有甚麼？請你給我五個餅或是可以找到的食物。」
1SAM|21|4|祭司對 大衛 說：「我手中沒有普通的餅，只有聖餅，只能給沒有親近婦人的年輕人。」
1SAM|21|5|大衛 回答祭司說：「我們確實沒有親近婦人，如同往常我出征的時候一樣。平常行路，僕人的身體 都還分別為聖，何況今日豈不更使自己分別為聖嗎？」
1SAM|21|6|祭司拿聖餅給他，因為在那裏沒有別的餅，只有那從耶和華面前撤下的供餅，就是換上熱餅的日子取下來的。
1SAM|21|7|當日，有 掃羅 的一個臣僕在那裏，他留在耶和華的面前，名叫 多益 ，是 以東 人，作 掃羅 的畜牧長。
1SAM|21|8|大衛 對 亞希米勒 說：「你手中有沒有槍或刀？因為王的事緊急，連刀劍兵器我都沒有帶。」
1SAM|21|9|祭司說：「你在 以拉谷 所殺的 非利士 人 歌利亞 的那刀，看哪，裹在布中，放在以弗得後邊。你若要可以拿去，除此以外，再沒有別的了。」 大衛 說：「沒有甚麼可以跟它比的了！請你給我。」
1SAM|21|10|那日 大衛 起來，躲避 掃羅 ，逃到 迦特 王 亞吉 那裏。
1SAM|21|11|亞吉 的臣僕對他說：「這不是那地的國王 大衛 嗎？那裏的人跳舞唱和： 『 掃羅 殺死千千， 大衛 殺死萬萬』， 不是指著他說的嗎？」
1SAM|21|12|大衛 把這些話放在心裏，就很懼怕 迦特 王 亞吉 。
1SAM|21|13|於是他在眾人眼前一反常態，在他們中間 裝瘋作癲，在城門的門扇上胡寫亂畫，任由唾沫流在鬍子上。
1SAM|21|14|亞吉 對臣僕說：「看哪，你們看這人瘋了，為甚麼帶他到我這裏來呢？
1SAM|21|15|我豈缺少瘋子，你們竟然帶這人到我面前瘋癲嗎？這個人可以進我的家嗎？」
1SAM|22|1|大衛 離開那裏，逃到 亞杜蘭 洞。他的兄弟和他父親全家聽見了，都下到他那裏去。
1SAM|22|2|凡生活窘迫的、欠債的、心裏苦惱的都聚集到 大衛 那裏，他就作他們的領袖，跟隨他的約有四百人。
1SAM|22|3|大衛 從那裏往 摩押 的 米斯巴 去，對 摩押 王說：「請你讓我父母搬來，跟你們在一起，等我知道上帝要為我怎樣做。」
1SAM|22|4|大衛 領他父母到 摩押 王面前。 大衛 住山寨一切的日子，他父母也都住在 摩押 王那裏。
1SAM|22|5|先知 迦得 對 大衛 說：「你不要住在山寨，要到 猶大 地去。」 大衛 就去，來到 哈列 的樹林。
1SAM|22|6|掃羅 聽見 大衛 和跟隨他之人的下落， 掃羅 正在 基比亞 ，坐在山頂 的柳樹下，手裏拿著槍，眾臣僕侍立在左右。
1SAM|22|7|掃羅 對左右侍立的臣僕說：「 便雅憫 人哪，聽著！ 耶西 的兒子也能把田地和葡萄園賜給你們各人嗎？他能立你們各人作千夫長和百夫長嗎？
1SAM|22|8|你們竟都結黨害我！我兒子與 耶西 的兒子立約的時候，無人告訴我；我兒子挑唆我的臣僕謀害我，像今日這樣，也無人告訴我，為我憂慮。」
1SAM|22|9|那時 以東 人 多益 站在 掃羅 的臣僕中，回答說：「我曾看見 耶西 的兒子往 挪伯 去，到了 亞希突 的兒子 亞希米勒 那裏。
1SAM|22|10|亞希米勒 為他求問耶和華，給他食物，又把 非利士 人 歌利亞 的刀給了他。」
1SAM|22|11|王就派人把 亞希突 的兒子 亞希米勒 祭司和他父親的全家，就是在 挪伯 的祭司都召了來，他們都來到王那裏。
1SAM|22|12|掃羅 說：「 亞希突 的兒子，聽著！」他說：「我主，我在這裏。」
1SAM|22|13|掃羅 對他說：「你為甚麼與 耶西 的兒子結黨害我，把食物和刀給他，又為他求問上帝，使他起來謀害我，像今日這樣？」
1SAM|22|14|亞希米勒 回答王說：「王的眾臣僕中有誰比 大衛 忠心呢？他是王的女婿，又是你的侍衛長 ，並且是你宮中受敬重的人。
1SAM|22|15|我今日才開始為他求問上帝嗎？絕非如此！王不要歸罪於我和我父全家，因為這事，無論大小，僕人都不知情。」
1SAM|22|16|王說：「 亞希米勒 ，你和你父全家都是該死的！」
1SAM|22|17|王吩咐左右的侍衛說：「你們轉身去殺耶和華的祭司吧！因為他們幫助 大衛 ，知道 大衛 逃跑卻不告訴我。」但王的臣僕都不願動手殺耶和華的祭司。
1SAM|22|18|王吩咐 多益 說：「你轉身去殺祭司吧！」 以東 人 多益 就轉身去殺祭司，那日殺了穿細麻布以弗得的，共八十五人，
1SAM|22|19|又用刀把祭司城 挪伯 中的男女、孩童和吃奶的都殺了，又用刀殺了牛、羊和驢子。
1SAM|22|20|亞希突 的兒子 亞希米勒 有一個兒子逃脫了；他名叫 亞比亞他 ，逃到 大衛 那裏。
1SAM|22|21|亞比亞他 把 掃羅 殺耶和華祭司的事告訴 大衛 。
1SAM|22|22|大衛 對 亞比亞他 說：「那日我見 以東 人 多益 在那裏，就知道他一定會告訴 掃羅 。你父的全家喪命，都是因我的緣故。
1SAM|22|23|你可以住在我這裏，不要懼怕。因為尋索你命的也要尋索我的命，你在我這裏可得保護。」
1SAM|23|1|有人告訴 大衛 說：「看哪， 非利士 人攻擊 基伊拉 ，搶奪禾場。」
1SAM|23|2|大衛 求問耶和華說：「我可以去嗎？我可以去攻打那些 非利士 人嗎？」耶和華對 大衛 說：「你可以去攻打 非利士 人，拯救 基伊拉 。」
1SAM|23|3|大衛 的人對他說：「看哪，我們在 猶大 這裏尚且懼怕，何況到 基伊拉 去攻打 非利士 人的軍隊呢？」
1SAM|23|4|大衛 又再求問耶和華，耶和華回答說：「你起身下 基伊拉 去，我必將 非利士 人交在你手裏。」
1SAM|23|5|於是 大衛 和他的人往 基伊拉 去，與 非利士 人打仗，大大擊敗他們，奪取他們的牲畜。這樣， 大衛 救了 基伊拉 的居民。
1SAM|23|6|亞希米勒 的兒子 亞比亞他 逃往 基伊拉 到 大衛 那裏的時候，手裏拿著以弗得。
1SAM|23|7|有人告訴 掃羅 ， 大衛 到了 基伊拉 。 掃羅 說：「上帝將他交在我手裏了，因為他進了有門有閂的城，把自己關起來了。」
1SAM|23|8|於是 掃羅 召集眾百姓，要下去攻打 基伊拉 ，圍困 大衛 和他的人。
1SAM|23|9|大衛 知道 掃羅 設計陷害他，就對 亞比亞他 祭司說：「把以弗得拿過來。」
1SAM|23|10|大衛 說：「耶和華－ 以色列 的上帝啊，你僕人確實聽見 掃羅 設法要到 基伊拉 來，為我的緣故毀滅這城。
1SAM|23|11|基伊拉 人會把我交在 掃羅 手裏嗎？ 掃羅 會下來，正如你僕人所聽見的嗎？耶和華－ 以色列 的上帝啊，求你指示僕人！」耶和華說：「他會下來。」
1SAM|23|12|大衛 又說：「 基伊拉 人會把我和我的人交在 掃羅 手裏嗎？」耶和華說：「他們會交出來。」
1SAM|23|13|於是 大衛 和他的人約有六百名起身離開 基伊拉 ，往他們所能去的地方去。有人告訴 掃羅 ， 大衛 離開 基伊拉 逃走了， 掃羅 就停止出發了。
1SAM|23|14|大衛 住在曠野的山寨裏，在 西弗 曠野的山區。 掃羅 天天尋索 大衛 ，上帝卻不將 大衛 交在他手裏。
1SAM|23|15|大衛 看到 掃羅 出來尋索他的命。那時，他住在 西弗 曠野的樹林裏 ；
1SAM|23|16|掃羅 的兒子 約拿單 起身，到樹林裏去見 大衛 ，使他的手倚靠上帝得以堅固，
1SAM|23|17|對他說：「不要懼怕！我父 掃羅 的手無法害你 ，你必作 以色列 的王，我必作你的宰相。我父 掃羅 也知道這事。」
1SAM|23|18|於是二人在耶和華面前立約。 大衛 仍住在樹林裏， 約拿單 就回家去了。
1SAM|23|19|西弗 人上 基比亞 到 掃羅 那裏，說：「 大衛 不是在我們那裏，在樹林裏的山寨中，在荒野 南邊的 哈基拉山 藏著嗎？
1SAM|23|20|現在，王啊，請隨你的心願要下來，就請下來；至於我們，一定會把他交在王的手裏。」
1SAM|23|21|掃羅 說：「願耶和華賜福給你們，因為你們體恤我。
1SAM|23|22|請你們回去，再確定一下，調查並看清楚他落腳的地方，是誰看見他在那裏 ，因為有人告訴我他很狡猾。
1SAM|23|23|你們要看清楚，調查他藏匿的每一個地方，回來給我確實的報告，我就與你們同去。他若在境內，我必從 猶大 的千門萬戶中搜出他來。」
1SAM|23|24|西弗 人動身，在 掃羅 以先往 西弗 去。 大衛 和他的人卻在 瑪雲 曠野，在荒野南邊的 亞拉巴 。
1SAM|23|25|掃羅 和他的人去尋索 大衛 。有人告訴 大衛 ，他就下到巖石那裏，留在 瑪雲 的曠野。 掃羅 聽見了，就在 瑪雲 的曠野追趕 大衛 。
1SAM|23|26|掃羅 在山的這一邊走， 大衛 和他的人在山的那一邊。 大衛 急忙躲避 掃羅 ， 掃羅 和他的人正四面圍住 大衛 和他的人，要捉拿他們。
1SAM|23|27|有使者來對 掃羅 說：「 非利士 人入境搶掠，請快快回去！」
1SAM|23|28|於是 掃羅 不再追趕 大衛 ，回去迎擊 非利士 人。因此那地方名叫 西拉‧哈瑪希羅結 。
1SAM|23|29|大衛 從那裏上去，住在 隱‧基底 的山寨裏。
1SAM|24|1|掃羅 追趕 非利士 人回來，有人告訴他說：「看哪， 大衛 在 隱‧基底 的曠野。」
1SAM|24|2|掃羅 就從全 以色列 中挑選三千精兵，往 野山羊磐石 的東邊 去，尋索 大衛 和他的人。
1SAM|24|3|到了路旁的羊圈，在那裏有個洞， 掃羅 進去大解。 大衛 和他的人正藏在洞裏的深處。
1SAM|24|4|大衛 的人對 大衛 說：「看哪，這日子到了！耶和華曾對你說：『看哪，我要將你的仇敵交在你手裏，你可以照你看為好的對待他。』」 大衛 就起來，悄悄地割下 掃羅 外袍的衣角。
1SAM|24|5|隨後 大衛 心中自責，因為他割下了 掃羅 的衣角。
1SAM|24|6|他對他的人說：「耶和華絕不允許我對我的主，耶和華的受膏者做這事，伸手害他，因為他是耶和華的受膏者。」
1SAM|24|7|大衛 用這話勸阻他的人，不許他們起來害 掃羅 。 掃羅 起來，從洞裏出去，預備上路。
1SAM|24|8|然後 大衛 也起來，從洞裏出去，呼喚 掃羅 說：「我主，我王！」 掃羅 回頭觀看， 大衛 就屈身，臉伏於地下拜。
1SAM|24|9|大衛 對 掃羅 說：「你為何聽信人的讒言，說『看哪， 大衛 想要害你』呢？
1SAM|24|10|看哪，今日你親眼看見，在洞中耶和華將你交在我手裏。有人要我殺你，我卻愛惜你，說：『我不敢伸手害我的主，因為他是耶和華的受膏者。』
1SAM|24|11|我父啊，請看，看你外袍的衣角在我手中。我割下你外袍的衣角，卻沒有殺你。你知道，並且看見我沒有惡意要悖逆你。你雖然要獵取我的命，我卻沒有得罪你。
1SAM|24|12|願耶和華在你我中間判斷，願耶和華在你身上為我伸冤，我卻不親手加害於你。
1SAM|24|13|古人有句俗語說：『惡事出於惡人。』我卻不親手加害於你。
1SAM|24|14|以色列 王出來要尋找誰呢？你要追趕誰呢？不過是一條死狗，一隻跳蚤而已。
1SAM|24|15|願耶和華作仲裁者，在你我中間判斷。願他鑒察，為我伸冤，救我脫離你的手。」
1SAM|24|16|大衛 向 掃羅 說完了這些話， 掃羅 說：「我兒 大衛 ，這是你的聲音嗎？」於是 掃羅 放聲大哭，
1SAM|24|17|對 大衛 說：「你比我公義，因為你以善待我，我卻以惡待你。
1SAM|24|18|今日你已顯明是以善待我，因為耶和華將我交在你手裏，你卻沒有殺我。
1SAM|24|19|人若遇見仇敵，豈肯放他平安上路呢？願耶和華因你今日向我所做的，以善回報你。
1SAM|24|20|現在，看哪，我知道你一定會作王， 以色列 的國必要堅立在你手裏。
1SAM|24|21|現在你要指著耶和華向我起誓，你必不剪除我的後裔，必不從我父家除去我的名。」
1SAM|24|22|於是 大衛 向 掃羅 起誓， 掃羅 就回家去， 大衛 和他的人也上山寨去了。
1SAM|25|1|撒母耳 死了， 以色列 眾人聚集，為他哀哭，把他葬在 拉瑪 他的家裏。 大衛 動身，下到 巴蘭 的曠野。
1SAM|25|2|在 瑪雲 有一個人，他的產業在 迦密 。這人是一個大富翁，有三千隻綿羊，一千隻山羊；他正在 迦密 剪羊毛。
1SAM|25|3|這人名叫 拿八 ，他的妻子名叫 亞比該 。 拿八 的妻子有美好的見識，又有美麗的容貌，但 拿八 為人剛愎兇惡，是 迦勒 族的人。
1SAM|25|4|大衛 在曠野聽見 拿八 正在剪羊毛，
1SAM|25|5|就派十個僕人，對他們說：「你們上 迦密 到 拿八 那裏，提我的名向他問安。
1SAM|25|6|你們要如此說：『願你來年平安 ，願你家平安，願你一切所有的都平安。
1SAM|25|7|現在我聽說你有剪羊毛的人，你的牧人和我們在一起，他們在 迦密 一切的日子，我們沒有欺負過他們，他們也未曾失去甚麼。
1SAM|25|8|你問你的僕人，他們會告訴你。願我的僕人在你眼前得歡心，因為我們是在好日子來的。請你隨手分點食物給僕人和你兒子 大衛 。』」
1SAM|25|9|大衛 的僕人到了，就提 大衛 的名，把這一切話告訴 拿八 ，他們就停頓下來。
1SAM|25|10|拿八 回答 大衛 的僕人說：「 大衛 是誰？ 耶西 的兒子是誰？今日悖逆主人奔逃的僕人很多。
1SAM|25|11|我豈可把飲食，以及我為剪羊毛的人所宰的肉給那些我不知道從哪裏來的人呢？」
1SAM|25|12|大衛 的僕人轉身從原路回去，照這一切的話告訴 大衛 。
1SAM|25|13|大衛 對他的人說：「你們各人都要佩上刀！」各人就都佩上刀， 大衛 也佩上刀。跟隨 大衛 上去的約有四百人，留下二百人看守物件。
1SAM|25|14|拿八 的一個僕人告訴 拿八 的妻子 亞比該 說：「看哪， 大衛 從曠野派使者來向我主人問安，主人卻辱罵他們。
1SAM|25|15|但是那些人待我們真好；我們在田野與他們一切來往的日子，沒有受他們欺負，也未曾失去甚麼。
1SAM|25|16|我們在他們那裏牧羊，一切的日子他們晝夜保護我們 。
1SAM|25|17|現在，你當知道，看怎樣做才好。不然，禍患必定臨到我主人和他全家。他性情兇暴，無人敢與他說話。」
1SAM|25|18|亞比該 急忙將二百個餅，兩皮袋酒，五隻宰好的羊，五細亞烘熟的穗子，一百個葡萄乾餅，二百個無花果餅，都馱在驢上，
1SAM|25|19|對僕人說：「你們在我前面走，看哪，我跟著你們去。」她卻沒有告訴丈夫 拿八 。
1SAM|25|20|亞比該 騎著驢，正下山坡，看哪， 大衛 和他的人正迎著 亞比該 下來，她就去迎接他們。
1SAM|25|21|大衛 曾說：「我在曠野為那人看守他一切所有的，以致他未失去任何一樣東西，實在是徒然了！他竟然向我以惡報善。
1SAM|25|22|凡屬 拿八 的男丁，我若留一個到明日早晨，願上帝重重懲罰 大衛 ！」
1SAM|25|23|亞比該 看見 大衛 ，就急忙下驢，在 大衛 面前臉伏於地叩拜。
1SAM|25|24|她俯伏在 大衛 的腳前，說：「我主啊，願這罪歸於我！求你容許使女向你進言，更求你聽使女的話。
1SAM|25|25|我主不必理會 拿八 這性情兇暴的人，他就像他的名字一樣；他名叫 拿八 ，為人也真是愚頑。至於我，你的使女並沒有看見我主所派來的僕人。
1SAM|25|26|現在，我主啊，耶和華既然阻止你親手報仇，避免流人的血，我指著永生的耶和華起誓，又指著你的性命起誓：『現在，願你的仇敵和謀害我主的人都像 拿八 一樣。』
1SAM|25|27|現在求我主把婢女送來的禮物給跟隨我主的僕人。
1SAM|25|28|求你原諒使女的冒犯。耶和華必為我主建立堅固的家，因為我主為耶和華爭戰，並且你一生的日子查不出有甚麼惡來。
1SAM|25|29|雖有人起來追逼你，要尋索你的性命，我主的性命在耶和華－你的上帝那裏，如同藏在生命的寶藏中。至於你仇敵的性命，耶和華必甩去，如用機弦甩石一樣。
1SAM|25|30|耶和華照所應許你的福氣賜給我主，立你作 以色列 王的時候，
1SAM|25|31|我主就不至於因為親手報仇，流了無辜人的血，而心裏不安，良心有虧了。耶和華賜福給我主的時候，求你記得你的使女。」
1SAM|25|32|大衛 對 亞比該 說：「耶和華－ 以色列 的上帝是應當稱頌的，因為他今日派你來迎接我。
1SAM|25|33|你和你的見識也配得稱讚，因為你今日攔阻我親手報仇、流人的血。
1SAM|25|34|我指著阻止我加害於你的耶和華－ 以色列 永生的上帝起誓，若不是你很快地來迎接我，到早晨天亮的時候，凡屬 拿八 的男丁，必定一個也不留。」
1SAM|25|35|大衛 從 亞比該 手中收了她帶來的禮物，對她說：「平平安安上你的家去吧！你看，我看了你的情面，聽了你的話。」
1SAM|25|36|亞比該 到 拿八 那裏，看哪，他在家裏擺設宴席，如同王的宴席。 拿八 心情舒暢，酩酊大醉。所以 亞比該 大小事都沒有告訴他，直等到早晨天亮的時候。
1SAM|25|37|到了早晨， 拿八 酒醒了，他的妻子把這些事都告訴他，他就發心臟病快死了，僵如石頭。
1SAM|25|38|過了十天，耶和華擊打 拿八 ，他就死了。
1SAM|25|39|大衛 聽見 拿八 死了，就說：「耶和華是應當稱頌的，因為我從 拿八 手中受了羞辱，他為我伸冤，又阻止他的僕人行惡；耶和華使 拿八 的惡歸到他自己頭上。」於是 大衛 派人去向 亞比該 說，要娶她為妻。
1SAM|25|40|大衛 的僕人來到 迦密 ，到 亞比該 那裏，對她說：「 大衛 派我們到你這裏，要娶你作他的妻子。」
1SAM|25|41|亞比該 起來叩拜，俯伏在地，說：「看哪，你的使女情願作婢女，為我主的僕人洗腳。」
1SAM|25|42|亞比該 立刻起身，騎上驢，五個女僕跟著她走。她跟從 大衛 的使者去，就作了 大衛 的妻子。
1SAM|25|43|大衛 先前娶了 耶斯列 人 亞希暖 ，她們二人都作了他的妻子。
1SAM|25|44|掃羅 已把他的女兒 米甲 ，就是 大衛 的妻子，給了 迦琳 人 拉億 的兒子 帕提 為妻。
1SAM|26|1|西弗 人來到 基比亞 ，到 掃羅 那裏，說：「 大衛 不是在荒野 東邊 的 哈基拉山 藏著嗎？」
1SAM|26|2|掃羅 動身，帶領 以色列 人中挑選的三千精兵下到 西弗 的曠野，要在那裏尋索 大衛 。
1SAM|26|3|掃羅 在荒野東邊的 哈基拉山 ，在路旁安營。那時 大衛 住在曠野，看見 掃羅 到曠野來追趕他，
1SAM|26|4|大衛 就派人去探聽，知道 掃羅 果然來了。
1SAM|26|5|大衛 起來，到 掃羅 安營的地方，看見 掃羅 和 尼珥 的兒子 押尼珥 元帥躺臥之處； 掃羅 睡在軍營裏，士兵安營在他周圍。
1SAM|26|6|大衛 對 赫 人 亞希米勒 和 洗魯雅 的兒子 約押 的兄弟 亞比篩 說：「誰同我下到 掃羅 營裏去？」 亞比篩 說：「我同你下去。」
1SAM|26|7|於是 大衛 和 亞比篩 夜間到了士兵那裏；看哪， 掃羅 睡在軍營裏，他的槍在頭旁，插在地上。 押尼珥 和士兵睡在他周圍。
1SAM|26|8|亞比篩 對 大衛 說：「上帝將你的仇敵交在你手裏，現在讓我拿槍把他刺透在地上，一刺就成，不用再刺他了。」
1SAM|26|9|大衛 對 亞比篩 說：「不可殺害他！有誰伸手害耶和華的受膏者而無罪呢？」
1SAM|26|10|大衛 又說：「我指著永生的耶和華起誓，他或被耶和華擊殺，或死期到了，或出戰陣亡，
1SAM|26|11|耶和華絕不允許我伸手害耶和華的受膏者。現在你可以把他頭旁的槍和水壺拿來，我們就走。」
1SAM|26|12|大衛 從 掃羅 的頭旁拿了槍和水壺，他們就走了。沒有人看見，沒有人知道，也沒有人醒過來。他們都睡著了，因為耶和華使他們沉睡了。
1SAM|26|13|大衛 過到另一邊去，遠遠地站在山頂上，與他們相離很遠。
1SAM|26|14|大衛 呼叫百姓和 尼珥 的兒子 押尼珥 說：「 押尼珥 ，你為何不回答呢？」 押尼珥 回答說：「你是誰？竟敢呼喚王呢？」
1SAM|26|15|大衛 對 押尼珥 說：「你不是個大丈夫嗎？ 以色列 中誰能比你呢？百姓中有一個人進來要害死你主你王，你為何沒有保護你主你王呢？
1SAM|26|16|你做的這件事不好！我指著永生的耶和華起誓，你們都是該死的，因為你們沒有保護你們的主，就是耶和華的受膏者。現在你看，王頭旁的槍和水壺在哪裏？」
1SAM|26|17|掃羅 認出 大衛 的聲音，就說：「我兒 大衛 ，這是你的聲音嗎？」 大衛 說：「我主我王啊，是我的聲音。」
1SAM|26|18|又說：「我主為何要追趕僕人呢？我做了甚麼？我手做了甚麼惡事呢？
1SAM|26|19|現在求我主我王聽僕人的話：若是耶和華激發你來攻擊我，願耶和華悅納供物；若是出於人，願他們在耶和華面前受詛咒，因為他們今日趕逐我，不讓我在耶和華的產業中有分，說：『你去事奉別神吧！』
1SAM|26|20|現在不要使我的血流在遠離耶和華面的地上。因為 以色列 王出來，只不過是尋找一隻跳蚤，如同人在山上獵取一隻鷓鴣。」
1SAM|26|21|掃羅 說：「我有罪了！我兒 大衛 ，回來吧！我必不再加害於你，因為你今日看我的性命為寶貴。看哪，我是個糊塗人，大大錯了。」
1SAM|26|22|大衛 回答說：「看哪，這是王的槍，可以吩咐一個僕人過來拿去。
1SAM|26|23|今日耶和華將王交在我手裏，我卻不肯伸手害耶和華的受膏者。耶和華必照各人的公義誠實報應他。
1SAM|26|24|看哪，我今日看重你的性命，願耶和華也照樣看重我的性命，並且拯救我脫離一切患難。」
1SAM|26|25|掃羅 對 大衛 說：「我兒 大衛 ，願你得福！你必做大事，也必得勝。」於是 大衛 上路， 掃羅 也回自己的地方去了。
1SAM|27|1|大衛 心裏說：「總有一天我會死在 掃羅 手裏，現在我最好逃到 非利士 人的地去， 掃羅 就會絕望，不會繼續在 以色列 全境內尋索我了。這樣，我才可以脫離他的手。」
1SAM|27|2|於是 大衛 動身，和跟隨他的六百人投奔 瑪俄 的兒子 迦特 王 亞吉 去了。
1SAM|27|3|大衛 和他的兩個妻子，就是 耶斯列 人 亞希暖 和作過 拿八 妻子的 迦密 人 亞比該 ，以及他的人，連同各人的眷屬，都住在 迦特 的 亞吉 那裏。
1SAM|27|4|有人告訴 掃羅 ：「 大衛 逃到 迦特 。」 掃羅 就不再尋索他了。
1SAM|27|5|大衛 對 亞吉 說：「我若蒙你看得起，求你在郊外的城鎮中賜我一個地方，讓我住在那裏。僕人何必與王同住京城呢？」
1SAM|27|6|當日 亞吉 把 洗革拉 賜給他，因此 洗革拉 屬於 猶大 王，直到今日。
1SAM|27|7|大衛 在 非利士 人的地，住的期間有一年四個月。
1SAM|27|8|大衛 和他的人上去，侵奪 基述 人、 基色 人、 亞瑪力 人，這些是從 帖蘭 經過 書珥 直到 埃及 地的居民 。
1SAM|27|9|大衛 攻擊那地，無論男女沒有留下一個活口，又奪獲牛、羊、驢、駱駝和衣服，回來到 亞吉 那裏。
1SAM|27|10|亞吉 說：「今日你們沒有去搶奪甚麼地方吧 ？」 大衛 說：「侵奪了 猶大 、 耶拉篾 、 基尼 等地的南方。」
1SAM|27|11|無論男女， 大衛 沒有留下一個活口帶到 迦特 來。他說：「恐怕他們把我們的事告訴人，說：『 大衛 如此做了。』」這是他住在 非利士 人之地一切日子的慣例。
1SAM|27|12|亞吉 信了 大衛 ，說：「 大衛 已經使本族 以色列 人憎惡他，所以他必永遠作我的僕人了。」
1SAM|28|1|那時， 非利士 人召集軍隊，要與 以色列 打仗。 亞吉 對 大衛 說：「你當知道，你和你的人都要隨我出征。」
1SAM|28|2|大衛 對 亞吉 說：「好，僕人所能做的事，王都知道。」 亞吉 對 大衛 說：「好，我立你終生作我 的侍衛。」
1SAM|28|3|那時 撒母耳 已經死了， 以色列 眾人為他哀哭，把他葬在他的本城 拉瑪 。 掃羅 曾在國內驅除招魂的和行巫術的人。
1SAM|28|4|非利士 人集合，來到 書念 安營； 掃羅 集合 以色列 眾人在 基利波 安營。
1SAM|28|5|掃羅 看見 非利士 的軍隊，就懼怕，心中大大戰兢。
1SAM|28|6|掃羅 求問耶和華，耶和華卻不藉夢，或烏陵，或先知回答他。
1SAM|28|7|掃羅 吩咐臣僕說：「為我找一個招魂的婦人，我好去問她。」臣僕對他說：「看哪，在 隱‧多珥 有一個招魂的婦人。」
1SAM|28|8|於是 掃羅 改了裝，穿上別的衣服，帶著兩個人，夜裏去見那婦人。 掃羅 說：「請你用招魂的法術，把我所告訴你的死人，為我招上來。」
1SAM|28|9|婦人對他說：「看哪，你知道 掃羅 所做的，他從國中剪除招魂的和行巫術的。你為何為我的性命設下羅網，要害死我呢？」
1SAM|28|10|掃羅 向婦人指著耶和華起誓說：「我指著永生的耶和華起誓，你必不因這事受罰。」
1SAM|28|11|婦人說：「我為你招誰上來呢？」他說：「為我招 撒母耳 上來。」
1SAM|28|12|婦人看見 撒母耳 ，就大聲喊叫。婦人對 掃羅 說：「你是 掃羅 ，為甚麼欺騙我呢？」
1SAM|28|13|王對婦人說：「不要懼怕，你看見甚麼呢？」婦人對 掃羅 說：「我看見有神明從地裏上來。」
1SAM|28|14|掃羅 說：「他是怎樣的形狀？」婦人說：「有一個老人上來，身穿長袍。」 掃羅 知道是 撒母耳 ，就屈身，臉伏於地下拜。
1SAM|28|15|撒母耳 對 掃羅 說：「你為甚麼攪擾我，招我上來呢？」 掃羅 說：「我十分為難，因為 非利士 人攻擊我，上帝離開我，不再藉先知或夢回答我。因此請你上來，好指示我應當怎樣做。」
1SAM|28|16|撒母耳 說：「耶和華已經離開你，與你為敵，你何必問我呢？
1SAM|28|17|耶和華照他藉我所說的話為他自己 實現了。耶和華已經從你手裏奪去國權，賜給別人，就是 大衛 。
1SAM|28|18|因為你沒有聽從耶和華的話，沒有執行他對 亞瑪力 人的惱怒，所以今日耶和華向你做這事。
1SAM|28|19|耶和華也必將你和 以色列 交在 非利士 人手裏。明日你和你兒子們必與我在一處了；耶和華也必將 以色列 的軍兵交在 非利士 人手裏。」
1SAM|28|20|掃羅 突然全身仆倒在地，因為 撒母耳 的話令他十分懼怕。他毫無氣力，因為他一日一夜都沒有吃甚麼。
1SAM|28|21|婦人到 掃羅 面前，見他極其驚恐，對他說：「看哪，婢女聽從了你，不顧惜自己的性命，遵從你吩咐我的話。
1SAM|28|22|現在求你也聽婢女的話，讓我在你面前擺上一點食物，你吃了才有氣力上路。」
1SAM|28|23|掃羅 不肯，說：「我不吃。」但他的僕人和那婦人再三勸他，他才聽他們的話，從地上起來，坐在床上。
1SAM|28|24|婦人急忙把家裏的一隻肥牛犢宰了，又拿麵來揉，烤成無酵餅，
1SAM|28|25|擺在 掃羅 和他僕人面前。他們吃了，當夜就起身走了。
1SAM|29|1|非利士 人聚集他們所有的軍隊到 亞弗 ； 以色列 人在 耶斯列 的泉旁安營。
1SAM|29|2|非利士 人的領袖各率隊伍，或百或千的前進； 大衛 和他的人同 亞吉 跟在後邊前進。
1SAM|29|3|非利士 人的領袖說：「這些 希伯來 人在這裏做甚麼呢？」 亞吉 對 非利士 人的領袖說：「這不是 以色列 王 掃羅 的臣僕 大衛 嗎？他在我這裏有些年日了。自從他投降直到今日，我未曾見他有甚麼過錯。」
1SAM|29|4|非利士 人的領袖向 亞吉 發怒，對他說：「叫這人回去！叫他回到你指派他的地方去，不可讓他同我們出征，免得他在陣上反成為我們的敵人。他用甚麼與他主人復和呢？豈不是用我們這些人的首級嗎？
1SAM|29|5|有人跳舞唱和說： 『 掃羅 殺死千千， 大衛 殺死萬萬』， 不就是這個 大衛 嗎？」
1SAM|29|6|亞吉 叫 大衛 來，對他說：「我指著永生的耶和華起誓，你是個正直人。你隨我在軍中出入，我也很滿意。自從你投奔我到如今，我未曾看見你有甚麼過失，但是眾領袖看你不順眼。
1SAM|29|7|現在你平平安安地回去，不要做 非利士 人領袖眼中看為惡的事。」
1SAM|29|8|大衛 對 亞吉 說：「但我做了甚麼呢？自從僕人到你面前，直到今日，你查出我有甚麼過錯，使我不去攻擊我主我王的仇敵呢？」
1SAM|29|9|亞吉 回答 大衛 說：「我知道你在我眼中是好人，如同上帝的使者一樣，只是 非利士 人的領袖說：『這人不可同我們上戰場。』
1SAM|29|10|現在，你和跟隨你來的，就是你主人的僕人，清晨要早早起來，回到我所指派你的地方去，不要把中傷的話放在心上，因為你在我面前很好 。你們清晨早早起來，天一亮就回去吧！」
1SAM|29|11|於是 大衛 和他的人清晨早早起來，回到 非利士 人的地去。 非利士 人也上 耶斯列 去了。
1SAM|30|1|第三日， 大衛 和他的人到了 洗革拉 。 亞瑪力 人已經侵奪 尼革夫 和 洗革拉 。他們攻破 洗革拉 ，用火焚燒。
1SAM|30|2|他們擄去城內的婦女和城中的大小人口，一個都沒有殺，全都帶走，他們就上路去了。
1SAM|30|3|大衛 和他的人到了那城，看哪，城已被火燒燬，他們的妻子兒女都被擄去了。
1SAM|30|4|大衛 和跟隨他的百姓就放聲大哭，直到沒有氣力再哭。
1SAM|30|5|大衛 的兩個妻子， 耶斯列 人 亞希暖 和作過 拿八 妻子的 迦密 人 亞比該 ，也被擄去了。
1SAM|30|6|大衛 非常焦急，因為眾百姓為自己的兒女痛心，說要用石頭打死他。 大衛 卻倚靠耶和華－他的上帝，堅定自己。
1SAM|30|7|大衛 對 亞希米勒 的兒子 亞比亞他 祭司說：「請你把以弗得拿來給我。」 亞比亞他 就把以弗得拿給 大衛 。
1SAM|30|8|大衛 求問耶和華說：「我追趕這群人，是否追得上呢？」耶和華對他說：「你可以追，一定追得上，也一定救得回來。」
1SAM|30|9|於是， 大衛 出發，他和跟隨他的六百人來到 比梭溪 ，那些不能前去的就留在那裏。
1SAM|30|10|大衛 帶著四百人往前追趕；有二百人疲乏，不能過 比梭溪 ，留在那裏。
1SAM|30|11|這四百人在田野遇見一個 埃及 人，就帶他到 大衛 面前，給他餅吃，給他水喝，
1SAM|30|12|又給他一塊無花果餅，兩個葡萄乾餅。他吃了，精神就恢復了，因為他三日三夜沒有吃餅，沒有喝水。
1SAM|30|13|大衛 對他說：「你是誰的人？你從哪裏來？」他說：「我是 埃及 的青年，是 亞瑪力 人的奴僕。因為我三天前生病，我主人就把我撇棄了。
1SAM|30|14|我們侵奪了 基利提 的南方和屬 猶大 的地，以及 迦勒 地的南方，又用火燒了 洗革拉 。」
1SAM|30|15|大衛 對他說：「你肯領我們下到那群人那裏嗎？」他說：「你要向我指著上帝起誓，你不殺我，也不把我交在我主人手裏，我就領你下到那群人那裏。」
1SAM|30|16|那人領 大衛 下去，看哪，他們分散在全地面，吃喝跳舞，因為他們從 非利士 人的地和 猶大 地擄來的財物非常多。
1SAM|30|17|大衛 擊殺他們，從黎明直到次日晚上，除了四百個騎駱駝逃走的青年之外，一個也沒有逃脫。
1SAM|30|18|亞瑪力 人所擄去的財物， 大衛 全都奪回，並救回他的兩個妻子。
1SAM|30|19|凡 亞瑪力 人所擄去的，無論大小、兒女、掠物和一切被擄去的， 大衛 全都奪回來。
1SAM|30|20|大衛 所奪來的牛群羊群，有人趕在群畜前面，說：「這是 大衛 的掠物。」
1SAM|30|21|大衛 到了那疲乏不能跟隨、留在 比梭溪 的二百人那裏。他們出來迎接 大衛 和跟隨他的百姓。 大衛 上前向他們問安。
1SAM|30|22|跟隨 大衛 去的人中，每一個惡人和無賴都說：「這些人既然沒有和我同去，我們所奪的財物就不分給他們，只把他們各人的妻子兒女給他們，讓他們帶回去就好了。」
1SAM|30|23|大衛 說：「我的弟兄，耶和華所賜給我們的，你們不可這麼做，因為他保佑了我們，把那群來攻擊我們的人交在我們手裏。
1SAM|30|24|誰肯在這事上聽你們呢？上陣的分得多少，留下看守物件的也分得多少，大家應當平分。」
1SAM|30|25|從那日起， 大衛 定此為 以色列 的律例典章，直到今日。
1SAM|30|26|大衛 到了 洗革拉 ，從掠物中取些送給他的朋友，就是 猶大 的長老，說：「看哪，這是從耶和華仇敵那裏奪來的，送給你們作禮物。」
1SAM|30|27|有在 伯特利 的， 尼革夫 之 拉末 的， 雅提珥 的，
1SAM|30|28|有在 亞羅珥 的， 息末 的， 以實提莫 的，
1SAM|30|29|有在 拉哈勒 的， 耶拉篾 各城的， 基尼 各城的，
1SAM|30|30|有在 何珥瑪 的， 坡拉珊 的， 亞撻 的，
1SAM|30|31|有在 希伯崙 的，以及 大衛 和跟隨他的人經常進出之處的。
1SAM|31|1|非利士 人攻打 以色列 。 以色列 人在 非利士 人面前逃跑，很多人 在 基利波山 被殺仆倒。
1SAM|31|2|非利士 人緊追 掃羅 和他的兒子，殺了 掃羅 的兒子 約拿單 、 亞比拿達 、 麥基‧舒亞 。
1SAM|31|3|攻擊 掃羅 的戰事激烈，弓箭手追上他，他被弓箭手射中，傷勢很重 。
1SAM|31|4|掃羅 吩咐拿他兵器的人說：「你拔出刀來，把我刺死，免得那些未受割禮的人來刺我，凌辱我。」但拿兵器的人不肯，因為他非常懼怕。於是 掃羅 拿起刀來，伏在刀上。
1SAM|31|5|拿兵器的人見 掃羅 已死，也伏在刀上跟他一起死。
1SAM|31|6|這樣， 掃羅 和他三個兒子，與拿他兵器的人，以及他所有的人 ，都在那日一起死了。
1SAM|31|7|住平原那邊和 約旦河 那邊的 以色列 人，見 以色列 軍兵逃跑， 掃羅 和他兒子都死了，就棄城逃跑。 非利士 人前來住在其中。
1SAM|31|8|次日， 非利士 人來剝那些被殺之人的衣服，看見 掃羅 和他三個兒子仆倒在 基利波山 。
1SAM|31|9|他們割下他的首級，剝了他的盔甲，派人到 非利士 人之地的四境，報信給他們廟裏的偶像和百姓。
1SAM|31|10|他們將 掃羅 的盔甲放在 亞斯她錄 廟裏，把他的屍身釘在 伯‧珊 的城牆上。
1SAM|31|11|基列 的 雅比 居民聽見 非利士 人向 掃羅 所行的事，
1SAM|31|12|他們所有的勇士就起身，走了一夜，把 掃羅 和他兒子的屍身從 伯‧珊 城牆上取下來，送到 雅比 ，在那裏用火燒了，
1SAM|31|13|把骸骨葬在 雅比 的柳樹下，並且禁食七日。
