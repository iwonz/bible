1TIM|1|1|Paul, an apostle of Christ Jesus by the command of God our Savior and of Christ Jesus our hope,
1TIM|1|2|To Timothy my true son in the faith: Grace, mercy and peace from God the Father and Christ Jesus our Lord.
1TIM|1|3|As I urged you when I went into Macedonia, stay there in Ephesus so that you may command certain men not to teach false doctrines any longer
1TIM|1|4|nor to devote themselves to myths and endless genealogies. These promote controversies rather than God's work--which is by faith.
1TIM|1|5|The goal of this command is love, which comes from a pure heart and a good conscience and a sincere faith.
1TIM|1|6|Some have wandered away from these and turned to meaningless talk.
1TIM|1|7|They want to be teachers of the law, but they do not know what they are talking about or what they so confidently affirm.
1TIM|1|8|We know that the law is good if one uses it properly.
1TIM|1|9|We also know that law is made not for the righteous but for lawbreakers and rebels, the ungodly and sinful, the unholy and irreligious; for those who kill their fathers or mothers, for murderers,
1TIM|1|10|for adulterers and perverts, for slave traders and liars and perjurers--and for whatever else is contrary to the sound doctrine
1TIM|1|11|that conforms to the glorious gospel of the blessed God, which he entrusted to me.
1TIM|1|12|I thank Christ Jesus our Lord, who has given me strength, that he considered me faithful, appointing me to his service.
1TIM|1|13|Even though I was once a blasphemer and a persecutor and a violent man, I was shown mercy because I acted in ignorance and unbelief.
1TIM|1|14|The grace of our Lord was poured out on me abundantly, along with the faith and love that are in Christ Jesus.
1TIM|1|15|Here is a trustworthy saying that deserves full acceptance: Christ Jesus came into the world to save sinners--of whom I am the worst.
1TIM|1|16|But for that very reason I was shown mercy so that in me, the worst of sinners, Christ Jesus might display his unlimited patience as an example for those who would believe on him and receive eternal life.
1TIM|1|17|Now to the King eternal, immortal, invisible, the only God, be honor and glory for ever and ever. Amen.
1TIM|1|18|Timothy, my son, I give you this instruction in keeping with the prophecies once made about you, so that by following them you may fight the good fight,
1TIM|1|19|holding on to faith and a good conscience. Some have rejected these and so have shipwrecked their faith.
1TIM|1|20|Among them are Hymenaeus and Alexander, whom I have handed over to Satan to be taught not to blaspheme.
1TIM|2|1|I urge, then, first of all, that requests, prayers, intercession and thanksgiving be made for everyone--
1TIM|2|2|for kings and all those in authority, that we may live peaceful and quiet lives in all godliness and holiness.
1TIM|2|3|This is good, and pleases God our Savior,
1TIM|2|4|who wants all men to be saved and to come to a knowledge of the truth.
1TIM|2|5|For there is one God and one mediator between God and men, the man Christ Jesus,
1TIM|2|6|who gave himself as a ransom for all men--the testimony given in its proper time.
1TIM|2|7|And for this purpose I was appointed a herald and an apostle--I am telling the truth, I am not lying--and a teacher of the true faith to the Gentiles.
1TIM|2|8|I want men everywhere to lift up holy hands in prayer, without anger or disputing.
1TIM|2|9|I also want women to dress modestly, with decency and propriety, not with braided hair or gold or pearls or expensive clothes,
1TIM|2|10|but with good deeds, appropriate for women who profess to worship God.
1TIM|2|11|A woman should learn in quietness and full submission.
1TIM|2|12|I do not permit a woman to teach or to have authority over a man; she must be silent.
1TIM|2|13|For Adam was formed first, then Eve.
1TIM|2|14|And Adam was not the one deceived; it was the woman who was deceived and became a sinner.
1TIM|2|15|But women will be saved through childbearing--if they continue in faith, love and holiness with propriety.
1TIM|3|1|Here is a trustworthy saying: If anyone sets his heart on being an overseer, he desires a noble task.
1TIM|3|2|Now the overseer must be above reproach, the husband of but one wife, temperate, self-controlled, respectable, hospitable, able to teach,
1TIM|3|3|not given to drunkenness, not violent but gentle, not quarrelsome, not a lover of money.
1TIM|3|4|He must manage his own family well and see that his children obey him with proper respect.
1TIM|3|5|(If anyone does not know how to manage his own family, how can he take care of God's church?)
1TIM|3|6|He must not be a recent convert, or he may become conceited and fall under the same judgment as the devil.
1TIM|3|7|He must also have a good reputation with outsiders, so that he will not fall into disgrace and into the devil's trap.
1TIM|3|8|Deacons, likewise, are to be men worthy of respect, sincere, not indulging in much wine, and not pursuing dishonest gain.
1TIM|3|9|They must keep hold of the deep truths of the faith with a clear conscience.
1TIM|3|10|They must first be tested; and then if there is nothing against them, let them serve as deacons.
1TIM|3|11|In the same way, their wives are to be women worthy of respect, not malicious talkers but temperate and trustworthy in everything.
1TIM|3|12|A deacon must be the husband of but one wife and must manage his children and his household well.
1TIM|3|13|Those who have served well gain an excellent standing and great assurance in their faith in Christ Jesus.
1TIM|3|14|Although I hope to come to you soon, I am writing you these instructions so that,
1TIM|3|15|if I am delayed, you will know how people ought to conduct themselves in God's household, which is the church of the living God, the pillar and foundation of the truth.
1TIM|3|16|Beyond all question, the mystery of godliness is great: He appeared in a body, was vindicated by the Spirit, was seen by angels, was preached among the nations, was believed on in the world, was taken up in glory.
1TIM|4|1|The Spirit clearly says that in later times some will abandon the faith and follow deceiving spirits and things taught by demons.
1TIM|4|2|Such teachings come through hypocritical liars, whose consciences have been seared as with a hot iron.
1TIM|4|3|They forbid people to marry and order them to abstain from certain foods, which God created to be received with thanksgiving by those who believe and who know the truth.
1TIM|4|4|For everything God created is good, and nothing is to be rejected if it is received with thanksgiving,
1TIM|4|5|because it is consecrated by the word of God and prayer.
1TIM|4|6|If you point these things out to the brothers, you will be a good minister of Christ Jesus, brought up in the truths of the faith and of the good teaching that you have followed.
1TIM|4|7|Have nothing to do with godless myths and old wives' tales; rather, train yourself to be godly.
1TIM|4|8|For physical training is of some value, but godliness has value for all things, holding promise for both the present life and the life to come.
1TIM|4|9|This is a trustworthy saying that deserves full acceptance
1TIM|4|10|(and for this we labor and strive), that we have put our hope in the living God, who is the Savior of all men, and especially of those who believe.
1TIM|4|11|Command and teach these things.
1TIM|4|12|Don't let anyone look down on you because you are young, but set an example for the believers in speech, in life, in love, in faith and in purity.
1TIM|4|13|Until I come, devote yourself to the public reading of Scripture, to preaching and to teaching.
1TIM|4|14|Do not neglect your gift, which was given you through a prophetic message when the body of elders laid their hands on you.
1TIM|4|15|Be diligent in these matters; give yourself wholly to them, so that everyone may see your progress.
1TIM|4|16|Watch your life and doctrine closely. Persevere in them, because if you do, you will save both yourself and your hearers.
1TIM|5|1|Do not rebuke an older man harshly, but exhort him as if he were your father. Treat younger men as brothers,
1TIM|5|2|older women as mothers, and younger women as sisters, with absolute purity.
1TIM|5|3|Give proper recognition to those widows who are really in need.
1TIM|5|4|But if a widow has children or grandchildren, these should learn first of all to put their religion into practice by caring for their own family and so repaying their parents and grandparents, for this is pleasing to God.
1TIM|5|5|The widow who is really in need and left all alone puts her hope in God and continues night and day to pray and to ask God for help.
1TIM|5|6|But the widow who lives for pleasure is dead even while she lives.
1TIM|5|7|Give the people these instructions, too, so that no one may be open to blame.
1TIM|5|8|If anyone does not provide for his relatives, and especially for his immediate family, he has denied the faith and is worse than an unbeliever.
1TIM|5|9|No widow may be put on the list of widows unless she is over sixty, has been faithful to her husband,
1TIM|5|10|and is well known for her good deeds, such as bringing up children, showing hospitality, washing the feet of the saints, helping those in trouble and devoting herself to all kinds of good deeds.
1TIM|5|11|As for younger widows, do not put them on such a list. For when their sensual desires overcome their dedication to Christ, they want to marry.
1TIM|5|12|Thus they bring judgment on themselves, because they have broken their first pledge.
1TIM|5|13|Besides, they get into the habit of being idle and going about from house to house. And not only do they become idlers, but also gossips and busybodies, saying things they ought not to.
1TIM|5|14|So I counsel younger widows to marry, to have children, to manage their homes and to give the enemy no opportunity for slander.
1TIM|5|15|Some have in fact already turned away to follow Satan.
1TIM|5|16|If any woman who is a believer has widows in her family, she should help them and not let the church be burdened with them, so that the church can help those widows who are really in need.
1TIM|5|17|The elders who direct the affairs of the church well are worthy of double honor, especially those whose work is preaching and teaching.
1TIM|5|18|For the Scripture says, "Do not muzzle the ox while it is treading out the grain," and "The worker deserves his wages."
1TIM|5|19|Do not entertain an accusation against an elder unless it is brought by two or three witnesses.
1TIM|5|20|Those who sin are to be rebuked publicly, so that the others may take warning.
1TIM|5|21|I charge you, in the sight of God and Christ Jesus and the elect angels, to keep these instructions without partiality, and to do nothing out of favoritism.
1TIM|5|22|Do not be hasty in the laying on of hands, and do not share in the sins of others. Keep yourself pure.
1TIM|5|23|Stop drinking only water, and use a little wine because of your stomach and your frequent illnesses.
1TIM|5|24|The sins of some men are obvious, reaching the place of judgment ahead of them; the sins of others trail behind them.
1TIM|5|25|In the same way, good deeds are obvious, and even those that are not cannot be hidden.
1TIM|6|1|All who are under the yoke of slavery should consider their masters worthy of full respect, so that God's name and our teaching may not be slandered.
1TIM|6|2|Those who have believing masters are not to show less respect for them because they are brothers. Instead, they are to serve them even better, because those who benefit from their service are believers, and dear to them. These are the things you are to teach and urge on them.
1TIM|6|3|If anyone teaches false doctrines and does not agree to the sound instruction of our Lord Jesus Christ and to godly teaching,
1TIM|6|4|he is conceited and understands nothing. He has an unhealthy interest in controversies and quarrels about words that result in envy, strife, malicious talk, evil suspicions
1TIM|6|5|and constant friction between men of corrupt mind, who have been robbed of the truth and who think that godliness is a means to financial gain.
1TIM|6|6|But godliness with contentment is great gain.
1TIM|6|7|For we brought nothing into the world, and we can take nothing out of it.
1TIM|6|8|But if we have food and clothing, we will be content with that.
1TIM|6|9|People who want to get rich fall into temptation and a trap and into many foolish and harmful desires that plunge men into ruin and destruction.
1TIM|6|10|For the love of money is a root of all kinds of evil. Some people, eager for money, have wandered from the faith and pierced themselves with many griefs.
1TIM|6|11|But you, man of God, flee from all this, and pursue righteousness, godliness, faith, love, endurance and gentleness.
1TIM|6|12|Fight the good fight of the faith. Take hold of the eternal life to which you were called when you made your good confession in the presence of many witnesses.
1TIM|6|13|In the sight of God, who gives life to everything, and of Christ Jesus, who while testifying before Pontius Pilate made the good confession, I charge you
1TIM|6|14|to keep this command without spot or blame until the appearing of our Lord Jesus Christ,
1TIM|6|15|which God will bring about in his own time--God, the blessed and only Ruler, the King of kings and Lord of lords,
1TIM|6|16|who alone is immortal and who lives in unapproachable light, whom no one has seen or can see. To him be honor and might forever. Amen.
1TIM|6|17|Command those who are rich in this present world not to be arrogant nor to put their hope in wealth, which is so uncertain, but to put their hope in God, who richly provides us with everything for our enjoyment.
1TIM|6|18|Command them to do good, to be rich in good deeds, and to be generous and willing to share.
1TIM|6|19|In this way they will lay up treasure for themselves as a firm foundation for the coming age, so that they may take hold of the life that is truly life.
1TIM|6|20|Timothy, guard what has been entrusted to your care. Turn away from godless chatter and the opposing ideas of what is falsely called knowledge,
1TIM|6|21|which some have professed and in so doing have wandered from the faith. Grace be with you.
