1JOHN|1|1|О том, что было от начала, что мы слышали, что видели своими очами, что рассматривали и что осязали руки наши, о Слове жизни, –
1JOHN|1|2|ибо жизнь явилась, и мы видели и свидетельствуем, и возвещаем вам сию вечную жизнь, которая была у Отца и явилась нам, –
1JOHN|1|3|о том, что мы видели и слышали, возвещаем вам, чтобы и вы имели общение с нами: а наше общение – с Отцем и Сыном Его, Иисусом Христом.
1JOHN|1|4|И сие пишем вам, чтобы радость ваша была совершенна.
1JOHN|1|5|И вот благовестие, которое мы слышали от Него и возвещаем вам: Бог есть свет, и нет в Нем никакой тьмы.
1JOHN|1|6|Если мы говорим, что имеем общение с Ним, а ходим во тьме, то мы лжем и не поступаем по истине;
1JOHN|1|7|если же ходим во свете, подобно как Он во свете, то имеем общение друг с другом, и Кровь Иисуса Христа, Сына Его, очищает нас от всякого греха.
1JOHN|1|8|Если говорим, что не имеем греха, – обманываем самих себя, и истины нет в нас.
1JOHN|1|9|Если исповедуем грехи наши, то Он, будучи верен и праведен, простит нам грехи наши и очистит нас от всякой неправды.
1JOHN|1|10|Если говорим, что мы не согрешили, то представляем Его лживым, и слова Его нет в нас.
1JOHN|2|1|Дети мои! сие пишу вам, чтобы вы не согрешали; а если бы кто согрешил, то мы имеем ходатая пред Отцем, Иисуса Христа, праведника;
1JOHN|2|2|Он есть умилостивление за грехи наши, и не только за наши, но и за [грехи] всего мира.
1JOHN|2|3|А что мы познали Его, узнаем из того, что соблюдаем Его заповеди.
1JOHN|2|4|Кто говорит: "я познал Его", но заповедей Его не соблюдает, тот лжец, и нет в нем истины;
1JOHN|2|5|а кто соблюдает слово Его, в том истинно любовь Божия совершилась: из сего узнаем, что мы в Нем.
1JOHN|2|6|Кто говорит, что пребывает в Нем, тот должен поступать так, как Он поступал.
1JOHN|2|7|Возлюбленные! пишу вам не новую заповедь, но заповедь древнюю, которую вы имели от начала. Заповедь древняя есть слово, которое вы слышали от начала.
1JOHN|2|8|Но притом и новую заповедь пишу вам, что есть истинно и в Нем и в вас: потому что тьма проходит и истинный свет уже светит.
1JOHN|2|9|Кто говорит, что он во свете, а ненавидит брата своего, тот еще во тьме.
1JOHN|2|10|Кто любит брата своего, тот пребывает во свете, и нет в нем соблазна.
1JOHN|2|11|А кто ненавидит брата своего, тот находится во тьме, и во тьме ходит, и не знает, куда идет, потому что тьма ослепила ему глаза.
1JOHN|2|12|Пишу вам, дети, потому что прощены вам грехи ради имени Его.
1JOHN|2|13|Пишу вам, отцы, потому что вы познали Сущего от начала. Пишу вам, юноши, потому что вы победили лукавого. Пишу вам, отроки, потому что вы познали Отца.
1JOHN|2|14|Я написал вам, отцы, потому что вы познали Безначального. Я написал вам, юноши, потому что вы сильны, и слово Божие пребывает в вас, и вы победили лукавого.
1JOHN|2|15|Не любите мира, ни того, что в мире: кто любит мир, в том нет любви Отчей.
1JOHN|2|16|Ибо все, что в мире: похоть плоти, похоть очей и гордость житейская, не есть от Отца, но от мира сего.
1JOHN|2|17|И мир проходит, и похоть его, а исполняющий волю Божию пребывает вовек.
1JOHN|2|18|Дети! последнее время. И как вы слышали, что придет антихрист, и теперь появилось много антихристов, то мы и познаем из того, что последнее время.
1JOHN|2|19|Они вышли от нас, но не были наши: ибо если бы они были наши, то остались бы с нами; но [они вышли, и] через то открылось, что не все наши.
1JOHN|2|20|Впрочем, вы имеете помазание от Святаго и знаете все.
1JOHN|2|21|Я написал вам не потому, чтобы вы не знали истины, но потому, что вы знаете ее, [равно как] и то, что всякая ложь не от истины.
1JOHN|2|22|Кто лжец, если не тот, кто отвергает, что Иисус есть Христос? Это антихрист, отвергающий Отца и Сына.
1JOHN|2|23|Всякий, отвергающий Сына, не имеет и Отца; а исповедующий Сына имеет и Отца.
1JOHN|2|24|Итак, что вы слышали от начала, то и да пребывает в вас; если пребудет в вас то, что вы слышали от начала, то и вы пребудете в Сыне и в Отце.
1JOHN|2|25|Обетование же, которое Он обещал нам, есть жизнь вечная.
1JOHN|2|26|Это я написал вам об обольщающих вас.
1JOHN|2|27|Впрочем, помазание, которое вы получили от Него, в вас пребывает, и вы не имеете нужды, чтобы кто учил вас; но как самое сие помазание учит вас всему, и оно истинно и неложно, то, чему оно научило вас, в том пребывайте.
1JOHN|2|28|Итак, дети, пребывайте в Нем, чтобы, когда Он явится, иметь нам дерзновение и не постыдиться пред Ним в пришествие Его.
1JOHN|2|29|Если вы знаете, что Он праведник, знайте и то, что всякий, делающий правду, рожден от Него.
1JOHN|3|1|Смотрите, какую любовь дал нам Отец, чтобы нам называться и быть детьми Божиими. Мир потому не знает нас, что не познал Его.
1JOHN|3|2|Возлюбленные! мы теперь дети Божии; но еще не открылось, что будем. Знаем только, что, когда откроется, будем подобны Ему, потому что увидим Его, как Он есть.
1JOHN|3|3|И всякий, имеющий сию надежду на Него, очищает себя так, как Он чист.
1JOHN|3|4|Всякий, делающий грех, делает и беззаконие; и грех есть беззаконие.
1JOHN|3|5|И вы знаете, что Он явился для того, чтобы взять грехи наши, и что в Нем нет греха.
1JOHN|3|6|Всякий, пребывающий в Нем, не согрешает; всякий согрешающий не видел Его и не познал Его.
1JOHN|3|7|Дети! да не обольщает вас никто. Кто делает правду, тот праведен, подобно как Он праведен.
1JOHN|3|8|Кто делает грех, тот от диавола, потому что сначала диавол согрешил. Для сего–то и явился Сын Божий, чтобы разрушить дела диавола.
1JOHN|3|9|Всякий, рожденный от Бога, не делает греха, потому что семя Его пребывает в нем; и он не может грешить, потому что рожден от Бога.
1JOHN|3|10|Дети Божии и дети диавола узнаются так: всякий, не делающий правды, не есть от Бога, равно и не любящий брата своего.
1JOHN|3|11|Ибо таково благовествование, которое вы слышали от начала, чтобы мы любили друг друга,
1JOHN|3|12|не так, как Каин, [который] был от лукавого и убил брата своего. А за что убил его? За то, что дела его были злы, а дела брата его праведны.
1JOHN|3|13|Не дивитесь, братия мои, если мир ненавидит вас.
1JOHN|3|14|Мы знаем, что мы перешли из смерти в жизнь, потому что любим братьев; не любящий брата пребывает в смерти.
1JOHN|3|15|Всякий, ненавидящий брата своего, есть человекоубийца; а вы знаете, что никакой человекоубийца не имеет жизни вечной, в нем пребывающей.
1JOHN|3|16|Любовь познали мы в том, что Он положил за нас душу Свою: и мы должны полагать души свои за братьев.
1JOHN|3|17|А кто имеет достаток в мире, но, видя брата своего в нужде, затворяет от него сердце свое, – как пребывает в том любовь Божия?
1JOHN|3|18|Дети мои! станем любить не словом или языком, но делом и истиною.
1JOHN|3|19|И вот по чему узнаем, что мы от истины, и успокаиваем пред Ним сердца наши;
1JOHN|3|20|ибо если сердце наше осуждает нас, то [кольми паче Бог], потому что Бог больше сердца нашего и знает все.
1JOHN|3|21|Возлюбленные! если сердце наше не осуждает нас, то мы имеем дерзновение к Богу,
1JOHN|3|22|и, чего ни попросим, получим от Него, потому что соблюдаем заповеди Его и делаем благоугодное пред Ним.
1JOHN|3|23|А заповедь Его та, чтобы мы веровали во имя Сына Его Иисуса Христа и любили друг друга, как Он заповедал нам.
1JOHN|3|24|И кто сохраняет заповеди Его, тот пребывает в Нем, и Он в том. А что Он пребывает в нас, узнаем по духу, который Он дал нам.
1JOHN|4|1|Возлюбленные! не всякому духу верьте, но испытывайте духов, от Бога ли они, потому что много лжепророков появилось в мире.
1JOHN|4|2|Духа Божия (и духа заблуждения) узнавайте так: всякий дух, который исповедует Иисуса Христа, пришедшего во плоти, есть от Бога;
1JOHN|4|3|а всякий дух, который не исповедует Иисуса Христа, пришедшего во плоти, не есть от Бога, но это дух антихриста, о котором вы слышали, что он придет и теперь есть уже в мире.
1JOHN|4|4|Дети! вы от Бога, и победили их; ибо Тот, Кто в вас, больше того, кто в мире.
1JOHN|4|5|Они от мира, потому и говорят по–мирски, и мир слушает их.
1JOHN|4|6|Мы от Бога; знающий Бога слушает нас; кто не от Бога, тот не слушает нас. По сему–то узнаем духа истины и духа заблуждения.
1JOHN|4|7|Возлюбленные! будем любить друг друга, потому что любовь от Бога, и всякий любящий рожден от Бога и знает Бога.
1JOHN|4|8|Кто не любит, тот не познал Бога, потому что Бог есть любовь.
1JOHN|4|9|Любовь Божия к нам открылась в том, что Бог послал в мир Единородного Сына Своего, чтобы мы получили жизнь через Него.
1JOHN|4|10|В том любовь, что не мы возлюбили Бога, но Он возлюбил нас и послал Сына Своего в умилостивление за грехи наши.
1JOHN|4|11|Возлюбленные! если так возлюбил нас Бог, то и мы должны любить друг друга.
1JOHN|4|12|Бога никто никогда не видел. Если мы любим друг друга, то Бог в нас пребывает, и любовь Его совершенна есть в нас.
1JOHN|4|13|Что мы пребываем в Нем и Он в нас, узнаем из того, что Он дал нам от Духа Своего.
1JOHN|4|14|И мы видели и свидетельствуем, что Отец послал Сына Спасителем миру.
1JOHN|4|15|Кто исповедует, что Иисус есть Сын Божий, в том пребывает Бог, и он в Боге.
1JOHN|4|16|И мы познали любовь, которую имеет к нам Бог, и уверовали в нее. Бог есть любовь, и пребывающий в любви пребывает в Боге, и Бог в нем.
1JOHN|4|17|Любовь до того совершенства достигает в нас, что мы имеем дерзновение в день суда, потому что поступаем в мире сем, как Он.
1JOHN|4|18|В любви нет страха, но совершенная любовь изгоняет страх, потому что в страхе есть мучение. Боящийся несовершен в любви.
1JOHN|4|19|Будем любить Его, потому что Он прежде возлюбил нас.
1JOHN|4|20|Кто говорит: "я люблю Бога", а брата своего ненавидит, тот лжец: ибо не любящий брата своего, которого видит, как может любить Бога, Которого не видит?
1JOHN|4|21|И мы имеем от Него такую заповедь, чтобы любящий Бога любил и брата своего.
1JOHN|5|1|Всякий верующий, что Иисус есть Христос, от Бога рожден, и всякий, любящий Родившего, любит и Рожденного от Него.
1JOHN|5|2|Что мы любим детей Божиих, узнаем из того, когда любим Бога и соблюдаем заповеди Его.
1JOHN|5|3|Ибо это есть любовь к Богу, чтобы мы соблюдали заповеди Его; и заповеди Его нетяжки.
1JOHN|5|4|Ибо всякий, рожденный от Бога, побеждает мир; и сия есть победа, победившая мир, вера наша.
1JOHN|5|5|Кто побеждает мир, как не тот, кто верует, что Иисус есть Сын Божий?
1JOHN|5|6|Сей есть Иисус Христос, пришедший водою и кровию и Духом, не водою только, но водою и кровию, и Дух свидетельствует о [Нем], потому что Дух есть истина.
1JOHN|5|7|Ибо три свидетельствуют на небе: Отец, Слово и Святый Дух; и Сии три суть едино.
1JOHN|5|8|И три свидетельствуют на земле: дух, вода и кровь; и сии три об одном.
1JOHN|5|9|Если мы принимаем свидетельство человеческое, свидетельство Божие – больше, ибо это есть свидетельство Божие, которым Бог свидетельствовал о Сыне Своем.
1JOHN|5|10|Верующий в Сына Божия имеет свидетельство в себе самом; не верующий Богу представляет Его лживым, потому что не верует в свидетельство, которым Бог свидетельствовал о Сыне Своем.
1JOHN|5|11|Свидетельство сие состоит в том, что Бог даровал нам жизнь вечную, и сия жизнь в Сыне Его.
1JOHN|5|12|Имеющий Сына (Божия) имеет жизнь; не имеющий Сына Божия не имеет жизни.
1JOHN|5|13|Сие написал я вам, верующим во имя Сына Божия, дабы вы знали, что вы, веруя в Сына Божия, имеете жизнь вечную.
1JOHN|5|14|И вот какое дерзновение мы имеем к Нему, что, когда просим чего по воле Его, Он слушает нас.
1JOHN|5|15|А когда мы знаем, что Он слушает нас во всем, чего бы мы ни просили, – знаем и то, что получаем просимое от Него.
1JOHN|5|16|Если кто видит брата своего согрешающего грехом не к смерти, то пусть молится, и [Бог] даст ему жизнь, [то есть] согрешающему [грехом] не к смерти. Есть грех к смерти: не о том говорю, чтобы он молился.
1JOHN|5|17|Всякая неправда есть грех; но есть грех не к смерти.
1JOHN|5|18|Мы знаем, что всякий, рожденный от Бога, не грешит; но рожденный от Бога хранит себя, и лукавый не прикасается к нему.
1JOHN|5|19|Мы знаем, что мы от Бога и что весь мир лежит во зле.
1JOHN|5|20|Знаем также, что Сын Божий пришел и дал нам свет и разум, да познаем Бога истинного и да будем в истинном Сыне Его Иисусе Христе. Сей есть истинный Бог и жизнь вечная.
1JOHN|5|21|Дети! храните себя от идолов. Аминь.
