RUTH|1|1|In diebus, quando iudices praeerant, facta est fames in ter ra. Abiitque homo de Bethlehem Iudae, ut peregrinaretur in regione Moabitide cum uxore sua ac duobus liberis.
RUTH|1|2|Ipse vocabatur Elimelech et uxor eius Noemi et duo filii alter Mahalon et alter Chelion Ephrathaei de Bethlehem Iudae. Ingressique regionem Moabitidem morabantur ibi.
RUTH|1|3|Et mortuus est Elimelech maritus Noemi, remansitque ipsa cum filiis,
RUTH|1|4|qui acceperunt uxores Moabitidas, quarum una vocabatur Orpha, altera Ruth; manseruntque ibi decem fere annis.
RUTH|1|5|Et ambo mortui sunt, Mahalon videlicet et Chelion; remansitque mulier orbata duobus liberis ac marito.
RUTH|1|6|Et surrexit, ut in patriam pergeret cum utraque nuru sua de regione Moabitide; audierat enim quod respexisset Dominus populum suum et dedisset eis escas.
RUTH|1|7|Egressa est itaque de loco peregrinationis suae cum utraque nuru et, iam in via posita revertendi in terram Iudae,
RUTH|1|8|dixit ad eas: " Ite in domum matris vestrae; faciat Dominus vobiscum misericordiam, sicut fecistis cum mortuis et mecum:
RUTH|1|9|det vobis invenire requiem in domibus virorum, quos sortiturae estis ". Et osculata est eas. Quae elevata voce flere coeperunt
RUTH|1|10|et dicere: " Tecum pergemus ad populum tuum ".
RUTH|1|11|Quibus illa respondit: " Revertimini, filiae meae; cur venitis mecum? Num ultra habeo filios in utero meo, ut viros ex me sperare possitis?
RUTH|1|12|Revertimini, filiae meae, abite; iam enim senectute confecta sum nec apta vinculo coniugali; etiamsi possem hac nocte concipere et parere filios,
RUTH|1|13|numquid exspectare velitis et abstinere vos a matrimonio, donec crescant et annos impleant pubertatis? Nolite, quaeso, filiae meae; quia amaritudo est mihi magis quam vobis, et egressa est manus Domini contra me.
RUTH|1|14|Elevata igitur voce, rursum flere coeperunt. Orpha osculata socrum est ac reversa; Ruth autem adhaesit socrui suae.
RUTH|1|15|Cui dixit Noemi: " En reversa est cognata tua ad populum suum et ad deos suos; vade cum ea".
RUTH|1|16|Quae respondit: "Noli instare mihi, ut relinquam te et abeam; quocumque perrexeris, pergam; ubi morata fueris, et ego pariter morabor: populus tuus populus meus et Deus tuus Deus meus.
RUTH|1|17|Quae te morientem terra susceperit, in ea moriar ibique locum accipiam sepulturae. Haec mihi faciat Dominus et haec addat, si non sola mors me et te separaverit ".
RUTH|1|18|Videns ergo Noemi quod obstinato Ruth animo decrevisset secum pergere, adversari noluit nec ultra ad suos reditum persuadere.
RUTH|1|19|Profectaeque sunt simul et venerunt in Bethlehem. Quibus urbem ingressis, tota urbs commota est super eas; dicebantque mulieres: "Haec est illa Noemi!".
RUTH|1|20|Quibus ait: "Ne vocetis me Noemi (id est Pulchram), sed vocate me Mara hoc est Amaram), quia valde me amaritudine replevit Omnipotens.
RUTH|1|21|Egressa sum plena, et vacuam reduxit me Dominus; cur igitur vocatis me Noemi, quam humiliavit Dominus, et afflixit Omnipotens? ".
RUTH|1|22|Venit ergo Noemi cum Ruth Moabitide nuru sua de terra peregrinationis suae ac reversa est in Bethlehem, quando hordea metere incipiebant.
RUTH|2|1|Erat autem Noemi consangui neus viri sui homo potens et for tis nomine Booz.
RUTH|2|2|Dixitque Ruth Moabitis ad socrum suam: " Si permittis, vadam in agrum et colligam spicas, quae fugerint manus metentium, ubicumque clementis in me patris familias repperero gratiam". Cui illa respondit: " Vade, filia mea.
RUTH|2|3|Abiit itaque et colligebat spicas post terga metentium. Accidit autem ut ager ille haberet dominum nomine Booz, qui erat de cognatione Elimelech.
RUTH|2|4|Et ecce ipse veniebat de Bethlehem dixitque messoribus: "Dominus vobiscum". Qui responderunt ei: " Benedicat tibi Dominus ".
RUTH|2|5|Dixitque Booz iuveni, qui messoribus praeerat: " Cuius est haec puella?.
RUTH|2|6|Qui respondit: " Haec est Moabitis, quae venit cum Noemi de regione Moabitide
RUTH|2|7|et rogavit, ut spicas colligeret remanentes sequens messorum vestigia; et de mane usque nunc stat in agro et nunc tantum ad momentum requievit ".
RUTH|2|8|Et ait Booz ad Ruth: " Audi, filia: ne vadas ad colligendum in alterum agrum nec recedas ab hoc loco, sed iungere puellis meis.
RUTH|2|9|Vide et, ubi messuerint, sequere eas; mandavi enim pueris, ut nemo tibi molestus sit; sed, si sitieris, vade ad sarcinulas et bibe de aqua, quam pueri hauserint ".
RUTH|2|10|Quae cadens in faciem suam et adorans super terram dixit ad eum: " Unde mihi hoc, ut invenirem gratiam ante oculos tuos, et nosse me dignareris peregrinam mulierem? ".
RUTH|2|11|Cui ille respondit: " Nuntiata sunt mihi omnia, quae feceris socrui tuae post mortem viri tui et quod dereliqueris parentes tuos et terram, in qua nata es, et veneris ad populum, quem ante nesciebas.
RUTH|2|12|Reddat tibi Dominus pro opere tuo, et plenam mercedem recipias a Domino, Deo Israel, ad quem venisti et sub cuius confugisti alas ".
RUTH|2|13|Quae ait: " Inveniam gratiam ante oculos tuos, domine mi, qui consolatus es me et locutus es ad cor ancillae tuae, quae non sum similis unius puellarum tuarum ".
RUTH|2|14|Dixitque ad eam Booz hora vescendi: "Veni huc et comede panem et intinge buccellam tuam in aceto ". Sedit itaque ad messorum latus, et porrexit ei polentam, comeditque et saturata est et tulit reliquias.
RUTH|2|15|Atque inde surrexit, ut spicas ex more colligeret. Praecepit autem Booz pueris suis dicens: "Etiam inter manipulos colligat, ne prohibeatis eam;
RUTH|2|16|quin et de fasciculis spicas proicite et remanere permittite, ut colligat, et colligentem nemo corripiat ".
RUTH|2|17|Collegit ergo in agro usque ad vesperam; et, quae collegerat virga excutiens, invenit hordei quasi ephi mensuram (id est tres modios).
RUTH|2|18|Quos portans reversa est in civitatem et ostendit socrui suae, quae collegerat; insuper protulit et dedit ei de reliquiis cibi sui, quo saturata fuerat.
RUTH|2|19|Dixitque ei socrus: " Ubi hodie collegisti et ubi fecisti opus? Sit benedictus, qui misertus est tui! ". Indicavitque ei apud quem esset operata et dixit: " Nomen viri est Booz ".
RUTH|2|20|Cui respondit Noemi: " Benedictus sit a Domino, quia non subtraxit gratiam suam nec vivis nec mortuis! ". Rursumque ait: " Propinquus noster est homo ex eis, qui pro nobis ius redemptionis habent ".
RUTH|2|21|Et Ruth: " Hoc quoque, inquit, praecepit mihi, ut tamdiu messoribus eius iungerer, donec omnes segetes meterentur ".
RUTH|2|22|Cui dixit socrus: " Melius est, filia mea, ut cum puellis eius exeas ad metendum, ne in alieno agro quispiam tibi molestus sit ".
RUTH|2|23|Iuncta est itaque puellis Booz usque ad finem messis hordei et tritici; et mansit cum socru sua.
RUTH|3|1|Et dixit ad eam Noemi socrus sua: " Filia mea, quaeram tibi requiem et providebo, ut bene sit tibi.
RUTH|3|2|Booz propinquus noster, cuius puellis in agro iuncta eras, ecce ipse hac nocte aream hordei ventilat.
RUTH|3|3|Lavare igitur, ungere et induere pallio tuo ac descende in aream; non te videat homo, donec esum potumque finierit.
RUTH|3|4|Quando autem ierit ad dormiendum, nota locum, in quo dormiat; veniesque et discooperies pallium, quo operitur a parte pedum, et ibi iacebis. Ipse autem dicet tibi quid agere debeas ".
RUTH|3|5|Quae respondit: " Quidquid praeceperis, faciam ".
RUTH|3|6|Descenditque in aream et fecit omnia, quae sibi imperaverat socrus.
RUTH|3|7|Cumque comedisset Booz et bibisset et factus esset hilarior issetque ad dormiendum in extrema parte acervi manipulorum, venit abscondite et, discooperto a pedibus eius pallio, se proiecit.
RUTH|3|8|Et ecce, nocte iam media, expavit homo et erexit se viditque mulierem iacentem ad pedes suos.
RUTH|3|9|Et ait illi: " Quae es? ". Illaque respondit: " Ego sum Ruth ancilla tua. Expande pallium tuum super famulam tuam, quia tibi est ius redemptionis ".
RUTH|3|10|Et ille: " Benedicta, inquit, es a Domino, filia; et priorem pietatem posteriore superasti, quia non es secuta iuvenes pauperes sive divites.
RUTH|3|11|Noli ergo metuere, sed, quidquid dixeris mihi, faciam tibi; scit enim omnis populus, qui habitat intra portas urbis meae, mulierem te esse fortem.
RUTH|3|12|Nec abnuo me propinquum, sed est alius me propinquior.
RUTH|3|13|Quiesce hac nocte et, facto mane, si te voluerit propinquitatis iure suscipere, bene, suscipiat; sin autem ille noluerit, vivit Dominus, ego te absque ulla dubitatione suscipiam! Dormi usque mane ".
RUTH|3|14|Dormivit itaque ad pedes eius usque ad noctis abscessum. Surrexitque, antequam homines se cognoscerent mutuo, et dixit Booz: " Cave, ne quis noverit quod huc veneris ".
RUTH|3|15|Et rursum: " Expande, inquit, palliolum tuum, quo operiris, et tene utraque manu ". Qua extendente et tenente, mensus est sex modios hordei et posuit super eam; quae portans ingressa est civitatem
RUTH|3|16|et venit ad socrum suam. Quae dixit ei: " Quid egisti, filia? ". Narravitque ei omnia, quae sibi fecisset homo,
RUTH|3|17|et ait: " Ecce sex modios hordei dedit mihi et ait: " Nolo vacuam te reverti ad socrum tuam ".
RUTH|3|18|Dixitque Noemi: " Exspecta, filia, donec videamus quem res exitum habeat; neque enim cessabit homo, nisi compleverit hodie, quod locutus est.
RUTH|4|1|Ascendit ergo Booz ad portam et sedit ibi. Cumque vidisset propinquum praeterire, de quo locutus erat, dixit ad eum: " Declina paulisper et sede hic ", vocans eum nomine suo. Qui divertit et sedit.
RUTH|4|2|Tollens autem Booz decem viros de senioribus civitatis dixit ad eos: " Sedete hic ".
RUTH|4|3|Quibus sedentibus, locutus est ad propinquum: " Partem agri fratris nostri Elimelech vendit Noemi, quae reversa est de regione Moabitide.
RUTH|4|4|Quod audire te volui et tibi dicere: Coram cunctis sedentibus et maioribus natu de populo meo, si vis possidere iure propinquitatis, eme et posside; sin autem tibi displicet, hoc ipsum indica mihi, ut sciam quid facere debeam. Nullus est enim propinquus, excepto te, qui prior es, et me, qui secundus sum ". At ille respondit: " Ego agrum emam ".
RUTH|4|5|Cui dixit Booz: " Quando emeris agrum de manu Noemi, Ruth quoque Moabitidem, quae uxor defuncti fuit, debes accipere, ut suscites nomen defuncti propinqui tui in hereditate sua ".
RUTH|4|6|Qui respondit: " Cedo iure propinquitatis; neque enim possessionem familiae meae delere debeo. Tu meo utere privilegio, quo me libenter carere profiteor ".
RUTH|4|7|Hic autem erat mos antiquitus in Israel pro redemptione et commutatione: ut esset firma concessio, solvebat homo calceamentum suum et dabat proximo suo. Hoc erat testimonium cessionis in Israel.
RUTH|4|8|Dixit ergo propinquus ad Booz: " Eme tibi ". Et solvit calceamentum suum de pede suo.
RUTH|4|9|Et Booz maioribus natu et universo populo: " Testes, inquit, vos estis hodie quod acquisierim omnia, quae fuerunt Elimelech et Chelion et Mahalon, tradente Noemi,
RUTH|4|10|et etiam Ruth Moabitidem uxorem Mahalon in coniugium sumpserim, ut suscitem nomen defuncti in hereditate sua, ne vocabulum eius de fratribus suis et de porta loci sui deleatur. Vos, inquam, huius rei hodie testes estis ".
RUTH|4|11|Respondit omnis populus, qui erat in porta, et maiores natu: " Nos testes sumus; faciat Dominus hanc mulierem, quae ingreditur domum tuam, sicut Rachel et Liam, quae aedificaverunt ambae domum Israel.Fortiter age in Ephrathaet fac tibi celebre nomen in Bethlehem!
RUTH|4|12|Fiatque domus tua sicut domus Phares, quem Thamar peperit Iudae, de semine, quod dederit Dominus tibi ex hac puella! ".
RUTH|4|13|Tulit itaque Booz Ruth et accepit uxorem; ingressusque est ad eam, et dedit illi Dominus, ut conciperet et pareret filium.
RUTH|4|14|Dixeruntque mulieres ad Noemi: " Benedictus Dominus, qui non est passus, ut deficeret tibi hodie, qui redimit familiam tuam, et vocetur nomen eius in Israel
RUTH|4|15|et consoletur animam tuam et enutriat senectutem; de nuru enim tua natus est, quae te diligit et multo tibi est melior quam septem filii ".
RUTH|4|16|Susceptumque Noemi puerum posuit in sinu suo et gerulae officio fungebatur.
RUTH|4|17|Vicinae autem mulieres congratulantes ei et dicentes: " Natus est filius Noemi! ", vocaverunt nomen eius Obed. Hic est pater Isai patris David.
RUTH|4|18|Hae sunt generationes Phares: Phares genuit Esrom,
RUTH|4|19|Esrom genuit Aram, Aram genuit Aminadab,
RUTH|4|20|Aminadab genuit Naasson, Naasson genuit Salmon,
RUTH|4|21|Salmon genuit Booz, Booz genuit Obed,
RUTH|4|22|Obed genuit Iesse, Iesse genuit David.
