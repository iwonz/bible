HOS|1|1|當 烏西雅 、 約坦 、 亞哈斯 、 希西家 作 猶大 王， 約阿施 的兒子 耶羅波安 作 以色列 王的時候，耶和華的話臨到 備利 的兒子 何西阿 。
HOS|1|2|耶和華初次向 何西阿 說話。耶和華對他說：「你去娶一個淫蕩的女子為妻，收那從淫亂所生的兒女；因為這地行大淫亂，離棄耶和華。」
HOS|1|3|於是， 何西阿 去娶了 滴拉音 的女兒 歌篾 。她就懷孕，為 何西阿 生了一個兒子。
HOS|1|4|耶和華對 何西阿 說：「給他起名叫 耶斯列 ；因為再過片時，我要懲罰 耶戶 家在 耶斯列 流人血的罪，也必終結 以色列 家的王朝。
HOS|1|5|到那日，我必在 耶斯列 平原折斷 以色列 的弓。」
HOS|1|6|歌篾 又懷孕，生了一個女兒，耶和華對 何西阿 說：「給她起名叫 羅‧路哈瑪 ；因為我必不再憐憫 以色列 家，絕不赦免他們。
HOS|1|7|我卻要憐憫 猶大 家，使他們靠耶和華－他們的上帝得救；我必不讓他們靠弓、刀、戰爭、馬匹與騎兵得救。」
HOS|1|8|歌篾 在 羅‧路哈瑪 斷奶以後，又懷孕生了一個兒子。
HOS|1|9|耶和華說：「給他起名叫 羅‧阿米 ；因為你們不是我的子民，我也不是你們的上帝 。」
HOS|1|10|然而， 以色列 的人數必多如海沙，不可量，不可數。從前在甚麼地方對他們說「你們不是我的子民」，將來就在那裏稱他們為「永生上帝的兒子」。
HOS|1|11|猶大 人和 以色列 人要一同聚集，為自己設立一個「頭」，從這地上來，因為 耶斯列 的日子必為大日。
HOS|2|1|你們要稱你們的眾弟兄 為 阿米 ，稱你們的眾姊妹 為 路哈瑪 。
HOS|2|2|要跟你們的母親理論，理論， ─因為她不是我的妻子， 我也不是她的丈夫─ 叫她除掉臉上的淫相 和胸間的淫態，
HOS|2|3|免得我剝光她，使她赤身， 如剛出生的時候一樣， 使她如曠野，如乾旱之地， 乾渴而死。
HOS|2|4|我必不憐憫她的兒女， 因為他們是從淫亂生的兒女。
HOS|2|5|他們的母親行了淫亂， 懷他們的做了可羞恥的事； 因為她說：「我要跟隨我所愛的， 我的餅、水、羊毛、麻、油、酒， 都是他們給的。」
HOS|2|6|因此，看哪，我要用荊棘堵塞她 的道， 築牆擋住她， 使她找不著路；
HOS|2|7|以致她追隨所愛的人，卻追不上， 尋找他們，卻尋不著， 就說：「我要回到前夫那裏去， 因我那時比現在還好。」
HOS|2|8|她不知道是我給她五穀、新酒和新的油， 又加添她的金銀； 他們卻用來供奉 巴力 。
HOS|2|9|因此，我要在收割的日子收回我的五穀， 在當令的季節收回我的新酒， 我要奪回她用以遮體的羊毛和麻。
HOS|2|10|如今我必在她所愛的人眼前顯露她的羞恥 ， 無人能救她脫離我的手。
HOS|2|11|我必使她的宴樂、節期、初一、安息日， 她一切的盛會都止息。
HOS|2|12|我要毀壞她的葡萄樹和無花果樹， 就是她所說「我所愛的給我為賞賜」的； 我要使它們變為荒林， 為野地的走獸所吞吃。
HOS|2|13|我要懲罰她素日給諸 巴力 燒香的罪； 那時她佩戴耳環和珠寶， 跟隨她所愛的，卻忘記我。 這是耶和華說的。
HOS|2|14|因此，看哪，我要誘導她，領她到曠野， 我要說動她的心。
HOS|2|15|在那裏，我必賜她葡萄園， 又賜她 亞割谷 作為指望的門。 她必在那裏回應， 像在年輕時從 埃及 地上來的時候一樣。
HOS|2|16|那日你必稱呼我 伊施 ，不再稱呼我 巴力 。這是耶和華說的。
HOS|2|17|因為我必從她口中除掉諸 巴力 的名號，不再有人提這名號。
HOS|2|18|當那日，我必為我的百姓，與野地的走獸、天空的飛鳥和地上爬行的動物立約；又要在國中折斷弓和刀，止息戰爭，使他們安然躺臥。
HOS|2|19|我必聘你永遠歸我為妻，以公義、公平、慈愛、憐憫聘你歸我；
HOS|2|20|又以信實聘你歸我，你就必認識耶和華。
HOS|2|21|耶和華說：那日我必應允， 我必應允天，天必應允地，
HOS|2|22|地必應允五穀、新酒和新的油； 這些都必應允在 耶斯列 身上。
HOS|2|23|我為自己必將她種在這地。 我必憐憫 羅‧路哈瑪 ； 對 羅‧阿米 說： 「你是我的子民」； 他必說：「我的上帝。」
HOS|3|1|耶和華又對我說：「你去愛那情人所愛卻犯姦淫的婦人，正如耶和華愛那偏向別神、喜愛葡萄餅 的 以色列 人。」
HOS|3|2|於是我用十五舍客勒銀子和一賀梅珥半大麥買她歸我。
HOS|3|3|我對她說：「你當多日與我同住，不可行淫，不可歸與別人，我對你也一樣。」
HOS|3|4|因為 以色列 人必多日過著無君王，無領袖，無祭祀，無柱像，無以弗得，無家中神像的生活。
HOS|3|5|後來 以色列 人必歸回 ，尋求耶和華─他們的上帝和他們的王 大衛 。在末後的日子，他們必敬畏耶和華，領受他的恩惠。
HOS|4|1|以色列 人哪，當聽耶和華的話。 耶和華指控這地的居民， 因為在這地上無誠信， 無慈愛，無人認識上帝；
HOS|4|2|惟起誓、欺騙、殺害、 偷盜、姦淫、殘暴、 流血又流血。
HOS|4|3|因此，這地悲哀， 其上的居民、野地的走獸、 天空的飛鳥都日趨衰微， 海中的魚也必消滅。
HOS|4|4|然而，人都不必爭辯，也不必指責。 你的百姓與抗拒祭司的人一樣。
HOS|4|5|日間你必跌倒， 夜間先知也要與你一同跌倒； 我要滅絕你的母親。
HOS|4|6|我的百姓因無知識而滅亡。 你拋棄知識， 我也必拋棄你， 使你不再作我的祭司。 你既忘了你上帝的律法， 我也必忘記你的兒女。
HOS|4|7|祭司越發增多，就越發得罪我； 我必使他們的榮耀變為羞辱。
HOS|4|8|他們吞吃我百姓的贖罪祭 ， 滿心願意我的子民犯罪。
HOS|4|9|將來百姓所受的， 祭司也必承受； 我必因他們所行的懲罰他們， 照他們所做的報應他們。
HOS|4|10|他們吃，卻不得飽足； 行淫，卻不繁衍； 因為他們離棄耶和華， 常行
HOS|4|11|淫亂。 酒和新酒奪去人的心。
HOS|4|12|我的百姓求問木頭， 以為木杖能指示他們； 淫亂的心使他們失迷， 以致行淫離棄他們的上帝，
HOS|4|13|在各山頂獻祭，在各高岡上燒香， 在橡樹、楊樹、大樹之下， 因為那裏樹影美好。 所以，你們的女兒行淫， 你們的媳婦 犯姦淫。
HOS|4|14|我不因你們的女兒行淫 或你們的媳婦犯姦淫懲罰她們； 因為人自己轉去與娼妓同居， 與神廟娼妓一同獻祭。 這無知的百姓必致傾倒。
HOS|4|15|以色列 啊，你雖然行淫， 猶大 卻不可犯罪； 不要往 吉甲 去， 不要上到 伯‧亞文 ， 也不要指著永生的耶和華起誓。
HOS|4|16|以色列 倔強， 猶如倔強的母牛； 現在耶和華能牧放他們， 如在寬闊之地牧放羔羊嗎？
HOS|4|17|以法蓮 親近偶像， 任憑他吧！
HOS|4|18|他們喝完了酒， 荒淫無度， 他們的官長甚愛羞恥的事。
HOS|4|19|風把他們捲在翅膀裏， 他們必因所獻的祭 蒙羞。
HOS|5|1|眾祭司啊，要聽這話！ 以色列 家啊，要留心聽！ 王室啊，要側耳而聽！ 審判將臨到你們， 因你們在 米斯巴 如羅網， 在 他泊山 如張開的網。
HOS|5|2|這些悖逆的人大行殺戮， 我要斥責他們眾人。
HOS|5|3|至於我，我認識 以法蓮 ， 以色列 不能向我隱藏。 以法蓮 哪，現在你竟然行淫 ， 以色列 竟然被污辱。
HOS|5|4|他們所做的使他們不能歸向上帝， 因有淫亂的心在他們裏面； 他們不認識耶和華。
HOS|5|5|以色列 的驕傲使自己臉面無光 ； 以色列 和 以法蓮 必因自己的罪孽跌倒， 猶大 也必與他們一同跌倒。
HOS|5|6|他們牽著牛羊去尋求耶和華， 卻尋不著； 因他已轉去離開他們。
HOS|5|7|他們不忠於耶和華， 生了私生子。 現在新月必吞滅他們和他們的地業。
HOS|5|8|你們當在 基比亞 吹角， 在 拉瑪 吹號， 在 伯‧亞文 發出警報； 便雅憫 哪，留意你的背後！
HOS|5|9|到了懲罰的日子， 以法蓮 必變為廢墟； 我在 以色列 眾支派中，已指示將來必成的事。
HOS|5|10|猶大 的領袖如同挪移地界的人， 我必把我的憤怒如水傾倒在他們身上。
HOS|5|11|以法蓮 因喜愛遵從荒謬的命令 就受欺壓，在審判中被壓碎。
HOS|5|12|我對 以法蓮 竟如蛀蟲， 向 猶大 家竟如朽爛。
HOS|5|13|以法蓮 見自己有病， 猶大 見自己有傷， 以法蓮 就前往 亞述 ， 差遣人去見大王 ； 他卻不能醫治你們， 不能治好你們的傷。
HOS|5|14|我必向 以法蓮 如獅子， 向 猶大 家如少壯獅子。 我要撕裂，並且離去， 我必奪去，無人搭救。
HOS|5|15|我要去，我要回到原處， 等他們自覺有罪，尋求我的面； 急難時他們必切切尋求我。
HOS|6|1|來，我們歸向耶和華吧！ 他撕裂我們，也必醫治； 打傷我們，也必包紮。
HOS|6|2|過兩天他必使我們甦醒， 第三天他必使我們興起， 我們就在他面前得以存活。
HOS|6|3|我們要認識，要追求認識耶和華。 他如黎明必然出現， 他必臨到我們像甘霖， 像滋潤土地的春雨。
HOS|6|4|以法蓮 哪，我可以向你怎樣行呢？ 猶大 啊，我可以向你怎樣做呢？ 因為你們的慈愛如同早晨的雲霧， 又如速散的露水。
HOS|6|5|因此，我藉先知砍伐他們， 以我口中的話殺戮他們； 對你的審判 如光發出。
HOS|6|6|我喜愛慈愛 ，不喜愛祭物； 喜愛人認識上帝，勝於燔祭。
HOS|6|7|他們卻如 亞當 背約， 在那裏向我行詭詐。
HOS|6|8|基列 是作惡之人的城， 被血沾染。
HOS|6|9|成群的祭司如強盜埋伏等候， 在 示劍 的路上殺戮， 行了邪惡。
HOS|6|10|在 以色列 家我看見可憎的事， 在 以法蓮 那裏有淫行， 以色列 被污辱了。
HOS|6|11|猶大 啊，我使被擄之民歸回的時候， 必有為你所預備的豐收。
HOS|7|1|我正要醫治 以色列 的時候， 以法蓮 的罪孽 和 撒瑪利亞 的邪惡就顯露出來。 他們行事虛謊， 內有賊人入侵， 外有群盜劫掠。
HOS|7|2|他們以為我不在意他們一切的惡行； 現在，他們所做的在我面前纏繞他們。
HOS|7|3|他們行惡使君王歡喜， 說謊使官長快樂。
HOS|7|4|他們全都犯姦淫， 如同烤熱的火爐， 師傅在揉麵到發麵時 暫時停止煽火。
HOS|7|5|在我們君王宴樂的日子， 官長因酒的烈性而生病 ， 王與褻慢的人握手。
HOS|7|6|他們臨近，心裏如火爐一般， 他們等待，如烤餅的整夜睡覺， 到了早晨卻如火焰熊熊。
HOS|7|7|他們全都熱如火爐， 吞滅他們的審判官。 他們的君王都仆倒， 他們中間無一人求告我。
HOS|7|8|以法蓮 混居在萬民中 ， 以法蓮 是沒有翻過的餅。
HOS|7|9|外邦人消耗他的力量，他卻不知道； 頭髮斑白，他也不覺得。
HOS|7|10|以色列 的驕傲使自己臉面無光。 他們雖遭遇這一切， 仍不歸向耶和華－他們的上帝， 也不尋求他。
HOS|7|11|以法蓮 好像鴿子愚蠢無知， 他們求告 埃及 ，投奔 亞述 。
HOS|7|12|他們去的時候，我要把我的網撒在他們身上； 我要捕獲他們如同空中的鳥。 我必按他們會眾所聽到的 懲罰他們。
HOS|7|13|他們因離棄我，必定有禍； 因違背我，必遭毀滅。 我雖想要救贖他們，他們卻向我說謊。
HOS|7|14|他們在床上呼號， 卻不誠心哀求我； 他們為求五穀新酒而聚集 ， 卻背叛我。
HOS|7|15|我雖管教他們，堅固他們的膀臂， 他們卻圖謀邪惡抗拒我。
HOS|7|16|他們歸向，但不是歸向至上者 ； 終究必如鬆弛的弓。 他們的領袖必因舌頭的狂傲倒在刀下， 這在 埃及 地必成為人的笑柄。
HOS|8|1|你用口吹角吧！ 敵人如鷹攻打耶和華的家； 因為他們違背了我的約， 干犯了我的律法。
HOS|8|2|他們必呼求我： 「我的上帝啊，我們 以色列 認識你了 。」
HOS|8|3|以色列 丟棄良善 ； 仇敵必追逼他。
HOS|8|4|他們立君王，並非出於我； 立官長，我卻不知道。 他們用金銀為自己製造偶像， 以致被剪除。
HOS|8|5|撒瑪利亞 啊，耶和華已拋棄你的牛犢； 我的怒氣向拜牛犢的人發作。 他們要到幾時方能無罪呢？
HOS|8|6|因這牛犢是出於 以色列 ， 是匠人所造的， 並不是上帝。 撒瑪利亞 的牛犢必被打碎。
HOS|8|7|他們所栽種的是風， 所收割的是暴風； 禾稼不長穗， 無以製成麵粉； 即便製成， 外邦人也必吞吃它。
HOS|8|8|以色列 被吞吃， 如今在列國中像人所不喜愛的器皿。
HOS|8|9|他們投奔 亞述 如獨行的野驢。 以法蓮 雇用情人，
HOS|8|10|他們雇用列國； 如今我要聚集他們， 他們必因君王和官長所加的重擔開始衰微 。
HOS|8|11|以法蓮 為贖罪增添許多祭壇， 這些祭壇卻使他犯罪。
HOS|8|12|我為他寫了許多條 律法， 他卻以為與他毫無關係。
HOS|8|13|他們獻祭物作為給我的供物， 卻自食其肉， 耶和華並不悅納他們。 現在他必記起他們的罪孽， 懲罰他們的罪惡； 他們必返回 埃及 。
HOS|8|14|以色列 忘記造他的主，建造宮殿， 猶大 增添許多堅固的城； 我卻要降火在他的城鎮， 吞滅其堡壘。
HOS|9|1|以色列 啊，不要歡喜， 像 萬民一樣快樂； 因為你行淫離棄你的上帝， 喜愛各禾場上賣淫所得的賞金。
HOS|9|2|禾場和壓酒池都不足以餵養他們， 它的新酒也必缺乏。
HOS|9|3|他們必不得住耶和華的地； 以法蓮 卻要返回 埃及 ， 在 亞述 吃不潔淨的食物。
HOS|9|4|他們必不得向耶和華獻澆酒祭， 所獻的祭也不蒙悅納。 他們的祭物如居喪者的食物， 凡吃的必使自己玷污； 因為他們的食物只為自己的口腹， 必不得入耶和華的殿。
HOS|9|5|到盛會的日子，在耶和華的節期， 你們要怎樣行呢？
HOS|9|6|看哪，他們要逃避災難； 埃及 人要收殮他們， 摩弗 人要埋葬他們。 蒺藜盤踞他們貴重的銀器， 荊棘必佔據他們的帳棚。
HOS|9|7|降罰的日子近了， 報應的時候已經來到。 以色列 必知道， 先知愚昧， 受靈感動的人狂妄， 皆因你多多作惡，大懷怨恨。
HOS|9|8|以法蓮 替我的上帝守望； 至於先知，他所到之處都有捕鳥人的羅網， 在他上帝的家中也遭人懷恨。
HOS|9|9|他們深深敗壞， 如在 基比亞 的日子一樣。 耶和華必記起他們的罪孽， 懲罰他們的罪惡。
HOS|9|10|我發現 以色列 ， 如在曠野的葡萄； 我看見你們的祖先， 如春季無花果樹上初熟的果子。 他們卻來到 巴力‧毗珥 ， 獻上自己做羞恥的事， 成為可憎惡的， 與他們所愛的一樣。
HOS|9|11|以法蓮 ，他們的榮耀如鳥飛去， 必不生產，不懷胎，不成孕；
HOS|9|12|他們縱然將兒女養大， 我卻要使他們喪子，一個也不留。 我離棄他們， 他們就有禍了。
HOS|9|13|我看 以法蓮 如 推羅 栽於美地。 以法蓮 卻要將自己的兒女帶出來， 交給行殺戮的人。
HOS|9|14|耶和華啊，求你加給他們， 加給他們甚麼呢？ 要使他們懷孕流產， 乳房枯乾。
HOS|9|15|因他們在 吉甲 的一切惡事， 我在那裏憎惡他們。 因他們所行的惡， 我必把他們趕出我的殿， 不再愛他們； 他們的領袖都是悖逆的。
HOS|9|16|以法蓮 受擊打， 其根枯乾，不能結果， 即或生產， 我也要殺他們所生的愛子。
HOS|9|17|我的上帝必棄絕他們， 因為他們不聽從他； 他們必飄流在列國中。
HOS|10|1|以色列 是茂盛的葡萄樹， 結果繁多。 果子越多， 就越增添祭壇； 土地越肥美， 就越建造美麗的柱像。
HOS|10|2|他們心懷二意， 現今要定為有罪。 耶和華必拆毀他們的祭壇， 粉碎他們的柱像。
HOS|10|3|現在他們要說： 「我們沒有王； 因為我們不敬畏耶和華， 王又能為我們做甚麼呢？」
HOS|10|4|他們講空話， 以假誓立約； 因此，懲罰如苦菜滋生 在田間的犁溝中。
HOS|10|5|撒瑪利亞 的居民必因 伯‧亞文 的牛犢驚恐； 它的百姓為它悲哀， 它的祭司為它戰兢， 因為榮耀已經離開它。
HOS|10|6|人必將牛犢帶到 亞述 ， 當作禮物獻給大王。 以法蓮 必蒙羞， 以色列 必因自己的計謀慚愧。
HOS|10|7|撒瑪利亞 的王要滅亡， 如水面上的泡沫一般。
HOS|10|8|亞文 的丘壇， 以色列 犯罪的地方必毀壞， 荊棘和蒺藜必長在他們的祭壇上。 他們要向大山說：遮蓋我們！ 向小山說：倒在我們身上！
HOS|10|9|以色列 啊， 你從 基比亞 的日子以來就時常犯罪， 他們仍停留在那裏。 攻擊罪孽之輩的戰事豈不會臨到 基比亞 嗎？
HOS|10|10|我必隨己意懲罰他們， 他們為雙重的罪所纏； 萬民必聚集攻擊他們。
HOS|10|11|以法蓮 是馴良的母牛犢，喜愛踹穀， 我要將軛套在牠肥美的頸項上， 我要使 以法蓮 被套住； 猶大 必耕田， 雅各 必耙地。
HOS|10|12|你們要為自己栽種公義， 收割慈愛。 你們要開墾荒地， 現今正是尋求耶和華的時候； 等他臨到，公義必如雨降給你們。
HOS|10|13|你們耕種奸惡， 收割罪孽， 吃的是謊言的果實。 因你倚靠自己的行為， 仰賴你眾多的勇士，
HOS|10|14|所以在你百姓中必掀起鬧鬨， 你一切的堡壘必被拆毀， 就如 沙勒幔 在爭戰的日子拆毀 伯‧亞比勒 ， 將城中的母子一同摔死。
HOS|10|15|伯特利 啊，因你們的大惡， 你們必遭遇如此。 黎明來臨， 以色列 的王必全然滅絕。
HOS|11|1|以色列 年幼的時候，我愛他， 就從 埃及 召我的兒子出來。
HOS|11|2|先知 越是呼喚他們， 他們越是遠離 ， 向諸 巴力 獻祭， 為雕刻的偶像燒香。
HOS|11|3|我曾教導 以法蓮 行走， 我用膀臂 抱起他們， 他們卻不知道是我醫治他們。
HOS|11|4|我用慈繩愛索牽引他們； 我待他們如人鬆開牛兩腮旁邊的軛， 彎下身來餵養他們。
HOS|11|5|他們必不返回 埃及 地； 然而 亞述 人要作他們的王， 因他們不肯歸向我。
HOS|11|6|刀劍必臨到他們的城鎮， 毀壞門閂，吞滅眾人， 都因他們自己的計謀。
HOS|11|7|我的百姓偏要背離我， 他們雖向至高者呼求， 他卻不抬舉他們 。
HOS|11|8|以法蓮 哪，我怎能捨棄你？ 以色列 啊，我怎能棄絕你？ 我怎能使你如 押瑪 ？ 怎能使你如 洗扁 ？ 我回心轉意， 我的憐憫燃了起來。
HOS|11|9|我必不發猛烈的怒氣， 也不再毀滅 以法蓮 。 因我是上帝，並非世人， 是你們中間的聖者； 我必不在怒中臨到你們。
HOS|11|10|耶和華如獅子吼叫， 他的兒女必跟隨他。 他一吼叫， 他們就從西方戰兢而來。
HOS|11|11|他們必如雀鳥從 埃及 戰兢而來， 又如鴿子從 亞述 地來到。 我必使他們住自己的房屋； 這是耶和華說的。
HOS|11|12|以法蓮 用謊言圍繞我， 以色列 家用詭計環繞我； 猶大 卻仍與上帝同行 ， 向聖者忠心。
HOS|12|1|以法蓮 以風為食物， 終日追逐東風， 增添虛謊和殘暴， 與 亞述 立約， 也把油送到 埃及 。
HOS|12|2|耶和華指控 猶大 ， 要照 雅各 所行的懲罰他， 按他所做的報應他。
HOS|12|3|他在腹中抓住哥哥的腳跟， 壯年的時候與上帝角力，
HOS|12|4|他與天使角力，並且得勝。 他曾哀哭，懇求施恩。 在 伯特利 遇見耶和華， 耶和華在那裏吩咐我們 ，
HOS|12|5|耶和華是萬軍之上帝， 耶和華是他可記念的名。
HOS|12|6|所以你當歸向你的上帝， 謹守慈愛和公平， 常常等候你的上帝。
HOS|12|7|商人 手持詭詐的天平， 喜愛欺壓。
HOS|12|8|以法蓮 說： 我果然富有，得了財寶； 我所勞碌得來的一切 人必找不到我有甚麼可算為有罪的惡。
HOS|12|9|自從你出 埃及 地以來， 我就是耶和華－你的上帝； 我必使你再住帳棚， 如同節期的日子一樣。
HOS|12|10|我已吩咐眾先知， 又增加異象， 藉先知設比喻。
HOS|12|11|基列 沒有罪孽嗎？ 他們誠然是虛假的， 在 吉甲 獻牛犢為祭； 他們的祭壇如同田間犁溝中的亂堆。
HOS|12|12|從前 雅各 逃到 亞蘭 地， 以色列 為娶妻子工作， 為娶妻子而牧放。
HOS|12|13|後來耶和華藉先知領 以色列 從 埃及 上來， 也藉先知看顧他們。
HOS|12|14|然而 以法蓮 大大惹動主怒， 他所流的血必歸到他身上。 主必使他的羞辱歸還給他。
HOS|13|1|從前 以法蓮 說話，人都戰兢， 他在 以色列 中居處高位； 但他因 巴力 犯罪就死了。
HOS|13|2|如今他們罪上加罪， 為自己鑄造偶像， 憑自己的聰明用銀子造偶像， 全都是匠人所製的。 論到它，有話說： 獻祭的人都要親吻牛犢。
HOS|13|3|因此，他們必如早晨的雲霧， 又如速散的露水， 如被狂風吹離禾場的糠秕， 又如煙囪冒出的煙。
HOS|13|4|自從你出 埃及 地以來， 我就是耶和華－你的上帝； 除了我上帝以外，你不認識別的， 在我以外，並沒有救主。
HOS|13|5|我曾在曠野， 就是那乾旱之地認識你。
HOS|13|6|他們得到餵養，就飽足； 既得飽足，就心高氣傲， 因而忘記了我。
HOS|13|7|因此我向他們如同獅子， 又如豹伏在道旁。
HOS|13|8|我如失去小熊的母熊，攻擊他們， 撕裂他們的胸膛。 在那裏我必如母獅吞吃他們， 如野獸撕開他們。
HOS|13|9|以色列 啊，你自取滅亡了 ， 因為我才是你的幫助。
HOS|13|10|現在，你的王在哪裏呢？ 讓他在你的各城中拯救你吧！ 你曾說「給我立君王和官長」， 那些治理你的又在哪裏呢？
HOS|13|11|我在怒氣中將王賜給你， 又在烈怒中將王廢去。
HOS|13|12|以法蓮 的罪孽被捲起來， 他的罪惡被收藏起來。
HOS|13|13|產婦的疼痛必臨到他身上； 他是無智慧之子， 如同臨盆時未出現的胎兒。
HOS|13|14|我必救贖他們脫離陰間， 救贖他們脫離死亡。 死亡啊，你的災害在哪裏？ 陰間哪，你的毀滅在哪裏？ 憐憫必從我眼前消逝。
HOS|13|15|他在弟兄中雖然旺盛， 卻有東風颳來， 就是耶和華的風從曠野上來。 他的泉源必乾涸， 他的源頭必枯竭， 這風必奪走他所積蓄的一切寶物。
HOS|13|16|撒瑪利亞 要擔當罪孽， 因為背叛自己的上帝。 他們必倒在刀下， 嬰孩必被摔死， 孕婦必被剖開。
HOS|14|1|以色列 啊，你要歸向耶和華－你的上帝， 你因自己的罪孽跌倒了。
HOS|14|2|當歸向耶和華， 用言語向他說： 「求你除盡罪孽，悅納善行， 我們就用嘴唇的祭代替牛犢獻上。
HOS|14|3|亞述 不能救我們， 我們不再騎馬， 也不再對我們手所造的偶像說： 『你是我們的上帝』； 孤兒在你那裏得蒙憐憫。」
HOS|14|4|我必醫治他們背道的病， 甘心愛他們， 因為我向他們所發的怒氣已轉消。
HOS|14|5|我必向 以色列 如甘露； 他必如百合花開放， 如 黎巴嫩 的樹扎根。
HOS|14|6|他的嫩枝必延伸， 他的榮華如橄欖樹， 香氣如 黎巴嫩 的香柏樹。
HOS|14|7|曾住在他蔭下的必歸回，使五穀生長 ， 他們要發旺如葡萄樹， 他的名氣 如 黎巴嫩 的酒。
HOS|14|8|以法蓮 說： 「我與偶像有何相干？」 我應允他，顧念他： 我如青翠的松樹， 你的果實從我而來。
HOS|14|9|智慧人必明白這些事， 聰明人必知道這一切。 耶和華的道是正直的， 義人行在其中， 罪人卻在其上跌倒。
