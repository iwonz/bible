1KGS|1|1|Now King David was old and advanced in years. And although they covered him with clothes, he could not get warm.
1KGS|1|2|Therefore his servants said to him, "Let a young woman be sought for my lord the king, and let her wait on the king and be in his service. Let her lie in your arms, that my lord the king may be warm."
1KGS|1|3|So they sought for a beautiful young woman throughout all the territory of Israel, and found Abishag the Shunammite, and brought her to the king.
1KGS|1|4|The young woman was very beautiful, and she was of service to the king and attended to him, but the king knew her not.
1KGS|1|5|Now Adonijah the son of Haggith exalted himself, saying, "I will be king." And he prepared for himself chariots and horsemen, and fifty men to run before him.
1KGS|1|6|His father had never at any time displeased him by asking, "Why have you done thus and so?" He was also a very handsome man, and he was born next after Absalom.
1KGS|1|7|He conferred with Joab the son of Zeruiah and with Abiathar the priest. And they followed Adonijah and helped him.
1KGS|1|8|But Zadok the priest and Benaiah the son of Jehoiada and Nathan the prophet and Shimei and Rei and David's mighty men were not with Adonijah.
1KGS|1|9|Adonijah sacrificed sheep, oxen, and fattened cattle by the Serpent's Stone, which is beside En-rogel, and he invited all his brothers, the king's sons, and all the royal officials of Judah,
1KGS|1|10|but he did not invite Nathan the prophet or Benaiah or the mighty men or Solomon his brother.
1KGS|1|11|Then Nathan said to Bathsheba the mother of Solomon, "Have you not heard that Adonijah the son of Haggith has become king and David our lord does not know it?
1KGS|1|12|Now therefore come, let me give you advice, that you may save your own life and the life of your son Solomon.
1KGS|1|13|Go in at once to King David, and say to him, 'Did you not, my lord the king, swear to your servant, saying, "Solomon your son shall reign after me, and he shall sit on my throne"? Why then is Adonijah king?'
1KGS|1|14|Then while you are still speaking with the king, I also will come in after you and confirm your words."
1KGS|1|15|So Bathsheba went to the king in his chamber (now the king was very old, and Abishag the Shunammite was attending to the king).
1KGS|1|16|Bathsheba bowed and paid homage to the king, and the king said, "What do you desire?"
1KGS|1|17|She said to him, "My lord, you swore to your servant by the LORD your God, saying, 'Solomon your son shall reign after me, and he shall sit on my throne.'
1KGS|1|18|And now, behold, Adonijah is king, although you, my lord the king, do not know it.
1KGS|1|19|He has sacrificed oxen, fattened cattle, and sheep in abundance, and has invited all the sons of the king, Abiathar the priest, and Joab the commander of the army, but Solomon your servant he has not invited.
1KGS|1|20|And now, my lord the king, the eyes of all Israel are on you, to tell them who shall sit on the throne of my lord the king after him.
1KGS|1|21|Otherwise it will come to pass, when my lord the king sleeps with his fathers, that I and my son Solomon will be counted offenders."
1KGS|1|22|While she was still speaking with the king, Nathan the prophet came in.
1KGS|1|23|And they told the king, "Here is Nathan the prophet." And when he came in before the king, he bowed before the king, with his face to the ground.
1KGS|1|24|And Nathan said, "My lord the king, have you said, 'Adonijah shall reign after me, and he shall sit on my throne'?
1KGS|1|25|For he has gone down this day and has sacrificed oxen, fattened cattle, and sheep in abundance, and has invited all the king's sons, the commanders of the army, and Abiathar the priest. And behold, they are eating and drinking before him, and saying, 'Long live King Adonijah!'
1KGS|1|26|But me, your servant, and Zadok the priest, and Benaiah the son of Jehoiada, and your servant Solomon he has not invited.
1KGS|1|27|Has this thing been brought about by my lord the king and you have not told your servants who should sit on the throne of my lord the king after him?"
1KGS|1|28|Then King David answered, "Call Bathsheba to me." So she came into the king's presence and stood before the king.
1KGS|1|29|And the king swore, saying, "As the LORD lives, who has redeemed my soul out of every adversity,
1KGS|1|30|as I swore to you by the LORD, the God of Israel, saying, 'Solomon your son shall reign after me, and he shall sit on my throne in my place,' even so will I do this day."
1KGS|1|31|Then Bathsheba bowed with her face to the ground and paid homage to the king and said, "May my lord King David live forever!"
1KGS|1|32|King David said, "Call to me Zadok the priest, Nathan the prophet, and Benaiah the son of Jehoiada." So they came before the king.
1KGS|1|33|And the king said to them, "Take with you the servants of your lord and have Solomon my son ride on my own mule, and bring him down to Gihon.
1KGS|1|34|And let Zadok the priest and Nathan the prophet there anoint him king over Israel. Then blow the trumpet and say, 'Long live King Solomon!'
1KGS|1|35|You shall then come up after him, and he shall come and sit on my throne, for he shall be king in my place. And I have appointed him to be ruler over Israel and over Judah."
1KGS|1|36|And Benaiah the son of Jehoiada answered the king, "Amen! May the LORD, the God of my lord the king, say so.
1KGS|1|37|As the LORD has been with my lord the king, even so may he be with Solomon, and make his throne greater than the throne of my lord King David."
1KGS|1|38|So Zadok the priest, Nathan the prophet, and Benaiah the son of Jehoiada, and the Cherethites and the Pelethites went down and had Solomon ride on King David's mule and brought him to Gihon.
1KGS|1|39|There Zadok the priest took the horn of oil from the tent and anointed Solomon. Then they blew the trumpet, and all the people said, "Long live King Solomon!"
1KGS|1|40|And all the people went up after him, playing on pipes, and rejoicing with great joy, so that the earth was split by their noise.
1KGS|1|41|Adonijah and all the guests who were with him heard it as they finished feasting. And when Joab heard the sound of the trumpet, he said, "What does this uproar in the city mean?"
1KGS|1|42|While he was still speaking, behold, Jonathan the son of Abiathar the priest came. And Adonijah said, "Come in, for you are a worthy man and bring good news."
1KGS|1|43|Jonathan answered Adonijah, "No, for our lord King David has made Solomon king,
1KGS|1|44|and the king has sent with him Zadok the priest, Nathan the prophet, and Benaiah the son of Jehoiada, and the Cherethites and the Pelethites. And they had him ride on the king's mule.
1KGS|1|45|And Zadok the priest and Nathan the prophet have anointed him king at Gihon, and they have gone up from there rejoicing, so that the city is in an uproar. This is the noise that you have heard.
1KGS|1|46|Solomon sits on the royal throne.
1KGS|1|47|Moreover, the king's servants came to congratulate our lord King David, saying, 'May your God make the name of Solomon more famous than yours, and make his throne greater than your throne.' And the king bowed himself on the bed.
1KGS|1|48|And the king also said, 'Blessed be the LORD, the God of Israel, who has granted someone to sit on my throne this day, my own eyes seeing it.'"
1KGS|1|49|Then all the guests of Adonijah trembled and rose, and each went his own way.
1KGS|1|50|And Adonijah feared Solomon. So he arose and went and took hold of the horns of the altar.
1KGS|1|51|Then it was told Solomon, "Behold, Adonijah fears King Solomon, for behold, he has laid hold of the horns of the altar, saying, 'Let King Solomon swear to me first that he will not put his servant to death with the sword.'"
1KGS|1|52|And Solomon said, "If he will show himself a worthy man, not one of his hairs shall fall to the earth, but if wickedness is found in him, he shall die."
1KGS|1|53|So King Solomon sent, and they brought him down from the altar. And he came and paid homage to King Solomon, and Solomon said to him, "Go to your house."
1KGS|2|1|When David's time to die drew near, he commanded Solomon his son, saying,
1KGS|2|2|"I am about to go the way of all the earth. Be strong, and show yourself a man,
1KGS|2|3|and keep the charge of the LORD your God, walking in his ways and keeping his statutes, his commandments, his rules, and his testimonies, as it is written in the Law of Moses, that you may prosper in all that you do and wherever you turn,
1KGS|2|4|that the LORD may establish his word that he spoke concerning me, saying, 'If your sons pay close attention to their way, to walk before me in faithfulness with all their heart and with all their soul, you shall not lack a man on the throne of Israel.'
1KGS|2|5|"Moreover, you also know what Joab the son of Zeruiah did to me, how he dealt with the two commanders of the armies of Israel, Abner the son of Ner, and Amasa the son of Jether, whom he killed, avenging in time of peace for blood that had been shed in war, and putting the blood of war on the belt around his waist and on the sandals on his feet.
1KGS|2|6|Act therefore according to your wisdom, but do not let his gray head go down to Sheol in peace.
1KGS|2|7|But deal loyally with the sons of Barzillai the Gileadite, and let them be among those who eat at your table, for with such loyalty they met me when I fled from Absalom your brother.
1KGS|2|8|And there is also with you Shimei the son of Gera, the Benjaminite from Bahurim, who cursed me with a grievous curse on the day when I went to Mahanaim. But when he came down to meet me at the Jordan, I swore to him by the LORD, saying, 'I will not put you to death with the sword.'
1KGS|2|9|Now therefore do not hold him guiltless, for you are a wise man. You will know what you ought to do to him, and you shall bring his gray head down with blood to Sheol."
1KGS|2|10|Then David slept with his fathers and was buried in the city of David.
1KGS|2|11|And the time that David reigned over Israel was forty years. He reigned seven years in Hebron and thirty-three years in Jerusalem.
1KGS|2|12|So Solomon sat on the throne of David his father, and his kingdom was firmly established.
1KGS|2|13|Then Adonijah the son of Haggith came to Bathsheba the mother of Solomon. And she said, "Do you come peacefully?" He said, "Peacefully."
1KGS|2|14|Then he said, "I have something to say to you." She said, "Speak."
1KGS|2|15|He said, "You know that the kingdom was mine, and that all Israel fully expected me to reign. However, the kingdom has turned about and become my brother's, for it was his from the LORD.
1KGS|2|16|And now I have one request to make of you; do not refuse me." She said to him, "Speak."
1KGS|2|17|And he said, "Please ask King Solomon- he will not refuse you- to give me Abishag the Shunammite as my wife."
1KGS|2|18|Bathsheba said, "Very well; I will speak for you to the king."
1KGS|2|19|So Bathsheba went to King Solomon to speak to him on behalf of Adonijah. And the king rose to meet her and bowed down to her. Then he sat on his throne and had a seat brought for the king's mother, and she sat on his right.
1KGS|2|20|Then she said, "I have one small request to make of you; do not refuse me." And the king said to her, "Make your request, my mother, for I will not refuse you."
1KGS|2|21|She said, "Let Abishag the Shunammite be given to Adonijah your brother as his wife."
1KGS|2|22|King Solomon answered his mother, "And why do you ask Abishag the Shunammite for Adonijah? Ask for him the kingdom also, for he is my older brother, and on his side are Abiathar the priest and Joab the son of Zeruiah."
1KGS|2|23|Then King Solomon swore by the LORD, saying, "God do so to me and more also if this word does not cost Adonijah his life!
1KGS|2|24|Now therefore as the LORD lives, who has established me and placed me on the throne of David my father, and who has made me a house, as he promised, Adonijah shall be put to death this day."
1KGS|2|25|So King Solomon sent Benaiah the son of Jehoiada, and he struck him down, and he died.
1KGS|2|26|And to Abiathar the priest the king said, "Go to Anathoth, to your estate, for you deserve death. But I will not at this time put you to death, because you carried the ark of the Lord GOD before David my father, and because you shared in all my father's affliction."
1KGS|2|27|So Solomon expelled Abiathar from being priest to the LORD, thus fulfilling the word of the LORD that he had spoken concerning the house of Eli in Shiloh.
1KGS|2|28|When the news came to Joab- for Joab had supported Adonijah although he had not supported Absalom- Joab fled to the tent of the LORD and caught hold of the horns of the altar.
1KGS|2|29|And when it was told King Solomon, "Joab has fled to the tent of the LORD, and behold, he is beside the altar," Solomon sent Benaiah the son of Jehoiada, saying, "Go, strike him down."
1KGS|2|30|So Benaiah came to the tent of the LORD and said to him, "The king commands, 'Come out.'"But he said, "No, I will die here." Then Benaiah brought the king word again, saying, "Thus said Joab, and thus he answered me."
1KGS|2|31|The king replied to him, "Do as he has said, strike him down and bury him, and thus take away from me and from my father's house the guilt for the blood that Joab shed without cause.
1KGS|2|32|The LORD will bring back his bloody deeds on his own head, because, without the knowledge of my father David, he attacked and killed with the sword two men more righteous and better than himself, Abner the son of Ner, commander of the army of Israel, and Amasa the son of Jether, commander of the army of Judah.
1KGS|2|33|So shall their blood come back on the head of Joab and on the head of his descendants forever. But for David and for his descendants and for his house and for his throne there shall be peace from the LORD forevermore."
1KGS|2|34|Then Benaiah the son of Jehoiada went up and struck him down and put him to death. And he was buried in his own house in the wilderness.
1KGS|2|35|The king put Benaiah the son of Jehoiada over the army in place of Joab, and the king put Zadok the priest in the place of Abiathar.
1KGS|2|36|Then the king sent and summoned Shimei and said to him, "Build yourself a house in Jerusalem and dwell there, and do not go out from there to any place whatever.
1KGS|2|37|For on the day you go out and cross the brook Kidron, know for certain that you shall die. Your blood shall be on your own head."
1KGS|2|38|And Shimei said to the king, "What you say is good; as my lord the king has said, so will your servant do." So Shimei lived in Jerusalem many days.
1KGS|2|39|But it happened at the end of three years that two of Shimei's servants ran away to Achish, son of Maacah, king of Gath. And when it was told Shimei, "Behold, your servants are in Gath,"
1KGS|2|40|Shimei arose and saddled a donkey and went to Gath to Achish to seek his servants. Shimei went and brought his servants from Gath.
1KGS|2|41|And when Solomon was told that Shimei had gone from Jerusalem to Gath and returned,
1KGS|2|42|the king sent and summoned Shimei and said to him, "Did I not make you swear by the LORD and solemnly warn you, saying, 'Know for certain that on the day you go out and go to any place whatever, you shall die'? And you said to me, 'What you say is good; I will obey.'
1KGS|2|43|Why then have you not kept your oath to the LORD and the commandment with which I commanded you?"
1KGS|2|44|The king also said to Shimei, "You know in your own heart all the harm that you did to David my father. So the LORD will bring back your harm on your own head.
1KGS|2|45|But King Solomon shall be blessed, and the throne of David shall be established before the LORD forever."
1KGS|2|46|Then the king commanded Benaiah the son of Jehoiada, and he went out and struck him down, and he died. So the kingdom was established in the hand of Solomon.
1KGS|3|1|Solomon made a marriage alliance with Pharaoh king of Egypt. He took Pharaoh's daughter and brought her into the city of David until he had finished building his own house and the house of the LORD and the wall around Jerusalem.
1KGS|3|2|The people were sacrificing at the high places, however, because no house had yet been built for the name of the LORD.
1KGS|3|3|Solomon loved the LORD, walking in the statutes of David his father, only he sacrificed and made offerings at the high places.
1KGS|3|4|And the king went to Gibeon to sacrifice there, for that was the great high place. Solomon used to offer a thousand burnt offerings on that altar.
1KGS|3|5|At Gibeon the LORD appeared to Solomon in a dream by night, and God said, "Ask what I shall give you."
1KGS|3|6|And Solomon said, "You have shown great and steadfast love to your servant David my father, because he walked before you in faithfulness, in righteousness, and in uprightness of heart toward you. And you have kept for him this great and steadfast love and have given him a son to sit on his throne this day.
1KGS|3|7|And now, O LORD my God, you have made your servant king in place of David my father, although I am but a little child. I do not know how to go out or come in.
1KGS|3|8|And your servant is in the midst of your people whom you have chosen, a great people, too many to be numbered or counted for multitude.
1KGS|3|9|Give your servant therefore an understanding mind to govern your people, that I may discern between good and evil, for who is able to govern this your great people?"
1KGS|3|10|It pleased the Lord that Solomon had asked this.
1KGS|3|11|And God said to him, "Because you have asked this, and have not asked for yourself long life or riches or the life of your enemies, but have asked for yourself understanding to discern what is right,
1KGS|3|12|behold, I now do according to your word. Behold, I give you a wise and discerning mind, so that none like you has been before you and none like you shall arise after you.
1KGS|3|13|I give you also what you have not asked, both riches and honor, so that no other king shall compare with you, all your days.
1KGS|3|14|And if you will walk in my ways, keeping my statutes and my commandments, as your father David walked, then I will lengthen your days."
1KGS|3|15|And Solomon awoke, and behold, it was a dream. Then he came to Jerusalem and stood before the ark of the covenant of the LORD, and offered up burnt offerings and peace offerings, and made a feast for all his servants.
1KGS|3|16|Then two prostitutes came to the king and stood before him.
1KGS|3|17|The one woman said, "Oh, my lord, this woman and I live in the same house, and I gave birth to a child while she was in the house.
1KGS|3|18|Then on the third day after I gave birth, this woman also gave birth. And we were alone. There was no one else with us in the house; only we two were in the house.
1KGS|3|19|And this woman's son died in the night, because she lay on him.
1KGS|3|20|And she arose at midnight and took my son from beside me, while your servant slept, and laid him at her breast, and laid her dead son at my breast.
1KGS|3|21|When I rose in the morning to nurse my child, behold, he was dead. But when I looked at him closely in the morning, behold, he was not the child that I had borne."
1KGS|3|22|But the other woman said, "No, the living child is mine, and the dead child is yours." The first said, "No, the dead child is yours, and the living child is mine." Thus they spoke before the king.
1KGS|3|23|Then the king said, "The one says, 'This is my son that is alive, and your son is dead'; and the other says, 'No; but your son is dead, and my son is the living one.'"
1KGS|3|24|And the king said, "Bring me a sword." So a sword was brought before the king.
1KGS|3|25|And the king said, "Divide the living child in two, and give half to the one and half to the other."
1KGS|3|26|Then the woman whose son was alive said to the king, because her heart yearned for her son, "Oh, my lord, give her the living child, and by no means put him to death." But the other said, "He shall be neither mine nor yours; divide him."
1KGS|3|27|Then the king answered and said, "Give the living child to the first woman, and by no means put him to death; she is his mother."
1KGS|3|28|And all Israel heard of the judgment that the king had rendered, and they stood in awe of the king, because they perceived that the wisdom of God was in him to do justice.
1KGS|4|1|King Solomon was king over all Israel,
1KGS|4|2|and these were his high officials: Azariah the son of Zadok was the priest;
1KGS|4|3|Elihoreph and Ahijah the sons of Shisha were secretaries; Jehoshaphat the son of Ahilud was recorder;
1KGS|4|4|Benaiah the son of Jehoiada was in command of the army; Zadok and Abiathar were priests;
1KGS|4|5|Azariah the son of Nathan was over the officers; Zabud the son of Nathan was priest and king's friend;
1KGS|4|6|Ahishar was in charge of the palace; and Adoniram the son of Abda was in charge of the forced labor.
1KGS|4|7|Solomon had twelve officers over all Israel, who provided food for the king and his household. Each man had to make provision for one month in the year.
1KGS|4|8|These were their names: Ben-hur, in the hill country of Ephraim;
1KGS|4|9|Ben-deker, in Makaz, Shaalbim, Beth-shemesh, and Elonbeth-hanan;
1KGS|4|10|Ben-hesed, in Arubboth (to him belonged Socoh and all the land of Hepher);
1KGS|4|11|Ben-abinadab, in all Naphath-dor (he had Taphath the daughter of Solomon as his wife);
1KGS|4|12|Baana the son of Ahilud, in Taanach, Megiddo, and all Beth-shean that is beside Zarethan below Jezreel, and from Beth-shean to Abel-meholah, as far as the other side of Jokmeam;
1KGS|4|13|Ben-geber, in Ramoth-gilead (he had the villages of Jair the son of Manasseh, which are in Gilead, and he had the region of Argob, which is in Bashan, sixty great cities with walls and bronze bars);
1KGS|4|14|Ahinadab the son of Iddo, in Mahanaim;
1KGS|4|15|Ahimaaz, in Naphtali (he had taken Basemath the daughter of Solomon as his wife);
1KGS|4|16|Baana the son of Hushai, in Asher and Bealoth;
1KGS|4|17|Jehoshaphat the son of Paruah, in Issachar;
1KGS|4|18|Shimei the son of Ela, in Benjamin;
1KGS|4|19|Geber the son of Uri, in the land of Gilead, the country of Sihon king of the Amorites and of Og king of Bashan. And there was one governor who was over the land.
1KGS|4|20|Judah and Israel were as many as the sand by the sea. They ate and drank and were happy.
1KGS|4|21|Solomon ruled over all the kingdoms from the Euphrates to the land of the Philistines and to the border of Egypt. They brought tribute and served Solomon all the days of his life.
1KGS|4|22|Solomon's provision for one day was thirty cors of fine flour and sixty cors of meal,
1KGS|4|23|ten fat oxen, and twenty pasture-fed cattle, a hundred sheep, besides deer, gazelles, roebucks, and fattened fowl.
1KGS|4|24|For he had dominion over all the region west of the Euphrates from Tiphsah to Gaza, over all the kings west of the Euphrates. And he had peace on all sides around him.
1KGS|4|25|And Judah and Israel lived in safety, from Dan even to Beersheba, every man under his vine and under his fig tree, all the days of Solomon.
1KGS|4|26|Solomon also had 40,000 stalls of horses for his chariots, and 12,000 horsemen.
1KGS|4|27|And those officers supplied provisions for King Solomon, and for all who came to King Solomon's table, each one in his month. They let nothing be lacking.
1KGS|4|28|Barley also and straw for the horses and swift steeds they brought to the place where it was required, each according to his duty.
1KGS|4|29|And God gave Solomon wisdom and understanding beyond measure, and breadth of mind like the sand on the seashore,
1KGS|4|30|so that Solomon's wisdom surpassed the wisdom of all the people of the east and all the wisdom of Egypt.
1KGS|4|31|For he was wiser than all other men, wiser than Ethan the Ezrahite, and Heman, Calcol, and Darda, the sons of Mahol, and his fame was in all the surrounding nations.
1KGS|4|32|He also spoke 3,000 proverbs, and his songs were 1,005.
1KGS|4|33|He spoke of trees, from the cedar that is in Lebanon to the hyssop that grows out of the wall. He spoke also of beasts, and of birds, and of reptiles, and of fish.
1KGS|4|34|And people of all nations came to hear the wisdom of Solomon, and from all the kings of the earth, who had heard of his wisdom.
1KGS|5|1|Now Hiram king of Tyre sent his servants to Solomon when he heard that they had anointed him king in place of his father, for Hiram always loved David.
1KGS|5|2|And Solomon sent word to Hiram,
1KGS|5|3|"You know that David my father could not build a house for the name of the LORD his God because of the warfare with which his enemies surrounded him, until the LORD put them under the soles of his feet.
1KGS|5|4|But now the LORD my God has given me rest on every side. There is neither adversary nor misfortune.
1KGS|5|5|And so I intend to build a house for the name of the LORD my God, as the LORD said to David my father, 'Your son, whom I will set on your throne in your place, shall build the house for my name.'
1KGS|5|6|Now therefore command that cedars of Lebanon be cut for me. And my servants will join your servants, and I will pay you for your servants such wages as you set, for you know that there is no one among us who knows how to cut timber like the Sidonians."
1KGS|5|7|As soon as Hiram heard the words of Solomon, he rejoiced greatly and said, "Blessed be the LORD this day, who has given to David a wise son to be over this great people."
1KGS|5|8|And Hiram sent to Solomon, saying, "I have heard the message that you have sent to me. I am ready to do all you desire in the matter of cedar and cypress timber.
1KGS|5|9|My servants shall bring it down to the sea from Lebanon, and I will make it into rafts to go by sea to the place you direct. And I will have them broken up there, and you shall receive it. And you shall meet my wishes by providing food for my household."
1KGS|5|10|So Hiram supplied Solomon with all the timber of cedar and cypress that he desired,
1KGS|5|11|while Solomon gave Hiram 20,000 cors of wheat as food for his household, and 20,000 cors of beaten oil. Solomon gave this to Hiram year by year.
1KGS|5|12|And the LORD gave Solomon wisdom, as he promised him. And there was peace between Hiram and Solomon, and the two of them made a treaty.
1KGS|5|13|King Solomon drafted forced labor out of all Israel, and the draft numbered 30,000 men.
1KGS|5|14|And he sent them to Lebanon, 10,000 a month in shifts. They would be a month in Lebanon and two months at home. Adoniram was in charge of the draft.
1KGS|5|15|Solomon also had 70,000 burden-bearers and 80,000 stonecutters in the hill country,
1KGS|5|16|besides Solomon's 3,300 chief officers who were over the work, who had charge of the people who carried on the work.
1KGS|5|17|At the king's command they quarried out great, costly stones in order to lay the foundation of the house with dressed stones.
1KGS|5|18|So Solomon's builders and Hiram's builders and the men of Gebal did the cutting and prepared the timber and the stone to build the house.
1KGS|6|1|In the four hundred and eightieth year after the people of Israel came out of the land of Egypt, in the fourth year of Solomon's reign over Israel, in the month of Ziv, which is the second month, he began to build the house of the LORD.
1KGS|6|2|The house that King Solomon built for the LORD was sixty cubits long, twenty cubits wide, and thirty cubits high.
1KGS|6|3|The vestibule in front of the nave of the house was twenty cubits long, equal to the width of the house, and ten cubits deep in front of the house.
1KGS|6|4|And he made for the house windows with recessed frames.
1KGS|6|5|He also built a structure against the wall of the house, running around the walls of the house, both the nave and the inner sanctuary. And he made side chambers all around.
1KGS|6|6|The lowest story was five cubits broad, the middle one was six cubits broad, and the third was seven cubits broad. For around the outside of the house he made offsets on the wall in order that the supporting beams should not be inserted into the walls of the house.
1KGS|6|7|When the house was built, it was with stone prepared at the quarry, so that neither hammer nor axe nor any tool of iron was heard in the temple while it was being built.
1KGS|6|8|The entrance for the lowest story was on the south side of the house, and one went up by stairs to the middle story, and from the middle story to the third.
1KGS|6|9|So he built the house and finished it, and he made the ceiling of the house of beams and planks of cedar.
1KGS|6|10|He built the structure against the whole house, five cubits high, and it was joined to the house with timbers of cedar.
1KGS|6|11|Now the word of the LORD came to Solomon,
1KGS|6|12|"Concerning this house that you are building, if you will walk in my statutes and obey my rules and keep all my commandments and walk in them, then I will establish my word with you, which I spoke to David your father.
1KGS|6|13|And I will dwell among the children of Israel and will not forsake my people Israel."
1KGS|6|14|So Solomon built the house and finished it.
1KGS|6|15|He lined the walls of the house on the inside with boards of cedar. From the floor of the house to the walls of the ceiling, he covered them on the inside with wood, and he covered the floor of the house with boards of cypress.
1KGS|6|16|He built twenty cubits of the rear of the house with boards of cedar from the floor to the walls, and he built this within as an inner sanctuary, as the Most Holy Place.
1KGS|6|17|The house, that is, the nave in front of the inner sanctuary, was forty cubits long.
1KGS|6|18|The cedar within the house was carved in the form of gourds and open flowers. All was cedar; no stone was seen.
1KGS|6|19|The inner sanctuary he prepared in the innermost part of the house, to set there the ark of the covenant of the LORD.
1KGS|6|20|The inner sanctuary was twenty cubits long, twenty cubits wide, and twenty cubits high, and he overlaid it with pure gold. He also overlaid an altar of cedar.
1KGS|6|21|And Solomon overlaid the inside of the house with pure gold, and he drew chains of gold across, in front of the inner sanctuary, and overlaid it with gold.
1KGS|6|22|And he overlaid the whole house with gold, until all the house was finished. Also the whole altar that belonged to the inner sanctuary he overlaid with gold.
1KGS|6|23|In the inner sanctuary he made two cherubim of olivewood, each ten cubits high.
1KGS|6|24|Five cubits was the length of one wing of the cherub, and five cubits the length of the other wing of the cherub; it was ten cubits from the tip of one wing to the tip of the other.
1KGS|6|25|The other cherub also measured ten cubits; both cherubim had the same measure and the same form.
1KGS|6|26|The height of one cherub was ten cubits, and so was that of the other cherub.
1KGS|6|27|He put the cherubim in the innermost part of the house. And the wings of the cherubim were spread out so that a wing of one touched the one wall, and a wing of the other cherub touched the other wall; their other wings touched each other in the middle of the house.
1KGS|6|28|And he overlaid the cherubim with gold.
1KGS|6|29|Around all the walls of the house he carved engraved figures of cherubim and palm trees and open flowers, in the inner and outer rooms.
1KGS|6|30|The floor of the house he overlaid with gold in the inner and outer rooms.
1KGS|6|31|For the entrance to the inner sanctuary he made doors of olivewood; the lintel and the doorposts were five-sided.
1KGS|6|32|He covered the two doors of olivewood with carvings of cherubim, palm trees, and open flowers. He overlaid them with gold and spread gold on the cherubim and on the palm trees.
1KGS|6|33|So also he made for the entrance to the nave doorposts of olivewood, in the form of a square,
1KGS|6|34|and two doors of cypress wood. The two leaves of the one door were folding, and the two leaves of the other door were folding.
1KGS|6|35|On them he carved cherubim and palm trees and open flowers, and he overlaid them with gold evenly applied on the carved work.
1KGS|6|36|He built the inner court with three courses of cut stone and one course of cedar beams.
1KGS|6|37|In the fourth year the foundation of the house of the LORD was laid, in the month of Ziv.
1KGS|6|38|And in the eleventh year, in the month of Bul, which is the eighth month, the house was finished in all its parts, and according to all its specifications. He was seven years in building it.
1KGS|7|1|Solomon was building his own house thirteen years, and he finished his entire house.
1KGS|7|2|He built the House of the Forest of Lebanon. Its length was a hundred cubits and its breadth fifty cubits and its height thirty cubits, and it was built on four rows of cedar pillars, with cedar beams on the pillars.
1KGS|7|3|And it was covered with cedar above the chambers that were on the forty-five pillars, fifteen in each row.
1KGS|7|4|There were window frames in three rows, and window opposite window in three tiers.
1KGS|7|5|All the doorways and windows had square frames, and window was opposite window in three tiers.
1KGS|7|6|And he made the Hall of Pillars; its length was fifty cubits, and its breadth thirty cubits. There was a porch in front with pillars, and a canopy in front of them.
1KGS|7|7|And he made the Hall of the Throne where he was to pronounce judgment, even the Hall of Judgment. It was finished with cedar from floor to rafters.
1KGS|7|8|His own house where he was to dwell, in the other court back of the hall, was of like workmanship. Solomon also made a house like this hall for Pharaoh's daughter whom he had taken in marriage.
1KGS|7|9|All these were made of costly stones, cut according to measure, sawed with saws, back and front, even from the foundation to the coping, and from the outside to the great court.
1KGS|7|10|The foundation was of costly stones, huge stones, stones of eight and ten cubits.
1KGS|7|11|And above were costly stones, cut according to measurement, and cedar.
1KGS|7|12|The great court had three courses of cut stone all around, and a course of cedar beams; so had the inner court of the house of the LORD and the vestibule of the house.
1KGS|7|13|And King Solomon sent and brought Hiram from Tyre.
1KGS|7|14|He was the son of a widow of the tribe of Naphtali, and his father was a man of Tyre, a worker in bronze. And he was full of wisdom, understanding, and skill for making any work in bronze. He came to King Solomon and did all his work.
1KGS|7|15|He cast two pillars of bronze. Eighteen cubits was the height of one pillar, and a line of twelve cubits measured its circumference. It was hollow, and its thickness was four fingers. The second pillar was the same.
1KGS|7|16|He also made two capitals of cast bronze to set on the tops of the pillars. The height of the one capital was five cubits, and the height of the other capital was five cubits.
1KGS|7|17|There were lattices of checker work with wreaths of chain work for the capitals on the tops of the pillars, a lattice for the one capital and a lattice for the other capital.
1KGS|7|18|Likewise he made pomegranates in two rows around the one latticework to cover the capital that was on the top of the pillar, and he did the same with the other capital.
1KGS|7|19|Now the capitals that were on the tops of the pillars in the vestibule were of lily-work, four cubits.
1KGS|7|20|The capitals were on the two pillars and also above the rounded projection which was beside the latticework. There were two hundred pomegranates in two rows all around, and so with the other capital.
1KGS|7|21|He set up the pillars at the vestibule of the temple. He set up the pillar on the south and called its name Jachin, and he set up the pillar on the north and called its name Boaz.
1KGS|7|22|And on the tops of the pillars was lily-work. Thus the work of the pillars was finished.
1KGS|7|23|Then he made the sea of cast metal. It was round, ten cubits from brim to brim, and five cubits high, and a line of thirty cubits measured its circumference.
1KGS|7|24|Under its brim were gourds, for ten cubits, compassing the sea all around. The gourds were in two rows, cast with it when it was cast.
1KGS|7|25|It stood on twelve oxen, three facing north, three facing west, three facing south, and three facing east. The sea was set on them, and all their rear parts were inward.
1KGS|7|26|Its thickness was a handbreadth, and its brim was made like the brim of a cup, like the flower of a lily. It held two thousand baths.
1KGS|7|27|He also made the ten stands of bronze. Each stand was four cubits long, four cubits wide, and three cubits high.
1KGS|7|28|This was the construction of the stands: they had panels, and the panels were set in the frames,
1KGS|7|29|and on the panels that were set in the frames were lions, oxen, and cherubim. On the frames, both above and below the lions and oxen, there were wreaths of beveled work.
1KGS|7|30|Moreover, each stand had four bronze wheels and axles of bronze, and at the four corners were supports for a basin. The supports were cast with wreaths at the side of each.
1KGS|7|31|Its opening was within a crown that projected upward one cubit. Its opening was round, as a pedestal is made, a cubit and a half deep. At its opening there were carvings, and its panels were square, not round.
1KGS|7|32|And the four wheels were underneath the panels. The axles of the wheels were of one piece with the stands, and the height of a wheel was a cubit and a half.
1KGS|7|33|The wheels were made like a chariot wheel; their axles, their rims, their spokes, and their hubs were all cast.
1KGS|7|34|There were four supports at the four corners of each stand. The supports were of one piece with the stands.
1KGS|7|35|And on the top of the stand there was a round band half a cubit high; and on the top of the stand its stays and its panels were of one piece with it.
1KGS|7|36|And on the surfaces of its stays and on its panels, he carved cherubim, lions, and palm trees, according to the space of each, with wreaths all around.
1KGS|7|37|After this manner he made the ten stands. All of them were cast alike, of the same measure and the same form.
1KGS|7|38|And he made ten basins of bronze. Each basin held forty baths, each basin measured four cubits, and there was a basin for each of the ten stands.
1KGS|7|39|And he set the stands, five on the south side of the house, and five on the north side of the house. And he set the sea at the southeast corner of the house.
1KGS|7|40|Hiram also made the pots, the shovels, and the basins. So Hiram finished all the work that he did for King Solomon on the house of the LORD:
1KGS|7|41|the two pillars, the two bowls of the capitals that were on the tops of the pillars, and the two latticeworks to cover the two bowls of the capitals that were on the tops of the pillars;
1KGS|7|42|and the four hundred pomegranates for the two latticeworks, two rows of pomegranates for each latticework, to cover the two bowls of the capitals that were on the pillars;
1KGS|7|43|the ten stands, and the ten basins on the stands;
1KGS|7|44|and the one sea, and the twelve oxen underneath the sea.
1KGS|7|45|Now the pots, the shovels, and the basins, all these vessels in the house of the LORD, which Hiram made for King Solomon, were of burnished bronze.
1KGS|7|46|In the plain of the Jordan the king cast them, in the clay ground between Succoth and Zarethan.
1KGS|7|47|And Solomon left all the vessels unweighed, because there were so many of them; the weight of the bronze was not ascertained.
1KGS|7|48|So Solomon made all the vessels that were in the house of the LORD: the golden altar, the golden table for the bread of the Presence,
1KGS|7|49|the lampstands of pure gold, five on the south side and five on the north, before the inner sanctuary; the flowers, the lamps, and the tongs, of gold;
1KGS|7|50|the cups, snuffers, basins, dishes for incense, and fire pans, of pure gold; and the sockets of gold, for the doors of the innermost part of the house, the Most Holy Place, and for the doors of the nave of the temple.
1KGS|7|51|Thus all the work that King Solomon did on the house of the LORD was finished. And Solomon brought in the things that David his father had dedicated, the silver, the gold, and the vessels, and stored them in the treasuries of the house of the LORD.
1KGS|8|1|Then Solomon assembled the elders of Israel and all the heads of the tribes, the leaders of the fathers' houses of the people of Israel, before King Solomon in Jerusalem, to bring up the ark of the covenant of the LORD out of the city of David, which is Zion.
1KGS|8|2|And all the men of Israel assembled to King Solomon at the feast in the month Ethanim, which is the seventh month.
1KGS|8|3|And all the elders of Israel came, and the priests took up the ark.
1KGS|8|4|And they brought up the ark of the LORD, the tent of meeting, and all the holy vessels that were in the tent; the priests and the Levites brought them up.
1KGS|8|5|And King Solomon and all the congregation of Israel, who had assembled before him, were with him before the ark, sacrificing so many sheep and oxen that they could not be counted or numbered.
1KGS|8|6|Then the priests brought the ark of the covenant of the LORD to its place in the inner sanctuary of the house, in the Most Holy Place, underneath the wings of the cherubim.
1KGS|8|7|For the cherubim spread out their wings over the place of the ark, so that the cherubim overshadowed the ark and its poles.
1KGS|8|8|And the poles were so long that the ends of the poles were seen from the Holy Place before the inner sanctuary; but they could not be seen from outside. And they are there to this day.
1KGS|8|9|There was nothing in the ark except the two tablets of stone that Moses put there at Horeb, where the LORD made a covenant with the people of Israel, when they came out of the land of Egypt.
1KGS|8|10|And when the priests came out of the Holy Place, a cloud filled the house of the LORD,
1KGS|8|11|so that the priests could not stand to minister because of the cloud, for the glory of the LORD filled the house of the LORD.
1KGS|8|12|Then Solomon said, "The LORD has said that he would dwell in thick darkness.
1KGS|8|13|I have indeed built you an exalted house, a place for you to dwell in forever."
1KGS|8|14|Then the king turned around and blessed all the assembly of Israel, while all the assembly of Israel stood.
1KGS|8|15|And he said, "Blessed be the LORD, the God of Israel, who with his hand has fulfilled what he promised with his mouth to David my father, saying,
1KGS|8|16|'Since the day that I brought my people Israel out of Egypt, I chose no city out of all the tribes of Israel in which to build a house, that my name might be there. But I chose David to be over my people Israel.'
1KGS|8|17|Now it was in the heart of David my father to build a house for the name of the LORD, the God of Israel.
1KGS|8|18|But the LORD said to David my father, 'Whereas it was in your heart to build a house for my name, you did well that it was in your heart.
1KGS|8|19|Nevertheless, you shall not build the house, but your son who shall be born to you shall build the house for my name.'
1KGS|8|20|Now the LORD has fulfilled his promise that he made. For I have risen in the place of David my father, and sit on the throne of Israel, as the LORD promised, and I have built the house for the name of the LORD, the God of Israel.
1KGS|8|21|And there I have provided a place for the ark, in which is the covenant of the LORD that he made with our fathers, when he brought them out of the land of Egypt."
1KGS|8|22|Then Solomon stood before the altar of the LORD in the presence of all the assembly of Israel and spread out his hands toward heaven,
1KGS|8|23|and said, "O LORD, God of Israel, there is no God like you, in heaven above or on earth beneath, keeping covenant and showing steadfast love to your servants who walk before you with all their heart,
1KGS|8|24|who have kept with your servant David my father what you declared to him. You spoke with your mouth, and with your hand have fulfilled it this day.
1KGS|8|25|Now therefore, O LORD, God of Israel, keep for your servant David my father what you have promised him, saying, 'You shall not lack a man to sit before me on the throne of Israel, if only your sons pay close attention to their way, to walk before me as you have walked before me.'
1KGS|8|26|Now therefore, O God of Israel, let your word be confirmed, which you have spoken to your servant David my father.
1KGS|8|27|"But will God indeed dwell on the earth? Behold, heaven and the highest heaven cannot contain you; how much less this house that I have built!
1KGS|8|28|Yet have regard to the prayer of your servant and to his plea, O LORD my God, listening to the cry and to the prayer that your servant prays before you this day,
1KGS|8|29|that your eyes may be open night and day toward this house, the place of which you have said, 'My name shall be there,' that you may listen to the prayer that your servant offers toward this place.
1KGS|8|30|And listen to the plea of your servant and of your people Israel, when they pray toward this place. And listen in heaven your dwelling place, and when you hear, forgive.
1KGS|8|31|"If a man sins against his neighbor and is made to take an oath and comes and swears his oath before your altar in this house,
1KGS|8|32|then hear in heaven and act and judge your servants, condemning the guilty by bringing his conduct on his own head, and vindicating the righteous by rewarding him according to his righteousness.
1KGS|8|33|"When your people Israel are defeated before the enemy because they have sinned against you, and if they turn again to you and acknowledge your name and pray and plead with you in this house,
1KGS|8|34|then hear in heaven and forgive the sin of your people Israel and bring them again to the land that you gave to their fathers.
1KGS|8|35|"When heaven is shut up and there is no rain because they have sinned against you, if they pray toward this place and acknowledge your name and turn from their sin, when you afflict them,
1KGS|8|36|then hear in heaven and forgive the sin of your servants, your people Israel, when you teach them the good way in which they should walk, and grant rain upon your land, which you have given to your people as an inheritance.
1KGS|8|37|"If there is famine in the land, if there is pestilence or blight or mildew or locust or caterpillar, if their enemy besieges them in the land at their gates, whatever plague, whatever sickness there is,
1KGS|8|38|whatever prayer, whatever plea is made by any man or by all your people Israel, each knowing the affliction of his own heart and stretching out his hands toward this house,
1KGS|8|39|then hear in heaven your dwelling place and forgive and act and render to each whose heart you know, according to all his ways (for you, you only, know the hearts of all the children of mankind),
1KGS|8|40|that they may fear you all the days that they live in the land that you gave to our fathers.
1KGS|8|41|"Likewise, when a foreigner, who is not of your people Israel, comes from a far country for your name's sake
1KGS|8|42|(for they shall hear of your great name and your mighty hand, and of your outstretched arm), when he comes and prays toward this house,
1KGS|8|43|hear in heaven your dwelling place and do according to all for which the foreigner calls to you, in order that all the peoples of the earth may know your name and fear you, as do your people Israel, and that they may know that this house that I have built is called by your name.
1KGS|8|44|"If your people go out to battle against their enemy, by whatever way you shall send them, and they pray to the LORD toward the city that you have chosen and the house that I have built for your name,
1KGS|8|45|then hear in heaven their prayer and their plea, and maintain their cause.
1KGS|8|46|"If they sin against you- for there is no one who does not sin- and you are angry with them and give them to an enemy, so that they are carried away captive to the land of the enemy, far off or near,
1KGS|8|47|yet if they turn their heart in the land to which they have been carried captive, and repent and plead with you in the land of their captors, saying, 'We have sinned and have acted perversely and wickedly,'
1KGS|8|48|if they repent with all their mind and with all their heart in the land of their enemies, who carried them captive, and pray to you toward their land, which you gave to their fathers, the city that you have chosen, and the house that I have built for your name,
1KGS|8|49|then hear in heaven your dwelling place their prayer and their plea, and maintain their cause
1KGS|8|50|and forgive your people who have sinned against you, and all their transgressions that they have committed against you, and grant them compassion in the sight of those who carried them captive, that they may have compassion on them
1KGS|8|51|(for they are your people, and your heritage, which you brought out of Egypt, from the midst of the iron furnace).
1KGS|8|52|Let your eyes be open to the plea of your servant and to the plea of your people Israel, giving ear to them whenever they call to you.
1KGS|8|53|For you separated them from among all the peoples of the earth to be your heritage, as you declared through Moses your servant, when you brought our fathers out of Egypt, O Lord GOD."
1KGS|8|54|Now as Solomon finished offering all this prayer and plea to the LORD, he arose from before the altar of the LORD, where he had knelt with hands outstretched toward heaven.
1KGS|8|55|And he stood and blessed all the assembly of Israel with a loud voice, saying,
1KGS|8|56|"Blessed be the LORD who has given rest to his people Israel, according to all that he promised. Not one word has failed of all his good promise, which he spoke by Moses his servant.
1KGS|8|57|The LORD our God be with us, as he was with our fathers. May he not leave us or forsake us,
1KGS|8|58|that he may incline our hearts to him, to walk in all his ways and to keep his commandments, his statutes, and his rules, which he commanded our fathers.
1KGS|8|59|Let these words of mine, with which I have pleaded before the LORD, be near to the LORD our God day and night, and may he maintain the cause of his servant and the cause of his people Israel, as each day requires,
1KGS|8|60|that all the peoples of the earth may know that the LORD is God; there is no other.
1KGS|8|61|Let your heart therefore be wholly true to the LORD our God, walking in his statutes and keeping his commandments, as at this day."
1KGS|8|62|Then the king, and all Israel with him, offered sacrifice before the LORD.
1KGS|8|63|Solomon offered as peace offerings to the LORD 22,000 oxen and 120,000 sheep. So the king and all the people of Israel dedicated the house of the LORD.
1KGS|8|64|The same day the king consecrated the middle of the court that was before the house of the LORD, for there he offered the burnt offering and the grain offering and the fat pieces of the peace offerings, because the bronze altar that was before the LORD was too small to receive the burnt offering and the grain offering and the fat pieces of the peace offerings.
1KGS|8|65|So Solomon held the feast at that time, and all Israel with him, a great assembly, from Lebo-hamath to the Brook of Egypt, before the LORD our God, seven days.
1KGS|8|66|On the eighth day he sent the people away, and they blessed the king and went to their homes joyful and glad of heart for all the goodness that the LORD had shown to David his servant and to Israel his people.
1KGS|9|1|As soon as Solomon had finished building the house of the LORD and the king's house and all that Solomon desired to build,
1KGS|9|2|the LORD appeared to Solomon a second time, as he had appeared to him at Gibeon.
1KGS|9|3|And the LORD said to him, "I have heard your prayer and your plea, which you have made before me. I have consecrated this house that you have built, by putting my name there forever. My eyes and my heart will be there for all time.
1KGS|9|4|And as for you, if you will walk before me, as David your father walked, with integrity of heart and uprightness, doing according to all that I have commanded you, and keeping my statutes and my rules,
1KGS|9|5|then I will establish your royal throne over Israel forever, as I promised David your father, saying, 'You shall not lack a man on the throne of Israel.'
1KGS|9|6|But if you turn aside from following me, you or your children, and do not keep my commandments and my statutes that I have set before you, but go and serve other gods and worship them,
1KGS|9|7|then I will cut off Israel from the land that I have given them, and the house that I have consecrated for my name I will cast out of my sight, and Israel will become a proverb and a byword among all peoples.
1KGS|9|8|And this house will become a heap of ruins. Everyone passing by it will be astonished and will hiss, and they will say, 'Why has the LORD done thus to this land and to this house?'
1KGS|9|9|Then they will say, 'Because they abandoned the LORD their God who brought their fathers out of the land of Egypt and laid hold on other gods and worshiped them and served them. Therefore the LORD has brought all this disaster on them.'"
1KGS|9|10|At the end of twenty years, in which Solomon had built the two houses, the house of the LORD and the king's house,
1KGS|9|11|and Hiram king of Tyre had supplied Solomon with cedar and cypress timber and gold, as much as he desired, King Solomon gave to Hiram twenty cities in the land of Galilee.
1KGS|9|12|But when Hiram came from Tyre to see the cities that Solomon had given him, they did not please him.
1KGS|9|13|Therefore he said, "What kind of cities are these that you have given me, my brother?" So they are called the land of Cabul to this day.
1KGS|9|14|Hiram had sent to the king 120 talents of gold.
1KGS|9|15|And this is the account of the forced labor that King Solomon drafted to build the house of the LORD and his own house and the Millo and the wall of Jerusalem and Hazor and Megiddo and Gezer
1KGS|9|16|(Pharaoh king of Egypt had gone up and captured Gezer and burned it with fire, and had killed the Canaanites who lived in the city, and had given it as dowry to his daughter, Solomon's wife;
1KGS|9|17|so Solomon rebuilt Gezer) and Lower Beth-horon
1KGS|9|18|and Baalath and Tamar in the wilderness, in the land of Judah,
1KGS|9|19|and all the store cities that Solomon had, and the cities for his chariots, and the cities for his horsemen, and whatever Solomon desired to build in Jerusalem, in Lebanon, and in all the land of his dominion.
1KGS|9|20|All the people who were left of the Amorites, the Hittites, the Perizzites, the Hivites, and the Jebusites, who were not of the people of Israel-
1KGS|9|21|their descendants who were left after them in the land, whom the people of Israel were unable to devote to destruction- these Solomon drafted to be slaves, and so they are to this day.
1KGS|9|22|But of the people of Israel Solomon made no slaves. They were the soldiers, they were his officials, his commanders, his captains, his chariot commanders and his horsemen.
1KGS|9|23|These were the chief officers who were over Solomon's work: 550 who had charge of the people who carried on the work.
1KGS|9|24|But Pharaoh's daughter went up from the city of David to her own house that Solomon had built for her. Then he built the Millo.
1KGS|9|25|Three times a year Solomon used to offer up burnt offerings and peace offerings on the altar that he built to the LORD, making offerings with it before the LORD. So he finished the house.
1KGS|9|26|King Solomon built a fleet of ships at Ezion-geber, which is near Eloth on the shore of the Red Sea, in the land of Edom.
1KGS|9|27|And Hiram sent with the fleet his servants, seamen who were familiar with the sea, together with the servants of Solomon.
1KGS|9|28|And they went to Ophir and brought from there gold, 420 talents, and they brought it to King Solomon.
1KGS|10|1|Now when the queen of Sheba heard of the fame of Solomon concerning the name of the LORD, she came to test him with hard questions.
1KGS|10|2|She came to Jerusalem with a very great retinue, with camels bearing spices and very much gold and precious stones. And when she came to Solomon, she told him all that was on her mind.
1KGS|10|3|And Solomon answered all her questions; there was nothing hidden from the king that he could not explain to her.
1KGS|10|4|And when the queen of Sheba had seen all the wisdom of Solomon, the house that he had built,
1KGS|10|5|the food of his table, the seating of his officials, and the attendance of his servants, their clothing, his cupbearers, and his burnt offerings that he offered at the house of the LORD, there was no more breath in her.
1KGS|10|6|And she said to the king, "The report was true that I heard in my own land of your words and of your wisdom,
1KGS|10|7|but I did not believe the reports until I came and my own eyes had seen it. And behold, the half was not told me. Your wisdom and prosperity surpass the report that I heard.
1KGS|10|8|Happy are your men! Happy are your servants, who continually stand before you and hear your wisdom!
1KGS|10|9|Blessed be the LORD your God, who has delighted in you and set you on the throne of Israel! Because the LORD loved Israel forever, he has made you king, that you may execute justice and righteousness."
1KGS|10|10|Then she gave the king 120 talents of gold, and a very great quantity of spices and precious stones. Never again came such an abundance of spices as these that the queen of Sheba gave to King Solomon.
1KGS|10|11|Moreover, the fleet of Hiram, which brought gold from Ophir, brought from Ophir a very great amount of almug wood and precious stones.
1KGS|10|12|And the king made of the almug wood supports for the house of the LORD and for the king's house, also lyres and harps for the singers. No such almug wood has come or been seen to this day.
1KGS|10|13|And King Solomon gave to the queen of Sheba all that she desired, whatever she asked besides what was given her by the bounty of King Solomon. So she turned and went back to her own land with her servants.
1KGS|10|14|Now the weight of gold that came to Solomon in one year was 666 talents of gold,
1KGS|10|15|besides that which came from the explorers and from the business of the merchants, and from all the kings of the west and from the governors of the land.
1KGS|10|16|King Solomon made 200 large shields of beaten gold; 600 shekels of gold went into each shield.
1KGS|10|17|And he made 300 shields of beaten gold; three minas of gold went into each shield. And the king put them in the House of the Forest of Lebanon.
1KGS|10|18|The king also made a great ivory throne and overlaid it with the finest gold.
1KGS|10|19|The throne had six steps, and at the back of the throne was a calf's head, and on each side of the seat were armrests and two lions standing beside the armrests,
1KGS|10|20|while twelve lions stood there, one on each end of a step on the six steps. The like of it was never made in any kingdom.
1KGS|10|21|All King Solomon's drinking vessels were of gold, and all the vessels of the House of the Forest of Lebanon were of pure gold. None were of silver; silver was not considered as anything in the days of Solomon.
1KGS|10|22|For the king had a fleet of ships of Tarshish at sea with the fleet of Hiram. Once every three years the fleet of ships of Tarshish used to come bringing gold, silver, ivory, apes, and peacocks.
1KGS|10|23|Thus King Solomon excelled all the kings of the earth in riches and in wisdom.
1KGS|10|24|And the whole earth sought the presence of Solomon to hear his wisdom, which God had put into his mind.
1KGS|10|25|Every one of them brought his present, articles of silver and gold, garments, myrrh, spices, horses, and mules, so much year by year.
1KGS|10|26|And Solomon gathered together chariots and horsemen. He had 1,400 chariots and 12,000 horsemen, whom he stationed in the chariot cities and with the king in Jerusalem.
1KGS|10|27|And the king made silver as common in Jerusalem as stone, and he made cedar as plentiful as the sycamore of the Shephelah.
1KGS|10|28|And Solomon's import of horses was from Egypt and Kue, and the king's traders received them from Kue at a price.
1KGS|10|29|A chariot could be imported from Egypt for 600 shekels of silver and a horse for 150, and so through the king's traders they were exported to all the kings of the Hittites and the kings of Syria.
1KGS|11|1|Now King Solomon loved many foreign women, along with the daughter of Pharaoh: Moabite, Ammonite, Edomite, Sidonian, and Hittite women,
1KGS|11|2|from the nations concerning which the LORD had said to the people of Israel, "You shall not enter into marriage with them, neither shall they with you, for surely they will turn away your heart after their gods." Solomon clung to these in love.
1KGS|11|3|He had 700 wives, princesses, and 300 concubines. And his wives turned away his heart.
1KGS|11|4|For when Solomon was old his wives turned away his heart after other gods, and his heart was not wholly true to the LORD his God, as was the heart of David his father.
1KGS|11|5|For Solomon went after Ashtoreth the goddess of the Sidonians, and after Milcom the abomination of the Ammonites.
1KGS|11|6|So Solomon did what was evil in the sight of the LORD and did not wholly follow the LORD, as David his father had done.
1KGS|11|7|Then Solomon built a high place for Chemosh the abomination of Moab, and for Molech the abomination of the Ammonites, on the mountain east of Jerusalem.
1KGS|11|8|And so he did for all his foreign wives, who made offerings and sacrificed to their gods.
1KGS|11|9|And the LORD was angry with Solomon, because his heart had turned away from the LORD, the God of Israel, who had appeared to him twice
1KGS|11|10|and had commanded him concerning this thing, that he should not go after other gods. But he did not keep what the LORD commanded.
1KGS|11|11|Therefore the LORD said to Solomon, "Since this has been your practice and you have not kept my covenant and my statutes that I have commanded you, I will surely tear the kingdom from you and will give it to your servant.
1KGS|11|12|Yet for the sake of David your father I will not do it in your days, but I will tear it out of the hand of your son.
1KGS|11|13|However, I will not tear away all the kingdom, but I will give one tribe to your son, for the sake of David my servant and for the sake of Jerusalem that I have chosen."
1KGS|11|14|And the LORD raised up an adversary against Solomon, Hadad the Edomite. He was of the royal house in Edom.
1KGS|11|15|For when David was in Edom, and Joab the commander of the army went up to bury the slain, he struck down every male in Edom
1KGS|11|16|(for Joab and all Israel remained there six months, until he had cut off every male in Edom).
1KGS|11|17|But Hadad fled to Egypt, together with certain Edomites of his father's servants, Hadad still being a little child.
1KGS|11|18|They set out from Midian and came to Paran and took men with them from Paran and came to Egypt, to Pharaoh king of Egypt, who gave him a house and assigned him an allowance of food and gave him land.
1KGS|11|19|And Hadad found great favor in the sight of Pharaoh, so that he gave him in marriage the sister of his own wife, the sister of Tahpenes the queen.
1KGS|11|20|And the sister of Tahpenes bore him Genubath his son, whom Tahpenes weaned in Pharaoh's house. And Genubath was in Pharaoh's house among the sons of Pharaoh.
1KGS|11|21|But when Hadad heard in Egypt that David slept with his fathers and that Joab the commander of the army was dead, Hadad said to Pharaoh, "Let me depart, that I may go to my own country."
1KGS|11|22|But Pharaoh said to him, "What have you lacked with me that you are now seeking to go to your own country?" And he said to him, "Only let me depart."
1KGS|11|23|God also raised up as an adversary to him, Rezon the son of Eliada, who had fled from his master Hadadezer king of Zobah.
1KGS|11|24|And he gathered men about him and became leader of a marauding band, after the killing by David. And they went to Damascus and lived there and made him king in Damascus.
1KGS|11|25|He was an adversary of Israel all the days of Solomon, doing harm as Hadad did. And he loathed Israel and reigned over Syria.
1KGS|11|26|Jeroboam the son of Nebat, an Ephraimite of Zeredah, a servant of Solomon, whose mother's name was Zeruah, a widow, also lifted up his hand against the king.
1KGS|11|27|And this was the reason why he lifted up his hand against the king. Solomon built the Millo, and closed up the breach of the city of David his father.
1KGS|11|28|The man Jeroboam was very able, and when Solomon saw that the young man was industrious he gave him charge over all the forced labor of the house of Joseph.
1KGS|11|29|And at that time, when Jeroboam went out of Jerusalem, the prophet Ahijah the Shilonite found him on the road. Now Ahijah had dressed himself in a new garment, and the two of them were alone in the open country.
1KGS|11|30|Then Ahijah laid hold of the new garment that was on him, and tore it into twelve pieces.
1KGS|11|31|And he said to Jeroboam, "Take for yourself ten pieces, for thus says the LORD, the God of Israel, 'Behold, I am about to tear the kingdom from the hand of Solomon and will give you ten tribes
1KGS|11|32|(but he shall have one tribe, for the sake of my servant David and for the sake of Jerusalem, the city that I have chosen out of all the tribes of Israel),
1KGS|11|33|because they have forsaken me and worshiped Ashtoreth the goddess of the Sidonians, Chemosh the god of Moab, and Milcom the god of the Ammonites, and they have not walked in my ways, doing what is right in my sight and keeping my statutes and my rules, as David his father did.
1KGS|11|34|Nevertheless, I will not take the whole kingdom out of his hand, but I will make him ruler all the days of his life, for the sake of David my servant whom I chose, who kept my commandments and my statutes.
1KGS|11|35|But I will take the kingdom out of his son's hand and will give it to you, ten tribes.
1KGS|11|36|Yet to his son I will give one tribe, that David my servant may always have a lamp before me in Jerusalem, the city where I have chosen to put my name.
1KGS|11|37|And I will take you, and you shall reign over all that your soul desires, and you shall be king over Israel.
1KGS|11|38|And if you will listen to all that I command you, and will walk in my ways, and do what is right in my eyes by keeping my statutes and my commandments, as David my servant did, I will be with you and will build you a sure house, as I built for David, and I will give Israel to you.
1KGS|11|39|And I will afflict the offspring of David because of this, but not forever.'"
1KGS|11|40|Solomon sought therefore to kill Jeroboam. But Jeroboam arose and fled into Egypt, to Shishak king of Egypt, and was in Egypt until the death of Solomon.
1KGS|11|41|Now the rest of the acts of Solomon, and all that he did, and his wisdom, are they not written in the Book of the Acts of Solomon?
1KGS|11|42|And the time that Solomon reigned in Jerusalem over all Israel was forty years.
1KGS|11|43|And Solomon slept with his fathers and was buried in the city of David his father. And Rehoboam his son reigned in his place.
1KGS|12|1|Rehoboam went to Shechem, for all Israel had come to Shechem to make him king.
1KGS|12|2|And as soon as Jeroboam the son of Nebat heard of it (for he was still in Egypt, where he had fled from King Solomon), then Jeroboam returned from Egypt.
1KGS|12|3|And they sent and called him, and Jeroboam and all the assembly of Israel came and said to Rehoboam,
1KGS|12|4|"Your father made our yoke heavy. Now therefore lighten the hard service of your father and his heavy yoke on us, and we will serve you."
1KGS|12|5|He said to them, "Go away for three days, then come again to me." So the people went away.
1KGS|12|6|Then King Rehoboam took counsel with the old men, who had stood before Solomon his father while he was yet alive, saying, "How do you advise me to answer this people?"
1KGS|12|7|And they said to him, "If you will be a servant to this people today and serve them, and speak good words to them when you answer them, then they will be your servants forever."
1KGS|12|8|But he abandoned the counsel that the old men gave him and took counsel with the young men who had grown up with him and stood before him.
1KGS|12|9|And he said to them, "What do you advise that we answer this people who have said to me, 'Lighten the yoke that your father put on us'?"
1KGS|12|10|And the young men who had grown up with him said to him, "Thus shall you speak to this people who said to you, 'Your father made our yoke heavy, but you lighten it for us,' thus shall you say to them, 'My little finger is thicker than my father's thighs.
1KGS|12|11|And now, whereas my father laid on you a heavy yoke, I will add to your yoke. My father disciplined you with whips, but I will discipline you with scorpions.'"
1KGS|12|12|So Jeroboam and all the people came to Rehoboam the third day, as the king said, "Come to me again the third day."
1KGS|12|13|And the king answered the people harshly, and forsaking the counsel that the old men had given him,
1KGS|12|14|he spoke to them according to the counsel of the young men, saying, "My father made your yoke heavy, but I will add to your yoke. My father disciplined you with whips, but I will discipline you with scorpions."
1KGS|12|15|So the king did not listen to the people, for it was a turn of affairs brought about by the LORD that he might fulfill his word, which the LORD spoke by Ahijah the Shilonite to Jeroboam the son of Nebat.
1KGS|12|16|And when all Israel saw that the king did not listen to them, the people answered the king, "What portion do we have in David? We have no inheritance in the son of Jesse. To your tents, O Israel! Look now to your own house, David." So Israel went to their tents.
1KGS|12|17|But Rehoboam reigned over the people of Israel who lived in the cities of Judah.
1KGS|12|18|Then King Rehoboam sent Adoram, who was taskmaster over the forced labor, and all Israel stoned him to death with stones. And King Rehoboam hurried to mount his chariot to flee to Jerusalem.
1KGS|12|19|So Israel has been in rebellion against the house of David to this day.
1KGS|12|20|And when all Israel heard that Jeroboam had returned, they sent and called him to the assembly and made him king over all Israel. There was none that followed the house of David but the tribe of Judah only.
1KGS|12|21|When Rehoboam came to Jerusalem, he assembled all the house of Judah and the tribe of Benjamin, 180,000 chosen warriors, to fight against the house of Israel, to restore the kingdom to Rehoboam the son of Solomon.
1KGS|12|22|But the word of God came to Shemaiah the man of God:
1KGS|12|23|"Say to Rehoboam the son of Solomon, king of Judah, and to all the house of Judah and Benjamin, and to the rest of the people,
1KGS|12|24|'Thus says the LORD, You shall not go up or fight against your relatives the people of Israel. Every man return to his home, for this thing is from me.'"So they listened to the word of the LORD and went home again, according to the word of the LORD.
1KGS|12|25|Then Jeroboam built Shechem in the hill country of Ephraim and lived there. And he went out from there and built Penuel.
1KGS|12|26|And Jeroboam said in his heart, "Now the kingdom will turn back to the house of David.
1KGS|12|27|If this people go up to offer sacrifices in the temple of the LORD at Jerusalem, then the heart of this people will turn again to their lord, to Rehoboam king of Judah, and they will kill me and return to Rehoboam king of Judah."
1KGS|12|28|So the king took counsel and made two calves of gold. And he said to the people, "You have gone up to Jerusalem long enough. Behold your gods, O Israel, who brought you up out of the land of Egypt."
1KGS|12|29|And he set one in Bethel, and the other he put in Dan.
1KGS|12|30|Then this thing became a sin, for the people went as far as Dan to be before one.
1KGS|12|31|He also made temples on high places and appointed priests from among all the people, who were not of the Levites.
1KGS|12|32|And Jeroboam appointed a feast on the fifteenth day of the eighth month like the feast that was in Judah, and he offered sacrifices on the altar. So he did in Bethel, sacrificing to the calves that he made. And he placed in Bethel the priests of the high places that he had made.
1KGS|12|33|He went up to the altar that he had made in Bethel on the fifteenth day in the eighth month, in the month that he had devised from his own heart. And he instituted a feast for the people of Israel and went up to the altar to make offerings.
1KGS|13|1|And behold, a man of God came out of Judah by the word of the LORD to Bethel. Jeroboam was standing by the altar to make offerings.
1KGS|13|2|And the man cried against the altar by the word of the LORD and said, "O altar, altar, thus says the LORD: 'Behold, a son shall be born to the house of David, Josiah by name, and he shall sacrifice on you the priests of the high places who make offerings on you, and human bones shall be burned on you.'"
1KGS|13|3|And he gave a sign the same day, saying, "This is the sign that the LORD has spoken: 'Behold, the altar shall be torn down, and the ashes that are on it shall be poured out.'"
1KGS|13|4|And when the king heard the saying of the man of God, which he cried against the altar at Bethel, Jeroboam stretched out his hand from the altar, saying, "Seize him." And his hand, which he stretched out against him, dried up, so that he could not draw it back to himself.
1KGS|13|5|The altar also was torn down, and the ashes poured out from the altar, according to the sign that the man of God had given by the word of the LORD.
1KGS|13|6|And the king said to the man of God, "Entreat now the favor of the LORD your God, and pray for me, that my hand may be restored to me." And the man of God entreated the LORD, and the king's hand was restored to him and became as it was before.
1KGS|13|7|And the king said to the man of God, "Come home with me, and refresh yourself, and I will give you a reward."
1KGS|13|8|And the man of God said to the king, "If you give me half your house, I will not go in with you. And I will not eat bread or drink water in this place,
1KGS|13|9|for so was it commanded me by the word of the LORD, saying, 'You shall neither eat bread nor drink water nor return by the way that you came.'"
1KGS|13|10|So he went another way and did not return by the way that he came to Bethel.
1KGS|13|11|Now an old prophet lived in Bethel. And his sons came and told him all that the man of God had done that day in Bethel. They also told to their father the words that he had spoken to the king.
1KGS|13|12|And their father said to them, "Which way did he go?" And his sons showed him the way that the man of God who came from Judah had gone.
1KGS|13|13|And he said to his sons, "Saddle the donkey for me." So they saddled the donkey for him and he mounted it.
1KGS|13|14|And he went after the man of God and found him sitting under an oak. And he said to him, "Are you the man of God who came from Judah?" And he said, "I am."
1KGS|13|15|Then he said to him, "Come home with me and eat bread."
1KGS|13|16|And he said, "I may not return with you, or go in with you, neither will I eat bread nor drink water with you in this place,
1KGS|13|17|for it was said to me by the word of the LORD, 'You shall neither eat bread nor drink water there, nor return by the way that you came.'"
1KGS|13|18|And he said to him, "I also am a prophet as you are, and an angel spoke to me by the word of the LORD, saying, 'Bring him back with you into your house that he may eat bread and drink water.'"But he lied to him.
1KGS|13|19|So he went back with him and ate bread in his house and drank water.
1KGS|13|20|And as they sat at the table, the word of the LORD came to the prophet who had brought him back.
1KGS|13|21|And he cried to the man of God who came from Judah, "Thus says the LORD, 'Because you have disobeyed the word of the LORD and have not kept the command that the LORD your God commanded you,
1KGS|13|22|but have come back and have eaten bread and drunk water in the place of which he said to you, "Eat no bread and drink no water," your body shall not come to the tomb of your fathers.'"
1KGS|13|23|And after he had eaten bread and drunk, he saddled the donkey for the prophet whom he had brought back.
1KGS|13|24|And as he went away a lion met him on the road and killed him. And his body was thrown in the road, and the donkey stood beside it; the lion also stood beside the body.
1KGS|13|25|And behold, men passed by and saw the body thrown in the road and the lion standing by the body. And they came and told it in the city where the old prophet lived.
1KGS|13|26|And when the prophet who had brought him back from the way heard of it, he said, "It is the man of God who disobeyed the word of the LORD; therefore the LORD has given him to the lion, which has torn him and killed him, according to the word that the LORD spoke to him."
1KGS|13|27|And he said to his sons, "Saddle the donkey for me." And they saddled it.
1KGS|13|28|And he went and found his body thrown in the road, and the donkey and the lion standing beside the body. The lion had not eaten the body or torn the donkey.
1KGS|13|29|And the prophet took up the body of the man of God and laid it on the donkey and brought it back to the city to mourn and to bury him.
1KGS|13|30|And he laid the body in his own grave. And they mourned over him, saying, "Alas, my brother!"
1KGS|13|31|And after he had buried him, he said to his sons, "When I die, bury me in the grave in which the man of God is buried; lay my bones beside his bones.
1KGS|13|32|For the saying that he called out by the word of the LORD against the altar in Bethel and against all the houses of the high places that are in the cities of Samaria shall surely come to pass."
1KGS|13|33|After this thing Jeroboam did not turn from his evil way, but made priests for the high places again from among all the people. Any who would, he ordained to be priests of the high places.
1KGS|13|34|And this thing became sin to the house of Jeroboam, so as to cut it off and to destroy it from the face of the earth.
1KGS|14|1|At that time Abijah the son of Jeroboam fell sick.
1KGS|14|2|And Jeroboam said to his wife, "Arise, and disguise yourself, that it not be known that you are the wife of Jeroboam, and go to Shiloh. Behold, Ahijah the prophet is there, who said of me that I should be king over this people.
1KGS|14|3|Take with you ten loaves, some cakes, and a jar of honey, and go to him. He will tell you what shall happen to the child."
1KGS|14|4|Jeroboam's wife did so. She arose and went to Shiloh and came to the house of Ahijah. Now Ahijah could not see, for his eyes were dim because of his age.
1KGS|14|5|And the LORD said to Ahijah, "Behold, the wife of Jeroboam is coming to inquire of you concerning her son, for he is sick. Thus and thus shall you say to her." When she came, she pretended to be another woman.
1KGS|14|6|But when Ahijah heard the sound of her feet, as she came in at the door, he said, "Come in, wife of Jeroboam. Why do you pretend to be another? For I am charged with unbearable news for you.
1KGS|14|7|Go, tell Jeroboam, 'Thus says the LORD, the God of Israel: "Because I exalted you from among the people and made you leader over my people Israel
1KGS|14|8|and tore the kingdom away from the house of David and gave it to you, and yet you have not been like my servant David, who kept my commandments and followed me with all his heart, doing only that which was right in my eyes,
1KGS|14|9|but you have done evil above all who were before you and have gone and made for yourself other gods and metal images, provoking me to anger, and have cast me behind your back,
1KGS|14|10|therefore behold, I will bring harm upon the house of Jeroboam and will cut off from Jeroboam every male, both bond and free in Israel, and will burn up the house of Jeroboam, as a man burns up dung until it is all gone.
1KGS|14|11|Anyone belonging to Jeroboam who dies in the city the dogs shall eat, and anyone who dies in the open country the birds of the heavens shall eat, for the LORD has spoken it."'
1KGS|14|12|Arise therefore, go to your house. When your feet enter the city, the child shall die.
1KGS|14|13|And all Israel shall mourn for him and bury him, for he only of Jeroboam shall come to the grave, because in him there is found something pleasing to the LORD, the God of Israel, in the house of Jeroboam.
1KGS|14|14|Moreover, the LORD will raise up for himself a king over Israel who shall cut off the house of Jeroboam today. And henceforth,
1KGS|14|15|the LORD will strike Israel as a reed is shaken in the water, and root up Israel out of this good land that he gave to their fathers and scatter them beyond the Euphrates, because they have made their Asherim, provoking the LORD to anger.
1KGS|14|16|And he will give Israel up because of the sins of Jeroboam, which he sinned and made Israel to sin."
1KGS|14|17|Then Jeroboam's wife arose and departed and came to Tirzah. And as she came to the threshold of the house, the child died.
1KGS|14|18|And all Israel buried him and mourned for him, according to the word of the LORD, which he spoke by his servant Ahijah the prophet.
1KGS|14|19|Now the rest of the acts of Jeroboam, how he warred and how he reigned, behold, they are written in the Book of the Chronicles of the Kings of Israel.
1KGS|14|20|And the time that Jeroboam reigned was twenty-two years. And he slept with his fathers, and Nadab his son reigned in his place.
1KGS|14|21|Now Rehoboam the son of Solomon reigned in Judah. Rehoboam was forty-one years old when he began to reign, and he reigned seventeen years in Jerusalem, the city that the LORD had chosen out of all the tribes of Israel, to put his name there. His mother's name was Naamah the Ammonite.
1KGS|14|22|And Judah did what was evil in the sight of the LORD, and they provoked him to jealousy with their sins that they committed, more than all that their fathers had done.
1KGS|14|23|For they also built for themselves high places and pillars and Asherim on every high hill and under every green tree,
1KGS|14|24|and there were also male cult prostitutes in the land. They did according to all the abominations of the nations that the LORD drove out before the people of Israel.
1KGS|14|25|In the fifth year of King Rehoboam, Shishak king of Egypt came up against Jerusalem.
1KGS|14|26|He took away the treasures of the house of the LORD and the treasures of the king's house. He took away everything. He also took away all the shields of gold that Solomon had made,
1KGS|14|27|and King Rehoboam made in their place shields of bronze, and committed them to the hands of the officers of the guard, who kept the door of the king's house.
1KGS|14|28|And as often as the king went into the house of the LORD, the guard carried them and brought them back to the guardroom.
1KGS|14|29|Now the rest of the acts of Rehoboam and all that he did, are they not written in the Book of the Chronicles of the Kings of Judah?
1KGS|14|30|And there was war between Rehoboam and Jeroboam continually.
1KGS|14|31|And Rehoboam slept with his fathers and was buried with his fathers in the city of David. His mother's name was Naamah the Ammonite. And Abijam his son reigned in his place.
1KGS|15|1|Now in the eighteenth year of King Jeroboam the son of Nebat, Abijam began to reign over Judah.
1KGS|15|2|He reigned for three years in Jerusalem. His mother's name was Maacah the daughter of Abishalom.
1KGS|15|3|And he walked in all the sins that his father did before him, and his heart was not wholly true to the LORD his God, as the heart of David his father.
1KGS|15|4|Nevertheless, for David's sake the LORD his God gave him a lamp in Jerusalem, setting up his son after him, and establishing Jerusalem,
1KGS|15|5|because David did what was right in the eyes of the LORD and did not turn aside from anything that he commanded him all the days of his life, except in the matter of Uriah the Hittite.
1KGS|15|6|Now there was war between Rehoboam and Jeroboam all the days of his life.
1KGS|15|7|The rest of the acts of Abijam and all that he did, are they not written in the Book of the Chronicles of the Kings of Judah? And there was war between Abijam and Jeroboam.
1KGS|15|8|And Abijam slept with his fathers, and they buried him in the city of David. And Asa his son reigned in his place.
1KGS|15|9|In the twentieth year of Jeroboam king of Israel, Asa began to reign over Judah,
1KGS|15|10|and he reigned forty-one years in Jerusalem. His mother's name was Maacah the daughter of Abishalom.
1KGS|15|11|And Asa did what was right in the eyes of the LORD, as David his father had done.
1KGS|15|12|He put away the male cult prostitutes out of the land and removed all the idols that his fathers had made.
1KGS|15|13|He also removed Maacah his mother from being queen mother because she had made an abominable image for Asherah. And Asa cut down her image and burned it at the brook Kidron.
1KGS|15|14|But the high places were not taken away. Nevertheless, the heart of Asa was wholly true to the LORD all his days.
1KGS|15|15|And he brought into the house of the LORD the sacred gifts of his father and his own sacred gifts, silver, and gold, and vessels.
1KGS|15|16|And there was war between Asa and Baasha king of Israel all their days.
1KGS|15|17|Baasha king of Israel went up against Judah and built Ramah, that he might permit no one to go out or come in to Asa king of Judah.
1KGS|15|18|Then Asa took all the silver and the gold that were left in the treasures of the house of the LORD and the treasures of the king's house and gave them into the hands of his servants. And King Asa sent them to Ben-hadad the son of Tabrimmon, the son of Hezion, king of Syria, who lived in Damascus, saying,
1KGS|15|19|"Let there be a covenant between me and you, as there was between my father and your father. Behold, I am sending to you a present of silver and gold. Go, break your covenant with Baasha king of Israel, that he may withdraw from me."
1KGS|15|20|And Ben-hadad listened to King Asa and sent the commanders of his armies against the cities of Israel and conquered Ijon, Dan, Abel-beth-maacah, and all Chinneroth, with all the land of Naphtali.
1KGS|15|21|And when Baasha heard of it, he stopped building Ramah, and he lived in Tirzah.
1KGS|15|22|Then King Asa made a proclamation to all Judah, none was exempt, and they carried away the stones of Ramah and its timber, with which Baasha had been building, and with them King Asa built Geba of Benjamin and Mizpah.
1KGS|15|23|Now the rest of all the acts of Asa, all his might, and all that he did, and the cities that he built, are they not written in the Book of the Chronicles of the Kings of Judah? But in his old age he was diseased in his feet.
1KGS|15|24|And Asa slept with his fathers and was buried with his fathers in the city of David his father, and Jehoshaphat his son reigned in his place.
1KGS|15|25|Nadab the son of Jeroboam began to reign over Israel in the second year of Asa king of Judah, and he reigned over Israel two years.
1KGS|15|26|He did what was evil in the sight of the LORD and walked in the way of his father, and in his sin which he made Israel to sin.
1KGS|15|27|Baasha the son of Ahijah, of the house of Issachar, conspired against him. And Baasha struck him down at Gibbethon, which belonged to the Philistines, for Nadab and all Israel were laying siege to Gibbethon.
1KGS|15|28|So Baasha killed him in the third year of Asa king of Judah and reigned in his place.
1KGS|15|29|And as soon as he was king, he killed all the house of Jeroboam. He left to the house of Jeroboam not one that breathed, until he had destroyed it, according to the word of the LORD that he spoke by his servant Ahijah the Shilonite.
1KGS|15|30|It was for the sins of Jeroboam that he sinned and that he made Israel to sin, and because of the anger to which he provoked the LORD, the God of Israel.
1KGS|15|31|Now the rest of the acts of Nadab and all that he did, are they not written in the Book of the Chronicles of the Kings of Israel?
1KGS|15|32|And there was war between Asa and Baasha king of Israel all their days.
1KGS|15|33|In the third year of Asa king of Judah, Baasha the son of Ahijah began to reign over all Israel at Tirzah, and he reigned twenty-four years.
1KGS|15|34|He did what was evil in the sight of the LORD and walked in the way of Jeroboam and in his sin which he made Israel to sin.
1KGS|16|1|And the word of the LORD came to Jehu the son of Hanani against Baasha, saying,
1KGS|16|2|"Since I exalted you out of the dust and made you leader over my people Israel, and you have walked in the way of Jeroboam and have made my people Israel to sin, provoking me to anger with their sins,
1KGS|16|3|behold, I will utterly sweep away Baasha and his house, and I will make your house like the house of Jeroboam the son of Nebat.
1KGS|16|4|Anyone belonging to Baasha who dies in the city the dogs shall eat, and anyone of his who dies in the field the birds of the heavens shall eat."
1KGS|16|5|Now the rest of the acts of Baasha and what he did, and his might, are they not written in the Book of the Chronicles of the Kings of Israel?
1KGS|16|6|And Baasha slept with his fathers and was buried at Tirzah, and Elah his son reigned in his place.
1KGS|16|7|Moreover, the word of the LORD came by the prophet Jehu the son of Hanani against Baasha and his house, both because of all the evil that he did in the sight of the LORD, provoking him to anger with the work of his hands, in being like the house of Jeroboam, and also because he destroyed it.
1KGS|16|8|In the twenty-sixth year of Asa king of Judah, Elah the son of Baasha began to reign over Israel in Tirzah, and he reigned two years.
1KGS|16|9|But his servant Zimri, commander of half his chariots, conspired against him. When he was at Tirzah, drinking himself drunk in the house of Arza, who was over the household in Tirzah,
1KGS|16|10|Zimri came in and struck him down and killed him, in the twenty-seventh year of Asa king of Judah, and reigned in his place.
1KGS|16|11|When he began to reign, as soon as he had seated himself on his throne, he struck down all the house of Baasha. He did not leave him a single male of his relatives or his friends.
1KGS|16|12|Thus Zimri destroyed all the house of Baasha, according to the word of the LORD, which he spoke against Baasha by Jehu the prophet,
1KGS|16|13|for all the sins of Baasha and the sins of Elah his son, which they sinned and which they made Israel to sin, provoking the LORD God of Israel to anger with their idols.
1KGS|16|14|Now the rest of the acts of Elah and all that he did, are they not written in the Book of the Chronicles of the Kings of Israel?
1KGS|16|15|In the twenty-seventh year of Asa king of Judah, Zimri reigned seven days in Tirzah. Now the troops were encamped against Gibbethon, which belonged to the Philistines,
1KGS|16|16|and the troops who were encamped heard it said, "Zimri has conspired, and he has killed the king." Therefore all Israel made Omri, the commander of the army, king over Israel that day in the camp.
1KGS|16|17|So Omri went up from Gibbethon, and all Israel with him, and they besieged Tirzah.
1KGS|16|18|And when Zimri saw that the city was taken, he went into the citadel of the king's house and burned the king's house over him with fire and died,
1KGS|16|19|because of his sins that he committed, doing evil in the sight of the LORD, walking in the way of Jeroboam, and for his sin which he committed, making Israel to sin.
1KGS|16|20|Now the rest of the acts of Zimri, and the conspiracy that he made, are they not written in the Book of the Chronicles of the Kings of Israel?
1KGS|16|21|Then the people of Israel were divided into two parts. Half of the people followed Tibni the son of Ginath, to make him king, and half followed Omri.
1KGS|16|22|But the people who followed Omri overcame the people who followed Tibni the son of Ginath. So Tibni died, and Omri became king.
1KGS|16|23|In the thirty-first year of Asa king of Judah, Omri began to reign over Israel, and he reigned for twelve years; six years he reigned in Tirzah.
1KGS|16|24|He bought the hill of Samaria from Shemer for two talents of silver, and he fortified the hill and called the name of the city that he built Samaria, after the name of Shemer, the owner of the hill.
1KGS|16|25|Omri did what was evil in the sight of the LORD, and did more evil than all who were before him.
1KGS|16|26|For he walked in all the way of Jeroboam the son of Nebat, and in the sins that he made Israel to sin, provoking the LORD, the God of Israel, to anger by their idols.
1KGS|16|27|Now the rest of the acts of Omri that he did, and the might that he showed, are they not written in the Book of the Chronicles of the Kings of Israel?
1KGS|16|28|And Omri slept with his fathers and was buried in Samaria, and Ahab his son reigned in his place.
1KGS|16|29|In the thirty-eighth year of Asa king of Judah, Ahab the son of Omri began to reign over Israel, and Ahab the son of Omri reigned over Israel in Samaria twenty-two years.
1KGS|16|30|And Ahab the son of Omri did evil in the sight of the LORD, more than all who were before him.
1KGS|16|31|And as if it had been a light thing for him to walk in the sins of Jeroboam the son of Nebat, he took for his wife Jezebel the daughter of Ethbaal king of the Sidonians, and went and served Baal and worshiped him.
1KGS|16|32|He erected an altar for Baal in the house of Baal, which he built in Samaria.
1KGS|16|33|And Ahab made an Asherah. Ahab did more to provoke the LORD, the God of Israel, to anger than all the kings of Israel who were before him.
1KGS|16|34|In his days Hiel of Bethel built Jericho. He laid its foundation at the cost of Abiram his firstborn, and set up its gates at the cost of his youngest son Segub, according to the word of the LORD, which he spoke by Joshua the son of Nun.
1KGS|17|1|Now Elijah the Tishbite, of Tishbe in Gilead, said to Ahab, "As the LORD the God of Israel lives, before whom I stand, there shall be neither dew nor rain these years, except by my word."
1KGS|17|2|And the word of the LORD came to him,
1KGS|17|3|"Depart from here and turn eastward and hide yourself by the brook Cherith, which is east of the Jordan.
1KGS|17|4|You shall drink from the brook, and I have commanded the ravens to feed you there."
1KGS|17|5|So he went and did according to the word of the LORD. He went and lived by the brook Cherith that is east of the Jordan.
1KGS|17|6|And the ravens brought him bread and meat in the morning, and bread and meat in the evening, and he drank from the brook.
1KGS|17|7|And after a while the brook dried up, because there was no rain in the land.
1KGS|17|8|Then the word of the LORD came to him,
1KGS|17|9|"Arise, go to Zarephath, which belongs to Sidon, and dwell there. Behold, I have commanded a widow there to feed you."
1KGS|17|10|So he arose and went to Zarephath. And when he came to the gate of the city, behold, a widow was there gathering sticks. And he called to her and said, "Bring me a little water in a vessel, that I may drink."
1KGS|17|11|And as she was going to bring it, he called to her and said, "Bring me a morsel of bread in your hand."
1KGS|17|12|And she said, "As the LORD your God lives, I have nothing baked, only a handful of flour in a jar and a little oil in a jug. And now I am gathering a couple of sticks that I may go in and prepare it for myself and my son, that we may eat it and die."
1KGS|17|13|And Elijah said to her, "Do not fear; go and do as you have said. But first make me a little cake of it and bring it to me, and afterward make something for yourself and your son.
1KGS|17|14|For thus says the LORD the God of Israel, 'The jar of flour shall not be spent, and the jug of oil shall not be empty, until the day that the LORD sends rain upon the earth.'"
1KGS|17|15|And she went and did as Elijah said. And she and he and her household ate for many days.
1KGS|17|16|The jar of flour was not spent, neither did the jug of oil become empty, according to the word of the LORD that he spoke by Elijah.
1KGS|17|17|After this the son of the woman, the mistress of the house, became ill. And his illness was so severe that there was no breath left in him.
1KGS|17|18|And she said to Elijah, "What have you against me, O man of God? You have come to me to bring my sin to remembrance and to cause the death of my son!"
1KGS|17|19|And he said to her, "Give me your son." And he took him from her arms and carried him up into the upper chamber where he lodged, and laid him on his own bed.
1KGS|17|20|And he cried to the LORD, "O LORD my God, have you brought calamity even upon the widow with whom I sojourn, by killing her son?"
1KGS|17|21|Then he stretched himself upon the child three times and cried to the LORD, "O LORD my God, let this child's life come into him again."
1KGS|17|22|And the LORD listened to the voice of Elijah. And the life of the child came into him again, and he revived.
1KGS|17|23|And Elijah took the child and brought him down from the upper chamber into the house and delivered him to his mother. And Elijah said, "See, your son lives."
1KGS|17|24|And the woman said to Elijah, "Now I know that you are a man of God, and that the word of the LORD in your mouth is truth."
1KGS|18|1|After many days the word of the LORD came to Elijah, in the third year, saying, "Go, show yourself to Ahab, and I will send rain upon the earth."
1KGS|18|2|So Elijah went to show himself to Ahab. Now the famine was severe in Samaria.
1KGS|18|3|And Ahab called Obadiah, who was over the household. (Now Obadiah feared the LORD greatly,
1KGS|18|4|and when Jezebel cut off the prophets of the LORD, Obadiah took a hundred prophets and hid them by fifties in a cave and fed them with bread and water.)
1KGS|18|5|And Ahab said to Obadiah, "Go through the land to all the springs of water and to all the valleys. Perhaps we may find grass and save the horses and mules alive, and not lose some of the animals."
1KGS|18|6|So they divided the land between them to pass through it. Ahab went in one direction by himself, and Obadiah went in another direction by himself.
1KGS|18|7|And as Obadiah was on the way, behold, Elijah met him. And Obadiah recognized him and fell on his face and said, "Is it you, my lord Elijah?"
1KGS|18|8|And he answered him, "It is I. Go, tell your lord, 'Behold, Elijah is here.'"
1KGS|18|9|And he said, "How have I sinned, that you would give your servant into the hand of Ahab, to kill me?
1KGS|18|10|As the LORD your God lives, there is no nation or kingdom where my lord has not sent to seek you. And when they would say, 'He is not here,' he would take an oath of the kingdom or nation, that they had not found you.
1KGS|18|11|And now you say, 'Go, tell your lord, "Behold, Elijah is here."'
1KGS|18|12|And as soon as I have gone from you, the Spirit of the LORD will carry you I know not where. And so, when I come and tell Ahab and he cannot find you, he will kill me, although I your servant have feared the LORD from my youth.
1KGS|18|13|Has it not been told my lord what I did when Jezebel killed the prophets of the LORD, how I hid a hundred men of the LORD's prophets by fifties in a cave and fed them with bread and water?
1KGS|18|14|And now you say, 'Go, tell your lord, "Behold, Elijah is here"'; and he will kill me."
1KGS|18|15|And Elijah said, "As the LORD of hosts lives, before whom I stand, I will surely show myself to him today."
1KGS|18|16|So Obadiah went to meet Ahab, and told him. And Ahab went to meet Elijah.
1KGS|18|17|When Ahab saw Elijah, Ahab said to him, "Is it you, you troubler of Israel?"
1KGS|18|18|And he answered, "I have not troubled Israel, but you have, and your father's house, because you have abandoned the commandments of the LORD and followed the Baals.
1KGS|18|19|Now therefore send and gather all Israel to me at Mount Carmel, and the 450 prophets of Baal and the 400 prophets of Asherah, who eat at Jezebel's table."
1KGS|18|20|So Ahab sent to all the people of Israel and gathered the prophets together at Mount Carmel.
1KGS|18|21|And Elijah came near to all the people and said, "How long will you go limping between two different opinions? If the LORD is God, follow him; but if Baal, then follow him." And the people did not answer him a word.
1KGS|18|22|Then Elijah said to the people, "I, even I only, am left a prophet of the LORD, but Baal's prophets are 450 men.
1KGS|18|23|Let two bulls be given to us, and let them choose one bull for themselves and cut it in pieces and lay it on the wood, but put no fire to it. And I will prepare the other bull and lay it on the wood and put no fire to it.
1KGS|18|24|And you call upon the name of your god, and I will call upon the name of the LORD, and the God who answers by fire, he is God." And all the people answered, "It is well spoken."
1KGS|18|25|Then Elijah said to the prophets of Baal, "Choose for yourselves one bull and prepare it first, for you are many, and call upon the name of your god, but put no fire to it."
1KGS|18|26|And they took the bull that was given them, and they prepared it and called upon the name of Baal from morning until noon, saying, "O Baal, answer us!" But there was no voice, and no one answered. And they limped around the altar that they had made.
1KGS|18|27|And at noon Elijah mocked them, saying, "Cry aloud, for he is a god. Either he is musing, or he is relieving himself, or he is on a journey, or perhaps he is asleep and must be awakened."
1KGS|18|28|And they cried aloud and cut themselves after their custom with swords and lances, until the blood gushed out upon them.
1KGS|18|29|And as midday passed, they raved on until the time of the offering of the oblation, but there was no voice. No one answered; no one paid attention.
1KGS|18|30|Then Elijah said to all the people, "Come near to me." And all the people came near to him. And he repaired the altar of the LORD that had been thrown down.
1KGS|18|31|Elijah took twelve stones, according to the number of the tribes of the sons of Jacob, to whom the word of the LORD came, saying, "Israel shall be your name,"
1KGS|18|32|and with the stones he built an altar in the name of the LORD. And he made a trench about the altar, as great as would contain two seahs of seed.
1KGS|18|33|And he put the wood in order and cut the bull in pieces and laid it on the wood. And he said, "Fill four jars with water and pour it on the burnt offering and on the wood."
1KGS|18|34|And he said, "Do it a second time." And they did it a second time. And he said, "Do it a third time." And they did it a third time.
1KGS|18|35|And the water ran around the altar and filled the trench also with water.
1KGS|18|36|And at the time of the offering of the oblation, Elijah the prophet came near and said, "O LORD, God of Abraham, Isaac, and Israel, let it be known this day that you are God in Israel, and that I am your servant, and that I have done all these things at your word.
1KGS|18|37|Answer me, O LORD, answer me, that this people may know that you, O LORD, are God, and that you have turned their hearts back."
1KGS|18|38|Then the fire of the LORD fell and consumed the burnt offering and the wood and the stones and the dust, and licked up the water that was in the trench.
1KGS|18|39|And when all the people saw it, they fell on their faces and said, "The LORD, he is God; the LORD, he is God."
1KGS|18|40|And Elijah said to them, "Seize the prophets of Baal; let not one of them escape." And they seized them. And Elijah brought them down to the brook Kishon and slaughtered them there.
1KGS|18|41|And Elijah said to Ahab, "Go up, eat and drink, for there is a sound of the rushing of rain."
1KGS|18|42|So Ahab went up to eat and to drink. And Elijah went up to the top of Mount Carmel. And he bowed himself down on the earth and put his face between his knees.
1KGS|18|43|And he said to his servant, "Go up now, look toward the sea." And he went up and looked and said, "There is nothing." And he said, "Go again," seven times.
1KGS|18|44|And at the seventh time he said, "Behold, a little cloud like a man's hand is rising from the sea." And he said, "Go up, say to Ahab, 'Prepare your chariot and go down, lest the rain stop you.'"
1KGS|18|45|And in a little while the heavens grew black with clouds and wind, and there was a great rain. And Ahab rode and went to Jezreel.
1KGS|18|46|And the hand of the LORD was on Elijah, and he gathered up his garment and ran before Ahab to the entrance of Jezreel.
1KGS|19|1|Ahab told Jezebel all that Elijah had done, and how he had killed all the prophets with the sword.
1KGS|19|2|Then Jezebel sent a messenger to Elijah, saying, "So may the gods do to me and more also, if I do not make your life as the life of one of them by this time tomorrow."
1KGS|19|3|Then he was afraid, and he arose and ran for his life and came to Beersheba, which belongs to Judah, and left his servant there.
1KGS|19|4|But he himself went a day's journey into the wilderness and came and sat down under a broom tree. And he asked that he might die, saying, "It is enough; now, O LORD, take away my life, for I am no better than my fathers."
1KGS|19|5|And he lay down and slept under a broom tree. And behold, an angel touched him and said to him, "Arise and eat."
1KGS|19|6|And he looked, and behold, there was at his head a cake baked on hot stones and a jar of water. And he ate and drank and lay down again.
1KGS|19|7|And the angel of the LORD came again a second time and touched him and said, "Arise and eat, for the journey is too great for you."
1KGS|19|8|And he arose and ate and drank, and went in the strength of that food forty days and forty nights to Horeb, the mount of God.
1KGS|19|9|There he came to a cave and lodged in it. And behold, the word of the LORD came to him, and he said to him, "What are you doing here, Elijah?"
1KGS|19|10|He said, "I have been very jealous for the LORD, the God of hosts. For the people of Israel have forsaken your covenant, thrown down your altars, and killed your prophets with the sword, and I, even I only, am left, and they seek my life, to take it away."
1KGS|19|11|And he said, "Go out and stand on the mount before the LORD." And behold, the LORD passed by, and a great and strong wind tore the mountains and broke in pieces the rocks before the LORD, but the LORD was not in the wind. And after the wind an earthquake, but the LORD was not in the earthquake.
1KGS|19|12|And after the earthquake a fire, but the LORD was not in the fire. And after the fire the sound of a low whisper.
1KGS|19|13|And when Elijah heard it, he wrapped his face in his cloak and went out and stood at the entrance of the cave. And behold, there came a voice to him and said, "What are you doing here, Elijah?"
1KGS|19|14|He said, "I have been very jealous for the LORD, the God of hosts. For the people of Israel have forsaken your covenant, thrown down your altars, and killed your prophets with the sword, and I, even I only, am left, and they seek my life, to take it away."
1KGS|19|15|And the LORD said to him, "Go, return on your way to the wilderness of Damascus. And when you arrive, you shall anoint Hazael to be king over Syria.
1KGS|19|16|And Jehu the son of Nimshi you shall anoint to be king over Israel, and Elisha the son of Shaphat of Abel-meholah you shall anoint to be prophet in your place.
1KGS|19|17|And the one who escapes from the sword of Hazael shall Jehu put to death, and the one who escapes from the sword of Jehu shall Elisha put to death.
1KGS|19|18|Yet I will leave seven thousand in Israel, all the knees that have not bowed to Baal, and every mouth that has not kissed him."
1KGS|19|19|So he departed from there and found Elisha the son of Shaphat, who was plowing with twelve yoke of oxen in front of him, and he was with the twelfth. Elijah passed by him and cast his cloak upon him.
1KGS|19|20|And he left the oxen and ran after Elijah and said, "Let me kiss my father and my mother, and then I will follow you." And he said to him, "Go back again, for what have I done to you?"
1KGS|19|21|And he returned from following him and took the yoke of oxen and sacrificed them and boiled their flesh with the yokes of the oxen and gave it to the people, and they ate. Then he arose and went after Elijah and assisted him.
1KGS|20|1|Ben-hadad the king of Syria gathered all his army together. Thirty-two kings were with him, and horses and chariots. And he went up and closed in on Samaria and fought against it.
1KGS|20|2|And he sent messengers into the city to Ahab king of Israel and said to him, "Thus says Ben-hadad:
1KGS|20|3|'Your silver and your gold are mine; your best wives and children also are mine.'"
1KGS|20|4|And the king of Israel answered, "As you say, my lord, O king, I am yours, and all that I have."
1KGS|20|5|The messengers came again and said, "Thus says Ben-hadad: 'I sent to you, saying, "Deliver to me your silver and your gold, your wives and your children."
1KGS|20|6|Nevertheless I will send my servants to you tomorrow about this time, and they shall search your house and the houses of your servants and lay hands on whatever pleases you and take it away.'"
1KGS|20|7|Then the king of Israel called all the elders of the land and said, "Mark, now, and see how this man is seeking trouble, for he sent to me for my wives and my children, and for my silver and my gold, and I did not refuse him."
1KGS|20|8|And all the elders and all the people said to him, "Do not listen or consent."
1KGS|20|9|So he said to the messengers of Ben-hadad, "Tell my lord the king, 'All that you first demanded of your servant I will do, but this thing I cannot do.'"And the messengers departed and brought him word again.
1KGS|20|10|Ben-hadad sent to him and said, "The gods do so to me and more also, if the dust of Samaria shall suffice for handfuls for all the people who follow me."
1KGS|20|11|And the king of Israel answered, "Tell him, 'Let not him who straps on his armor boast himself like he who takes it off.'"
1KGS|20|12|When Ben-hadad heard this message as he was drinking with the kings in the booths, he said to his men, "Take your positions." And they took their positions against the city.
1KGS|20|13|And behold, a prophet came near to Ahab king of Israel and said, "Thus says the LORD, Have you seen all this great multitude? Behold, I will give it into your hand this day, and you shall know that I am the LORD."
1KGS|20|14|And Ahab said, "By whom?" He said, "Thus says the LORD, By the servants of the governors of the districts." Then he said, "Who shall begin the battle?" He answered, "You."
1KGS|20|15|Then he mustered the servants of the governors of the districts, and they were 232. And after them he mustered all the people of Israel, seven thousand.
1KGS|20|16|And they went out at noon, while Ben-hadad was drinking himself drunk in the booths, he and the thirty-two kings who helped him.
1KGS|20|17|The servants of the governors of the districts went out first. And Ben-hadad sent out scouts, and they reported to him, "Men are coming out from Samaria."
1KGS|20|18|He said, "If they have come out for peace, take them alive. Or if they have come out for war, take them alive."
1KGS|20|19|So these went out of the city, the servants of the governors of the districts and the army that followed them.
1KGS|20|20|And each struck down his man. The Syrians fled, and Israel pursued them, but Ben-hadad king of Syria escaped on a horse with horsemen.
1KGS|20|21|And the king of Israel went out and struck the horses and chariots, and struck the Syrians with a great blow.
1KGS|20|22|Then the prophet came near to the king of Israel and said to him, "Come, strengthen yourself, and consider well what you have to do, for in the spring the king of Syria will come up against you."
1KGS|20|23|And the servants of the king of Syria said to him, "Their gods are gods of the hills, and so they were stronger than we. But let us fight against them in the plain, and surely we shall be stronger than they.
1KGS|20|24|And do this: remove the kings, each from his post, and put commanders in their places,
1KGS|20|25|and muster an army like the army that you have lost, horse for horse, and chariot for chariot. Then we will fight against them in the plain, and surely we shall be stronger than they." And he listened to their voice and did so.
1KGS|20|26|In the spring, Ben-hadad mustered the Syrians and went up to Aphek to fight against Israel.
1KGS|20|27|And the people of Israel were mustered and were provisioned and went against them. The people of Israel encamped before them like two little flocks of goats, but the Syrians filled the country.
1KGS|20|28|And a man of God came near and said to the king of Israel, "Thus says the LORD, 'Because the Syrians have said, "The LORD is a god of the hills but he is not a god of the valleys," therefore I will give all this great multitude into your hand, and you shall know that I am the LORD.'"
1KGS|20|29|And they encamped opposite one another seven days. Then on the seventh day the battle was joined. And the people of Israel struck down of the Syrians 100,000 foot soldiers in one day.
1KGS|20|30|And the rest fled into the city of Aphek, and the wall fell upon 27,000 men who were left. Ben-hadad also fled and entered an inner chamber in the city.
1KGS|20|31|And his servants said to him, "Behold now, we have heard that the kings of the house of Israel are merciful kings. Let us put sackcloth around our waists and ropes on our heads and go out to the king of Israel. Perhaps he will spare your life."
1KGS|20|32|So they tied sackcloth around their waists and put ropes on their heads and went to the king of Israel and said, "Your servant Ben-hadad says, 'Please, let me live.'"And he said, "Does he still live? He is my brother."
1KGS|20|33|Now the men were watching for a sign, and they quickly took it up from him and said, "Yes, your brother Ben-hadad." Then he said, "Go and bring him." Then Ben-hadad came out to him, and he caused him to come up into the chariot.
1KGS|20|34|And Ben-hadad said to him, "The cities that my father took from your father I will restore, and you may establish bazaars for yourself in Damascus, as my father did in Samaria." And Ahab said, "I will let you go on these terms." So he made a covenant with him and let him go.
1KGS|20|35|And a certain man of the sons of the prophets said to his fellow at the command of the LORD, "Strike me, please." But the man refused to strike him.
1KGS|20|36|Then he said to him, "Because you have not obeyed the voice of the LORD, behold, as soon as you have gone from me, a lion shall strike you down." And as soon as he had departed from him, a lion met him and struck him down.
1KGS|20|37|Then he found another man and said, "Strike me, please." And the man struck him- struck him and wounded him.
1KGS|20|38|So the prophet departed and waited for the king by the way, disguising himself with a bandage over his eyes.
1KGS|20|39|And as the king passed, he cried to the king and said, "Your servant went out into the midst of the battle, and behold, a soldier turned and brought a man to me and said, 'Guard this man; if by any means he is missing, your life shall be for his life, or else you shall pay a talent of silver.'
1KGS|20|40|And as your servant was busy here and there, he was gone." The king of Israel said to him, "So shall your judgment be; you yourself have decided it."
1KGS|20|41|Then he hurried to take the bandage away from his eyes, and the king of Israel recognized him as one of the prophets.
1KGS|20|42|And he said to him, "Thus says the LORD, 'Because you have let go out of your hand the man whom I had devoted to destruction, therefore your life shall be for his life, and your people for his people.'"
1KGS|20|43|And the king of Israel went to his house vexed and sullen and came to Samaria.
1KGS|21|1|Now Naboth the Jezreelite had a vineyard in Jezreel, beside the palace of Ahab king of Samaria.
1KGS|21|2|And after this Ahab said to Naboth, "Give me your vineyard, that I may have it for a vegetable garden, because it is near my house, and I will give you a better vineyard for it; or, if it seems good to you, I will give you its value in money."
1KGS|21|3|But Naboth said to Ahab, "The LORD forbid that I should give you the inheritance of my fathers."
1KGS|21|4|And Ahab went into his house vexed and sullen because of what Naboth the Jezreelite had said to him, for he had said, "I will not give you the inheritance of my fathers." And he lay down on his bed and turned away his face and would eat no food.
1KGS|21|5|But Jezebel his wife came to him and said to him, "Why is your spirit so vexed that you eat no food?"
1KGS|21|6|And he said to her, "Because I spoke to Naboth the Jezreelite and said to him, 'Give me your vineyard for money, or else, if it please you, I will give you another vineyard for it.' And he answered, 'I will not give you my vineyard.'"
1KGS|21|7|And Jezebel his wife said to him, "Do you now govern Israel? Arise and eat bread and let your heart be cheerful; I will give you the vineyard of Naboth the Jezreelite."
1KGS|21|8|So she wrote letters in Ahab's name and sealed them with his seal, and she sent the letters to the elders and the leaders who lived with Naboth in his city.
1KGS|21|9|And she wrote in the letters, "Proclaim a fast, and set Naboth at the head of the people.
1KGS|21|10|And set two worthless men opposite him, and let them bring a charge against him, saying, 'You have cursed God and the king.' Then take him out and stone him to death."
1KGS|21|11|And the men of his city, the elders and the leaders who lived in his city, did as Jezebel had sent word to them. As it was written in the letters that she had sent to them,
1KGS|21|12|they proclaimed a fast and set Naboth at the head of the people.
1KGS|21|13|And the two worthless men came in and sat opposite him. And the worthless men brought a charge against Naboth in the presence of the people, saying, "Naboth cursed God and the king." So they took him outside the city and stoned him to death with stones.
1KGS|21|14|Then they sent to Jezebel, saying, "Naboth has been stoned; he is dead."
1KGS|21|15|As soon as Jezebel heard that Naboth had been stoned and was dead, Jezebel said to Ahab, "Arise, take possession of the vineyard of Naboth the Jezreelite, which he refused to give you for money, for Naboth is not alive, but dead."
1KGS|21|16|And as soon as Ahab heard that Naboth was dead, Ahab arose to go down to the vineyard of Naboth the Jezreelite, to take possession of it.
1KGS|21|17|Then the word of the LORD came to Elijah the Tishbite, saying,
1KGS|21|18|"Arise, go down to meet Ahab king of Israel, who is in Samaria; behold, he is in the vineyard of Naboth, where he has gone to take possession.
1KGS|21|19|And you shall say to him, 'Thus says the LORD, "Have you killed and also taken possession?"'And you shall say to him, 'Thus says the LORD: "In the place where dogs licked up the blood of Naboth shall dogs lick your own blood."'"
1KGS|21|20|Ahab said to Elijah, "Have you found me, O my enemy?" He answered, "I have found you, because you have sold yourself to do what is evil in the sight of the LORD.
1KGS|21|21|Behold, I will bring disaster upon you. I will utterly burn you up, and will cut off from Ahab every male, bond or free, in Israel.
1KGS|21|22|And I will make your house like the house of Jeroboam the son of Nebat, and like the house of Baasha the son of Ahijah, for the anger to which you have provoked me, and because you have made Israel to sin.
1KGS|21|23|And of Jezebel the LORD also said, 'The dogs shall eat Jezebel within the walls of Jezreel.'
1KGS|21|24|Anyone belonging to Ahab who dies in the city the dogs shall eat, and anyone of his who dies in the open country the birds of the heavens shall eat."
1KGS|21|25|(There was none who sold himself to do what was evil in the sight of the LORD like Ahab, whom Jezebel his wife incited.
1KGS|21|26|He acted very abominably in going after idols, as the Amorites had done, whom the LORD cast out before the people of Israel.)
1KGS|21|27|And when Ahab heard those words, he tore his clothes and put sackcloth on his flesh and fasted and lay in sackcloth and went about dejectedly.
1KGS|21|28|And the word of the LORD came to Elijah the Tishbite, saying,
1KGS|21|29|"Have you seen how Ahab has humbled himself before me? Because he has humbled himself before me, I will not bring the disaster in his days; but in his son's days I will bring the disaster upon his house."
1KGS|22|1|For three years Syria and Israel continued without war.
1KGS|22|2|But in the third year Jehoshaphat the king of Judah came down to the king of Israel.
1KGS|22|3|And the king of Israel said to his servants, "Do you know that Ramoth-gilead belongs to us, and we keep quiet and do not take it out of the hand of the king of Syria?"
1KGS|22|4|And he said to Jehoshaphat, "Will you go with me to battle at Ramoth-gilead?" And Jehoshaphat said to the king of Israel, "I am as you are, my people as your people, my horses as your horses."
1KGS|22|5|And Jehoshaphat said to the king of Israel, "Inquire first for the word of the LORD."
1KGS|22|6|Then the king of Israel gathered the prophets together, about four hundred men, and said to them, "Shall I go to battle against Ramoth-gilead, or shall I refrain?" And they said, "Go up, for the Lord will give it into the hand of the king."
1KGS|22|7|But Jehoshaphat said, "Is there not here another prophet of the LORD of whom we may inquire?"
1KGS|22|8|And the king of Israel said to Jehoshaphat, "There is yet one man by whom we may inquire of the LORD, Micaiah the son of Imlah, but I hate him, for he never prophesies good concerning me, but evil." And Jehoshaphat said, "Let not the king say so."
1KGS|22|9|Then the king of Israel summoned an officer and said, "Bring quickly Micaiah the son of Imlah."
1KGS|22|10|Now the king of Israel and Jehoshaphat the king of Judah were sitting on their thrones, arrayed in their robes, at the threshing floor at the entrance of the gate of Samaria, and all the prophets were prophesying before them.
1KGS|22|11|And Zedekiah the son of Chenaanah made for himself horns of iron and said, "Thus says the LORD, 'With these you shall push the Syrians until they are destroyed.'"
1KGS|22|12|And all the prophets prophesied so and said, "Go up to Ramoth-gilead and triumph; the LORD will give it into the hand of the king."
1KGS|22|13|And the messenger who went to summon Micaiah said to him, "Behold, the words of the prophets with one accord are favorable to the king. Let your word be like the word of one of them, and speak favorably."
1KGS|22|14|But Micaiah said, "As the LORD lives, what the LORD says to me, that I will speak."
1KGS|22|15|And when he had come to the king, the king said to him, "Micaiah, shall we go to Ramoth-gilead to battle, or shall we refrain?" And he answered him, "Go up and triumph; the LORD will give it into the hand of the king."
1KGS|22|16|But the king said to him, "How many times shall I make you swear that you speak to me nothing but the truth in the name of the LORD?"
1KGS|22|17|And he said, "I saw all Israel scattered on the mountains, as sheep that have no shepherd. And the LORD said, 'These have no master; let each return to his home in peace.'"
1KGS|22|18|And the king of Israel said to Jehoshaphat, "Did I not tell you that he would not prophesy good concerning me, but evil?"
1KGS|22|19|And Micaiah said, "Therefore hear the word of the LORD: I saw the LORD sitting on his throne, and all the host of heaven standing beside him on his right hand and on his left;
1KGS|22|20|and the LORD said, 'Who will entice Ahab, that he may go up and fall at Ramoth-gilead?' And one said one thing, and another said another.
1KGS|22|21|Then a spirit came forward and stood before the LORD, saying, 'I will entice him.'
1KGS|22|22|And the LORD said to him, 'By what means?' And he said, 'I will go out, and will be a lying spirit in the mouth of all his prophets.' And he said, 'You are to entice him, and you shall succeed; go out and do so.'
1KGS|22|23|Now therefore behold, the LORD has put a lying spirit in the mouth of all these your prophets; the LORD has declared disaster for you."
1KGS|22|24|Then Zedekiah the son of Chenaanah came near and struck Micaiah on the cheek and said, "How did the Spirit of the LORD go from me to speak to you?"
1KGS|22|25|And Micaiah said, "Behold, you shall see on that day when you go into an inner chamber to hide yourself."
1KGS|22|26|And the king of Israel said, "Seize Micaiah, and take him back to Amon the governor of the city and to Joash the king's son,
1KGS|22|27|and say, 'Thus says the king, "Put this fellow in prison and feed him meager rations of bread and water, until I come in peace."'"
1KGS|22|28|And Micaiah said, "If you return in peace, the LORD has not spoken by me." And he said, "Hear, all you peoples!"
1KGS|22|29|So the king of Israel and Jehoshaphat the king of Judah went up to Ramoth-gilead.
1KGS|22|30|And the king of Israel said to Jehoshaphat, "I will disguise myself and go into battle, but you wear your robes." And the king of Israel disguised himself and went into battle.
1KGS|22|31|Now the king of Syria had commanded the thirty-two captains of his chariots, "Fight with neither small nor great, but only with the king of Israel."
1KGS|22|32|And when the captains of the chariots saw Jehoshaphat, they said, "It is surely the king of Israel." So they turned to fight against him. And Jehoshaphat cried out.
1KGS|22|33|And when the captains of the chariots saw that it was not the king of Israel, they turned back from pursuing him.
1KGS|22|34|But a certain man drew his bow at random and struck the king of Israel between the scale armor and the breastplate. Therefore he said to the driver of his chariot, "Turn around and carry me out of the battle, for I am wounded."
1KGS|22|35|And the battle continued that day, and the king was propped up in his chariot facing the Syrians, until at evening he died. And the blood of the wound flowed into the bottom of the chariot.
1KGS|22|36|And about sunset a cry went through the army, "Every man to his city, and every man to his country!"
1KGS|22|37|So the king died, and was brought to Samaria. And they buried the king in Samaria.
1KGS|22|38|And they washed the chariot by the pool of Samaria, and the dogs licked up his blood, and the prostitutes washed themselves in it, according to the word of the LORD that he had spoken.
1KGS|22|39|Now the rest of the acts of Ahab and all that he did, and the ivory house that he built and all the cities that he built, are they not written in the Book of the Chronicles of the Kings of Israel?
1KGS|22|40|So Ahab slept with his fathers, and Ahaziah his son reigned in his place.
1KGS|22|41|Jehoshaphat the son of Asa began to reign over Judah in the fourth year of Ahab king of Israel.
1KGS|22|42|Jehoshaphat was thirty-five years old when he began to reign, and he reigned twenty-five years in Jerusalem. His mother's name was Azubah the daughter of Shilhi.
1KGS|22|43|He walked in all the way of Asa his father. He did not turn aside from it, doing what was right in the sight of the LORD. Yet the high places were not taken away, and the people still sacrificed and made offerings on the high places.
1KGS|22|44|Jehoshaphat also made peace with the king of Israel.
1KGS|22|45|Now the rest of the acts of Jehoshaphat, and his might that he showed, and how he warred, are they not written in the Book of the Chronicles of the Kings of Judah?
1KGS|22|46|And from the land he exterminated the remnant of the male cult prostitutes who remained in the days of his father Asa.
1KGS|22|47|There was no king in Edom; a deputy was king.
1KGS|22|48|Jehoshaphat made ships of Tarshish to go to Ophir for gold, but they did not go, for the ships were wrecked at Ezion-geber.
1KGS|22|49|Then Ahaziah the son of Ahab said to Jehoshaphat, "Let my servants go with your servants in the ships," but Jehoshaphat was not willing.
1KGS|22|50|And Jehoshaphat slept with his fathers and was buried with his fathers in the city of David his father, and Jehoram his son reigned in his place.
1KGS|22|51|Ahaziah the son of Ahab began to reign over Israel in Samaria in the seventeenth year of Jehoshaphat king of Judah, and he reigned two years over Israel.
1KGS|22|52|He did what was evil in the sight of the LORD and walked in the way of his father and in the way of his mother and in the way of Jeroboam the son of Nebat, who made Israel to sin.
1KGS|22|53|He served Baal and worshiped him and provoked the LORD, the God of Israel, to anger in every way that his father had done.
