JUDE|1|1|Jude, a servant of Jesus Christ and brother of James, To those who are called, beloved in God the Father and kept for Jesus Christ:
JUDE|1|2|May mercy, peace, and love be multiplied to you.
JUDE|1|3|Beloved, although I was very eager to write to you about our common salvation, I found it necessary to write appealing to you to contend for the faith that was once for all delivered to the saints.
JUDE|1|4|For certain people have crept in unnoticed who long ago were designated for this condemnation, ungodly people, who pervert the grace of our God into sensuality and deny our only Master and Lord, Jesus Christ.
JUDE|1|5|Now I want to remind you, although you once fully knew it, that Jesus, who saved a people out of the land of Egypt, afterward destroyed those who did not believe.
JUDE|1|6|And the angels who did not stay within their own position of authority, but left their proper dwelling, he has kept in eternal chains under gloomy darkness until the judgment of the great day-
JUDE|1|7|just as Sodom and Gomorrah and the surrounding cities, which likewise indulged in sexual immorality and pursued unnatural desire, serve as an example by undergoing a punishment of eternal fire.
JUDE|1|8|Yet in like manner these people also, relying on their dreams, defile the flesh, reject authority, and blaspheme the glorious ones.
JUDE|1|9|But when the archangel Michael, contending with the devil, was disputing about the body of Moses, he did not presume to pronounce a blasphemous judgment, but said, "The Lord rebuke you."
JUDE|1|10|But these people blaspheme all that they do not understand, and they are destroyed by all that they, like unreasoning animals, understand instinctively.
JUDE|1|11|Woe to them! For they walked in the way of Cain and abandoned themselves for the sake of gain to Balaam's error and perished in Korah's rebellion.
JUDE|1|12|These are blemishes on your love feasts, as they feast with you without fear, looking after themselves; waterless clouds, swept along by winds; fruitless trees in late autumn, twice dead, uprooted;
JUDE|1|13|wild waves of the sea, casting up the foam of their own shame; wandering stars, for whom the gloom of utter darkness has been reserved forever.
JUDE|1|14|It was also about these that Enoch, the seventh from Adam, prophesied, saying, "Behold, the Lord came with ten thousands of his holy ones,
JUDE|1|15|to execute judgment on all and to convict all the ungodly of all their deeds of ungodliness that they have committed in such an ungodly way, and of all the harsh things that ungodly sinners have spoken against him."
JUDE|1|16|These are grumblers, malcontents, following their own sinful desires; they are loud-mouthed boasters, showing favoritism to gain advantage.
JUDE|1|17|But you must remember, beloved, the predictions of the apostles of our Lord Jesus Christ.
JUDE|1|18|They said to you, "In the last time there will be scoffers, following their own ungodly passions."
JUDE|1|19|It is these who cause divisions, worldly people, devoid of the Spirit.
JUDE|1|20|But you, beloved, build yourselves up in your most holy faith; pray in the Holy Spirit;
JUDE|1|21|keep yourselves in the love of God, waiting for the mercy of our Lord Jesus Christ that leads to eternal life.
JUDE|1|22|And have mercy on those who doubt;
JUDE|1|23|save others by snatching them out of the fire; to others show mercy with fear, hating even the garment stained by the flesh.
JUDE|1|24|Now to him who is able to keep you from stumbling and to present you blameless before the presence of his glory with great joy,
JUDE|1|25|to the only God, our Savior, through Jesus Christ our Lord, be glory, majesty, dominion, and authority, before all time and now and forever. Amen.
