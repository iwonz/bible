1PET|1|1|耶穌基督的使徒 彼得 寫信給那些被揀選，分散在 本都 、 加拉太 、 加帕多家 、 亞細亞 、 庇推尼 寄居的人，
1PET|1|2|就是照父上帝的預知，藉著聖靈得以成聖，以致順服耶穌基督，又蒙他血所灑的人。願恩惠、平安 多多地賜給你們！
1PET|1|3|願頌讚歸於我們主耶穌基督的父上帝！他曾照自己的大憐憫，藉著耶穌基督從死人中復活，重生了我們，使我們有活的盼望，
1PET|1|4|好得到不朽壞、不玷污、不衰殘、為你們存留在天上的基業，
1PET|1|5|就是為你們這些藉著信、蒙上帝大能保守的人，能獲得他所預備、到末世要顯現的救恩。
1PET|1|6|雖然你們必須在百般試煉中暫時憂愁，你們要為此喜樂 ，
1PET|1|7|使你們的信心既被考驗，就比那被火試煉仍然能壞的金子更顯寶貴，可以在耶穌基督顯現的時候得著稱讚、榮耀、尊貴。
1PET|1|8|雖然你們沒有見過他，卻是愛他；如今雖看不見，你們卻因信他而有說不出來、滿有榮光的喜樂，
1PET|1|9|因為你們 得到信心的效果，就是靈魂的得救。
1PET|1|10|論到這救恩，那預先說你們要得恩典的眾先知已經詳細地搜索查考過，
1PET|1|11|查考在他們心裏的基督的靈預先證明基督受苦難，後來得榮耀，是指甚麼時候，甚麼樣的情況。
1PET|1|12|他們得了啟示，知道他們所服事的不是自己，而是你們。那藉著從天上差來的聖靈傳福音給你們的人，現在將這些事傳給你們；這些事連天使也都切望察看呢！
1PET|1|13|所以，要準備 好你們的心，謹慎自守，專心盼望耶穌基督顯現的時候帶給你們的恩惠。
1PET|1|14|作為順服的兒女，就不要效法從前蒙昧無知的時候那放縱私慾的樣子。
1PET|1|15|但那召你們的既是聖潔，你們在一切所行的事上也要聖潔；
1PET|1|16|因為經上記著：「你們要成為聖，因為我是神聖的。」
1PET|1|17|既然你們稱那不偏待人、按各人行為審判人的主為父 ，就當存敬畏的心，度你們在世寄居的日子。
1PET|1|18|你們知道，你們得以從你們祖先傳下來虛妄的行為中救贖出來，不是靠著會朽壞的金銀等物，
1PET|1|19|而是憑著基督的寶血，如同無瑕疵、無玷污的羔羊的血。
1PET|1|20|基督是上帝在創世以前所預知，而在這末世才為你們顯現的。
1PET|1|21|你們也因著他而信那使他從死人中復活、又給他榮耀的上帝，好讓你們的信心和盼望都在於上帝。
1PET|1|22|既然你們因順從真理而潔淨了自己的心靈，能真誠愛弟兄，就該以清潔的心 彼此切實相愛。
1PET|1|23|你們蒙了重生，不是由於會朽壞的種子，而是由於不會朽壞的種子，是藉著上帝永活常存的道。
1PET|1|24|因為 「凡血肉之軀的盡都如草， 他的一切榮美像草上的花； 草必枯乾，花必凋謝，
1PET|1|25|惟有主的道永遠常存。」 這話就是傳給你們的福音。
1PET|2|1|所以，你們要除去一切的惡毒，一切詭詐、假善、嫉妒，和一切毀謗的話。
1PET|2|2|要愛慕那純淨的靈奶，像初生的嬰孩愛慕奶一樣，好使你們藉著它成長，以致得救，
1PET|2|3|因為你們已經嘗過主恩的滋味。
1PET|2|4|要親近主，他是活石，雖然被人所丟棄，卻是上帝所揀選、所珍貴的。
1PET|2|5|你們作為活石，要被建造成屬靈的殿，成為聖潔的祭司，藉著耶穌基督獻上蒙上帝悅納的屬靈祭物。
1PET|2|6|因為經上說： 「看哪，我把一塊石頭放在 錫安 — 一塊蒙揀選、珍貴的房角石； 信靠他的人必不蒙羞。」
1PET|2|7|所以，這石頭在你們信的人是珍貴的；在那不信的人卻有話說： 「匠人所丟棄的石頭 已作了房角的頭塊石頭。」
1PET|2|8|又說： 「作了絆腳的石頭， 使人跌倒的磐石。」 他們絆跌，因為不順從這道，這也是預定的。
1PET|2|9|不過，你們是被揀選的一族，是君尊的祭司，是神聖的國度，是屬上帝的子民，要使你們宣揚那召你們出黑暗入奇妙光明者的美德。
1PET|2|10|「你們從前不是子民， 現在卻成了上帝的子民； 從前未曾蒙憐憫， 現在卻蒙了憐憫。」
1PET|2|11|親愛的，你們是客旅，是寄居的，我勸你們要禁戒肉體的情慾；這情慾是與靈魂爭戰的。
1PET|2|12|你們在外邦人中要品行端正，好讓那些人，雖然毀謗你們是作惡的，會因看見你們的好行為而在鑒察 的日子歸榮耀給上帝。
1PET|2|13|你們為主的緣故要順服人的一切制度，或是在上的君王，
1PET|2|14|或是君王所派懲惡賞善的官員。
1PET|2|15|因為上帝的旨意原是要你們以行善來堵住糊塗無知人的口。
1PET|2|16|雖然你們是自由的，卻不可藉著自由遮蓋惡毒，總要作上帝的僕人。
1PET|2|17|務要尊重眾人；要敬愛教中的弟兄姊妹；要敬畏上帝；要尊敬君王。
1PET|2|18|你們作奴僕的，凡事要存敬畏的心順服主人；不但順服善良溫和的，就是乖僻的也要順服。
1PET|2|19|倘若你們為使良心對得起上帝，忍受冤屈的痛苦，這是可讚許的。
1PET|2|20|你們若因犯罪受責打而忍耐，有甚麼可稱讚的呢？但你們若因行善受苦而忍耐，這在上帝看來是可讚許的。
1PET|2|21|你們蒙召就是為此，因為基督也為你們受過苦，給你們留下榜樣，為要使你們跟隨他的腳蹤。
1PET|2|22|「他並沒有犯罪， 口裏也沒有詭詐。」
1PET|2|23|他被辱罵不還口，受害也不說威嚇的話，只將自己交託給公義的審判者。
1PET|2|24|他被掛在木頭上，親身擔當了我們的罪，使我們既然在罪上死，就得以在義上活。因他受的鞭傷，你們得了醫治。
1PET|2|25|你們從前好像迷路的羊，如今卻歸回你們靈魂的牧人和監督了。
1PET|3|1|同樣，你們作妻子的，要順服自己的丈夫，這樣，即使有不信從道理的丈夫，也會因妻子的品行，並非言語，而感化過來，
1PET|3|2|因為看見了你們敬虔純潔的品行。
1PET|3|3|你們不要藉外表來妝飾自己，如編頭髮，戴金飾，穿美麗的衣裳等，
1PET|3|4|而要有蘊藏在人內心不衰退的美，以溫柔嫻靜的心妝飾自己；這在上帝面前是極寶貴的。
1PET|3|5|因為古時仰賴上帝的聖潔婦人正是以此為妝飾，順服自己的丈夫。
1PET|3|6|就如 撒拉 聽從 亞伯拉罕 ，稱他為主。你們只要行善，不怕任何恐嚇，就成為 撒拉 的女兒了。
1PET|3|7|同樣，你們作丈夫的，要按情理 跟妻子共同生活，體貼女性是比較軟弱的器皿；要尊重她，因為她也與你一同承受生命之恩。這樣，你們的禱告就不會受阻礙。
1PET|3|8|總而言之，你們都要同心，彼此體恤，相愛如弟兄，存憐憫和謙卑的心。
1PET|3|9|不要以惡報惡，以辱罵還辱罵，倒要祝福，因為你們正是為此蒙召的，好使你們承受福氣。
1PET|3|10|因為經上說： 「凡要愛惜生命、 享受好日子的人， 要禁止舌頭不出惡言， 嘴唇不說詭詐的話。
1PET|3|11|也要棄惡行善， 尋求和睦，一心追求。
1PET|3|12|因為主的眼看顧義人， 他的耳聽他們的祈禱； 但主向行惡的人變臉。」
1PET|3|13|你們若熱心行善，有誰會害你們呢？
1PET|3|14|即使你們為義受苦，也是有福的。不要怕人的威嚇，也不要驚慌；
1PET|3|15|只要心裏奉主基督為聖，尊他為主。有人問你們心中盼望的理由，要隨時準備答覆；
1PET|3|16|不過，要以溫柔、敬畏的心回答。要存無虧的良心，使你們在何事上被毀謗，就在何事上使那些凌辱你們在基督裏有好品行的人自覺羞愧。
1PET|3|17|上帝的旨意若是要你們因行善受苦，這總比因行惡受苦好。
1PET|3|18|因為基督也曾一次為罪受苦 ， 就是義的代替不義的， 為要引領你們 到上帝面前。 在肉體裏，他被治死； 但在靈裏，他復活了。
1PET|3|19|他藉這靈也曾去向那些在監獄裏的靈傳道，
1PET|3|20|就是那些從前在 挪亞 預備方舟、上帝容忍等待的時候不信從的人。當時進入方舟，藉著水得救的不多，只有八個人。
1PET|3|21|這水所預表的洗禮，現在藉著耶穌基督的復活拯救你們，不是除掉肉體的污穢，而是向上帝懇求有無虧的良心。
1PET|3|22|耶穌已經到天上去，在上帝的右邊，眾天使、有權柄的、有權能的都服從了他。
1PET|4|1|既然基督在肉身受苦，你們也該將這樣的心志作為兵器，因為在肉身受過苦的已經與罪斷絕了，
1PET|4|2|使你們從今以後不再隨從人的情慾，只順從上帝的旨意，在世度餘下的光陰。
1PET|4|3|因為你們從前隨從外邦人的心意，生活在淫蕩、情慾、醉酒、荒宴、狂飲和可憎的偶像崇拜中，時候已經夠了。
1PET|4|4|在這些事上，他們見你們不與他們同奔放蕩無度的路就以為怪，毀謗你們。
1PET|4|5|他們必須在那位將要審判活人死人的主面前交賬。
1PET|4|6|為此，死人也曾有福音傳給他們，要使他們的肉體按著人受審判，他們的靈卻靠上帝活著。
1PET|4|7|萬物的結局近了。所以你們要謹慎自守，要警醒禱告。
1PET|4|8|最要緊的是彼此切實相愛，因為愛能遮掩許多的罪。
1PET|4|9|你們要互相款待，不發怨言。
1PET|4|10|人人要照自己所得的恩賜彼此服事，作上帝各種恩賜的好管家。
1PET|4|11|若有人講道，他要按著上帝的聖言講；若有人服事，他要按著上帝所賜的力量服事，好讓上帝在凡事上因耶穌基督得榮耀。願榮耀和權能都歸給他，直到永永遠遠。阿們！
1PET|4|12|親愛的，有火一般的考驗臨到你們，不要奇怪，似乎是遭遇非常的事；
1PET|4|13|倒要歡喜，因為你們是與基督一同受苦，使你們在他榮耀顯現的時候也可以歡喜快樂。
1PET|4|14|你們若為基督的名受辱罵是有福的，因為榮耀的靈，就是上帝的靈，在你們身上。
1PET|4|15|你們中間，不可有人因為殺人、偷竊、作惡、好管閒事而受苦。
1PET|4|16|若有人因是基督徒而受苦，不要引以為恥，倒要因這名而歸榮耀給上帝。
1PET|4|17|因為時候到了，審判要從上帝的家開始；若是先從我們開始，那麼，不信從上帝福音的人將有何等的結局呢？
1PET|4|18|「若是義人還僅僅得救， 不虔敬和犯罪的人將有何地可站呢？」
1PET|4|19|所以，照上帝旨意受苦的人要一心為善，將自己的靈魂交給那信實的造物主。
1PET|5|1|所以，我這同作長老，作基督受苦的證人和分享將來所要顯現的榮耀的人，勉勵在你們中間的長老們：
1PET|5|2|務要牧養在你們當中上帝的群羊，按著上帝的旨意照顧他們 ，不是出於勉強，而是出於甘心；也不是因為貪財，而是出於樂意。
1PET|5|3|不要轄制所託付你們的群羊，而是要作他們的榜樣。
1PET|5|4|到了大牧人顯現的時候，你們必得到那永不衰殘、榮耀的冠冕。
1PET|5|5|同樣，你們年輕的，要順服年長的。你們大家都要以謙卑當衣服穿上，彼此順服，因為 「上帝抵擋驕傲的人， 但賜恩給謙卑的人。」
1PET|5|6|所以，你們要謙卑服在上帝大能的手下，這樣，到了適當的時候，他必使你們升高。
1PET|5|7|你們要將一切的憂慮卸給上帝，因為他顧念你們。
1PET|5|8|務要謹慎，要警醒。因為你們的仇敵魔鬼，如同咆哮的獅子，走來走去，尋找可吞吃的人。
1PET|5|9|你們要用堅固的信心抵擋他，因為知道你們在世上的眾弟兄也正在經歷這樣的苦難。
1PET|5|10|那賜一切恩典的上帝曾在基督 裏召了你們，得享他永遠的榮耀，在你們暫受苦難之後，必要親自成全你們，堅固你們，賜力量給你們，建立你們 。
1PET|5|11|願權能歸給他，直到永永遠遠。阿們！
1PET|5|12|我簡單地寫了這信，託我所看為忠心的弟兄 西拉 交給你們，勸勉你們，又證明這恩是上帝真實的恩典；你們務要在這恩上站立得住。
1PET|5|13|在 巴比倫 與你們同蒙揀選的教會向你們問安。我兒子 馬可 也向你們問安。
1PET|5|14|你們要用愛心彼此親吻問安。願平安 歸給你們所有在基督裏的人！
