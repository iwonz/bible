LAM|1|1|How doth the city sit solitary, that was full of people! how is she become as a widow! she that was great among the nations, and princess among the provinces, how is she become tributary!
LAM|1|2|She weepeth sore in the night, and her tears are on her cheeks: among all her lovers she hath none to comfort her: all her friends have dealt treacherously with her, they are become her enemies.
LAM|1|3|Judah is gone into captivity because of affliction, and because of great servitude: she dwelleth among the heathen, she findeth no rest: all her persecutors overtook her between the straits.
LAM|1|4|The ways of Zion do mourn, because none come to the solemn feasts: all her gates are desolate: her priests sigh, her virgins are afflicted, and she is in bitterness.
LAM|1|5|Her adversaries are the chief, her enemies prosper; for the LORD hath afflicted her for the multitude of her transgressions: her children are gone into captivity before the enemy.
LAM|1|6|And from the daughter of Zion all her beauty is departed: her princes are become like harts that find no pasture, and they are gone without strength before the pursuer.
LAM|1|7|Jerusalem remembered in the days of her affliction and of her miseries all her pleasant things that she had in the days of old, when her people fell into the hand of the enemy, and none did help her: the adversaries saw her, and did mock at her sabbaths.
LAM|1|8|Jerusalem hath grievously sinned; therefore she is removed: all that honoured her despise her, because they have seen her nakedness: yea, she sigheth, and turneth backward.
LAM|1|9|Her filthiness is in her skirts; she remembereth not her last end; therefore she came down wonderfully: she had no comforter. O LORD, behold my affliction: for the enemy hath magnified himself.
LAM|1|10|The adversary hath spread out his hand upon all her pleasant things: for she hath seen that the heathen entered into her sanctuary, whom thou didst command that they should not enter into thy congregation.
LAM|1|11|All her people sigh, they seek bread; they have given their pleasant things for meat to relieve the soul: see, O LORD, and consider; for I am become vile.
LAM|1|12|Is it nothing to you, all ye that pass by? behold, and see if there be any sorrow like unto my sorrow, which is done unto me, wherewith the LORD hath afflicted me in the day of his fierce anger.
LAM|1|13|From above hath he sent fire into my bones, and it prevaileth against them: he hath spread a net for my feet, he hath turned me back: he hath made me desolate and faint all the day.
LAM|1|14|The yoke of my transgressions is bound by his hand: they are wreathed, and come up upon my neck: he hath made my strength to fall, the LORD hath delivered me into their hands, from whom I am not able to rise up.
LAM|1|15|The LORD hath trodden under foot all my mighty men in the midst of me: he hath called an assembly against me to crush my young men: the LORD hath trodden the virgin, the daughter of Judah, as in a winepress.
LAM|1|16|For these things I weep; mine eye, mine eye runneth down with water, because the comforter that should relieve my soul is far from me: my children are desolate, because the enemy prevailed.
LAM|1|17|Zion spreadeth forth her hands, and there is none to comfort her: the LORD hath commanded concerning Jacob, that his adversaries should be round about him: Jerusalem is as a menstruous woman among them.
LAM|1|18|The LORD is righteous; for I have rebelled against his commandment: hear, I pray you, all people, and behold my sorrow: my virgins and my young men are gone into captivity.
LAM|1|19|I called for my lovers, but they deceived me: my priests and mine elders gave up the ghost in the city, while they sought their meat to relieve their souls.
LAM|1|20|Behold, O LORD; for I am in distress: my bowels are troubled; mine heart is turned within me; for I have grievously rebelled: abroad the sword bereaveth, at home there is as death.
LAM|1|21|They have heard that I sigh: there is none to comfort me: all mine enemies have heard of my trouble; they are glad that thou hast done it: thou wilt bring the day that thou hast called, and they shall be like unto me.
LAM|1|22|Let all their wickedness come before thee; and do unto them, as thou hast done unto me for all my transgressions: for my sighs are many, and my heart is faint.
LAM|2|1|How hath the LORD covered the daughter of Zion with a cloud in his anger, and cast down from heaven unto the earth the beauty of Israel, and remembered not his footstool in the day of his anger!
LAM|2|2|The LORD hath swallowed up all the habitations of Jacob, and hath not pitied: he hath thrown down in his wrath the strong holds of the daughter of Judah; he hath brought them down to the ground: he hath polluted the kingdom and the princes thereof.
LAM|2|3|He hath cut off in his fierce anger all the horn of Israel: he hath drawn back his right hand from before the enemy, and he burned against Jacob like a flaming fire, which devoureth round about.
LAM|2|4|He hath bent his bow like an enemy: he stood with his right hand as an adversary, and slew all that were pleasant to the eye in the tabernacle of the daughter of Zion: he poured out his fury like fire.
LAM|2|5|The LORD was as an enemy: he hath swallowed up Israel, he hath swallowed up all her palaces: he hath destroyed his strong holds, and hath increased in the daughter of Judah mourning and lamentation.
LAM|2|6|And he hath violently taken away his tabernacle, as if it were of a garden: he hath destroyed his places of the assembly: the LORD hath caused the solemn feasts and sabbaths to be forgotten in Zion, and hath despised in the indignation of his anger the king and the priest.
LAM|2|7|The LORD hath cast off his altar, he hath abhorred his sanctuary, he hath given up into the hand of the enemy the walls of her palaces; they have made a noise in the house of the LORD, as in the day of a solemn feast.
LAM|2|8|The LORD hath purposed to destroy the wall of the daughter of Zion: he hath stretched out a line, he hath not withdrawn his hand from destroying: therefore he made the rampart and the wall to lament; they languished together.
LAM|2|9|Her gates are sunk into the ground; he hath destroyed and broken her bars: her king and her princes are among the Gentiles: the law is no more; her prophets also find no vision from the LORD.
LAM|2|10|The elders of the daughter of Zion sit upon the ground, and keep silence: they have cast up dust upon their heads; they have girded themselves with sackcloth: the virgins of Jerusalem hang down their heads to the ground.
LAM|2|11|Mine eyes do fail with tears, my bowels are troubled, my liver is poured upon the earth, for the destruction of the daughter of my people; because the children and the sucklings swoon in the streets of the city.
LAM|2|12|They say to their mothers, Where is corn and wine? when they swooned as the wounded in the streets of the city, when their soul was poured out into their mothers' bosom.
LAM|2|13|What thing shall I take to witness for thee? what thing shall I liken to thee, O daughter of Jerusalem? what shall I equal to thee, that I may comfort thee, O virgin daughter of Zion? for thy breach is great like the sea: who can heal thee?
LAM|2|14|Thy prophets have seen vain and foolish things for thee: and they have not discovered thine iniquity, to turn away thy captivity; but have seen for thee false burdens and causes of banishment.
LAM|2|15|All that pass by clap their hands at thee; they hiss and wag their head at the daughter of Jerusalem, saying, Is this the city that men call The perfection of beauty, The joy of the whole earth?
LAM|2|16|All thine enemies have opened their mouth against thee: they hiss and gnash the teeth: they say, We have swallowed her up: certainly this is the day that we looked for; we have found, we have seen it.
LAM|2|17|The LORD hath done that which he had devised; he hath fulfilled his word that he had commanded in the days of old: he hath thrown down, and hath not pitied: and he hath caused thine enemy to rejoice over thee, he hath set up the horn of thine adversaries.
LAM|2|18|Their heart cried unto the LORD, O wall of the daughter of Zion, let tears run down like a river day and night: give thyself no rest; let not the apple of thine eye cease.
LAM|2|19|Arise, cry out in the night: in the beginning of the watches pour out thine heart like water before the face of the LORD: lift up thy hands toward him for the life of thy young children, that faint for hunger in the top of every street.
LAM|2|20|Behold, O LORD, and consider to whom thou hast done this. Shall the women eat their fruit, and children of a span long? shall the priest and the prophet be slain in the sanctuary of the Lord?
LAM|2|21|The young and the old lie on the ground in the streets: my virgins and my young men are fallen by the sword; thou hast slain them in the day of thine anger; thou hast killed, and not pitied.
LAM|2|22|Thou hast called as in a solemn day my terrors round about, so that in the day of the LORD's anger none escaped nor remained: those that I have swaddled and brought up hath mine enemy consumed.
LAM|3|1|I AM the man that hath seen affliction by the rod of his wrath.
LAM|3|2|He hath led me, and brought me into darkness, but not into light.
LAM|3|3|Surely against me is he turned; he turneth his hand against me all the day.
LAM|3|4|My flesh and my skin hath he made old; he hath broken my bones.
LAM|3|5|He hath builded against me, and compassed me with gall and travail.
LAM|3|6|He hath set me in dark places, as they that be dead of old.
LAM|3|7|He hath hedged me about, that I cannot get out: he hath made my chain heavy.
LAM|3|8|Also when I cry and shout, he shutteth out my prayer.
LAM|3|9|He hath inclosed my ways with hewn stone, he hath made my paths crooked.
LAM|3|10|He was unto me as a bear lying in wait, and as a lion in secret places.
LAM|3|11|He hath turned aside my ways, and pulled me in pieces: he hath made me desolate.
LAM|3|12|He hath bent his bow, and set me as a mark for the arrow.
LAM|3|13|He hath caused the arrows of his quiver to enter into my reins.
LAM|3|14|I was a derision to all my people; and their song all the day.
LAM|3|15|He hath filled me with bitterness, he hath made me drunken with wormwood.
LAM|3|16|He hath also broken my teeth with gravel stones, he hath covered me with ashes.
LAM|3|17|And thou hast removed my soul far off from peace: I forgat prosperity.
LAM|3|18|And I said, My strength and my hope is perished from the LORD:
LAM|3|19|Remembering mine affliction and my misery, the wormwood and the gall.
LAM|3|20|My soul hath them still in remembrance, and is humbled in me.
LAM|3|21|This I recall to my mind, therefore have I hope.
LAM|3|22|It is of the LORD's mercies that we are not consumed, because his compassions fail not.
LAM|3|23|They are new every morning: great is thy faithfulness.
LAM|3|24|The LORD is my portion, saith my soul; therefore will I hope in him.
LAM|3|25|The LORD is good unto them that wait for him, to the soul that seeketh him.
LAM|3|26|It is good that a man should both hope and quietly wait for the salvation of the LORD.
LAM|3|27|It is good for a man that he bear the yoke of his youth.
LAM|3|28|He sitteth alone and keepeth silence, because he hath borne it upon him.
LAM|3|29|He putteth his mouth in the dust; if so be there may be hope.
LAM|3|30|He giveth his cheek to him that smiteth him: he is filled full with reproach.
LAM|3|31|For the LORD will not cast off for ever:
LAM|3|32|But though he cause grief, yet will he have compassion according to the multitude of his mercies.
LAM|3|33|For he doth not afflict willingly nor grieve the children of men.
LAM|3|34|To crush under his feet all the prisoners of the earth.
LAM|3|35|To turn aside the right of a man before the face of the most High,
LAM|3|36|To subvert a man in his cause, the LORD approveth not.
LAM|3|37|Who is he that saith, and it cometh to pass, when the Lord commandeth it not?
LAM|3|38|Out of the mouth of the most High proceedeth not evil and good?
LAM|3|39|Wherefore doth a living man complain, a man for the punishment of his sins?
LAM|3|40|Let us search and try our ways, and turn again to the LORD.
LAM|3|41|Let us lift up our heart with our hands unto God in the heavens.
LAM|3|42|We have transgressed and have rebelled: thou hast not pardoned.
LAM|3|43|Thou hast covered with anger, and persecuted us: thou hast slain, thou hast not pitied.
LAM|3|44|Thou hast covered thyself with a cloud, that our prayer should not pass through.
LAM|3|45|Thou hast made us as the offscouring and refuse in the midst of the people.
LAM|3|46|All our enemies have opened their mouths against us.
LAM|3|47|Fear and a snare is come upon us, desolation and destruction.
LAM|3|48|Mine eye runneth down with rivers of water for the destruction of the daughter of my people.
LAM|3|49|Mine eye trickleth down, and ceaseth not, without any intermission.
LAM|3|50|Till the LORD look down, and behold from heaven.
LAM|3|51|Mine eye affecteth mine heart because of all the daughters of my city.
LAM|3|52|Mine enemies chased me sore, like a bird, without cause.
LAM|3|53|They have cut off my life in the dungeon, and cast a stone upon me.
LAM|3|54|Waters flowed over mine head; then I said, I am cut off.
LAM|3|55|I called upon thy name, O LORD, out of the low dungeon.
LAM|3|56|Thou hast heard my voice: hide not thine ear at my breathing, at my cry.
LAM|3|57|Thou drewest near in the day that I called upon thee: thou saidst, Fear not.
LAM|3|58|O LORD, thou hast pleaded the causes of my soul; thou hast redeemed my life.
LAM|3|59|O LORD, thou hast seen my wrong: judge thou my cause.
LAM|3|60|Thou hast seen all their vengeance and all their imaginations against me.
LAM|3|61|Thou hast heard their reproach, O LORD, and all their imaginations against me;
LAM|3|62|The lips of those that rose up against me, and their device against me all the day.
LAM|3|63|Behold their sitting down, and their rising up; I am their musick.
LAM|3|64|Render unto them a recompence, O LORD, according to the work of their hands.
LAM|3|65|Give them sorrow of heart, thy curse unto them.
LAM|3|66|Persecute and destroy them in anger from under the heavens of the LORD.
LAM|4|1|How is the gold become dim! how is the most fine gold changed! the stones of the sanctuary are poured out in the top of every street.
LAM|4|2|The precious sons of Zion, comparable to fine gold, how are they esteemed as earthen pitchers, the work of the hands of the potter!
LAM|4|3|Even the sea monsters draw out the breast, they give suck to their young ones: the daughter of my people is become cruel, like the ostriches in the wilderness.
LAM|4|4|The tongue of the sucking child cleaveth to the roof of his mouth for thirst: the young children ask bread, and no man breaketh it unto them.
LAM|4|5|They that did feed delicately are desolate in the streets: they that were brought up in scarlet embrace dunghills.
LAM|4|6|For the punishment of the iniquity of the daughter of my people is greater than the punishment of the sin of Sodom, that was overthrown as in a moment, and no hands stayed on her.
LAM|4|7|Her Nazarites were purer than snow, they were whiter than milk, they were more ruddy in body than rubies, their polishing was of sapphire:
LAM|4|8|Their visage is blacker than a coal; they are not known in the streets: their skin cleaveth to their bones; it is withered, it is become like a stick.
LAM|4|9|They that be slain with the sword are better than they that be slain with hunger: for these pine away, stricken through for want of the fruits of the field.
LAM|4|10|The hands of the pitiful women have sodden their own children: they were their meat in the destruction of the daughter of my people.
LAM|4|11|The LORD hath accomplished his fury; he hath poured out his fierce anger, and hath kindled a fire in Zion, and it hath devoured the foundations thereof.
LAM|4|12|The kings of the earth, and all the inhabitants of the world, would not have believed that the adversary and the enemy should have entered into the gates of Jerusalem.
LAM|4|13|For the sins of her prophets, and the iniquities of her priests, that have shed the blood of the just in the midst of her,
LAM|4|14|They have wandered as blind men in the streets, they have polluted themselves with blood, so that men could not touch their garments.
LAM|4|15|They cried unto them, Depart ye; it is unclean; depart, depart, touch not: when they fled away and wandered, they said among the heathen, They shall no more sojourn there.
LAM|4|16|The anger of the LORD hath divided them; he will no more regard them: they respected not the persons of the priests, they favoured not the elders.
LAM|4|17|As for us, our eyes as yet failed for our vain help: in our watching we have watched for a nation that could not save us.
LAM|4|18|They hunt our steps, that we cannot go in our streets: our end is near, our days are fulfilled; for our end is come.
LAM|4|19|Our persecutors are swifter than the eagles of the heaven: they pursued us upon the mountains, they laid wait for us in the wilderness.
LAM|4|20|The breath of our nostrils, the anointed of the LORD, was taken in their pits, of whom we said, Under his shadow we shall live among the heathen.
LAM|4|21|Rejoice and be glad, O daughter of Edom, that dwellest in the land of Uz; the cup also shall pass through unto thee: thou shalt be drunken, and shalt make thyself naked.
LAM|4|22|The punishment of thine iniquity is accomplished, O daughter of Zion; he will no more carry thee away into captivity: he will visit thine iniquity, O daughter of Edom; he will discover thy sins.
LAM|5|1|Remember, O LORD, what is come upon us: consider, and behold our reproach.
LAM|5|2|Our inheritance is turned to strangers, our houses to aliens.
LAM|5|3|We are orphans and fatherless, our mothers are as widows.
LAM|5|4|We have drunken our water for money; our wood is sold unto us.
LAM|5|5|Our necks are under persecution: we labour, and have no rest.
LAM|5|6|We have given the hand to the Egyptians, and to the Assyrians, to be satisfied with bread.
LAM|5|7|Our fathers have sinned, and are not; and we have borne their iniquities.
LAM|5|8|Servants have ruled over us: there is none that doth deliver us out of their hand.
LAM|5|9|We gat our bread with the peril of our lives because of the sword of the wilderness.
LAM|5|10|Our skin was black like an oven because of the terrible famine.
LAM|5|11|They ravished the women in Zion, and the maids in the cities of Judah.
LAM|5|12|Princes are hanged up by their hand: the faces of elders were not honoured.
LAM|5|13|They took the young men to grind, and the children fell under the wood.
LAM|5|14|The elders have ceased from the gate, the young men from their musick.
LAM|5|15|The joy of our heart is ceased; our dance is turned into mourning.
LAM|5|16|The crown is fallen from our head: woe unto us, that we have sinned!
LAM|5|17|For this our heart is faint; for these things our eyes are dim.
LAM|5|18|Because of the mountain of Zion, which is desolate, the foxes walk upon it.
LAM|5|19|Thou, O LORD, remainest for ever; thy throne from generation to generation.
LAM|5|20|Wherefore dost thou forget us for ever, and forsake us so long time?
LAM|5|21|Turn thou us unto thee, O LORD, and we shall be turned; renew our days as of old.
LAM|5|22|But thou hast utterly rejected us; thou art very wroth against us.
