ACTS|1|1|In the first book, O Theophilus, I have dealt with all that Jesus began to do and teach,
ACTS|1|2|until the day when he was taken up, after he had given commands through the Holy Spirit to the apostles whom he had chosen.
ACTS|1|3|To them he presented himself alive after his suffering by many proofs, appearing to them during forty days and speaking about the kingdom of God.
ACTS|1|4|And while staying with them he ordered them not to depart from Jerusalem, but to wait for the promise of the Father, which, he said, "you heard from me;
ACTS|1|5|for John baptized with water, but you will be baptized with the Holy Spirit not many days from now."
ACTS|1|6|So when they had come together, they asked him, "Lord, will you at this time restore the kingdom to Israel?"
ACTS|1|7|He said to them, "It is not for you to know times or seasons that the Father has fixed by his own authority.
ACTS|1|8|But you will receive power when the Holy Spirit has come upon you, and you will be my witnesses in Jerusalem and in all Judea and Samaria, and to the end of the earth."
ACTS|1|9|And when he had said these things, as they were looking on, he was lifted up, and a cloud took him out of their sight.
ACTS|1|10|And while they were gazing into heaven as he went, behold, two men stood by them in white robes,
ACTS|1|11|and said, "Men of Galilee, why do you stand looking into heaven? This Jesus, who was taken up from you into heaven, will come in the same way as you saw him go into heaven."
ACTS|1|12|Then they returned to Jerusalem from the mount called Olivet, which is near Jerusalem, a Sabbath day's journey away.
ACTS|1|13|And when they had entered, they went up to the upper room, where they were staying, Peter and John and James and Andrew, Philip and Thomas, Bartholomew and Matthew, James the son of Alphaeus and Simon the Zealot and Judas the son of James.
ACTS|1|14|All these with one accord were devoting themselves to prayer, together with the women and Mary the mother of Jesus, and his brothers.
ACTS|1|15|In those days Peter stood up among the brothers (the company of persons was in all about 120) and said,
ACTS|1|16|"Brothers, the Scripture had to be fulfilled, which the Holy Spirit spoke beforehand by the mouth of David concerning Judas, who became a guide to those who arrested Jesus.
ACTS|1|17|For he was numbered among us and was allotted his share in this ministry."
ACTS|1|18|(Now this man bought a field with the reward of his wickedness, and falling headlong he burst open in the middle and all his bowels gushed out.
ACTS|1|19|And it became known to all the inhabitants of Jerusalem, so that the field was called in their own language Akeldama, that is, Field of Blood.)
ACTS|1|20|"For it is written in the Book of Psalms, "' May his camp become desolate, and let there be no one to dwell in it'; and "'Let another take his office.'
ACTS|1|21|So one of the men who have accompanied us during all the time that the Lord Jesus went in and out among us,
ACTS|1|22|beginning from the baptism of John until the day when he was taken up from us- one of these men must become with us a witness to his resurrection."
ACTS|1|23|And they put forward two, Joseph called Barsabbas, who was also called Justus, and Matthias.
ACTS|1|24|And they prayed and said, "You, Lord, who know the hearts of all, show which one of these two you have chosen
ACTS|1|25|to take the place in this ministry and apostleship from which Judas turned aside to go to his own place."
ACTS|1|26|And they cast lots for them, and the lot fell on Matthias, and he was numbered with the eleven apostles.
ACTS|2|1|When the day of Pentecost arrived, they were all together in one place.
ACTS|2|2|And suddenly there came from heaven a sound like a mighty rushing wind, and it filled the entire house where they were sitting.
ACTS|2|3|And divided tongues as of fire appeared to them and rested on each one of them.
ACTS|2|4|And they were all filled with the Holy Spirit and began to speak in other tongues as the Spirit gave them utterance.
ACTS|2|5|Now there were dwelling in Jerusalem Jews, devout men from every nation under heaven.
ACTS|2|6|And at this sound the multitude came together, and they were bewildered, because each one was hearing them speak in his own language.
ACTS|2|7|And they were amazed and astonished, saying, "Are not all these who are speaking Galileans?
ACTS|2|8|And how is it that we hear, each of us in his own native language?
ACTS|2|9|Parthians and Medes and Elamites and residents of Mesopotamia, Judea and Cappadocia, Pontus and Asia,
ACTS|2|10|Phrygia and Pamphylia, Egypt and the parts of Libya belonging to Cyrene, and visitors from Rome,
ACTS|2|11|both Jews and proselytes, Cretans and Arabians- we hear them telling in our own tongues the mighty works of God."
ACTS|2|12|And all were amazed and perplexed, saying to one another, "What does this mean?"
ACTS|2|13|But others mocking said, "They are filled with new wine."
ACTS|2|14|But Peter, standing with the eleven, lifted up his voice and addressed them, "Men of Judea and all who dwell in Jerusalem, let this be known to you, and give ear to my words.
ACTS|2|15|For these men are not drunk, as you suppose, since it is only the third hour of the day.
ACTS|2|16|But this is what was uttered through the prophet Joel:
ACTS|2|17|"'And in the last days it shall be, God declares, that I will pour out my Spirit on all flesh, and your sons and your daughters shall prophesy, and your young men shall see visions, and your old men shall dream dreams;
ACTS|2|18|even on my male servants and female servants in those days I will pour out my Spirit, and they shall prophesy.
ACTS|2|19|And I will show wonders in the heavens above and signs on the earth below, blood, and fire, and vapor of smoke;
ACTS|2|20|the sun shall be turned to darkness and the moon to blood, before the day of the Lord comes, the great and magnificent day.
ACTS|2|21|And it shall come to pass that everyone who calls upon the name of the Lord shall be saved.'
ACTS|2|22|"Men of Israel, hear these words: Jesus of Nazareth, a man attested to you by God with mighty works and wonders and signs that God did through him in your midst, as you yourselves know-
ACTS|2|23|this Jesus, delivered up according to the definite plan and foreknowledge of God, you crucified and killed by the hands of lawless men.
ACTS|2|24|God raised him up, loosing the pangs of death, because it was not possible for him to be held by it.
ACTS|2|25|For David says concerning him, "' I saw the Lord always before me, for he is at my right hand that I may not be shaken;
ACTS|2|26|therefore my heart was glad, and my tongue rejoiced; my flesh also will dwell in hope.
ACTS|2|27|For you will not abandon my soul to Hades, or let your Holy One see corruption.
ACTS|2|28|You have made known to me the paths of life; you will make me full of gladness with your presence.'
ACTS|2|29|"Brothers, I may say to you with confidence about the patriarch David that he both died and was buried, and his tomb is with us to this day.
ACTS|2|30|Being therefore a prophet, and knowing that God had sworn with an oath to him that he would set one of his descendants on his throne,
ACTS|2|31|he foresaw and spoke about the resurrection of the Christ, that he was not abandoned to Hades, nor did his flesh see corruption.
ACTS|2|32|This Jesus God raised up, and of that we all are witnesses.
ACTS|2|33|Being therefore exalted at the right hand of God, and having received from the Father the promise of the Holy Spirit, he has poured out this that you yourselves are seeing and hearing.
ACTS|2|34|For David did not ascend into the heavens, but he himself says, "' The Lord said to my Lord, Sit at my right hand,
ACTS|2|35|until I make your enemies your footstool.'
ACTS|2|36|Let all the house of Israel therefore know for certain that God has made him both Lord and Christ, this Jesus whom you crucified."
ACTS|2|37|Now when they heard this they were cut to the heart, and said to Peter and the rest of the apostles, "Brothers, what shall we do?"
ACTS|2|38|And Peter said to them, "Repent and be baptized every one of you in the name of Jesus Christ for the forgiveness of your sins, and you will receive the gift of the Holy Spirit.
ACTS|2|39|For the promise is for you and for your children and for all who are far off, everyone whom the Lord our God calls to himself."
ACTS|2|40|And with many other words he bore witness and continued to exhort them, saying, "Save yourselves from this crooked generation."
ACTS|2|41|So those who received his word were baptized, and there were added that day about three thousand souls.
ACTS|2|42|And they devoted themselves to the apostles' teaching and fellowship, to the breaking of bread and the prayers.
ACTS|2|43|And awe came upon every soul, and many wonders and signs were being done through the apostles.
ACTS|2|44|And all who believed were together and had all things in common.
ACTS|2|45|And they were selling their possessions and belongings and distributing the proceeds to all, as any had need.
ACTS|2|46|And day by day, attending the temple together and breaking bread in their homes, they received their food with glad and generous hearts,
ACTS|2|47|praising God and having favor with all the people. And the Lord added to their number day by day those who were being saved.
ACTS|3|1|Now Peter and John were going up to the temple at the hour of prayer, the ninth hour.
ACTS|3|2|And a man lame from birth was being carried, whom they laid daily at the gate of the temple that is called the Beautiful Gate to ask alms of those entering the temple.
ACTS|3|3|Seeing Peter and John about to go into the temple, he asked to receive alms.
ACTS|3|4|And Peter directed his gaze at him, as did John, and said, "Look at us."
ACTS|3|5|And he fixed his attention on them, expecting to receive something from them.
ACTS|3|6|But Peter said, "I have no silver and gold, but what I do have I give to you. In the name of Jesus Christ of Nazareth, rise up and walk!"
ACTS|3|7|And he took him by the right hand and raised him up, and immediately his feet and ankles were made strong.
ACTS|3|8|And leaping up he stood and began to walk, and entered the temple with them, walking and leaping and praising God.
ACTS|3|9|And all the people saw him walking and praising God,
ACTS|3|10|and recognized him as the one who sat at the Beautiful Gate of the temple, asking for alms. And they were filled with wonder and amazement at what had happened to him.
ACTS|3|11|While he clung to Peter and John, all the people ran together to them in the portico called Solomon's, astounded.
ACTS|3|12|And when Peter saw it he addressed the people: "Men of Israel, why do you wonder at this, or why do you stare at us, as though by our own power or piety we have made him walk?
ACTS|3|13|The God of Abraham, the God of Isaac, and the God of Jacob, the God of our fathers, glorified his servant Jesus, whom you delivered over and denied in the presence of Pilate, when he had decided to release him.
ACTS|3|14|But you denied the Holy and Righteous One, and asked for a murderer to be granted to you,
ACTS|3|15|and you killed the Author of life, whom God raised from the dead. To this we are witnesses.
ACTS|3|16|And his name- by faith in his name- has made this man strong whom you see and know, and the faith that is through Jesus has given the man this perfect health in the presence of you all.
ACTS|3|17|"And now, brothers, I know that you acted in ignorance, as did also your rulers.
ACTS|3|18|But what God foretold by the mouth of all the prophets, that his Christ would suffer, he thus fulfilled.
ACTS|3|19|Repent therefore, and turn again, that your sins may be blotted out,
ACTS|3|20|that times of refreshing may come from the presence of the Lord, and that he may send the Christ appointed for you, Jesus,
ACTS|3|21|whom heaven must receive until the time for restoring all the things about which God spoke by the mouth of his holy prophets long ago.
ACTS|3|22|Moses said, 'The Lord God will raise up for you a prophet like me from your brothers. You shall listen to him in whatever he tells you.
ACTS|3|23|And it shall be that every soul who does not listen to that prophet shall be destroyed from the people.'
ACTS|3|24|And all the prophets who have spoken, from Samuel and those who came after him, also proclaimed these days.
ACTS|3|25|You are the sons of the prophets and of the covenant that God made with your fathers, saying to Abraham, 'And in your offspring shall all the families of the earth be blessed.'
ACTS|3|26|God, having raised up his servant, sent him to you first, to bless you by turning every one of you from your wickedness."
ACTS|4|1|And as they were speaking to the people, the priests and the captain of the temple and the Sadducees came upon them,
ACTS|4|2|greatly annoyed because they were teaching the people and proclaiming in Jesus the resurrection from the dead.
ACTS|4|3|And they arrested them and put them in custody until the next day, for it was already evening.
ACTS|4|4|But many of those who had heard the word believed, and the number of the men came to about five thousand.
ACTS|4|5|On the next day their rulers and elders and scribes gathered together in Jerusalem,
ACTS|4|6|with Annas the high priest and Caiaphas and John and Alexander, and all who were of the high-priestly family.
ACTS|4|7|And when they had set them in the midst, they inquired, "By what power or by what name did you do this?"
ACTS|4|8|Then Peter, filled with the Holy Spirit, said to them, "Rulers of the people and elders,
ACTS|4|9|if we are being examined today concerning a good deed done to a crippled man, by what means this man has been healed,
ACTS|4|10|let it be known to all of you and to all the people of Israel that by the name of Jesus Christ of Nazareth, whom you crucified, whom God raised from the dead- by him this man is standing before you well.
ACTS|4|11|This Jesus is the stone that was rejected by you, the builders, which has become the cornerstone.
ACTS|4|12|And there is salvation in no one else, for there is no other name under heaven given among men by which we must be saved."
ACTS|4|13|Now when they saw the boldness of Peter and John, and perceived that they were uneducated, common men, they were astonished. And they recognized that they had been with Jesus.
ACTS|4|14|But seeing the man who was healed standing beside them, they had nothing to say in opposition.
ACTS|4|15|But when they had commanded them to leave the council, they conferred with one another,
ACTS|4|16|saying, "What shall we do with these men? For that a notable sign has been performed through them is evident to all the inhabitants of Jerusalem, and we cannot deny it.
ACTS|4|17|But in order that it may spread no further among the people, let us warn them to speak no more to anyone in this name."
ACTS|4|18|So they called them and charged them not to speak or teach at all in the name of Jesus.
ACTS|4|19|But Peter and John answered them, "Whether it is right in the sight of God to listen to you rather than to God, you must judge,
ACTS|4|20|for we cannot but speak of what we have seen and heard."
ACTS|4|21|And when they had further threatened them, they let them go, finding no way to punish them, because of the people, for all were praising God for what had happened.
ACTS|4|22|For the man on whom this sign of healing was performed was more than forty years old.
ACTS|4|23|When they were released, they went to their friends and reported what the chief priests and the elders had said to them.
ACTS|4|24|And when they heard it, they lifted their voices together to God and said, "Sovereign Lord, who made the heaven and the earth and the sea and everything in them,
ACTS|4|25|who through the mouth of our father David, your servant, said by the Holy Spirit, "' Why did the Gentiles rage, and the peoples plot in vain?
ACTS|4|26|The kings of the earth set themselves, and the rulers were gathered together, against the Lord and against his Anointed'-
ACTS|4|27|for truly in this city there were gathered together against your holy servant Jesus, whom you anointed, both Herod and Pontius Pilate, along with the Gentiles and the peoples of Israel,
ACTS|4|28|to do whatever your hand and your plan had predestined to take place.
ACTS|4|29|And now, Lord, look upon their threats and grant to your servants to continue to speak your word with all boldness,
ACTS|4|30|while you stretch out your hand to heal, and signs and wonders are performed through the name of your holy servant Jesus."
ACTS|4|31|And when they had prayed, the place in which they were gathered together was shaken, and they were all filled with the Holy Spirit and continued to speak the word of God with boldness.
ACTS|4|32|Now the full number of those who believed were of one heart and soul, and no one said that any of the things that belonged to him was his own, but they had everything in common.
ACTS|4|33|And with great power the apostles were giving their testimony to the resurrection of the Lord Jesus, and great grace was upon them all.
ACTS|4|34|There was not a needy person among them, for as many as were owners of lands or houses sold them and brought the proceeds of what was sold
ACTS|4|35|and laid it at the apostles' feet, and it was distributed to each as any had need.
ACTS|4|36|Thus Joseph, who was also called by the apostles Barnabas (which means son of encouragement), a Levite, a native of Cyprus,
ACTS|4|37|sold a field that belonged to him and brought the money and laid it at the apostles' feet.
ACTS|5|1|But a man named Ananias, with his wife Sapphira, sold a piece of property,
ACTS|5|2|and with his wife's knowledge he kept back for himself some of the proceeds and brought only a part of it and laid it at the apostles' feet.
ACTS|5|3|But Peter said, "Ananias, why has Satan filled your heart to lie to the Holy Spirit and to keep back for yourself part of the proceeds of the land?
ACTS|5|4|While it remained unsold, did it not remain your own? And after it was sold, was it not at your disposal? Why is it that you have contrived this deed in your heart? You have not lied to men but to God."
ACTS|5|5|When Ananias heard these words, he fell down and breathed his last. And great fear came upon all who heard of it.
ACTS|5|6|The young men rose and wrapped him up and carried him out and buried him.
ACTS|5|7|After an interval of about three hours his wife came in, not knowing what had happened.
ACTS|5|8|And Peter said to her, "Tell me whether you sold the land for so much." And she said, "Yes, for so much."
ACTS|5|9|But Peter said to her, "How is it that you have agreed together to test the Spirit of the Lord? Behold, the feet of those who have buried your husband are at the door, and they will carry you out."
ACTS|5|10|Immediately she fell down at his feet and breathed her last. When the young men came in they found her dead, and they carried her out and buried her beside her husband.
ACTS|5|11|And great fear came upon the whole church and upon all who heard of these things.
ACTS|5|12|Now many signs and wonders were regularly done among the people by the hands of the apostles. And they were all together in Solomon's Portico.
ACTS|5|13|None of the rest dared join them, but the people held them in high esteem.
ACTS|5|14|And more than ever believers were added to the Lord, multitudes of both men and women,
ACTS|5|15|so that they even carried out the sick into the streets and laid them on cots and mats, that as Peter came by at least his shadow might fall on some of them.
ACTS|5|16|The people also gathered from the towns around Jerusalem, bringing the sick and those afflicted with unclean spirits, and they were all healed.
ACTS|5|17|But the high priest rose up, and all who were with him (that is, the party of the Sadducees), and filled with jealousy
ACTS|5|18|they arrested the apostles and put them in the public prison.
ACTS|5|19|But during the night an angel of the Lord opened the prison doors and brought them out, and said,
ACTS|5|20|"Go and stand in the temple and speak to the people all the words of this Life."
ACTS|5|21|And when they heard this, they entered the temple at daybreak and began to teach. Now when the high priest came, and those who were with him, they called together the council and all the senate of Israel and sent to the prison to have them brought.
ACTS|5|22|But when the officers came, they did not find them in the prison, so they returned and reported,
ACTS|5|23|"We found the prison securely locked and the guards standing at the doors, but when we opened them we found no one inside."
ACTS|5|24|Now when the captain of the temple and the chief priests heard these words, they were greatly perplexed about them, wondering what this would come to.
ACTS|5|25|And someone came and told them, "Look! The men whom you put in prison are standing in the temple and teaching the people."
ACTS|5|26|Then the captain with the officers went and brought them, but not by force, for they were afraid of being stoned by the people.
ACTS|5|27|And when they had brought them, they set them before the council. And the high priest questioned them,
ACTS|5|28|saying, "We strictly charged you not to teach in this name, yet here you have filled Jerusalem with your teaching, and you intend to bring this man's blood upon us."
ACTS|5|29|But Peter and the apostles answered, "We must obey God rather than men.
ACTS|5|30|The God of our fathers raised Jesus, whom you killed by hanging him on a tree.
ACTS|5|31|God exalted him at his right hand as Leader and Savior, to give repentance to Israel and forgiveness of sins.
ACTS|5|32|And we are witnesses to these things, and so is the Holy Spirit, whom God has given to those who obey him."
ACTS|5|33|When they heard this, they were enraged and wanted to kill them.
ACTS|5|34|But a Pharisee in the council named Gamaliel, a teacher of the law held in honor by all the people, stood up and gave orders to put the men outside for a little while.
ACTS|5|35|And he said to them, "Men of Israel, take care what you are about to do with these men.
ACTS|5|36|For before these days Theudas rose up, claiming to be somebody, and a number of men, about four hundred, joined him. He was killed, and all who followed him were dispersed and came to nothing.
ACTS|5|37|After him Judas the Galilean rose up in the days of the census and drew away some of the people after him. He too perished, and all who followed him were scattered.
ACTS|5|38|So in the present case I tell you, keep away from these men and let them alone, for if this plan or this undertaking is of man, it will fail;
ACTS|5|39|but if it is of God, you will not be able to overthrow them. You might even be found opposing God!" So they took his advice,
ACTS|5|40|and when they had called in the apostles, they beat them and charged them not to speak in the name of Jesus, and let them go.
ACTS|5|41|Then they left the presence of the council, rejoicing that they were counted worthy to suffer dishonor for the name.
ACTS|5|42|And every day, in the temple and from house to house, they did not cease teaching and preaching Jesus as the Christ.
ACTS|6|1|Now in these days when the disciples were increasing in number, a complaint by the Hellenists arose against the Hebrews because their widows were being neglected in the daily distribution.
ACTS|6|2|And the twelve summoned the full number of the disciples and said, "It is not right that we should give up preaching the word of God to serve tables.
ACTS|6|3|Therefore, brothers, pick out from among you seven men of good repute, full of the Spirit and of wisdom, whom we will appoint to this duty.
ACTS|6|4|But we will devote ourselves to prayer and to the ministry of the word."
ACTS|6|5|And what they said pleased the whole gathering, and they chose Stephen, a man full of faith and of the Holy Spirit, and Philip, and Prochorus, and Nicanor, and Timon, and Parmenas, and Nicolaus, a proselyte of Antioch.
ACTS|6|6|These they set before the apostles, and they prayed and laid their hands on them.
ACTS|6|7|And the word of God continued to increase, and the number of the disciples multiplied greatly in Jerusalem, and a great many of the priests became obedient to the faith.
ACTS|6|8|And Stephen, full of grace and power, was doing great wonders and signs among the people.
ACTS|6|9|Then some of those who belonged to the synagogue of the Freedmen (as it was called), and of the Cyrenians, and of the Alexandrians, and of those from Cilicia and Asia, rose up and disputed with Stephen.
ACTS|6|10|But they could not withstand the wisdom and the Spirit with which he was speaking.
ACTS|6|11|Then they secretly instigated men who said, "We have heard him speak blasphemous words against Moses and God."
ACTS|6|12|And they stirred up the people and the elders and the scribes, and they came upon him and seized him and brought him before the council,
ACTS|6|13|and they set up false witnesses who said, "This man never ceases to speak words against this holy place and the law,
ACTS|6|14|for we have heard him say that this Jesus of Nazareth will destroy this place and will change the customs that Moses delivered to us."
ACTS|6|15|And gazing at him, all who sat in the council saw that his face was like the face of an angel.
ACTS|7|1|And the high priest said, "Are these things so?"
ACTS|7|2|And Stephen said: "Brothers and fathers, hear me. The God of glory appeared to our father Abraham when he was in Mesopotamia, before he lived in Haran,
ACTS|7|3|and said to him, 'Go out from your land and from your kindred and go into the land that I will show you.'
ACTS|7|4|Then he went out from the land of the Chaldeans and lived in Haran. And after his father died, God removed him from there into this land in which you are now living.
ACTS|7|5|Yet he gave him no inheritance in it, not even a foot's length, but promised to give it to him as a possession and to his offspring after him, though he had no child.
ACTS|7|6|And God spoke to this effect- that his offspring would be sojourners in a land belonging to others, who would enslave them and afflict them four hundred years.
ACTS|7|7|'But I will judge the nation that they serve,' said God, 'and after that they shall come out and worship me in this place.'
ACTS|7|8|And he gave him the covenant of circumcision. And so Abraham became the father of Isaac, and circumcised him on the eighth day, and Isaac became the father of Jacob, and Jacob of the twelve patriarchs.
ACTS|7|9|"And the patriarchs, jealous of Joseph, sold him into Egypt; but God was with him
ACTS|7|10|and rescued him out of all his afflictions and gave him favor and wisdom before Pharaoh, king of Egypt, who made him ruler over Egypt and over all his household.
ACTS|7|11|Now there came a famine throughout all Egypt and Canaan, and great affliction, and our fathers could find no food.
ACTS|7|12|But when Jacob heard that there was grain in Egypt, he sent out our fathers on their first visit.
ACTS|7|13|And on the second visit Joseph made himself known to his brothers, and Joseph's family became known to Pharaoh.
ACTS|7|14|And Joseph sent and summoned Jacob his father and all his kindred, seventy-five persons in all.
ACTS|7|15|And Jacob went down into Egypt, and he died, he and our fathers,
ACTS|7|16|and they were carried back to Shechem and laid in the tomb that Abraham had bought for a sum of silver from the sons of Hamor in Shechem.
ACTS|7|17|"But as the time of the promise drew near, which God had granted to Abraham, the people increased and multiplied in Egypt
ACTS|7|18|until there arose over Egypt another king who did not know Joseph.
ACTS|7|19|He dealt shrewdly with our race and forced our fathers to expose their infants, so that they would not be kept alive.
ACTS|7|20|At this time Moses was born; and he was beautiful in God's sight. And he was brought up for three months in his father's house,
ACTS|7|21|and when he was exposed, Pharaoh's daughter adopted him and brought him up as her own son.
ACTS|7|22|And Moses was instructed in all the wisdom of the Egyptians, and he was mighty in his words and deeds.
ACTS|7|23|"When he was forty years old, it came into his heart to visit his brothers, the children of Israel.
ACTS|7|24|And seeing one of them being wronged, he defended the oppressed man and avenged him by striking down the Egyptian.
ACTS|7|25|He supposed that his brothers would understand that God was giving them salvation by his hand, but they did not understand.
ACTS|7|26|And on the following day he appeared to them as they were quarreling and tried to reconcile them, saying, 'Men, you are brothers. Why do you wrong each other?'
ACTS|7|27|But the man who was wronging his neighbor thrust him aside, saying, 'Who made you a ruler and a judge over us?
ACTS|7|28|Do you want to kill me as you killed the Egyptian yesterday?'
ACTS|7|29|At this retort Moses fled and became an exile in the land of Midian, where he became the father of two sons.
ACTS|7|30|"Now when forty years had passed, an angel appeared to him in the wilderness of Mount Sinai, in a flame of fire in a bush.
ACTS|7|31|When Moses saw it, he was amazed at the sight, and as he drew near to look, there came the voice of the Lord:
ACTS|7|32|'I am the God of your fathers, the God of Abraham and of Isaac and of Jacob.' And Moses trembled and did not dare to look.
ACTS|7|33|Then the Lord said to him, 'Take off the sandals from your feet, for the place where you are standing is holy ground.
ACTS|7|34|I have surely seen the affliction of my people who are in Egypt, and have heard their groaning, and I have come down to deliver them. And now come, I will send you to Egypt.'
ACTS|7|35|"This Moses, whom they rejected, saying, 'Who made you a ruler and a judge?'- this man God sent as both ruler and redeemer by the hand of the angel who appeared to him in the bush.
ACTS|7|36|This man led them out, performing wonders and signs in Egypt and at the Red Sea and in the wilderness for forty years.
ACTS|7|37|This is the Moses who said to the Israelites, 'God will raise up for you a prophet like me from your brothers.'
ACTS|7|38|This is the one who was in the congregation in the wilderness with the angel who spoke to him at Mount Sinai, and with our fathers. He received living oracles to give to us.
ACTS|7|39|Our fathers refused to obey him, but thrust him aside, and in their hearts they turned to Egypt,
ACTS|7|40|saying to Aaron, 'Make for us gods who will go before us. As for this Moses who led us out from the land of Egypt, we do not know what has become of him.'
ACTS|7|41|And they made a calf in those days, and offered a sacrifice to the idol and were rejoicing in the works of their hands.
ACTS|7|42|But God turned away and gave them over to worship the host of heaven, as it is written in the book of the prophets: "' Did you bring to me slain beasts and sacrifices, during the forty years in the wilderness, O house of Israel?
ACTS|7|43|You took up the tent of Moloch and the star of your god Rephan, the images that you made to worship; and I will send you into exile beyond Babylon.'
ACTS|7|44|"Our fathers had the tent of witness in the wilderness, just as he who spoke to Moses directed him to make it, according to the pattern that he had seen.
ACTS|7|45|Our fathers in turn brought it in with Joshua when they dispossessed the nations that God drove out before our fathers. So it was until the days of David,
ACTS|7|46|who found favor in the sight of God and asked to find a dwelling place for the God of Jacob.
ACTS|7|47|But it was Solomon who built a house for him.
ACTS|7|48|Yet the Most High does not dwell in houses made by hands, as the prophet says,
ACTS|7|49|"'Heaven is my throne, and the earth is my footstool. What kind of house will you build for me, says the Lord, or what is the place of my rest?
ACTS|7|50|Did not my hand make all these things?'
ACTS|7|51|"You stiff-necked people, uncircumcised in heart and ears, you always resist the Holy Spirit. As your fathers did, so do you.
ACTS|7|52|Which of the prophets did not your fathers persecute? And they killed those who announced beforehand the coming of the Righteous One, whom you have now betrayed and murdered,
ACTS|7|53|you who received the law as delivered by angels and did not keep it."
ACTS|7|54|Now when they heard these things they were enraged, and they ground their teeth at him.
ACTS|7|55|But he, full of the Holy Spirit, gazed into heaven and saw the glory of God, and Jesus standing at the right hand of God.
ACTS|7|56|And he said, "Behold, I see the heavens opened, and the Son of Man standing at the right hand of God."
ACTS|7|57|But they cried out with a loud voice and stopped their ears and rushed together at him.
ACTS|7|58|Then they cast him out of the city and stoned him. And the witnesses laid down their garments at the feet of a young man named Saul.
ACTS|7|59|And as they were stoning Stephen, he called out, "Lord Jesus, receive my spirit."
ACTS|7|60|And falling to his knees he cried out with a loud voice, "Lord, do not hold this sin against them." And when he had said this, he fell asleep.
ACTS|8|1|And Saul approved of his execution. And there arose on that day a great persecution against the church in Jerusalem, and they were all scattered throughout the regions of Judea and Samaria, except the apostles.
ACTS|8|2|Devout men buried Stephen and made great lamentation over him.
ACTS|8|3|But Saul was ravaging the church, and entering house after house, he dragged off men and women and committed them to prison.
ACTS|8|4|Now those who were scattered went about preaching the word.
ACTS|8|5|Philip went down to the city of Samaria and proclaimed to them the Christ.
ACTS|8|6|And the crowds with one accord paid attention to what was being said by Philip when they heard him and saw the signs that he did.
ACTS|8|7|For unclean spirits came out of many who were possessed, crying with a loud voice, and many who were paralyzed or lame were healed.
ACTS|8|8|So there was much joy in that city.
ACTS|8|9|But there was a man named Simon, who had previously practiced magic in the city and amazed the people of Samaria, saying that he himself was somebody great.
ACTS|8|10|They all paid attention to him, from the least to the greatest, saying, "This man is the power of God that is called Great."
ACTS|8|11|And they paid attention to him because for a long time he had amazed them with his magic.
ACTS|8|12|But when they believed Philip as he preached good news about the kingdom of God and the name of Jesus Christ, they were baptized, both men and women.
ACTS|8|13|Even Simon himself believed, and after being baptized he continued with Philip. And seeing signs and great miracles performed, he was amazed.
ACTS|8|14|Now when the apostles at Jerusalem heard that Samaria had received the word of God, they sent to them Peter and John,
ACTS|8|15|who came down and prayed for them that they might receive the Holy Spirit,
ACTS|8|16|for he had not yet fallen on any of them, but they had only been baptized in the name of the Lord Jesus.
ACTS|8|17|Then they laid their hands on them and they received the Holy Spirit.
ACTS|8|18|Now when Simon saw that the Spirit was given through the laying on of the apostles' hands, he offered them money,
ACTS|8|19|saying, "Give me this power also, so that anyone on whom I lay my hands may receive the Holy Spirit."
ACTS|8|20|But Peter said to him, "May your silver perish with you, because you thought you could obtain the gift of God with money!
ACTS|8|21|You have neither part nor lot in this matter, for your heart is not right before God.
ACTS|8|22|Repent, therefore, of this wickedness of yours, and pray to the Lord that, if possible, the intent of your heart may be forgiven you.
ACTS|8|23|For I see that you are in the gall of bitterness and in the bond of iniquity."
ACTS|8|24|And Simon answered, "Pray for me to the Lord, that nothing of what you have said may come upon me."
ACTS|8|25|Now when they had testified and spoken the word of the Lord, they returned to Jerusalem, preaching the gospel to many villages of the Samaritans.
ACTS|8|26|Now an angel of the Lord said to Philip, "Rise and go toward the south to the road that goes down from Jerusalem to Gaza." This is a desert place.
ACTS|8|27|And he rose and went. And there was an Ethiopian, a eunuch, a court official of Candace, queen of the Ethiopians, who was in charge of all her treasure. He had come to Jerusalem to worship
ACTS|8|28|and was returning, seated in his chariot, and he was reading the prophet Isaiah.
ACTS|8|29|And the Spirit said to Philip, "Go over and join this chariot."
ACTS|8|30|So Philip ran to him and heard him reading Isaiah the prophet and asked, "Do you understand what you are reading?"
ACTS|8|31|And he said, "How can I, unless someone guides me?" And he invited Philip to come up and sit with him.
ACTS|8|32|Now the passage of the Scripture that he was reading was this: "Like a sheep he was led to the slaughter and like a lamb before its shearer is silent, so he opens not his mouth.
ACTS|8|33|In his humiliation justice was denied him. Who can describe his generation? For his life is taken away from the earth."
ACTS|8|34|And the eunuch said to Philip, "About whom, I ask you, does the prophet say this, about himself or about someone else?"
ACTS|8|35|Then Philip opened his mouth, and beginning with this Scripture he told him the good news about Jesus.
ACTS|8|36|And as they were going along the road they came to some water, and the eunuch said, "See, here is water! What prevents me from being baptized?"
ACTS|8|37|***
ACTS|8|38|And he commanded the chariot to stop, and they both went down into the water, Philip and the eunuch, and he baptized him.
ACTS|8|39|And when they came up out of the water, the Spirit of the Lord carried Philip away, and the eunuch saw him no more, and went on his way rejoicing.
ACTS|8|40|But Philip found himself at Azotus, and as he passed through he preached the gospel to all the towns until he came to Caesarea.
ACTS|9|1|But Saul, still breathing threats and murder against the disciples of the Lord, went to the high priest
ACTS|9|2|and asked him for letters to the synagogues at Damascus, so that if he found any belonging to the Way, men or women, he might bring them bound to Jerusalem.
ACTS|9|3|Now as he went on his way, he approached Damascus, and suddenly a light from heaven flashed around him.
ACTS|9|4|And falling to the ground he heard a voice saying to him, "Saul, Saul, why are you persecuting me?"
ACTS|9|5|And he said, "Who are you, Lord?" And he said, "I am Jesus, whom you are persecuting.
ACTS|9|6|But rise and enter the city, and you will be told what you are to do."
ACTS|9|7|The men who were traveling with him stood speechless, hearing the voice but seeing no one.
ACTS|9|8|Saul rose from the ground, and although his eyes were opened, he saw nothing. So they led him by the hand and brought him into Damascus.
ACTS|9|9|And for three days he was without sight, and neither ate nor drank.
ACTS|9|10|Now there was a disciple at Damascus named Ananias. The Lord said to him in a vision, "Ananias." And he said, "Here I am, Lord."
ACTS|9|11|And the Lord said to him, "Rise and go to the street called Straight, and at the house of Judas look for a man of Tarsus named Saul, for behold, he is praying,
ACTS|9|12|and he has seen in a vision a man named Ananias come in and lay his hands on him so that he might regain his sight."
ACTS|9|13|But Ananias answered, "Lord, I have heard from many about this man, how much evil he has done to your saints at Jerusalem.
ACTS|9|14|And here he has authority from the chief priests to bind all who call on your name."
ACTS|9|15|But the Lord said to him, "Go, for he is a chosen instrument of mine to carry my name before the Gentiles and kings and the children of Israel.
ACTS|9|16|For I will show him how much he must suffer for the sake of my name."
ACTS|9|17|So Ananias departed and entered the house. And laying his hands on him he said, "Brother Saul, the Lord Jesus who appeared to you on the road by which you came has sent me so that you may regain your sight and be filled with the Holy Spirit."
ACTS|9|18|And immediately something like scales fell from his eyes, and he regained his sight. Then he rose and was baptized;
ACTS|9|19|and taking food, he was strengthened. For some days he was with the disciples at Damascus.
ACTS|9|20|And immediately he proclaimed Jesus in the synagogues, saying, "He is the Son of God."
ACTS|9|21|And all who heard him were amazed and said, "Is not this the man who made havoc in Jerusalem of those who called upon this name? And has he not come here for this purpose, to bring them bound before the chief priests?"
ACTS|9|22|But Saul increased all the more in strength, and confounded the Jews who lived in Damascus by proving that Jesus was the Christ.
ACTS|9|23|When many days had passed, the Jews plotted to kill him,
ACTS|9|24|but their plot became known to Saul. They were watching the gates day and night in order to kill him,
ACTS|9|25|but his disciples took him by night and let him down through an opening in the wall, lowering him in a basket.
ACTS|9|26|And when he had come to Jerusalem, he attempted to join the disciples. And they were all afraid of him, for they did not believe that he was a disciple.
ACTS|9|27|But Barnabas took him and brought him to the apostles and declared to them how on the road he had seen the Lord, who spoke to him, and how at Damascus he had preached boldly in the name of Jesus.
ACTS|9|28|So he went in and out among them at Jerusalem, preaching boldly in the name of the Lord.
ACTS|9|29|And he spoke and disputed against the Hellenists. But they were seeking to kill him.
ACTS|9|30|And when the brothers learned this, they brought him down to Caesarea and sent him off to Tarsus.
ACTS|9|31|So the church throughout all Judea and Galilee and Samaria had peace and was being built up. And walking in the fear of the Lord and in the comfort of the Holy Spirit, it multiplied.
ACTS|9|32|Now as Peter went here and there among them all, he came down also to the saints who lived at Lydda.
ACTS|9|33|There he found a man named Aeneas, bedridden for eight years, who was paralyzed.
ACTS|9|34|And Peter said to him, "Aeneas, Jesus Christ heals you; rise and make your bed." And immediately he rose.
ACTS|9|35|And all the residents of Lydda and Sharon saw him, and they turned to the Lord.
ACTS|9|36|Now there was in Joppa a disciple named Tabitha, which, translated, means Dorcas. She was full of good works and acts of charity.
ACTS|9|37|In those days she became ill and died, and when they had washed her, they laid her in an upper room.
ACTS|9|38|Since Lydda was near Joppa, the disciples, hearing that Peter was there, sent two men to him, urging him, "Please come to us without delay."
ACTS|9|39|So Peter rose and went with them. And when he arrived, they took him to the upper room. All the widows stood beside him weeping and showing tunics and other garments that Dorcas made while she was with them.
ACTS|9|40|But Peter put them all outside, and knelt down and prayed; and turning to the body he said, "Tabitha, arise." And she opened her eyes, and when she saw Peter she sat up.
ACTS|9|41|And he gave her his hand and raised her up. Then calling the saints and widows, he presented her alive.
ACTS|9|42|And it became known throughout all Joppa, and many believed in the Lord.
ACTS|9|43|And he stayed in Joppa for many days with one Simon, a tanner.
ACTS|10|1|At Caesarea there was a man named Cornelius, a centurion of what was known as the Italian Cohort,
ACTS|10|2|a devout man who feared God with all his household, gave alms generously to the people, and prayed continually to God.
ACTS|10|3|About the ninth hour of the day he saw clearly in a vision an angel of God come in and say to him, "Cornelius."
ACTS|10|4|And he stared at him in terror and said, "What is it, Lord?" And he said to him, "Your prayers and your alms have ascended as a memorial before God.
ACTS|10|5|And now send men to Joppa and bring one Simon who is called Peter.
ACTS|10|6|He is lodging with one Simon, a tanner, whose house is by the seaside."
ACTS|10|7|When the angel who spoke to him had departed, he called two of his servants and a devout soldier from among those who attended him,
ACTS|10|8|and having related everything to them, he sent them to Joppa.
ACTS|10|9|The next day, as they were on their journey and approaching the city, Peter went up on the housetop about the sixth hour to pray.
ACTS|10|10|And he became hungry and wanted something to eat, but while they were preparing it, he fell into a trance
ACTS|10|11|and saw the heavens opened and something like a great sheet descending, being let down by its four corners upon the earth.
ACTS|10|12|In it were all kinds of animals and reptiles and birds of the air.
ACTS|10|13|And there came a voice to him: "Rise, Peter; kill and eat."
ACTS|10|14|But Peter said, "By no means, Lord; for I have never eaten anything that is common or unclean."
ACTS|10|15|And the voice came to him again a second time, "What God has made clean, do not call common."
ACTS|10|16|This happened three times, and the thing was taken up at once to heaven.
ACTS|10|17|Now while Peter was inwardly perplexed as to what the vision that he had seen might mean, behold, the men who were sent by Cornelius, having made inquiry for Simon's house, stood at the gate
ACTS|10|18|and called out to ask whether Simon who was called Peter was lodging there.
ACTS|10|19|And while Peter was pondering the vision, the Spirit said to him, "Behold, three men are looking for you.
ACTS|10|20|Rise and go down and accompany them without hesitation, for I have sent them."
ACTS|10|21|And Peter went down to the men and said, "I am the one you are looking for. What is the reason for your coming?"
ACTS|10|22|And they said, "Cornelius, a centurion, an upright and God-fearing man, who is well spoken of by the whole Jewish nation, was directed by a holy angel to send for you to come to his house and to hear what you have to say."
ACTS|10|23|So he invited them in to be his guests. The next day he rose and went away with them, and some of the brothers from Joppa accompanied him.
ACTS|10|24|And on the following day they entered Caesarea. Cornelius was expecting them and had called together his relatives and close friends.
ACTS|10|25|When Peter entered, Cornelius met him and fell down at his feet and worshiped him.
ACTS|10|26|But Peter lifted him up, saying, "Stand up; I too am a man."
ACTS|10|27|And as he talked with him, he went in and found many persons gathered.
ACTS|10|28|And he said to them, "You yourselves know how unlawful it is for a Jew to associate with or to visit anyone of another nation, but God has shown me that I should not call any person common or unclean.
ACTS|10|29|So when I was sent for, I came without objection. I ask then why you sent for me."
ACTS|10|30|And Cornelius said, "Four days ago, about this hour, I was praying in my house at the ninth hour, and behold, a man stood before me in bright clothing
ACTS|10|31|and said, 'Cornelius, your prayer has been heard and your alms have been remembered before God.
ACTS|10|32|Send therefore to Joppa and ask for Simon who is called Peter. He is lodging in the house of Simon, a tanner, by the sea.'
ACTS|10|33|So I sent for you at once, and you have been kind enough to come. Now therefore we are all here in the presence of God to hear all that you have been commanded by the Lord."
ACTS|10|34|So Peter opened his mouth and said: "Truly I understand that God shows no partiality,
ACTS|10|35|but in every nation anyone who fears him and does what is right is acceptable to him.
ACTS|10|36|As for the word that he sent to Israel, preaching good news of peace through Jesus Christ (he is Lord of all),
ACTS|10|37|you yourselves know what happened throughout all Judea, beginning from Galilee after the baptism that John proclaimed:
ACTS|10|38|how God anointed Jesus of Nazareth with the Holy Spirit and with power. He went about doing good and healing all who were oppressed by the devil, for God was with him.
ACTS|10|39|And we are witnesses of all that he did both in the country of the Jews and in Jerusalem. They put him to death by hanging him on a tree,
ACTS|10|40|but God raised him on the third day and made him to appear,
ACTS|10|41|not to all the people but to us who had been chosen by God as witnesses, who ate and drank with him after he rose from the dead.
ACTS|10|42|And he commanded us to preach to the people and to testify that he is the one appointed by God to be judge of the living and the dead.
ACTS|10|43|To him all the prophets bear witness that everyone who believes in him receives forgiveness of sins through his name."
ACTS|10|44|While Peter was still saying these things, the Holy Spirit fell on all who heard the word.
ACTS|10|45|And the believers from among the circumcised who had come with Peter were amazed, because the gift of the Holy Spirit was poured out even on the Gentiles.
ACTS|10|46|For they were hearing them speaking in tongues and extolling God. Then Peter declared,
ACTS|10|47|"Can anyone withhold water for baptizing these people, who have received the Holy Spirit just as we have?"
ACTS|10|48|And he commanded them to be baptized in the name of Jesus Christ. Then they asked him to remain for some days.
ACTS|11|1|Now the apostles and the brothers who were throughout Judea heard that the Gentiles also had received the word of God.
ACTS|11|2|So when Peter went up to Jerusalem, the circumcision party criticized him, saying,
ACTS|11|3|"You went to uncircumcised men and ate with them."
ACTS|11|4|But Peter began and explained it to them in order:
ACTS|11|5|"I was in the city of Joppa praying, and in a trance I saw a vision, something like a great sheet descending, being let down from heaven by its four corners, and it came down to me.
ACTS|11|6|Looking at it closely, I observed animals and beasts of prey and reptiles and birds of the air.
ACTS|11|7|And I heard a voice saying to me, 'Rise, Peter; kill and eat.'
ACTS|11|8|But I said, 'By no means, Lord; for nothing common or unclean has ever entered my mouth.'
ACTS|11|9|But the voice answered a second time from heaven, 'What God has made clean, do not call common.'
ACTS|11|10|This happened three times, and all was drawn up again into heaven.
ACTS|11|11|And behold, at that very moment three men arrived at the house in which we were, sent to me from Caesarea.
ACTS|11|12|And the Spirit told me to go with them, making no distinction. These six brothers also accompanied me, and we entered the man's house.
ACTS|11|13|And he told us how he had seen the angel stand in his house and say, 'Send to Joppa and bring Simon who is called Peter;
ACTS|11|14|he will declare to you a message by which you will be saved, you and all your household.'
ACTS|11|15|As I began to speak, the Holy Spirit fell on them just as on us at the beginning.
ACTS|11|16|And I remembered the word of the Lord, how he said, 'John baptized with water, but you will be baptized with the Holy Spirit.'
ACTS|11|17|If then God gave the same gift to them as he gave to us when we believed in the Lord Jesus Christ, who was I that I could stand in God's way?"
ACTS|11|18|When they heard these things they fell silent. And they glorified God, saying, "Then to the Gentiles also God has granted repentance that leads to life."
ACTS|11|19|Now those who were scattered because of the persecution that arose over Stephen traveled as far as Phoenicia and Cyprus and Antioch, speaking the word to no one except Jews.
ACTS|11|20|But there were some of them, men of Cyprus and Cyrene, who on coming to Antioch spoke to the Hellenists also, preaching the Lord Jesus.
ACTS|11|21|And the hand of the Lord was with them, and a great number who believed turned to the Lord.
ACTS|11|22|The report of this came to the ears of the church in Jerusalem, and they sent Barnabas to Antioch.
ACTS|11|23|When he came and saw the grace of God, he was glad, and he exhorted them all to remain faithful to the Lord with steadfast purpose,
ACTS|11|24|for he was a good man, full of the Holy Spirit and of faith. And a great many people were added to the Lord.
ACTS|11|25|So Barnabas went to Tarsus to look for Saul,
ACTS|11|26|and when he had found him, he brought him to Antioch. For a whole year they met with the church and taught a great many people. And in Antioch the disciples were first called Christians.
ACTS|11|27|Now in these days prophets came down from Jerusalem to Antioch.
ACTS|11|28|And one of them named Agabus stood up and foretold by the Spirit that there would be a great famine over all the world (this took place in the days of Claudius).
ACTS|11|29|So the disciples determined, everyone according to his ability, to send relief to the brothers living in Judea.
ACTS|11|30|And they did so, sending it to the elders by the hand of Barnabas and Saul.
ACTS|12|1|About that time Herod the king laid violent hands on some who belonged to the church.
ACTS|12|2|He killed James the brother of John with the sword,
ACTS|12|3|and when he saw that it pleased the Jews, he proceeded to arrest Peter also. This was during the days of Unleavened Bread.
ACTS|12|4|And when he had seized him, he put him in prison, delivering him over to four squads of soldiers to guard him, intending after the Passover to bring him out to the people.
ACTS|12|5|So Peter was kept in prison, but earnest prayer for him was made to God by the church.
ACTS|12|6|Now when Herod was about to bring him out, on that very night, Peter was sleeping between two soldiers, bound with two chains, and sentries before the door were guarding the prison.
ACTS|12|7|And behold, an angel of the Lord stood next to him, and a light shone in the cell. He struck Peter on the side and woke him, saying, "Get up quickly." And the chains fell off his hands.
ACTS|12|8|And the angel said to him, "Dress yourself and put on your sandals." And he did so. And he said to him, "Wrap your cloak around you and follow me."
ACTS|12|9|And he went out and followed him. He did not know that what was being done by the angel was real, but thought he was seeing a vision.
ACTS|12|10|When they had passed the first and the second guard, they came to the iron gate leading into the city. It opened for them of its own accord, and they went out and went along one street, and immediately the angel left him.
ACTS|12|11|When Peter came to himself, he said, "Now I am sure that the Lord has sent his angel and rescued me from the hand of Herod and from all that the Jewish people were expecting."
ACTS|12|12|When he realized this, he went to the house of Mary, the mother of John whose other name was Mark, where many were gathered together and were praying.
ACTS|12|13|And when he knocked at the door of the gateway, a servant girl named Rhoda came to answer.
ACTS|12|14|Recognizing Peter's voice, in her joy she did not open the gate but ran in and reported that Peter was standing at the gate.
ACTS|12|15|They said to her, "You are out of your mind." But she kept insisting that it was so, and they kept saying, "It is his angel!"
ACTS|12|16|But Peter continued knocking, and when they opened, they saw him and were amazed.
ACTS|12|17|But motioning to them with his hand to be silent, he described to them how the Lord had brought him out of the prison. And he said, "Tell these things to James and to the brothers." Then he departed and went to another place.
ACTS|12|18|Now when day came, there was no little disturbance among the soldiers over what had become of Peter.
ACTS|12|19|And after Herod searched for him and did not find him, he examined the sentries and ordered that they should be put to death. Then he went down from Judea to Caesarea and spent time there.
ACTS|12|20|Now Herod was angry with the people of Tyre and Sidon, and they came to him with one accord, and having persuaded Blastus, the king's chamberlain, they asked for peace, because their country depended on the king's country for food.
ACTS|12|21|On an appointed day Herod put on his royal robes, took his seat upon the throne, and delivered an oration to them.
ACTS|12|22|And the people were shouting, "The voice of a god, and not of a man!"
ACTS|12|23|Immediately an angel of the Lord struck him down, because he did not give God the glory, and he was eaten by worms and breathed his last.
ACTS|12|24|But the word of God increased and multiplied.
ACTS|12|25|And Barnabas and Saul returned from Jerusalem when they had completed their service, bringing with them John, whose other name was Mark.
ACTS|13|1|Now there were in the church at Antioch prophets and teachers, Barnabas, Simeon who was called Niger, Lucius of Cyrene, Manaen a member of the court of Herod the tetrarch, and Saul.
ACTS|13|2|While they were worshiping the Lord and fasting, the Holy Spirit said, "Set apart for me Barnabas and Saul for the work to which I have called them."
ACTS|13|3|Then after fasting and praying they laid their hands on them and sent them off.
ACTS|13|4|So, being sent out by the Holy Spirit, they went down to Seleucia, and from there they sailed to Cyprus.
ACTS|13|5|When they arrived at Salamis, they proclaimed the word of God in the synagogues of the Jews. And they had John to assist them.
ACTS|13|6|When they had gone through the whole island as far as Paphos, they came upon a certain magician, a Jewish false prophet named Bar-Jesus.
ACTS|13|7|He was with the proconsul, Sergius Paulus, a man of intelligence, who summoned Barnabas and Saul and sought to hear the word of God.
ACTS|13|8|But Elymas the magician (for that is the meaning of his name) opposed them, seeking to turn the proconsul away from the faith.
ACTS|13|9|But Saul, who was also called Paul, filled with the Holy Spirit, looked intently at him
ACTS|13|10|and said, "You son of the devil, you enemy of all righteousness, full of all deceit and villainy, will you not stop making crooked the straight paths of the Lord?
ACTS|13|11|And now, behold, the hand of the Lord is upon you, and you will be blind and unable to see the sun for a time." Immediately mist and darkness fell upon him, and he went about seeking people to lead him by the hand.
ACTS|13|12|Then the proconsul believed, when he saw what had occurred, for he was astonished at the teaching of the Lord.
ACTS|13|13|Now Paul and his companions set sail from Paphos and came to Perga in Pamphylia. And John left them and returned to Jerusalem,
ACTS|13|14|but they went on from Perga and came to Antioch in Pisidia. And on the Sabbath day they went into the synagogue and sat down.
ACTS|13|15|After the reading from the Law and the Prophets, the rulers of the synagogue sent a message to them, saying, "Brothers, if you have any word of exhortation for the people, say it."
ACTS|13|16|So Paul stood up, and motioning with his hand said: "Men of Israel and you who fear God, listen.
ACTS|13|17|The God of this people Israel chose our fathers and made the people great during their stay in the land of Egypt, and with uplifted arm he led them out of it.
ACTS|13|18|And for about forty years he put up with them in the wilderness.
ACTS|13|19|And after destroying seven nations in the land of Canaan, he gave them their land as an inheritance.
ACTS|13|20|All this took about 450 years. And after that he gave them judges until Samuel the prophet.
ACTS|13|21|Then they asked for a king, and God gave them Saul the son of Kish, a man of the tribe of Benjamin, for forty years.
ACTS|13|22|And when he had removed him, he raised up David to be their king, of whom he testified and said, 'I have found in David the son of Jesse a man after my heart, who will do all my will.'
ACTS|13|23|Of this man's offspring God has brought to Israel a Savior, Jesus, as he promised.
ACTS|13|24|Before his coming, John had proclaimed a baptism of repentance to all the people of Israel.
ACTS|13|25|And as John was finishing his course, he said, 'What do you suppose that I am? I am not he. No, but behold, after me one is coming, the sandals of whose feet I am not worthy to untie.'
ACTS|13|26|"Brothers, sons of the family of Abraham, and those among you who fear God, to us has been sent the message of this salvation.
ACTS|13|27|For those who live in Jerusalem and their rulers, because they did not recognize him nor understand the utterances of the prophets, which are read every Sabbath, fulfilled them by condemning him.
ACTS|13|28|And though they found in him no guilt worthy of death, they asked Pilate to have him executed.
ACTS|13|29|And when they had carried out all that was written of him, they took him down from the tree and laid him in a tomb.
ACTS|13|30|But God raised him from the dead,
ACTS|13|31|and for many days he appeared to those who had come up with him from Galilee to Jerusalem, who are now his witnesses to the people.
ACTS|13|32|And we bring you the good news that what God promised to the fathers,
ACTS|13|33|this he has fulfilled to us their children by raising Jesus, as also it is written in the second Psalm, "' You are my Son, today I have begotten you.'
ACTS|13|34|And as for the fact that he raised him from the dead, no more to return to corruption, he has spoken in this way, "' I will give you the holy and sure blessings of David.'
ACTS|13|35|Therefore he says also in another psalm, "' You will not let your Holy One see corruption.'
ACTS|13|36|For David, after he had served the purpose of God in his own generation, fell asleep and was laid with his fathers and saw corruption,
ACTS|13|37|but he whom God raised up did not see corruption.
ACTS|13|38|Let it be known to you therefore, brothers, that through this man forgiveness of sins is proclaimed to you, and by him everyone who believes is freed from everything
ACTS|13|39|from which you could not be freed by the law of Moses.
ACTS|13|40|Beware, therefore, lest what is said in the Prophets should come about:
ACTS|13|41|"'Look, you scoffers, be astounded and perish; for I am doing a work in your days, a work that you will not believe, even if one tells it to you.'"
ACTS|13|42|As they went out, the people begged that these things might be told them the next Sabbath.
ACTS|13|43|And after the meeting of the synagogue broke up, many Jews and devout converts to Judaism followed Paul and Barnabas, who, as they spoke with them, urged them to continue in the grace of God.
ACTS|13|44|The next Sabbath almost the whole city gathered to hear the word of the Lord.
ACTS|13|45|But when the Jews saw the crowds, they were filled with jealousy and began to contradict what was spoken by Paul, reviling him.
ACTS|13|46|And Paul and Barnabas spoke out boldly, saying, "It was necessary that the word of God be spoken first to you. Since you thrust it aside and judge yourselves unworthy of eternal life, behold, we are turning to the Gentiles.
ACTS|13|47|For so the Lord has commanded us, saying, "' I have made you a light for the Gentiles, that you may bring salvation to the ends of the earth.'"
ACTS|13|48|And when the Gentiles heard this, they began rejoicing and glorifying the word of the Lord, and as many as were appointed to eternal life believed.
ACTS|13|49|And the word of the Lord was spreading throughout the whole region.
ACTS|13|50|But the Jews incited the devout women of high standing and the leading men of the city, stirred up persecution against Paul and Barnabas, and drove them out of their district.
ACTS|13|51|But they shook off the dust from their feet against them and went to Iconium.
ACTS|13|52|And the disciples were filled with joy and with the Holy Spirit.
ACTS|14|1|Now at Iconium they entered together into the Jewish synagogue and spoke in such a way that a great number of both Jews and Greeks believed.
ACTS|14|2|But the unbelieving Jews stirred up the Gentiles and poisoned their minds against the brothers.
ACTS|14|3|So they remained for a long time, speaking boldly for the Lord, who bore witness to the word of his grace, granting signs and wonders to be done by their hands.
ACTS|14|4|But the people of the city were divided; some sided with the Jews and some with the apostles.
ACTS|14|5|When an attempt was made by both Gentiles and Jews, with their rulers, to mistreat them and to stone them,
ACTS|14|6|they learned of it and fled to Lystra and Derbe, cities of Lycaonia, and to the surrounding country,
ACTS|14|7|and there they continued to preach the gospel.
ACTS|14|8|Now at Lystra there was a man sitting who could not use his feet. He was crippled from birth and had never walked.
ACTS|14|9|He listened to Paul speaking. And Paul, looking intently at him and seeing that he had faith to be made well,
ACTS|14|10|said in a loud voice, "Stand upright on your feet." And he sprang up and began walking.
ACTS|14|11|And when the crowds saw what Paul had done, they lifted up their voices, saying in Lycaonian, "The gods have come down to us in the likeness of men!"
ACTS|14|12|Barnabas they called Zeus, and Paul, Hermes, because he was the chief speaker.
ACTS|14|13|And the priest of Zeus, whose temple was at the entrance to the city, brought oxen and garlands to the gates and wanted to offer sacrifice with the crowds.
ACTS|14|14|But when the apostles Barnabas and Paul heard of it, they tore their garments and rushed out into the crowd, crying out,
ACTS|14|15|"Men, why are you doing these things? We also are men, of like nature with you, and we bring you good news, that you should turn from these vain things to a living God, who made the heaven and the earth and the sea and all that is in them.
ACTS|14|16|In past generations he allowed all the nations to walk in their own ways.
ACTS|14|17|Yet he did not leave himself without witness, for he did good by giving you rains from heaven and fruitful seasons, satisfying your hearts with food and gladness."
ACTS|14|18|Even with these words they scarcely restrained the people from offering sacrifice to them.
ACTS|14|19|But Jews came from Antioch and Iconium, and having persuaded the crowds, they stoned Paul and dragged him out of the city, supposing that he was dead.
ACTS|14|20|But when the disciples gathered about him, he rose up and entered the city, and on the next day he went on with Barnabas to Derbe.
ACTS|14|21|When they had preached the gospel to that city and had made many disciples, they returned to Lystra and to Iconium and to Antioch,
ACTS|14|22|strengthening the souls of the disciples, encouraging them to continue in the faith, and saying that through many tribulations we must enter the kingdom of God.
ACTS|14|23|And when they had appointed elders for them in every church, with prayer and fasting they committed them to the Lord in whom they had believed.
ACTS|14|24|Then they passed through Pisidia and came to Pamphylia.
ACTS|14|25|And when they had spoken the word in Perga, they went down to Attalia,
ACTS|14|26|and from there they sailed to Antioch, where they had been commended to the grace of God for the work that they had fulfilled.
ACTS|14|27|And when they arrived and gathered the church together, they declared all that God had done with them, and how he had opened a door of faith to the Gentiles.
ACTS|14|28|And they remained no little time with the disciples.
ACTS|15|1|But some men came down from Judea and were teaching the brothers, "Unless you are circumcised according to the custom of Moses, you cannot be saved."
ACTS|15|2|And after Paul and Barnabas had no small dissension and debate with them, Paul and Barnabas and some of the others were appointed to go up to Jerusalem to the apostles and the elders about this question.
ACTS|15|3|So, being sent on their way by the church, they passed through both Phoenicia and Samaria, describing in detail the conversion of the Gentiles, and brought great joy to all the brothers.
ACTS|15|4|When they came to Jerusalem, they were welcomed by the church and the apostles and the elders, and they declared all that God had done with them.
ACTS|15|5|But some believers who belonged to the party of the Pharisees rose up and said, "It is necessary to circumcise them and to order them to keep the law of Moses."
ACTS|15|6|The apostles and the elders were gathered together to consider this matter.
ACTS|15|7|And after there had been much debate, Peter stood up and said to them, "Brothers, you know that in the early days God made a choice among you, that by my mouth the Gentiles should hear the word of the gospel and believe.
ACTS|15|8|And God, who knows the heart, bore witness to them, by giving them the Holy Spirit just as he did to us,
ACTS|15|9|and he made no distinction between us and them, having cleansed their hearts by faith.
ACTS|15|10|Now, therefore, why are you putting God to the test by placing a yoke on the neck of the disciples that neither our fathers nor we have been able to bear?
ACTS|15|11|But we believe that we will be saved through the grace of the Lord Jesus, just as they will."
ACTS|15|12|And all the assembly fell silent, and they listened to Barnabas and Paul as they related what signs and wonders God had done through them among the Gentiles.
ACTS|15|13|After they finished speaking, James replied, "Brothers, listen to me.
ACTS|15|14|Simeon has related how God first visited the Gentiles, to take from them a people for his name.
ACTS|15|15|And with this the words of the prophets agree, just as it is written,
ACTS|15|16|"'After this I will return, and I will rebuild the tent of David that has fallen; I will rebuild its ruins, and I will restore it,
ACTS|15|17|that the remnant of mankind may seek the Lord, and all the Gentiles who are called by my name, says the Lord, who makes these things
ACTS|15|18|known from of old.'
ACTS|15|19|Therefore my judgment is that we should not trouble those of the Gentiles who turn to God,
ACTS|15|20|but should write to them to abstain from the things polluted by idols, and from sexual immorality, and from what has been strangled, and from blood.
ACTS|15|21|For from ancient generations Moses has had in every city those who proclaim him, for he is read every Sabbath in the synagogues."
ACTS|15|22|Then it seemed good to the apostles and the elders, with the whole church, to choose men from among them and send them to Antioch with Paul and Barnabas. They sent Judas called Barsabbas, and Silas, leading men among the brothers,
ACTS|15|23|with the following letter: "The brothers, both the apostles and the elders, to the brothers who are of the Gentiles in Antioch and Syria and Cilicia, greetings.
ACTS|15|24|Since we have heard that some persons have gone out from us and troubled you with words, unsettling your minds, although we gave them no instructions,
ACTS|15|25|it has seemed good to us, having come to one accord, to choose men and send them to you with our beloved Barnabas and Paul,
ACTS|15|26|men who have risked their lives for the sake of our Lord Jesus Christ.
ACTS|15|27|We have therefore sent Judas and Silas, who themselves will tell you the same things by word of mouth.
ACTS|15|28|For it has seemed good to the Holy Spirit and to us to lay on you no greater burden than these requirements:
ACTS|15|29|that you abstain from what has been sacrificed to idols, and from blood, and from what has been strangled, and from sexual immorality. If you keep yourselves from these, you will do well. Farewell."
ACTS|15|30|So when they were sent off, they went down to Antioch, and having gathered the congregation together, they delivered the letter.
ACTS|15|31|And when they had read it, they rejoiced because of its encouragement.
ACTS|15|32|And Judas and Silas, who were themselves prophets, encouraged and strengthened the brothers with many words.
ACTS|15|33|And after they had spent some time, they were sent off in peace by the brothers to those who had sent them.
ACTS|15|34|***
ACTS|15|35|But Paul and Barnabas remained in Antioch, teaching and preaching the word of the Lord, with many others also.
ACTS|15|36|And after some days Paul said to Barnabas, "Let us return and visit the brothers in every city where we proclaimed the word of the Lord, and see how they are."
ACTS|15|37|Now Barnabas wanted to take with them John called Mark.
ACTS|15|38|But Paul thought best not to take with them one who had withdrawn from them in Pamphylia and had not gone with them to the work.
ACTS|15|39|And there arose a sharp disagreement, so that they separated from each other. Barnabas took Mark with him and sailed away to Cyprus,
ACTS|15|40|but Paul chose Silas and departed, having been commended by the brothers to the grace of the Lord.
ACTS|15|41|And he went through Syria and Cilicia, strengthening the churches.
ACTS|16|1|Paul came also to Derbe and to Lystra. A disciple was there, named Timothy, the son of a Jewish woman who was a believer, but his father was a Greek.
ACTS|16|2|He was well spoken of by the brothers at Lystra and Iconium.
ACTS|16|3|Paul wanted Timothy to accompany him, and he took him and circumcised him because of the Jews who were in those places, for they all knew that his father was a Greek.
ACTS|16|4|As they went on their way through the cities, they delivered to them for observance the decisions that had been reached by the apostles and elders who were in Jerusalem.
ACTS|16|5|So the churches were strengthened in the faith, and they increased in numbers daily.
ACTS|16|6|And they went through the region of Phrygia and Galatia, having been forbidden by the Holy Spirit to speak the word in Asia.
ACTS|16|7|And when they had come up to Mysia, they attempted to go into Bithynia, but the Spirit of Jesus did not allow them.
ACTS|16|8|So, passing by Mysia, they went down to Troas.
ACTS|16|9|And a vision appeared to Paul in the night: a man of Macedonia was standing there, urging him and saying, "Come over to Macedonia and help us."
ACTS|16|10|And when Paul had seen the vision, immediately we sought to go on into Macedonia, concluding that God had called us to preach the gospel to them.
ACTS|16|11|So, setting sail from Troas, we made a direct voyage to Samothrace, and the following day to Neapolis,
ACTS|16|12|and from there to Philippi, which is a leading city of the district of Macedonia and a Roman colony. We remained in this city some days.
ACTS|16|13|And on the Sabbath day we went outside the gate to the riverside, where we supposed there was a place of prayer, and we sat down and spoke to the women who had come together.
ACTS|16|14|One who heard us was a woman named Lydia, from the city of Thyatira, a seller of purple goods, who was a worshiper of God. The Lord opened her heart to pay attention to what was said by Paul.
ACTS|16|15|And after she was baptized, and her household as well, she urged us, saying, "If you have judged me to be faithful to the Lord, come to my house and stay." And she prevailed upon us.
ACTS|16|16|As we were going to the place of prayer, we were met by a slave girl who had a spirit of divination and brought her owners much gain by fortune-telling.
ACTS|16|17|She followed Paul and us, crying out, "These men are servants of the Most High God, who proclaim to you the way of salvation."
ACTS|16|18|And this she kept doing for many days. Paul, having become greatly annoyed, turned and said to the spirit, "I command you in the name of Jesus Christ to come out of her." And it came out that very hour.
ACTS|16|19|But when her owners saw that their hope of gain was gone, they seized Paul and Silas and dragged them into the marketplace before the rulers.
ACTS|16|20|And when they had brought them to the magistrates, they said, "These men are Jews, and they are disturbing our city.
ACTS|16|21|They advocate customs that are not lawful for us as Romans to accept or practice."
ACTS|16|22|The crowd joined in attacking them, and the magistrates tore the garments off them and gave orders to beat them with rods.
ACTS|16|23|And when they had inflicted many blows upon them, they threw them into prison, ordering the jailer to keep them safely.
ACTS|16|24|Having received this order, he put them into the inner prison and fastened their feet in the stocks.
ACTS|16|25|About midnight Paul and Silas were praying and singing hymns to God, and the prisoners were listening to them,
ACTS|16|26|and suddenly there was a great earthquake, so that the foundations of the prison were shaken. And immediately all the doors were opened, and everyone's bonds were unfastened.
ACTS|16|27|When the jailer woke and saw that the prison doors were open, he drew his sword and was about to kill himself, supposing that the prisoners had escaped.
ACTS|16|28|But Paul cried with a loud voice, "Do not harm yourself, for we are all here."
ACTS|16|29|And the jailer called for lights and rushed in, and trembling with fear he fell down before Paul and Silas.
ACTS|16|30|Then he brought them out and said, "Sirs, what must I do to be saved?"
ACTS|16|31|And they said, "Believe in the Lord Jesus, and you will be saved, you and your household."
ACTS|16|32|And they spoke the word of the Lord to him and to all who were in his house.
ACTS|16|33|And he took them the same hour of the night and washed their wounds; and he was baptized at once, he and all his family.
ACTS|16|34|Then he brought them up into his house and set food before them. And he rejoiced along with his entire household that he had believed in God.
ACTS|16|35|But when it was day, the magistrates sent the police, saying, "Let those men go."
ACTS|16|36|And the jailer reported these words to Paul, saying, "The magistrates have sent to let you go. Therefore come out now and go in peace."
ACTS|16|37|But Paul said to them, "They have beaten us publicly, uncondemned, men who are Roman citizens, and have thrown us into prison; and do they now throw us out secretly? No! Let them come themselves and take us out."
ACTS|16|38|The police reported these words to the magistrates, and they were afraid when they heard that they were Roman citizens.
ACTS|16|39|So they came and apologized to them. And they took them out and asked them to leave the city.
ACTS|16|40|So they went out of the prison and visited Lydia. And when they had seen the brothers, they encouraged them and departed.
ACTS|17|1|Now when they had passed through Amphipolis and Apollonia, they came to Thessalonica, where there was a synagogue of the Jews.
ACTS|17|2|And Paul went in, as was his custom, and on three Sabbath days he reasoned with them from the Scriptures,
ACTS|17|3|explaining and proving that it was necessary for the Christ to suffer and to rise from the dead, and saying, "This Jesus, whom I proclaim to you, is the Christ."
ACTS|17|4|And some of them were persuaded and joined Paul and Silas, as did a great many of the devout Greeks and not a few of the leading women.
ACTS|17|5|But the Jews were jealous, and taking some wicked men of the rabble, they formed a mob, set the city in an uproar, and attacked the house of Jason, seeking to bring them out to the crowd.
ACTS|17|6|And when they could not find them, they dragged Jason and some of the brothers before the city authorities, shouting, "These men who have turned the world upside down have come here also,
ACTS|17|7|and Jason has received them, and they are all acting against the decrees of Caesar, saying that there is another king, Jesus."
ACTS|17|8|And the people and the city authorities were disturbed when they heard these things.
ACTS|17|9|And when they had taken money as security from Jason and the rest, they let them go.
ACTS|17|10|The brothers immediately sent Paul and Silas away by night to Berea, and when they arrived they went into the Jewish synagogue.
ACTS|17|11|Now these Jews were more noble than those in Thessalonica; they received the word with all eagerness, examining the Scriptures daily to see if these things were so.
ACTS|17|12|Many of them therefore believed, with not a few Greek women of high standing as well as men.
ACTS|17|13|But when the Jews from Thessalonica learned that the word of God was proclaimed by Paul at Berea also, they came there too, agitating and stirring up the crowds.
ACTS|17|14|Then the brothers immediately sent Paul off on his way to the sea, but Silas and Timothy remained there.
ACTS|17|15|Those who conducted Paul brought him as far as Athens, and after receiving a command for Silas and Timothy to come to him as soon as possible, they departed.
ACTS|17|16|Now while Paul was waiting for them at Athens, his spirit was provoked within him as he saw that the city was full of idols.
ACTS|17|17|So he reasoned in the synagogue with the Jews and the devout persons, and in the marketplace every day with those who happened to be there.
ACTS|17|18|Some of the Epicurean and Stoic philosophers also conversed with him. And some said, "What does this babbler wish to say?" Others said, "He seems to be a preacher of foreign divinities"- because he was preaching Jesus and the resurrection.
ACTS|17|19|And they took hold of him and brought him to the Areopagus, saying, "May we know what this new teaching is that you are presenting?
ACTS|17|20|For you bring some strange things to our ears. We wish to know therefore what these things mean."
ACTS|17|21|Now all the Athenians and the foreigners who lived there would spend their time in nothing except telling or hearing something new.
ACTS|17|22|So Paul, standing in the midst of the Areopagus, said: "Men of Athens, I perceive that in every way you are very religious.
ACTS|17|23|For as I passed along and observed the objects of your worship, I found also an altar with this inscription, 'To the unknown god.' What therefore you worship as unknown, this I proclaim to you.
ACTS|17|24|The God who made the world and everything in it, being Lord of heaven and earth, does not live in temples made by man,
ACTS|17|25|nor is he served by human hands, as though he needed anything, since he himself gives to all mankind life and breath and everything.
ACTS|17|26|And he made from one man every nation of mankind to live on all the face of the earth, having determined allotted periods and the boundaries of their dwelling place,
ACTS|17|27|that they should seek God, in the hope that they might feel their way toward him and find him. Yet he is actually not far from each one of us,
ACTS|17|28|for "'In him we live and move and have our being'; as even some of your own poets have said, "' For we are indeed his offspring.'
ACTS|17|29|Being then God's offspring, we ought not to think that the divine being is like gold or silver or stone, an image formed by the art and imagination of man.
ACTS|17|30|The times of ignorance God overlooked, but now he commands all people everywhere to repent,
ACTS|17|31|because he has fixed a day on which he will judge the world in righteousness by a man whom he has appointed; and of this he has given assurance to all by raising him from the dead."
ACTS|17|32|Now when they heard of the resurrection of the dead, some mocked. But others said, "We will hear you again about this."
ACTS|17|33|So Paul went out from their midst.
ACTS|17|34|But some men joined him and believed, among them Dionysius the Areopagite and a woman named Damaris and others with them.
ACTS|18|1|After this Paul left Athens and went to Corinth.
ACTS|18|2|And he found a Jew named Aquila, a native of Pontus, recently come from Italy with his wife Priscilla, because Claudius had commanded all the Jews to leave Rome. And he went to see them,
ACTS|18|3|and because he was of the same trade he stayed with them and worked, for they were tentmakers by trade.
ACTS|18|4|And he reasoned in the synagogue every Sabbath, and tried to persuade Jews and Greeks.
ACTS|18|5|When Silas and Timothy arrived from Macedonia, Paul was occupied with the word, testifying to the Jews that the Christ was Jesus.
ACTS|18|6|And when they opposed and reviled him, he shook out his garments and said to them, "Your blood be on your own heads! I am innocent. From now on I will go to the Gentiles."
ACTS|18|7|And he left there and went to the house of a man named Titius Justus, a worshiper of God. His house was next door to the synagogue.
ACTS|18|8|Crispus, the ruler of the synagogue, believed in the Lord, together with his entire household. And many of the Corinthians hearing Paul believed and were baptized.
ACTS|18|9|And the Lord said to Paul one night in a vision, "Do not be afraid, but go on speaking and do not be silent,
ACTS|18|10|for I am with you, and no one will attack you to harm you, for I have many in this city who are my people."
ACTS|18|11|And he stayed a year and six months, teaching the word of God among them.
ACTS|18|12|But when Gallio was proconsul of Achaia, the Jews made a united attack on Paul and brought him before the tribunal,
ACTS|18|13|saying, "This man is persuading people to worship God contrary to the law."
ACTS|18|14|But when Paul was about to open his mouth, Gallio said to the Jews, "If it were a matter of wrongdoing or vicious crime, O Jews, I would have reason to accept your complaint.
ACTS|18|15|But since it is a matter of questions about words and names and your own law, see to it yourselves. I refuse to be a judge of these things."
ACTS|18|16|And he drove them from the tribunal.
ACTS|18|17|And they all seized Sosthenes, the ruler of the synagogue, and beat him in front of the tribunal. But Gallio paid no attention to any of this.
ACTS|18|18|After this, Paul stayed many days longer and then took leave of the brothers and set sail for Syria, and with him Priscilla and Aquila. At Cenchreae he had cut his hair, for he was under a vow.
ACTS|18|19|And they came to Ephesus, and he left them there, but he himself went into the synagogue and reasoned with the Jews.
ACTS|18|20|When they asked him to stay for a longer period, he declined.
ACTS|18|21|But on taking leave of them he said, "I will return to you if God wills," and he set sail from Ephesus.
ACTS|18|22|When he had landed at Caesarea, he went up and greeted the church, and then went down to Antioch.
ACTS|18|23|After spending some time there, he departed and went from one place to the next through the region of Galatia and Phrygia, strengthening all the disciples.
ACTS|18|24|Now a Jew named Apollos, a native of Alexandria, came to Ephesus. He was an eloquent man, competent in the Scriptures.
ACTS|18|25|He had been instructed in the way of the Lord. And being fervent in spirit, he spoke and taught accurately the things concerning Jesus, though he knew only the baptism of John.
ACTS|18|26|He began to speak boldly in the synagogue, but when Priscilla and Aquila heard him, they took him and explained to him the way of God more accurately.
ACTS|18|27|And when he wished to cross to Achaia, the brothers encouraged him and wrote to the disciples to welcome him. When he arrived, he greatly helped those who through grace had believed,
ACTS|18|28|for he powerfully refuted the Jews in public, showing by the Scriptures that the Christ was Jesus.
ACTS|19|1|And it happened that while Apollos was at Corinth, Paul passed through the inland country and came to Ephesus. There he found some disciples.
ACTS|19|2|And he said to them, "Did you receive the Holy Spirit when you believed?" And they said, "No, we have not even heard that there is a Holy Spirit."
ACTS|19|3|And he said, "Into what then were you baptized?" They said, "Into John's baptism."
ACTS|19|4|And Paul said, "John baptized with the baptism of repentance, telling the people to believe in the one who was to come after him, that is, Jesus."
ACTS|19|5|On hearing this, they were baptized in the name of the Lord Jesus.
ACTS|19|6|And when Paul had laid his hands on them, the Holy Spirit came on them, and they began speaking in tongues and prophesying.
ACTS|19|7|There were about twelve men in all.
ACTS|19|8|And he entered the synagogue and for three months spoke boldly, reasoning and persuading them about the kingdom of God.
ACTS|19|9|But when some became stubborn and continued in unbelief, speaking evil of the Way before the congregation, he withdrew from them and took the disciples with him, reasoning daily in the hall of Tyrannus.
ACTS|19|10|This continued for two years, so that all the residents of Asia heard the word of the Lord, both Jews and Greeks.
ACTS|19|11|And God was doing extraordinary miracles by the hands of Paul,
ACTS|19|12|so that even handkerchiefs or aprons that had touched his skin were carried away to the sick, and their diseases left them and the evil spirits came out of them.
ACTS|19|13|Then some of the itinerant Jewish exorcists undertook to invoke the name of the Lord Jesus over those who had evil spirits, saying, "I adjure you by the Jesus, whom Paul proclaims."
ACTS|19|14|Seven sons of a Jewish high priest named Sceva were doing this.
ACTS|19|15|But the evil spirit answered them, "Jesus I know, and Paul I recognize, but who are you?"
ACTS|19|16|And the man in whom was the evil spirit leaped on them, mastered all of them and overpowered them, so that they fled out of that house naked and wounded.
ACTS|19|17|And this became known to all the residents of Ephesus, both Jews and Greeks. And fear fell upon them all, and the name of the Lord Jesus was extolled.
ACTS|19|18|Also many of those who were now believers came, confessing and divulging their practices.
ACTS|19|19|And a number of those who had practiced magic arts brought their books together and burned them in the sight of all. And they counted the value of them and found it came to fifty thousand pieces of silver.
ACTS|19|20|So the word of the Lord continued to increase and prevail mightily.
ACTS|19|21|Now after these events Paul resolved in the Spirit to pass through Macedonia and Achaia and go to Jerusalem, saying, "After I have been there, I must also see Rome."
ACTS|19|22|And having sent into Macedonia two of his helpers, Timothy and Erastus, he himself stayed in Asia for a while.
ACTS|19|23|About that time there arose no little disturbance concerning the Way.
ACTS|19|24|For a man named Demetrius, a silversmith, who made silver shrines of Artemis, brought no little business to the craftsmen.
ACTS|19|25|These he gathered together, with the workmen in similar trades, and said, "Men, you know that from this business we have our wealth.
ACTS|19|26|And you see and hear that not only in Ephesus but in almost all of Asia this Paul has persuaded and turned away a great many people, saying that gods made with hands are not gods.
ACTS|19|27|And there is danger not only that this trade of ours may come into disrepute but also that the temple of the great goddess Artemis may be counted as nothing, and that she may even be deposed from her magnificence, she whom all Asia and the world worship."
ACTS|19|28|When they heard this they were enraged and were crying out, "Great is Artemis of the Ephesians!"
ACTS|19|29|So the city was filled with the confusion, and they rushed together into the theater, dragging with them Gaius and Aristarchus, Macedonians who were Paul's companions in travel.
ACTS|19|30|But when Paul wished to go in among the crowd, the disciples would not let him.
ACTS|19|31|And even some of the Asiarchs, who were friends of his, sent to him and were urging him not to venture into the theater.
ACTS|19|32|Now some cried out one thing, some another, for the assembly was in confusion, and most of them did not know why they had come together.
ACTS|19|33|Some of the crowd prompted Alexander, whom the Jews had put forward. And Alexander, motioning with his hand, wanted to make a defense to the crowd.
ACTS|19|34|But when they recognized that he was a Jew, for about two hours they all cried out with one voice, "Great is Artemis of the Ephesians!"
ACTS|19|35|And when the town clerk had quieted the crowd, he said, "Men of Ephesus, who is there who does not know that the city of the Ephesians is temple keeper of the great Artemis, and of the sacred stone that fell from the sky?
ACTS|19|36|Seeing then that these things cannot be denied, you ought to be quiet and do nothing rash.
ACTS|19|37|For you have brought these men here who are neither sacrilegious nor blasphemers of our goddess.
ACTS|19|38|If therefore Demetrius and the craftsmen with him have a complaint against anyone, the courts are open, and there are proconsuls. Let them bring charges against one another.
ACTS|19|39|But if you seek anything further, it shall be settled in the regular assembly.
ACTS|19|40|For we really are in danger of being charged with rioting today, since there is no cause that we can give to justify this commotion."
ACTS|19|41|And when he had said these things, he dismissed the assembly.
ACTS|20|1|After the uproar ceased, Paul sent for the disciples, and after encouraging them, he said farewell and departed for Macedonia.
ACTS|20|2|When he had gone through those regions and had given them much encouragement, he came to Greece.
ACTS|20|3|There he spent three months, and when a plot was made against him by the Jews as he was about to set sail for Syria, he decided to return through Macedonia.
ACTS|20|4|Sopater of Berea, the son of Pyrrhus from Berea, accompanied him; and of the Thessalonians, Aristarchus and Secundus; and Gaius of Derbe, and Timothy; and the Asians, Tychicus and Trophimus.
ACTS|20|5|These went on ahead and were waiting for us at Troas,
ACTS|20|6|but we sailed away from Philippi after the days of Unleavened Bread, and in five days we came to them at Troas, where we stayed for seven days.
ACTS|20|7|On the first day of the week, when we were gathered together to break bread, Paul talked with them, intending to depart on the next day, and he prolonged his speech until midnight.
ACTS|20|8|There were many lamps in the upper room where we were gathered.
ACTS|20|9|And a young man named Eutychus, sitting at the window, sank into a deep sleep as Paul talked still longer. And being overcome by sleep, he fell down from the third story and was taken up dead.
ACTS|20|10|But Paul went down and bent over him, and taking him in his arms, said, "Do not be alarmed, for his life is in him."
ACTS|20|11|And when Paul had gone up and had broken bread and eaten, he conversed with them a long while, until daybreak, and so departed.
ACTS|20|12|And they took the youth away alive, and were not a little comforted.
ACTS|20|13|But going ahead to the ship, we set sail for Assos, intending to take Paul aboard there, for so he had arranged, intending himself to go by land.
ACTS|20|14|And when he met us at Assos, we took him on board and went to Mitylene.
ACTS|20|15|And sailing from there we came the following day opposite Chios; the next day we touched at Samos; and the day after that we went to Miletus.
ACTS|20|16|For Paul had decided to sail past Ephesus, so that he might not have to spend time in Asia, for he was hastening to be at Jerusalem, if possible, on the day of Pentecost.
ACTS|20|17|Now from Miletus he sent to Ephesus and called the elders of the church to come to him.
ACTS|20|18|And when they came to him, he said to them: "You yourselves know how I lived among you the whole time from the first day that I set foot in Asia,
ACTS|20|19|serving the Lord with all humility and with tears and with trials that happened to me through the plots of the Jews;
ACTS|20|20|how I did not shrink from declaring to you anything that was profitable, and teaching you in public and from house to house,
ACTS|20|21|testifying both to Jews and to Greeks of repentance toward God and of faith in our Lord Jesus Christ.
ACTS|20|22|And now, behold, I am going to Jerusalem, constrained by the Spirit, not knowing what will happen to me there,
ACTS|20|23|except that the Holy Spirit testifies to me in every city that imprisonment and afflictions await me.
ACTS|20|24|But I do not account my life of any value nor as precious to myself, if only I may finish my course and the ministry that I received from the Lord Jesus, to testify to the gospel of the grace of God.
ACTS|20|25|And now, behold, I know that none of you among whom I have gone about proclaiming the kingdom will see my face again.
ACTS|20|26|Therefore I testify to you this day that I am innocent of the blood of all of you,
ACTS|20|27|for I did not shrink from declaring to you the whole counsel of God.
ACTS|20|28|Pay careful attention to yourselves and to all the flock, in which the Holy Spirit has made you overseers, to care for the church of God, which he obtained with his own blood.
ACTS|20|29|I know that after my departure fierce wolves will come in among you, not sparing the flock;
ACTS|20|30|and from among your own selves will arise men speaking twisted things, to draw away the disciples after them.
ACTS|20|31|Therefore be alert, remembering that for three years I did not cease night or day to admonish everyone with tears.
ACTS|20|32|And now I commend you to God and to the word of his grace, which is able to build you up and to give you the inheritance among all those who are sanctified.
ACTS|20|33|I coveted no one's silver or gold or apparel.
ACTS|20|34|You yourselves know that these hands ministered to my necessities and to those who were with me.
ACTS|20|35|In all things I have shown you that by working hard in this way we must help the weak and remember the words of the Lord Jesus, how he himself said, 'It is more blessed to give than to receive.'"
ACTS|20|36|And when he had said these things, he knelt down and prayed with them all.
ACTS|20|37|And there was much weeping on the part of all; they embraced Paul and kissed him,
ACTS|20|38|being sorrowful most of all because of the word he had spoken, that they would not see his face again. And they accompanied him to the ship.
ACTS|21|1|And when we had parted from them and set sail, we came by a straight course to Cos, and the next day to Rhodes, and from there to Patara.
ACTS|21|2|And having found a ship crossing to Phoenicia, we went aboard and set sail.
ACTS|21|3|When we had come in sight of Cyprus, leaving it on the left we sailed to Syria and landed at Tyre, for there the ship was to unload its cargo.
ACTS|21|4|And having sought out the disciples, we stayed there for seven days. And through the Spirit they were telling Paul not to go on to Jerusalem.
ACTS|21|5|When our days there were ended, we departed and went on our journey, and they all, with wives and children, accompanied us until we were outside the city. And kneeling down on the beach, we prayed
ACTS|21|6|and said farewell to one another. Then we went on board the ship, and they returned home.
ACTS|21|7|When we had finished the voyage from Tyre, we arrived at Ptolemais, and we greeted the brothers and stayed with them for one day.
ACTS|21|8|On the next day we departed and came to Caesarea, and we entered the house of Philip the evangelist, who was one of the seven, and stayed with him.
ACTS|21|9|He had four unmarried daughters, who prophesied.
ACTS|21|10|While we were staying for many days, a prophet named Agabus came down from Judea.
ACTS|21|11|And coming to us, he took Paul's belt and bound his own feet and hands and said, "Thus says the Holy Spirit, 'This is how the Jews at Jerusalem will bind the man who owns this belt and deliver him into the hands of the Gentiles.'"
ACTS|21|12|When we heard this, we and the people there urged him not to go up to Jerusalem.
ACTS|21|13|Then Paul answered, "What are you doing, weeping and breaking my heart? For I am ready not only to be imprisoned but even to die in Jerusalem for the name of the Lord Jesus."
ACTS|21|14|And since he would not be persuaded, we ceased and said, "Let the will of the Lord be done."
ACTS|21|15|After these days we got ready and went up to Jerusalem.
ACTS|21|16|And some of the disciples from Caesarea went with us, bringing us to the house of Mnason of Cyprus, an early disciple, with whom we should lodge.
ACTS|21|17|When we had come to Jerusalem, the brothers received us gladly.
ACTS|21|18|On the following day Paul went in with us to James, and all the elders were present.
ACTS|21|19|After greeting them, he related one by one the things that God had done among the Gentiles through his ministry.
ACTS|21|20|And when they heard it, they glorified God. And they said to him, "You see, brother, how many thousands there are among the Jews of those who have believed. They are all zealous for the law,
ACTS|21|21|and they have been told about you that you teach all the Jews who are among the Gentiles to forsake Moses, telling them not to circumcise their children or walk according to our customs.
ACTS|21|22|What then is to be done? They will certainly hear that you have come.
ACTS|21|23|Do therefore what we tell you. We have four men who are under a vow;
ACTS|21|24|take these men and purify yourself along with them and pay their expenses, so that they may shave their heads. Thus all will know that there is nothing in what they have been told about you, but that you yourself also live in observance of the law.
ACTS|21|25|But as for the Gentiles who have believed, we have sent a letter with our judgment that they should abstain from what has been sacrificed to idols, and from blood, and from what has been strangled, and from sexual immorality."
ACTS|21|26|Then Paul took the men, and the next day he purified himself along with them and went into the temple, giving notice when the days of purification would be fulfilled and the offering presented for each one of them.
ACTS|21|27|When the seven days were almost completed, the Jews from Asia, seeing him in the temple, stirred up the whole crowd and laid hands on him,
ACTS|21|28|crying out, "Men of Israel, help! This is the man who is teaching everyone everywhere against the people and the law and this place. Moreover, he even brought Greeks into the temple and has defiled this holy place."
ACTS|21|29|For they had previously seen Trophimus the Ephesian with him in the city, and they supposed that Paul had brought him into the temple.
ACTS|21|30|Then all the city was stirred up, and the people ran together. They seized Paul and dragged him out of the temple, and at once the gates were shut.
ACTS|21|31|And as they were seeking to kill him, word came to the tribune of the cohort that all Jerusalem was in confusion.
ACTS|21|32|He at once took soldiers and centurions and ran down to them. And when they saw the tribune and the soldiers, they stopped beating Paul.
ACTS|21|33|Then the tribune came up and arrested him and ordered him to be bound with two chains. He inquired who he was and what he had done.
ACTS|21|34|Some in the crowd were shouting one thing, some another. And as he could not learn the facts because of the uproar, he ordered him to be brought into the barracks.
ACTS|21|35|And when he came to the steps, he was actually carried by the soldiers because of the violence of the crowd,
ACTS|21|36|for the mob of the people followed, crying out, "Away with him!"
ACTS|21|37|As Paul was about to be brought into the barracks, he said to the tribune, "May I say something to you?" And he said, "Do you know Greek?
ACTS|21|38|Are you not the Egyptian, then, who recently stirred up a revolt and led the four thousand men of the Assassins out into the wilderness?"
ACTS|21|39|Paul replied, "I am a Jew, from Tarsus in Cilicia, a citizen of no obscure city. I beg you, permit me to speak to the people."
ACTS|21|40|And when he had given him permission, Paul, standing on the steps, motioned with his hand to the people. And when there was a great hush, he addressed them in the Hebrew language, saying:
ACTS|22|1|"Brothers and fathers, hear the defense that I now make before you."
ACTS|22|2|And when they heard that he was addressing them in the Hebrew language, they became even more quiet. And he said:
ACTS|22|3|"I am a Jew, born in Tarsus in Cilicia, but brought up in this city, educated at the feet of Gamaliel according to the strict manner of the law of our fathers, being zealous for God as all of you are this day.
ACTS|22|4|I persecuted this Way to the death, binding and delivering to prison both men and women,
ACTS|22|5|as the high priest and the whole council of elders can bear me witness. From them I received letters to the brothers, and I journeyed toward Damascus to take those also who were there and bring them in bonds to Jerusalem to be punished.
ACTS|22|6|"As I was on my way and drew near to Damascus, about noon a great light from heaven suddenly shone around me.
ACTS|22|7|And I fell to the ground and heard a voice saying to me, 'Saul, Saul, why are you persecuting me?'
ACTS|22|8|And I answered, 'Who are you, Lord?' And he said to me, 'I am Jesus of Nazareth, whom you are persecuting.'
ACTS|22|9|Now those who were with me saw the light but did not understand the voice of the one who was speaking to me.
ACTS|22|10|And I said, 'What shall I do, Lord?' And the Lord said to me, 'Rise, and go into Damascus, and there you will be told all that is appointed for you to do.'
ACTS|22|11|And since I could not see because of the brightness of that light, I was led by the hand by those who were with me, and came into Damascus.
ACTS|22|12|"And one Ananias, a devout man according to the law, well spoken of by all the Jews who lived there,
ACTS|22|13|came to me, and standing by me said to me, 'Brother Saul, receive your sight.' And at that very hour I received my sight and saw him.
ACTS|22|14|And he said, 'The God of our fathers appointed you to know his will, to see the Righteous One and to hear a voice from his mouth;
ACTS|22|15|for you will be a witness for him to everyone of what you have seen and heard.
ACTS|22|16|And now why do you wait? Rise and be baptized and wash away your sins, calling on his name.'
ACTS|22|17|"When I had returned to Jerusalem and was praying in the temple, I fell into a trance
ACTS|22|18|and saw him saying to me, 'Make haste and get out of Jerusalem quickly, because they will not accept your testimony about me.'
ACTS|22|19|And I said, 'Lord, they themselves know that in one synagogue after another I imprisoned and beat those who believed in you.
ACTS|22|20|And when the blood of Stephen your witness was being shed, I myself was standing by and approving and watching over the garments of those who killed him.'
ACTS|22|21|And he said to me, 'Go, for I will send you far away to the Gentiles.'"
ACTS|22|22|Up to this word they listened to him. Then they raised their voices and said, "Away with such a fellow from the earth! For he should not be allowed to live."
ACTS|22|23|And as they were shouting and throwing off their cloaks and flinging dust into the air,
ACTS|22|24|the tribune ordered him to be brought into the barracks, saying that he should be examined by flogging, to find out why they were shouting against him like this.
ACTS|22|25|But when they had stretched him out for the whips, Paul said to the centurion who was standing by, "Is it lawful for you to flog a man who is a Roman citizen and uncondemned?"
ACTS|22|26|When the centurion heard this, he went to the tribune and said to him, "What are you about to do? For this man is a Roman citizen."
ACTS|22|27|So the tribune came and said to him, "Tell me, are you a Roman citizen?" And he said, "Yes."
ACTS|22|28|The tribune answered, "I bought this citizenship for a large sum." Paul said, "But I am a citizen by birth."
ACTS|22|29|So those who were about to examine him withdrew from him immediately, and the tribune also was afraid, for he realized that Paul was a Roman citizen and that he had bound him.
ACTS|22|30|But on the next day, desiring to know the real reason why he was being accused by the Jews, he unbound him and commanded the chief priests and all the council to meet, and he brought Paul down and set him before them.
ACTS|23|1|And looking intently at the council, Paul said, "Brothers, I have lived my life before God in all good conscience up to this day."
ACTS|23|2|And the high priest Ananias commanded those who stood by him to strike him on the mouth.
ACTS|23|3|Then Paul said to him, "God is going to strike you, you whitewashed wall! Are you sitting to judge me according to the law, and yet contrary to the law you order me to be struck?"
ACTS|23|4|Those who stood by said, "Would you revile God's high priest?"
ACTS|23|5|And Paul said, "I did not know, brothers, that he was the high priest, for it is written, 'You shall not speak evil of a ruler of your people.'"
ACTS|23|6|Now when Paul perceived that one part were Sadducees and the other Pharisees, he cried out in the council, "Brothers, I am a Pharisee, a son of Pharisees. It is with respect to the hope and the resurrection of the dead that I am on trial."
ACTS|23|7|And when he had said this, a dissension arose between the Pharisees and the Sadducees, and the assembly was divided.
ACTS|23|8|For the Sadducees say that there is no resurrection, nor angel, nor spirit, but the Pharisees acknowledge them all.
ACTS|23|9|Then a great clamor arose, and some of the scribes of the Pharisees' party stood up and contended sharply, "We find nothing wrong in this man. What if a spirit or an angel spoke to him?"
ACTS|23|10|And when the dissension became violent, the tribune, afraid that Paul would be torn to pieces by them, commanded the soldiers to go down and take him away from among them by force and bring him into the barracks.
ACTS|23|11|The following night the Lord stood by him and said, "Take courage, for as you have testified to the facts about me in Jerusalem, so you must testify also in Rome."
ACTS|23|12|When it was day, the Jews made a plot and bound themselves by an oath neither to eat nor drink till they had killed Paul.
ACTS|23|13|There were more than forty who made this conspiracy.
ACTS|23|14|They went to the chief priests and elders and said, "We have strictly bound ourselves by an oath to taste no food till we have killed Paul.
ACTS|23|15|Now therefore you, along with the council, give notice to the tribune to bring him down to you, as though you were going to determine his case more exactly. And we are ready to kill him before he comes near."
ACTS|23|16|Now the son of Paul's sister heard of their ambush, so he went and entered the barracks and told Paul.
ACTS|23|17|Paul called one of the centurions and said, "Take this young man to the tribune, for he has something to tell him."
ACTS|23|18|So he took him and brought him to the tribune and said, "Paul the prisoner called me and asked me to bring this young man to you, as he has something to say to you."
ACTS|23|19|The tribune took him by the hand, and going aside asked him privately, "What is it that you have to tell me?"
ACTS|23|20|And he said, "The Jews have agreed to ask you to bring Paul down to the council tomorrow, as though they were going to inquire somewhat more closely about him.
ACTS|23|21|But do not be persuaded by them, for more than forty of their men are lying in ambush for him, who have bound themselves by an oath neither to eat nor drink till they have killed him. And now they are ready, waiting for your consent."
ACTS|23|22|So the tribune dismissed the young man, charging him, "Tell no one that you have informed me of these things."
ACTS|23|23|Then he called two of the centurions and said, "Get ready two hundred soldiers, with seventy horsemen and two hundred spearmen to go as far as Caesarea at the third hour of the night.
ACTS|23|24|Also provide mounts for Paul to ride and bring him safely to Felix the governor."
ACTS|23|25|And he wrote a letter to this effect:
ACTS|23|26|"Claudius Lysias, to his Excellency the governor Felix, greetings.
ACTS|23|27|This man was seized by the Jews and was about to be killed by them when I came upon them with the soldiers and rescued him, having learned that he was a Roman citizen.
ACTS|23|28|And desiring to know the charge for which they were accusing him, I brought him down to their council.
ACTS|23|29|I found that he was being accused about questions of their law, but charged with nothing deserving death or imprisonment.
ACTS|23|30|And when it was disclosed to me that there would be a plot against the man, I sent him to you at once, ordering his accusers also to state before you what they have against him."
ACTS|23|31|So the soldiers, according to their instructions, took Paul and brought him by night to Antipatris.
ACTS|23|32|And on the next day they returned to the barracks, letting the horsemen go on with him.
ACTS|23|33|When they had come to Caesarea and delivered the letter to the governor, they presented Paul also before him.
ACTS|23|34|On reading the letter, he asked what province he was from. And when he learned that he was from Cilicia,
ACTS|23|35|he said, "I will give you a hearing when your accusers arrive." And he commanded him to be guarded in Herod's praetorium.
ACTS|24|1|And after five days the high priest Ananias came down with some elders and a spokesman, one Tertullus. They laid before the governor their case against Paul.
ACTS|24|2|And when he had been summoned, Tertullus began to accuse him, saying: "Since through you we enjoy much peace, and since by your foresight, most excellent Felix, reforms are being made for this nation,
ACTS|24|3|in every way and everywhere we accept this with all gratitude.
ACTS|24|4|But, to detain you no further, I beg you in your kindness to hear us briefly.
ACTS|24|5|For we have found this man a plague, one who stirs up riots among all the Jews throughout the world and is a ringleader of the sect of the Nazarenes.
ACTS|24|6|He even tried to profane the temple, but we seized him.
ACTS|24|7|***
ACTS|24|8|By examining him yourself you will be able to find out from him about everything of which we accuse him."
ACTS|24|9|The Jews also joined in the charge, affirming that all these things were so.
ACTS|24|10|And when the governor had nodded to him to speak, Paul replied: "Knowing that for many years you have been a judge over this nation, I cheerfully make my defense.
ACTS|24|11|You can verify that it is not more than twelve days since I went up to worship in Jerusalem,
ACTS|24|12|and they did not find me disputing with anyone or stirring up a crowd, either in the temple or in the synagogues or in the city.
ACTS|24|13|Neither can they prove to you what they now bring up against me.
ACTS|24|14|But this I confess to you, that according to the Way, which they call a sect, I worship the God of our fathers, believing everything laid down by the Law and written in the Prophets,
ACTS|24|15|having a hope in God, which these men themselves accept, that there will be a resurrection of both the just and the unjust.
ACTS|24|16|So I always take pains to have a clear conscience toward both God and man.
ACTS|24|17|Now after several years I came to bring alms to my nation and to present offerings.
ACTS|24|18|While I was doing this, they found me purified in the temple, without any crowd or tumult. But some Jews from Asia-
ACTS|24|19|they ought to be here before you and to make an accusation, should they have anything against me.
ACTS|24|20|Or else let these men themselves say what wrongdoing they found when I stood before the council,
ACTS|24|21|other than this one thing that I cried out while standing among them: 'It is with respect to the resurrection of the dead that I am on trial before you this day.'"
ACTS|24|22|But Felix, having a rather accurate knowledge of the Way, put them off, saying, "When Lysias the tribune comes down, I will decide your case."
ACTS|24|23|Then he gave orders to the centurion that he should be kept in custody but have some liberty, and that none of his friends should be prevented from attending to his needs.
ACTS|24|24|After some days Felix came with his wife Drusilla, who was Jewish, and he sent for Paul and heard him speak about faith in Christ Jesus.
ACTS|24|25|And as he reasoned about righteousness and self-control and the coming judgment, Felix was alarmed and said, "Go away for the present. When I get an opportunity I will summon you."
ACTS|24|26|At the same time he hoped that money would be given him by Paul. So he sent for him often and conversed with him.
ACTS|24|27|When two years had elapsed, Felix was succeeded by Porcius Festus. And desiring to do the Jews a favor, Felix left Paul in prison.
ACTS|25|1|Now three days after Festus had arrived in the province, he went up to Jerusalem from Caesarea.
ACTS|25|2|And the chief priests and the principal men of the Jews laid out their case against Paul, and they urged him,
ACTS|25|3|asking as a favor against Paul that he summon him to Jerusalem- because they were planning an ambush to kill him on the way.
ACTS|25|4|Festus replied that Paul was being kept at Caesarea and that he himself intended to go there shortly.
ACTS|25|5|"So," said he, "let the men of authority among you go down with me, and if there is anything wrong about the man, let them bring charges against him."
ACTS|25|6|After he stayed among them not more than eight or ten days, he went down to Caesarea. And the next day he took his seat on the tribunal and ordered Paul to be brought.
ACTS|25|7|When he had arrived, the Jews who had come down from Jerusalem stood around him, bringing many and serious charges against him that they could not prove.
ACTS|25|8|Paul argued in his defense, "Neither against the law of the Jews, nor against the temple, nor against Caesar have I committed any offense."
ACTS|25|9|But Festus, wishing to do the Jews a favor, said to Paul, "Do you wish to go up to Jerusalem and there be tried on these charges before me?"
ACTS|25|10|But Paul said, "I am standing before Caesar's tribunal, where I ought to be tried. To the Jews I have done no wrong, as you yourselves know very well.
ACTS|25|11|If then I am a wrongdoer and have committed anything for which I deserve to die, I do not seek to escape death. But if there is nothing to their charges against me, no one can give me up to them. I appeal to Caesar."
ACTS|25|12|Then Festus, when he had conferred with his council, answered, "To Caesar you have appealed; to Caesar you shall go."
ACTS|25|13|Now when some days had passed, Agrippa the king and Bernice arrived at Caesarea and greeted Festus.
ACTS|25|14|And as they stayed there many days, Festus laid Paul's case before the king, saying, "There is a man left prisoner by Felix,
ACTS|25|15|and when I was at Jerusalem, the chief priests and the elders of the Jews laid out their case against him, asking for a sentence of condemnation against him.
ACTS|25|16|I answered them that it was not the custom of the Romans to give up anyone before the accused met the accusers face to face and had opportunity to make his defense concerning the charge laid against him.
ACTS|25|17|So when they came together here, I made no delay, but on the next day took my seat on the tribunal and ordered the man to be brought.
ACTS|25|18|When the accusers stood up, they brought no charge in his case of such evils as I supposed.
ACTS|25|19|Rather they had certain points of dispute with him about their own religion and about a certain Jesus, who was dead, but whom Paul asserted to be alive.
ACTS|25|20|Being at a loss how to investigate these questions, I asked whether he wanted to go to Jerusalem and be tried there regarding them.
ACTS|25|21|But when Paul had appealed to be kept in custody for the decision of the emperor, I ordered him to be held until I could send him to Caesar."
ACTS|25|22|Then Agrippa said to Festus, "I would like to hear the man myself." "Tomorrow," said he, "you will hear him."
ACTS|25|23|So on the next day Agrippa and Bernice came with great pomp, and they entered the audience hall with the military tribunes and the prominent men of the city. Then, at the command of Festus, Paul was brought in.
ACTS|25|24|And Festus said, "King Agrippa and all who are present with us, you see this man about whom the whole Jewish people petitioned me, both in Jerusalem and here, shouting that he ought not to live any longer.
ACTS|25|25|But I found that he had done nothing deserving death. And as he himself appealed to the emperor, I decided to go ahead and send him.
ACTS|25|26|But I have nothing definite to write to my lord about him. Therefore I have brought him before you all, and especially before you, King Agrippa, so that, after we have examined him, I may have something to write.
ACTS|25|27|For it seems to me unreasonable, in sending a prisoner, not to indicate the charges against him."
ACTS|26|1|So Agrippa said to Paul, "You have permission to speak for yourself." Then Paul stretched out his hand and made his defense:
ACTS|26|2|"I consider myself fortunate that it is before you, King Agrippa, I am going to make my defense today against all the accusations of the Jews,
ACTS|26|3|especially because you are familiar with all the customs and controversies of the Jews. Therefore I beg you to listen to me patiently.
ACTS|26|4|"My manner of life from my youth, spent from the beginning among my own nation and in Jerusalem, is known by all the Jews.
ACTS|26|5|They have known for a long time, if they are willing to testify, that according to the strictest party of our religion I have lived as a Pharisee.
ACTS|26|6|And now I stand here on trial because of my hope in the promise made by God to our fathers,
ACTS|26|7|to which our twelve tribes hope to attain, as they earnestly worship night and day. And for this hope I am accused by Jews, O king!
ACTS|26|8|Why is it thought incredible by any of you that God raises the dead?
ACTS|26|9|"I myself was convinced that I ought to do many things in opposing the name of Jesus of Nazareth.
ACTS|26|10|And I did so in Jerusalem. I not only locked up many of the saints in prison after receiving authority from the chief priests, but when they were put to death I cast my vote against them.
ACTS|26|11|And I punished them often in all the synagogues and tried to make them blaspheme, and in raging fury against them I persecuted them even to foreign cities.
ACTS|26|12|"In this connection I journeyed to Damascus with the authority and commission of the chief priests.
ACTS|26|13|At midday, O king, I saw on the way a light from heaven, brighter than the sun, that shone around me and those who journeyed with me.
ACTS|26|14|And when we had all fallen to the ground, I heard a voice saying to me in the Hebrew language, 'Saul, Saul, why are you persecuting me? It is hard for you to kick against the goads.'
ACTS|26|15|And I said, 'Who are you, Lord?' And the Lord said, 'I am Jesus whom you are persecuting.
ACTS|26|16|But rise and stand upon your feet, for I have appeared to you for this purpose, to appoint you as a servant and witness to the things in which you have seen me and to those in which I will appear to you,
ACTS|26|17|delivering you from your people and from the Gentiles- to whom I am sending you
ACTS|26|18|to open their eyes, so that they may turn from darkness to light and from the power of Satan to God, that they may receive forgiveness of sins and a place among those who are sanctified by faith in me.'
ACTS|26|19|"Therefore, O King Agrippa, I was not disobedient to the heavenly vision,
ACTS|26|20|but declared first to those in Damascus, then in Jerusalem and throughout all the region of Judea, and also to the Gentiles, that they should repent and turn to God, performing deeds in keeping with their repentance.
ACTS|26|21|For this reason the Jews seized me in the temple and tried to kill me.
ACTS|26|22|To this day I have had the help that comes from God, and so I stand here testifying both to small and great, saying nothing but what the prophets and Moses said would come to pass:
ACTS|26|23|that the Christ must suffer and that, by being the first to rise from the dead, he would proclaim light both to our people and to the Gentiles."
ACTS|26|24|And as he was saying these things in his defense, Festus said with a loud voice, "Paul, you are out of your mind; your great learning is driving you out of your mind."
ACTS|26|25|But Paul said, "I am not out of my mind, most excellent Festus, but I am speaking true and rational words.
ACTS|26|26|For the king knows about these things, and to him I speak boldly. For I am persuaded that none of these things has escaped his notice, for this has not been done in a corner.
ACTS|26|27|King Agrippa, do you believe the prophets? I know that you believe."
ACTS|26|28|And Agrippa said to Paul, "In a short time would you persuade me to be a Christian?"
ACTS|26|29|And Paul said, "Whether short or long, I would to God that not only you but also all who hear me this day might become such as I am- except for these chains."
ACTS|26|30|Then the king rose, and the governor and Bernice and those who were sitting with them.
ACTS|26|31|And when they had withdrawn, they said to one another, "This man is doing nothing to deserve death or imprisonment."
ACTS|26|32|And Agrippa said to Festus, "This man could have been set free if he had not appealed to Caesar."
ACTS|27|1|And when it was decided that we should sail for Italy, they delivered Paul and some other prisoners to a centurion of the Augustan Cohort named Julius.
ACTS|27|2|And embarking in a ship of Adramyttium, which was about to sail to the ports along the coast of Asia, we put to sea, accompanied by Aristarchus, a Macedonian from Thessalonica.
ACTS|27|3|The next day we put in at Sidon. And Julius treated Paul kindly and gave him leave to go to his friends and be cared for.
ACTS|27|4|And putting out to sea from there we sailed under the lee of Cyprus, because the winds were against us.
ACTS|27|5|And when we had sailed across the open sea along the coast of Cilicia and Pamphylia, we came to Myra in Lycia.
ACTS|27|6|There the centurion found a ship of Alexandria sailing for Italy and put us on board.
ACTS|27|7|We sailed slowly for a number of days and arrived with difficulty off Cnidus, and as the wind did not allow us to go farther, we sailed under the lee of Crete off Salmone.
ACTS|27|8|Coasting along it with difficulty, we came to a place called Fair Havens, near which was the city of Lasea.
ACTS|27|9|Since much time had passed, and the voyage was now dangerous because even the Fast was already over, Paul advised them,
ACTS|27|10|saying, "Sirs, I perceive that the voyage will be with injury and much loss, not only of the cargo and the ship, but also of our lives."
ACTS|27|11|But the centurion paid more attention to the pilot and to the owner of the ship than to what Paul said.
ACTS|27|12|And because the harbor was not suitable to spend the winter in, the majority decided to put out to sea from there, on the chance that somehow they could reach Phoenix, a harbor of Crete, facing both southwest and northwest, and spend the winter there.
ACTS|27|13|Now when the south wind blew gently, supposing that they had obtained their purpose, they weighed anchor and sailed along Crete, close to the shore.
ACTS|27|14|But soon a tempestuous wind, called the northeaster, struck down from the land.
ACTS|27|15|And when the ship was caught and could not face the wind, we gave way to it and were driven along.
ACTS|27|16|Running under the lee of a small island called Cauda, we managed with difficulty to secure the ship's boat.
ACTS|27|17|After hoisting it up, they used supports to undergird the ship. Then, fearing that they would run aground on the Syrtis, they lowered the gear, and thus they were driven along.
ACTS|27|18|Since we were violently storm-tossed, they began the next day to jettison the cargo.
ACTS|27|19|And on the third day they threw the ship's tackle overboard with their own hands.
ACTS|27|20|When neither sun nor stars appeared for many days, and no small tempest lay on us, all hope of our being saved was at last abandoned.
ACTS|27|21|Since they had been without food for a long time, Paul stood up among them and said, "Men, you should have listened to me and not have set sail from Crete and incurred this injury and loss.
ACTS|27|22|Yet now I urge you to take heart, for there will be no loss of life among you, but only of the ship.
ACTS|27|23|For this very night there stood before me an angel of the God to whom I belong and whom I worship,
ACTS|27|24|and he said, 'Do not be afraid, Paul; you must stand before Caesar. And behold, God has granted you all those who sail with you.'
ACTS|27|25|So take heart, men, for I have faith in God that it will be exactly as I have been told.
ACTS|27|26|But we must run aground on some island."
ACTS|27|27|When the fourteenth night had come, as we were being driven across the Adriatic Sea, about midnight the sailors suspected that they were nearing land.
ACTS|27|28|So they took a sounding and found twenty fathoms. A little farther on they took a sounding again and found fifteen fathoms.
ACTS|27|29|And fearing that we might run on the rocks, they let down four anchors from the stern and prayed for day to come.
ACTS|27|30|And as the sailors were seeking to escape from the ship, and had lowered the ship's boat into the sea under pretense of laying out anchors from the bow,
ACTS|27|31|Paul said to the centurion and the soldiers, "Unless these men stay in the ship, you cannot be saved."
ACTS|27|32|Then the soldiers cut away the ropes of the ship's boat and let it go.
ACTS|27|33|As day was about to dawn, Paul urged them all to take some food, saying, "Today is the fourteenth day that you have continued in suspense and without food, having taken nothing.
ACTS|27|34|Therefore I urge you to take some food. It will give you strength, for not a hair is to perish from the head of any of you."
ACTS|27|35|And when he had said these things, he took bread, and giving thanks to God in the presence of all he broke it and began to eat.
ACTS|27|36|Then they all were encouraged and ate some food themselves.
ACTS|27|37|(We were in all 276 persons in the ship.)
ACTS|27|38|And when they had eaten enough, they lightened the ship, throwing out the wheat into the sea.
ACTS|27|39|Now when it was day, they did not recognize the land, but they noticed a bay with a beach, on which they planned if possible to run the ship ashore.
ACTS|27|40|So they cast off the anchors and left them in the sea, at the same time loosening the ropes that tied the rudders. Then hoisting the foresail to the wind they made for the beach.
ACTS|27|41|But striking a reef, they ran the vessel aground. The bow stuck and remained immovable, and the stern was being broken up by the surf.
ACTS|27|42|The soldiers' plan was to kill the prisoners, lest any should swim away and escape.
ACTS|27|43|But the centurion, wishing to save Paul, kept them from carrying out their plan. He ordered those who could swim to jump overboard first and make for the land,
ACTS|27|44|and the rest on planks or on pieces of the ship. And so it was that all were brought safely to land.
ACTS|28|1|After we were brought safely through, we then learned that the island was called Malta.
ACTS|28|2|The native people showed us unusual kindness, for they kindled a fire and welcomed us all, because it had begun to rain and was cold.
ACTS|28|3|When Paul had gathered a bundle of sticks and put them on the fire, a viper came out because of the heat and fastened on his hand.
ACTS|28|4|When the native people saw the creature hanging from his hand, they said to one another, "No doubt this man is a murderer. Though he has escaped from the sea, Justice has not allowed him to live."
ACTS|28|5|He, however, shook off the creature into the fire and suffered no harm.
ACTS|28|6|They were waiting for him to swell up or suddenly fall down dead. But when they had waited a long time and saw no misfortune come to him, they changed their minds and said that he was a god.
ACTS|28|7|Now in the neighborhood of that place were lands belonging to the chief man of the island, named Publius, who received us and entertained us hospitably for three days.
ACTS|28|8|It happened that the father of Publius lay sick with fever and dysentery. And Paul visited him and prayed, and putting his hands on him healed him.
ACTS|28|9|And when this had taken place, the rest of the people on the island who had diseases also came and were cured.
ACTS|28|10|They also honored us greatly, and when we were about to sail, they put on board whatever we needed.
ACTS|28|11|After three months we set sail in a ship that had wintered in the island, a ship of Alexandria, with the twin gods as a figurehead.
ACTS|28|12|Putting in at Syracuse, we stayed there for three days.
ACTS|28|13|And from there we made a circuit and arrived at Rhegium. And after one day a south wind sprang up, and on the second day we came to Puteoli.
ACTS|28|14|There we found brothers and were invited to stay with them for seven days. And so we came to Rome.
ACTS|28|15|And the brothers there, when they heard about us, came as far as the Forum of Appius and Three Taverns to meet us. On seeing them, Paul thanked God and took courage.
ACTS|28|16|And when we came into Rome, Paul was allowed to stay by himself, with the soldier that guarded him.
ACTS|28|17|After three days he called together the local leaders of the Jews, and when they had gathered, he said to them, "Brothers, though I had done nothing against our people or the customs of our fathers, yet I was delivered as a prisoner from Jerusalem into the hands of the Romans.
ACTS|28|18|When they had examined me, they wished to set me at liberty, because there was no reason for the death penalty in my case.
ACTS|28|19|But because the Jews objected, I was compelled to appeal to Caesar- though I had no charge to bring against my nation.
ACTS|28|20|For this reason, therefore, I have asked to see you and speak with you, since it is because of the hope of Israel that I am wearing this chain."
ACTS|28|21|And they said to him, "We have received no letters from Judea about you, and none of the brothers coming here has reported or spoken any evil about you.
ACTS|28|22|But we desire to hear from you what your views are, for with regard to this sect we know that everywhere it is spoken against."
ACTS|28|23|When they had appointed a day for him, they came to him at his lodging in greater numbers. From morning till evening he expounded to them, testifying to the kingdom of God and trying to convince them about Jesus both from the Law of Moses and from the Prophets.
ACTS|28|24|And some were convinced by what he said, but others disbelieved.
ACTS|28|25|And disagreeing among themselves, they departed after Paul had made one statement: "The Holy Spirit was right in saying to your fathers through Isaiah the prophet:
ACTS|28|26|"'Go to this people, and say, You will indeed hear but never understand, and you will indeed see but never perceive.
ACTS|28|27|For this people's heart has grown dull, and with their ears they can barely hear, and their eyes they have closed; lest they should see with their eyes and hear with their ears and understand with their heart and turn, and I would heal them.'
ACTS|28|28|Therefore let it be known to you that this salvation of God has been sent to the Gentiles; they will listen."
ACTS|28|29|***
ACTS|28|30|He lived there two whole years at his own expense, and welcomed all who came to him,
ACTS|28|31|proclaiming the kingdom of God and teaching about the Lord Jesus Christ with all boldness and without hindrance.
