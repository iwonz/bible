ZEPH|1|1|当 亚们 的儿子 犹大 王 约西亚 在位的时候，耶和华的话临到 希西家 的玄孙， 亚玛利雅 的曾孙， 基大利 的孙子， 古示 的儿子 西番雅 。
ZEPH|1|2|耶和华说： “我必从地面上彻底除灭万物。
ZEPH|1|3|我必除灭人与牲畜， 除灭空中的鸟、海里的鱼、 绊脚石和恶人； 我必把人从地面上剪除， 这是耶和华说的。
ZEPH|1|4|我必伸手攻击 犹大 和 耶路撒冷 所有的居民； 从这地方剪除剩下的 巴力 、 事奉偶像之祭司的名字与祭司；
ZEPH|1|5|还有那些在屋顶拜天上万象的， 那些敬拜耶和华指着他起誓， 却又指着 米勒公 起誓的；
ZEPH|1|6|并那些转去不跟从耶和华， 不寻求耶和华，也不求问他的。”
ZEPH|1|7|在主耶和华面前要静默无声， 因为耶和华的日子快到了。 耶和华已经预备祭物， 将召来的人分别为圣。
ZEPH|1|8|“到了献祭给耶和华的日子， 我要惩罚领袖和王子， 及所有穿外邦衣服的人。
ZEPH|1|9|到那日，我必惩罚所有跳过门槛， 以残暴和诡诈塞满主人房屋的人。
ZEPH|1|10|“当那日，从 鱼门 必发出悲哀的声音， 从第二城区发出哀号的声音， 从山间发出破裂的大响声。 这是耶和华说的。
ZEPH|1|11|玛革提施 的居民哪，你们要哀号， 因为所有的商人 都灭亡了， 满载银子的人都被剪除。
ZEPH|1|12|那时，我必用灯巡查 耶路撒冷 ， 惩罚那些沉湎在酒渣上的人； 他们心里说： ‘耶和华必不降福，也不降祸。’
ZEPH|1|13|他们的财宝成为掠物， 房屋变为废墟。 他们建造房屋，却不得住在其内； 栽葡萄园，却不得喝其中所出的酒。”
ZEPH|1|14|耶和华的大日临近， 临近而且甚快； 那是耶和华日子的风声， 勇士必在那里痛痛地哭号。
ZEPH|1|15|那日是愤怒的日子， 急难困苦的日子， 荒废凄凉的日子， 黑暗幽冥的日子， 乌云密布的日子，
ZEPH|1|16|是吹角呐喊的日子， 要攻击坚固的城， 攻击高大的城楼。
ZEPH|1|17|我必使灾祸临到人身上， 使他们行走如同盲人， 因为他们得罪了耶和华； 他们的血必倒出如灰尘， 肉身抛弃如粪土。
ZEPH|1|18|当耶和华发怒的日子， 他们的金银不能救自己； 耶和华妒忌的火必烧灭全地， 要向地上所有的居民施行可怕的毁灭。
ZEPH|2|1|不知羞耻的国民哪， 趁命令尚未发出， 日子流逝如糠秕， 耶和华的烈怒尚未临到你们， 他发怒的日子未到以先， 你们应当聚集，聚集起来。
ZEPH|2|2|
ZEPH|2|3|世上遵守耶和华典章的谦卑人哪， 你们都当寻求耶和华， 寻求公义，寻求谦卑； 或许在耶和华发怒的日子得以隐藏。
ZEPH|2|4|迦萨 必遭遗弃 ， 亚实基伦 必然荒凉； 亚实突 人必在正午被赶出， 以革伦 也要连根拔除 。
ZEPH|2|5|祸哉，住沿海之地的 基利提 人！ 迦南 、 非利士 人之地啊，耶和华的话攻击你们： 我必毁灭你，以致无人居住。
ZEPH|2|6|沿海之地要变为草场， 牧人的住处 和羊群的圈。
ZEPH|2|7|这地必为 犹大 家的余民所得； 他们要在那里放牧， 晚上躺卧在 亚实基伦 的房屋中； 因为耶和华－他们的上帝必眷顾他们， 使被掳的人归回。
ZEPH|2|8|我听见 摩押 毁谤， 亚扪 人辱骂； 他们辱骂我的百姓， 自夸自大，侵犯他们的疆土。”
ZEPH|2|9|万军之耶和华－ 以色列 的上帝说： 因此，我指着我的永生起誓： 摩押 必如 所多玛 ， 亚扪 人必像 蛾摩拉 ， 都变为刺草、盐坑、永远荒废之地。 我百姓中剩余的必掳掠他们， 我国中的幸存者必得他们的地。
ZEPH|2|10|这事临到他们是因他们的骄傲， 他们自夸自大， 辱骂万军之耶和华的百姓。
ZEPH|2|11|耶和华必向他们显为可畏， 因他使地上的众神衰微； 列国的海岛各在自己的地方敬拜他。
ZEPH|2|12|你们 古实 人， 也是被我的刀所杀的。
ZEPH|2|13|耶和华要伸手攻击北方， 毁灭 亚述 ， 使 尼尼微 荒凉， 干旱如同旷野。
ZEPH|2|14|群畜，就是各类 的走兽必卧在其中， 鹈鹕和豪猪要宿在柱顶； 窗户有鸣叫的声音， 门槛毁坏 ， 他要毁坏香柏木板 。
ZEPH|2|15|这素来欢乐、安然居住的城， 心里说：“惟有我，除我以外再没有别的”， 现在竟然荒凉，成为野兽躺卧之处！ 凡经过的人都必摇着手嗤笑它。
ZEPH|3|1|祸哉，这欺压的城！ 悖逆，污秽，
ZEPH|3|2|不听从命令， 不领受训诲， 不倚靠耶和华， 不亲近它的上帝。
ZEPH|3|3|其中的领袖是咆哮的狮子， 审判官是晚上 的野狼， 不留一点到早晨。
ZEPH|3|4|它的先知是虚浮诡诈的人， 祭司亵渎圣所，强解律法。
ZEPH|3|5|耶和华在它中间行公义， 断不做非义的事， 每早晨显明他的公义，无日不然； 只是不义的人不知羞耻。
ZEPH|3|6|“我已经除灭列国， 使他们的城楼荒废。 我使他们街道荒凉， 无人经过； 他们的城镇毁坏， 没有人，没有居民。
ZEPH|3|7|我说：‘只要你敬畏我， 领受训诲； 其住处就不会照我原先所定的被剪除 。’ 然而，他们从早起来就在各样事上败坏自己。
ZEPH|3|8|“你们要等候我， 直到我兴起掳掠 的日子； 因为我已定意招聚列邦，聚集列国， 将我的恼怒，我一切的烈怒，都倾倒在它们身上。 我妒忌的火必烧灭全地。 这是耶和华说的。
ZEPH|3|9|“那时，我要改变万民， 使他们有清洁的嘴唇， 好求告耶和华的名， 同心合意事奉我。
ZEPH|3|10|那些向我祈求的， 我所分散的子民 ， 必从 古实河 的那一边， 献供物给我。
ZEPH|3|11|“当那日，你必不再因一切得罪我的事蒙羞， 因为那时我必从你中间除掉狂喜高傲的人， 在我的圣山上你也不再狂傲。
ZEPH|3|12|我却要在你中间留下困苦贫寒的百姓， 他们必投靠耶和华的名。
ZEPH|3|13|以色列 的余民必不行恶， 不说谎，口中没有诡诈的舌头； 他们吃喝躺卧， 无人使他们惊吓。”
ZEPH|3|14|锡安 哪，应当歌唱！ 以色列 啊，应当欢呼！ 耶路撒冷 啊，应当满心欢喜快乐！
ZEPH|3|15|耶和华已经免去对你的审判， 赶出你的仇敌。 以色列 的王－耶和华在你中间； 你必不再惧怕灾祸。
ZEPH|3|16|当那日，必有话对 耶路撒冷 说： “不要惧怕！ 锡安 哪，不要手软！
ZEPH|3|17|耶和华－你的上帝在你中间 大有能力，施行拯救。 他必因你欢欣喜乐， 他在爱中静默， 且因你而喜乐欢呼。
ZEPH|3|18|我要聚集那些因无节期而愁烦的人， 他们曾远离你， 是你的重担和羞辱 。
ZEPH|3|19|那时，看哪，我必对付所有苦待你的人， 拯救瘸腿的，召集被赶出的； 那些在全地受羞辱的， 我必使他们得称赞，享名声。
ZEPH|3|20|那时，我必领你们回来，召集你们； 我使你们被掳之人归回的时候， 我必使你们在地上的万民中享名声，得称赞； 这是耶和华说的。”
