2PET|1|1|耶稣基督的仆人和使徒 西门．彼得 写信给那因我们的上帝和 救主耶稣基督的义，与我们同得一样宝贵信心的人。
2PET|1|2|愿恩惠、平安 ，因你们认识上帝和我们的主耶稣，多多加给你们！
2PET|1|3|上帝的神能已把一切关乎生命和虔敬的事赐给我们，因我们认识那用自己荣耀和美德召我们的上帝。
2PET|1|4|因此，他已把又宝贵又极大的应许赐给我们，使我们既脱离世上从情欲来的败坏，就得分享上帝的本性。
2PET|1|5|正因这缘故，你们要分外地努力。有了信心，又要加上德行；有了德行，又要加上知识；
2PET|1|6|有了知识，又要加上节制；有了节制，又要加上忍耐；有了忍耐，又要加上虔敬；
2PET|1|7|有了虔敬，又要加上爱弟兄的心；有了爱弟兄的心，又要加上爱众人的心。
2PET|1|8|你们有了这几样，再继续增长，就必使你们在认识我们的主耶稣基督上，不至于懒散和不结果子了。
2PET|1|9|没有这几样的人就是瞎眼，是短视，忘了他过去的罪已经得了洁净。
2PET|1|10|所以，弟兄们，要更加努力，使你们的蒙召和被选坚定不移。你们实行这几样，就永不失脚。
2PET|1|11|这样，必叫你们丰丰富富地得以进入我们主－救主耶稣基督永远的国度。
2PET|1|12|虽然你们已经知道这些事，并且在你们已有的真道上得到坚固，我还是要常常提醒你们这些事。
2PET|1|13|我认为趁我还在这帐棚的时候，应该激发你们的记忆，
2PET|1|14|因为知道我脱离这帐棚的时候快到了，正如我们的主耶稣基督所指示我的。
2PET|1|15|我也要尽心竭力，使你们在我去世以后时常记念这些事。
2PET|1|16|我们从前把我们主耶稣基督的大能和他来临的事告诉你们，并不是随从一些捏造出来的无稽传说，我们是曾经亲眼见过他的威荣的人。
2PET|1|17|他从父上帝得尊贵荣耀的时候，从至高无上的荣耀有声音出来，对他说：“这是我的爱子，我所喜悦的。”
2PET|1|18|我们同他在圣山的时候，亲自听见这声音从天上出来。
2PET|1|19|我们有先知更确实的信息，你们要好好地留意这信息，如同留意照耀在暗处的明灯，直等到天亮，晨星在你们心里升起的时候。
2PET|1|20|第一要紧的，你们要知道，经上所有的预言是不可随私意解释的，
2PET|1|21|因为预言从来没有出于人意的，而是人被圣灵感动说出上帝的话来。
2PET|2|1|从前在民间有假先知起来；同样，将来在你们中间也会有假教师，偷偷地引进使人灭亡的异端。他们甚至不认买他们的主人，自取迅速灭亡。
2PET|2|2|许多人会随从他们淫荡的行为，以致真理之道因他们的缘故被毁谤。
2PET|2|3|他们因贪婪，要用捏造的言语在你们身上取得利益。他们的惩罚，自古以来并不迟延；他们的灭亡也必迅速来到。
2PET|2|4|既然上帝没有宽容犯了罪的天使，反而把他们丢在地狱里，囚禁在幽暗中等候审判；
2PET|2|5|既然上帝也没有宽容上古的世界，曾叫洪水临到那不敬虔的世界，只保护了报公义信息的 挪亚 一家八口；
2PET|2|6|既然上帝判决了 所多玛 和 蛾摩拉 ，将二城倾覆 ，焚烧成灰，作为后世不敬虔人的鉴戒，
2PET|2|7|只搭救了那常为恶人的淫荡忧伤的义人 罗得 —
2PET|2|8|因为那义人住在他们当中，他正义的心因天天看见和听见他们不法的事而伤痛；
2PET|2|9|那么，主知道搭救敬虔的人脱离试炼，把不义的人留在惩罚之下等候审判的日子，
2PET|2|10|尤其那些随从肉体、放纵污秽的情欲、藐视主的权威的人更是如此。 他们胆大任性，无惧地毁谤众尊荣者；
2PET|2|11|就是天使，虽然力量权能更大，在对他们宣告从主来的审判的时候还不用毁谤的话 。
2PET|2|12|但这些人好像没有理性的牲畜，生来就是要被捉拿宰杀的。他们毁谤自己所不知道的事，正在败坏人的时候，自己也遭遇败坏，
2PET|2|13|为所行的不义受不义的工钱。他们喜爱白昼狂欢，他们已被玷污，又有瑕疵，正与你们一同欢宴，以自己的诡诈为乐。
2PET|2|14|他们满眼是淫色，是止不住的罪，引诱心不坚定的人，心中习惯了贪婪，正是被诅咒的种类。
2PET|2|15|他们离弃了正路，走入歧途，随从 比珥 的儿子 巴兰 的路； 巴兰 就是那贪爱不义的工钱的人，
2PET|2|16|他却为自己的过犯受了责备，而那不能说话的驴以人的声音阻止了先知的狂妄。
2PET|2|17|这些人是无水的泉源，是狂风催逼的雾气，有漆黑的幽暗为他们存留。
2PET|2|18|他们说虚妄夸大的话，用肉体的情欲和淫荡的事引诱那些刚脱离错谬生活的人。
2PET|2|19|他们应许人自由，自己却作了腐败的奴隶，因为人被谁制伏就是谁的奴隶。
2PET|2|20|倘若他们因认识我们的主和救主耶稣基督而得以脱离世上的污秽，后来又被污秽缠住，被制伏，他们末后的景况就比先前更不好了。
2PET|2|21|他们知道义路，竟背弃了传授给他们那神圣的诫命，倒不如不知道为妙。
2PET|2|22|俗语说得好，这话正印证在他们身上了： “狗转过来吃自己所吐的；” 又说： “猪洗净了，又回到烂泥里打滚。”
2PET|3|1|亲爱的，我现在写给你们的是第二封信。在这两封信里，我都提醒你们，激发你们真诚的心，
2PET|3|2|要你们记得圣先知预先所说的话和主—救主的命令，就是使徒所传给你们的。
2PET|3|3|第一要紧的，你们要知道，在末世必有好讥诮的人随从自己的私欲出来讥诮，
2PET|3|4|说：“他要来临的应许在哪里呢？因为从列祖长眠以来，万物与起初创造的时候仍是一样啊！”
2PET|3|5|他们故意忘记这事，就是从太古凭上帝的话有了天，并由水而出和藉着水而成的地；
2PET|3|6|藉着水，当时的世界被水淹没而消灭了。
2PET|3|7|但现在的天地还是凭着上帝的话存留，直留到不敬虔之人受审判遭沉沦的日子，用火焚烧。
2PET|3|8|亲爱的，有一件事你们不可忘记，就是：主看一日如千年，千年如一日。
2PET|3|9|主没有迟延他的应许，就如有人以为他是迟延，其实他是宽容你们，不愿一人沉沦，而是人人都来悔改。
2PET|3|10|但主的日子要像贼一样来到；那日，天必在轰然一声中消失，天体都要被烈火熔化，地和地上的万物都要烧尽 。
2PET|3|11|既然这一切都要如此消失，你们 处世为人必须圣洁敬虔，
2PET|3|12|等候并催促上帝的日子来到。因为在那日，天要被火烧而消灭，天体都要被烈火熔化。
2PET|3|13|但照他的应许，我们等候新天新地，其中有正义常住。
2PET|3|14|所以，亲爱的，既然你们等候这些事，就要竭力使自己没有玷污，无可指责，在主前和睦；
2PET|3|15|并且要以我们主的容忍作为你们得救的机会，就如我们所亲爱的弟兄 保罗 ，照着所赐给他的智慧写信给你们。
2PET|3|16|他一切的信上都谈到这事。信中有些难明白的，那无学问、不坚定的人加以曲解，如曲解别的经书一样，自取灭亡。
2PET|3|17|所以，亲爱的，既然你们预先知道这事，就当防备，免得被恶人的错谬诱惑，从自己稳定的立场上坠落。
2PET|3|18|你们倒要在我们的主和救主耶稣基督的恩典和知识上有长进。愿荣耀归给他，从今直到永远之日。阿们！
