MAL|1|1|Пророческое слово Господа к Израилю через Малахию.
MAL|1|2|Я возлюбил вас, говорит Господь. А вы говорите: "в чем явил Ты любовь к нам?" – Не брат ли Исав Иакову? говорит Господь; и однако же Я возлюбил Иакова,
MAL|1|3|а Исава возненавидел и предал горы его опустошению, и владения его – шакалам пустыни.
MAL|1|4|Если Едом скажет: "мы разорены, но мы восстановим разрушенное", то Господь Саваоф говорит: они построят, а Я разрушу, и прозовут их областью нечестивою, народом, на который Господь прогневался навсегда.
MAL|1|5|И увидят это глаза ваши, и вы скажете: "возвеличился Господь над пределами Израиля!"
MAL|1|6|Сын чтит отца и раб – господина своего; если Я отец, то где почтение ко Мне? и если Я Господь, то где благоговение предо Мною? говорит Господь Саваоф вам, священники, бесславящие имя Мое. Вы говорите: "чем мы бесславим имя Твое?"
MAL|1|7|Вы приносите на жертвенник Мой нечистый хлеб, и говорите: "чем мы бесславим Тебя?" – Тем, что говорите: "трапеза Господня не стоит уважения".
MAL|1|8|И когда приносите в жертву слепое, не худо ли это? или когда приносите хромое и больное, не худо ли это? Поднеси это твоему князю; будет ли он доволен тобою и благосклонно ли примет тебя? говорит Господь Саваоф.
MAL|1|9|Итак молитесь Богу, чтобы помиловал нас; а когда такое исходит из рук ваших, то может ли Он милостиво принимать вас? говорит Господь Саваоф.
MAL|1|10|Лучше кто–нибудь из вас запер бы двери, чтобы напрасно не держали огня на жертвеннике Моем. Нет Моего благоволения к вам, говорит Господь Саваоф, и приношение из рук ваших неблагоугодно Мне.
MAL|1|11|Ибо от востока солнца до запада велико будет имя Мое между народами, и на всяком месте будут приносить фимиам имени Моему, чистую жертву; велико будет имя Мое между народами, говорит Господь Саваоф.
MAL|1|12|А вы хулите его тем, что говорите: "трапеза Господня не стоит уважения, и доход от нее – пища ничтожная".
MAL|1|13|Притом говорите: "вот сколько труда!" и пренебрегаете ею, говорит Господь Саваоф, и приносите украденное, хромое и больное, и такого же свойства приносите хлебный дар: могу ли с благоволением принимать это из рук ваших? говорит Господь.
MAL|1|14|Проклят лживый, у которого в стаде есть неиспорченный самец, и он дал обет, а приносит в жертву Господу поврежденное: ибо Я Царь великий, и имя Мое страшно у народов.
MAL|2|1|Итак для вас, священники, эта заповедь:
MAL|2|2|если вы не послушаетесь и если не примете к сердцу, чтобы воздавать славу имени Моему, говорит Господь Саваоф, то Я пошлю на вас проклятие и прокляну ваши благословения, и уже проклинаю, потому что вы не хотите приложить к тому сердца.
MAL|2|3|Вот, Я отниму у вас плечо, и помет раскидаю на лица ваши, помет праздничных жертв ваших, и выбросят вас вместе с ним.
MAL|2|4|И вы узнаете, что Я дал эту заповедь для сохранения завета Моего с Левием, говорит Господь Саваоф.
MAL|2|5|Завет Мой с ним был [завет] жизни и мира, и Я дал его ему для страха, и он боялся Меня и благоговел пред именем Моим.
MAL|2|6|Закон истины был в устах его, и неправды не обреталось на языке его; в мире и правде он ходил со Мною и многих отвратил от греха.
MAL|2|7|Ибо уста священника должны хранить ведение, и закона ищут от уст его, потому что он вестник Господа Саваофа.
MAL|2|8|Но вы уклонились от пути сего, для многих послужили соблазном в законе, разрушили завет Левия, говорит Господь Саваоф.
MAL|2|9|За то и Я сделаю вас презренными и униженными перед всем народом, так как вы не соблюдаете путей Моих, лицеприятствуете в делах закона.
MAL|2|10|Не один ли у всех нас Отец? Не один ли Бог сотворил нас? Почему же мы вероломно поступаем друг против друга, нарушая тем завет отцов наших?
MAL|2|11|Вероломно поступает Иуда, и мерзость совершается в Израиле и в Иерусалиме; ибо унизил Иуда святыню Господню, которую любил, и женился на дочери чужого бога.
MAL|2|12|У того, кто делает это, истребит Господь из шатров Иаковлевых бдящего на страже и отвечающего, и приносящего жертву Господу Саваофу.
MAL|2|13|И вот еще что вы делаете: вы заставляете обливать слезами жертвенник Господа с рыданием и воплем, так что Он уже не призирает более на приношение и не принимает умилоствительной жертвы из рук ваших.
MAL|2|14|Вы скажете: "за что?" За то, что Господь был свидетелем между тобою и женою юности твоей, против которой ты поступил вероломно, между тем как она подруга твоя и законная жена твоя.
MAL|2|15|Но не сделал ли того же один, и в нем пребывал превосходный дух? что же сделал этот один? он желал получить от Бога потомство. Итак берегите дух ваш, и никто не поступай вероломно против жены юности своей.
MAL|2|16|Если ты ненавидишь ее, отпусти, говорит Господь Бог Израилев; обида покроет одежду его, говорит Господь Саваоф; посему наблюдайте за духом вашим и не поступайте вероломно.
MAL|2|17|Вы прогневляете Господа словами вашими и говорите: "чем прогневляем мы Его?" Тем, что говорите: "всякий, делающий зло, хорош пред очами Господа, и к таким Он благоволит", или: "где Бог правосудия?"
MAL|3|1|Вот, Я посылаю Ангела Моего, и он приготовит путь предо Мною, и внезапно придет в храм Свой Господь, Которого вы ищете, и Ангел завета, Которого вы желаете; вот, Он идет, говорит Господь Саваоф.
MAL|3|2|И кто выдержит день пришествия Его, и кто устоит, когда Он явится? Ибо Он – как огонь расплавляющий и как щелок очищающий,
MAL|3|3|и сядет переплавлять и очищать серебро, и очистит сынов Левия и переплавит их, как золото и как серебро, чтобы приносили жертву Господу в правде.
MAL|3|4|Тогда благоприятна будет Господу жертва Иуды и Иерусалима, как во дни древние и как в лета прежние.
MAL|3|5|И приду к вам для суда и буду скорым обличителем чародеев и прелюбодеев и тех, которые клянутся ложно и удерживают плату у наемника, притесняют вдову и сироту, и отталкивают пришельца, и Меня не боятся, говорит Господь Саваоф.
MAL|3|6|Ибо Я – Господь, Я не изменяюсь; посему вы, сыны Иакова, не уничтожились.
MAL|3|7|Со дней отцов ваших вы отступили от уставов Моих и не соблюдаете их; обратитесь ко Мне, и я обращусь к вам, говорит Господь Саваоф. Вы скажете: "как нам обратиться?"
MAL|3|8|Можно ли человеку обкрадывать Бога? А вы обкрадываете Меня. Скажете: "чем обкрадываем мы Тебя?" Десятиною и приношениями.
MAL|3|9|Проклятием вы прокляты, потому что вы – весь народ – обкрадываете Меня.
MAL|3|10|Принесите все десятины в дом хранилища, чтобы в доме Моем была пища, и хотя в этом испытайте Меня, говорит Господь Саваоф: не открою ли Я для вас отверстий небесных и не изолью ли на вас благословения до избытка?
MAL|3|11|Я для вас запрещу пожирающим истреблять у вас плоды земные, и виноградная лоза на поле у вас не лишится плодов своих, говорит Господь Саваоф.
MAL|3|12|И блаженными называть будут вас все народы, потому что вы будете землею вожделенною, говорит Господь Саваоф.
MAL|3|13|Дерзостны предо Мною слова ваши, говорит Господь. Вы скажете: "что мы говорим против Тебя?"
MAL|3|14|Вы говорите: "тщетно служение Богу, и что пользы, что мы соблюдали постановления Его и ходили в печальной одежде пред лицем Господа Саваофа?
MAL|3|15|И ныне мы считаем надменных счастливыми: лучше устраивают себя делающие беззакония, и хотя искушают Бога, но остаются целы".
MAL|3|16|Но боящиеся Бога говорят друг другу: "внимает Господь и слышит это, и пред лицем Его пишется памятная книга о боящихся Господа и чтущих имя Его".
MAL|3|17|И они будут Моими, говорит Господь Саваоф, собственностью Моею в тот день, который Я соделаю, и буду миловать их, как милует человек сына своего, служащего ему.
MAL|3|18|И тогда снова увидите различие между праведником и нечестивым, между служащим Богу и не служащим Ему.
MAL|4|1|Ибо вот, придет день, пылающий как печь; тогда все надменные и поступающие нечестиво будут как солома, и попалит их грядущий день, говорит Господь Саваоф, так что не оставит у них ни корня, ни ветвей.
MAL|4|2|А для вас, благоговеющие пред именем Моим, взойдет Солнце правды и исцеление в лучах Его, и вы выйдете и взыграете, как тельцы упитанные;
MAL|4|3|и будете попирать нечестивых, ибо они будут прахом под стопами ног ваших в тот день, который Я соделаю, говорит Господь Саваоф.
MAL|4|4|Помните закон Моисея, раба Моего, который Я заповедал ему на Хориве для всего Израиля, равно как и правила и уставы.
MAL|4|5|Вот, Я пошлю к вам Илию пророка пред наступлением дня Господня, великого и страшного.
MAL|4|6|И он обратит сердца отцов к детям и сердца детей к отцам их, чтобы Я, придя, не поразил земли проклятием.
