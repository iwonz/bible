2CHR|1|1|Solomon son of David established himself firmly over his kingdom, for the LORD his God was with him and made him exceedingly great.
2CHR|1|2|Then Solomon spoke to all Israel-to the commanders of thousands and commanders of hundreds, to the judges and to all the leaders in Israel, the heads of families-
2CHR|1|3|and Solomon and the whole assembly went to the high place at Gibeon, for God's Tent of Meeting was there, which Moses the LORD's servant had made in the desert.
2CHR|1|4|Now David had brought up the ark of God from Kiriath Jearim to the place he had prepared for it, because he had pitched a tent for it in Jerusalem.
2CHR|1|5|But the bronze altar that Bezalel son of Uri, the son of Hur, had made was in Gibeon in front of the tabernacle of the LORD; so Solomon and the assembly inquired of him there.
2CHR|1|6|Solomon went up to the bronze altar before the LORD in the Tent of Meeting and offered a thousand burnt offerings on it.
2CHR|1|7|That night God appeared to Solomon and said to him, "Ask for whatever you want me to give you."
2CHR|1|8|Solomon answered God, "You have shown great kindness to David my father and have made me king in his place.
2CHR|1|9|Now, LORD God, let your promise to my father David be confirmed, for you have made me king over a people who are as numerous as the dust of the earth.
2CHR|1|10|Give me wisdom and knowledge, that I may lead this people, for who is able to govern this great people of yours?"
2CHR|1|11|God said to Solomon, "Since this is your heart's desire and you have not asked for wealth, riches or honor, nor for the death of your enemies, and since you have not asked for a long life but for wisdom and knowledge to govern my people over whom I have made you king,
2CHR|1|12|therefore wisdom and knowledge will be given you. And I will also give you wealth, riches and honor, such as no king who was before you ever had and none after you will have."
2CHR|1|13|Then Solomon went to Jerusalem from the high place at Gibeon, from before the Tent of Meeting. And he reigned over Israel.
2CHR|1|14|Solomon accumulated chariots and horses; he had fourteen hundred chariots and twelve thousand horses, which he kept in the chariot cities and also with him in Jerusalem.
2CHR|1|15|The king made silver and gold as common in Jerusalem as stones, and cedar as plentiful as sycamore-fig trees in the foothills.
2CHR|1|16|Solomon's horses were imported from Egypt and from Kue - the royal merchants purchased them from Kue.
2CHR|1|17|They imported a chariot from Egypt for six hundred shekels of silver, and a horse for a hundred and fifty. They also exported them to all the kings of the Hittites and of the Arameans.
2CHR|2|1|Solomon gave orders to build a temple for the Name of the LORD and a royal palace for himself.
2CHR|2|2|He conscripted seventy thousand men as carriers and eighty thousand as stonecutters in the hills and thirty-six hundred as foremen over them.
2CHR|2|3|Solomon sent this message to Hiram king of Tyre: "Send me cedar logs as you did for my father David when you sent him cedar to build a palace to live in.
2CHR|2|4|Now I am about to build a temple for the Name of the LORD my God and to dedicate it to him for burning fragrant incense before him, for setting out the consecrated bread regularly, and for making burnt offerings every morning and evening and on Sabbaths and New Moons and at the appointed feasts of the LORD our God. This is a lasting ordinance for Israel.
2CHR|2|5|"The temple I am going to build will be great, because our God is greater than all other gods.
2CHR|2|6|But who is able to build a temple for him, since the heavens, even the highest heavens, cannot contain him? Who then am I to build a temple for him, except as a place to burn sacrifices before him?
2CHR|2|7|"Send me, therefore, a man skilled to work in gold and silver, bronze and iron, and in purple, crimson and blue yarn, and experienced in the art of engraving, to work in Judah and Jerusalem with my skilled craftsmen, whom my father David provided.
2CHR|2|8|"Send me also cedar, pine and algum logs from Lebanon, for I know that your men are skilled in cutting timber there. My men will work with yours
2CHR|2|9|to provide me with plenty of lumber, because the temple I build must be large and magnificent.
2CHR|2|10|I will give your servants, the woodsmen who cut the timber, twenty thousand cors of ground wheat, twenty thousand cors of barley, twenty thousand baths of wine and twenty thousand baths of olive oil."
2CHR|2|11|Hiram king of Tyre replied by letter to Solomon: "Because the LORD loves his people, he has made you their king."
2CHR|2|12|And Hiram added: "Praise be to the LORD, the God of Israel, who made heaven and earth! He has given King David a wise son, endowed with intelligence and discernment, who will build a temple for the LORD and a palace for himself.
2CHR|2|13|"I am sending you Huram-Abi, a man of great skill,
2CHR|2|14|whose mother was from Dan and whose father was from Tyre. He is trained to work in gold and silver, bronze and iron, stone and wood, and with purple and blue and crimson yarn and fine linen. He is experienced in all kinds of engraving and can execute any design given to him. He will work with your craftsmen and with those of my Lord, David your father.
2CHR|2|15|"Now let my Lord send his servants the wheat and barley and the olive oil and wine he promised,
2CHR|2|16|and we will cut all the logs from Lebanon that you need and will float them in rafts by sea down to Joppa. You can then take them up to Jerusalem."
2CHR|2|17|Solomon took a census of all the aliens who were in Israel, after the census his father David had taken; and they were found to be 153,600.
2CHR|2|18|He assigned 70,000 of them to be carriers and 80,000 to be stonecutters in the hills, with 3,600 foremen over them to keep the people working.
2CHR|3|1|Then Solomon began to build the temple of the LORD in Jerusalem on Mount Moriah, where the LORD had appeared to his father David. It was on the threshing floor of Araunah the Jebusite, the place provided by David.
2CHR|3|2|He began building on the second day of the second month in the fourth year of his reign.
2CHR|3|3|The foundation Solomon laid for building the temple of God was sixty cubits long and twenty cubits wide (using the cubit of the old standard).
2CHR|3|4|The portico at the front of the temple was twenty cubits long across the width of the building and twenty cubits high. He overlaid the inside with pure gold.
2CHR|3|5|He paneled the main hall with pine and covered it with fine gold and decorated it with palm tree and chain designs.
2CHR|3|6|He adorned the temple with precious stones. And the gold he used was gold of Parvaim.
2CHR|3|7|He overlaid the ceiling beams, doorframes, walls and doors of the temple with gold, and he carved cherubim on the walls.
2CHR|3|8|He built the Most Holy Place, its length corresponding to the width of the temple-twenty cubits long and twenty cubits wide. He overlaid the inside with six hundred talents of fine gold.
2CHR|3|9|The gold nails weighed fifty shekels. He also overlaid the upper parts with gold.
2CHR|3|10|In the Most Holy Place he made a pair of sculptured cherubim and overlaid them with gold.
2CHR|3|11|The total wingspan of the cherubim was twenty cubits. One wing of the first cherub was five cubits long and touched the temple wall, while its other wing, also five cubits long, touched the wing of the other cherub.
2CHR|3|12|Similarly one wing of the second cherub was five cubits long and touched the other temple wall, and its other wing, also five cubits long, touched the wing of the first cherub.
2CHR|3|13|The wings of these cherubim extended twenty cubits. They stood on their feet, facing the main hall.
2CHR|3|14|He made the curtain of blue, purple and crimson yarn and fine linen, with cherubim worked into it.
2CHR|3|15|In the front of the temple he made two pillars, which together were thirty-five cubits long, each with a capital on top measuring five cubits.
2CHR|3|16|He made interwoven chains and put them on top of the pillars. He also made a hundred pomegranates and attached them to the chains.
2CHR|3|17|He erected the pillars in the front of the temple, one to the south and one to the north. The one to the south he named Jakin and the one to the north Boaz.
2CHR|4|1|He made a bronze altar twenty cubits long, twenty cubits wide and ten cubits high.
2CHR|4|2|He made the Sea of cast metal, circular in shape, measuring ten cubits from rim to rim and five cubits high. It took a line of thirty cubits to measure around it.
2CHR|4|3|Below the rim, figures of bulls encircled it-ten to a cubit. The bulls were cast in two rows in one piece with the Sea.
2CHR|4|4|The Sea stood on twelve bulls, three facing north, three facing west, three facing south and three facing east. The Sea rested on top of them, and their hindquarters were toward the center.
2CHR|4|5|It was a handbreadth in thickness, and its rim was like the rim of a cup, like a lily blossom. It held three thousand baths.
2CHR|4|6|He then made ten basins for washing and placed five on the south side and five on the north. In them the things to be used for the burnt offerings were rinsed, but the Sea was to be used by the priests for washing.
2CHR|4|7|He made ten gold lampstands according to the specifications for them and placed them in the temple, five on the south side and five on the north.
2CHR|4|8|He made ten tables and placed them in the temple, five on the south side and five on the north. He also made a hundred gold sprinkling bowls.
2CHR|4|9|He made the courtyard of the priests, and the large court and the doors for the court, and overlaid the doors with bronze.
2CHR|4|10|He placed the Sea on the south side, at the southeast corner.
2CHR|4|11|He also made the pots and shovels and sprinkling bowls. So Huram finished the work he had undertaken for King Solomon in the temple of God:
2CHR|4|12|the two pillars; the two bowl-shaped capitals on top of the pillars; the two sets of network decorating the two bowl-shaped capitals on top of the pillars;
2CHR|4|13|the four hundred pomegranates for the two sets of network (two rows of pomegranates for each network, decorating the bowl-shaped capitals on top of the pillars);
2CHR|4|14|the stands with their basins;
2CHR|4|15|the Sea and the twelve bulls under it;
2CHR|4|16|the pots, shovels, meat forks and all related articles. All the objects that Huram-Abi made for King Solomon for the temple of the LORD were of polished bronze.
2CHR|4|17|The king had them cast in clay molds in the plain of the Jordan between Succoth and Zarethan.
2CHR|4|18|All these things that Solomon made amounted to so much that the weight of the bronze was not determined.
2CHR|4|19|Solomon also made all the furnishings that were in God's temple: the golden altar; the tables on which was the bread of the Presence;
2CHR|4|20|the lampstands of pure gold with their lamps, to burn in front of the inner sanctuary as prescribed;
2CHR|4|21|the gold floral work and lamps and tongs (they were solid gold);
2CHR|4|22|the pure gold wick trimmers, sprinkling bowls, dishes and censers; and the gold doors of the temple: the inner doors to the Most Holy Place and the doors of the main hall.
2CHR|5|1|When all the work Solomon had done for the temple of the LORD was finished, he brought in the things his father David had dedicated-the silver and gold and all the furnishings-and he placed them in the treasuries of God's temple.
2CHR|5|2|Then Solomon summoned to Jerusalem the elders of Israel, all the heads of the tribes and the chiefs of the Israelite families, to bring up the ark of the LORD's covenant from Zion, the City of David.
2CHR|5|3|And all the men of Israel came together to the king at the time of the festival in the seventh month.
2CHR|5|4|When all the elders of Israel had arrived, the Levites took up the ark,
2CHR|5|5|and they brought up the ark and the Tent of Meeting and all the sacred furnishings in it. The priests, who were Levites, carried them up;
2CHR|5|6|and King Solomon and the entire assembly of Israel that had gathered about him were before the ark, sacrificing so many sheep and cattle that they could not be recorded or counted.
2CHR|5|7|The priests then brought the ark of the LORD's covenant to its place in the inner sanctuary of the temple, the Most Holy Place, and put it beneath the wings of the cherubim.
2CHR|5|8|The cherubim spread their wings over the place of the ark and covered the ark and its carrying poles.
2CHR|5|9|These poles were so long that their ends, extending from the ark, could be seen from in front of the inner sanctuary, but not from outside the Holy Place; and they are still there today.
2CHR|5|10|There was nothing in the ark except the two tablets that Moses had placed in it at Horeb, where the LORD made a covenant with the Israelites after they came out of Egypt.
2CHR|5|11|The priests then withdrew from the Holy Place. All the priests who were there had consecrated themselves, regardless of their divisions.
2CHR|5|12|All the Levites who were musicians-Asaph, Heman, Jeduthun and their sons and relatives-stood on the east side of the altar, dressed in fine linen and playing cymbals, harps and lyres. They were accompanied by 120 priests sounding trumpets.
2CHR|5|13|The trumpeters and singers joined in unison, as with one voice, to give praise and thanks to the LORD. Accompanied by trumpets, cymbals and other instruments, they raised their voices in praise to the LORD and sang: "He is good; his love endures forever." Then the temple of the LORD was filled with a cloud,
2CHR|5|14|and the priests could not perform their service because of the cloud, for the glory of the LORD filled the temple of God.
2CHR|6|1|Then Solomon said, "The LORD has said that he would dwell in a dark cloud;
2CHR|6|2|I have built a magnificent temple for you, a place for you to dwell forever."
2CHR|6|3|While the whole assembly of Israel was standing there, the king turned around and blessed them.
2CHR|6|4|Then he said: "Praise be to the LORD, the God of Israel, who with his hands has fulfilled what he promised with his mouth to my father David. For he said,
2CHR|6|5|'Since the day I brought my people out of Egypt, I have not chosen a city in any tribe of Israel to have a temple built for my Name to be there, nor have I chosen anyone to be the leader over my people Israel.
2CHR|6|6|But now I have chosen Jerusalem for my Name to be there, and I have chosen David to rule my people Israel.'
2CHR|6|7|"My father David had it in his heart to build a temple for the Name of the LORD, the God of Israel.
2CHR|6|8|But the LORD said to my father David, 'Because it was in your heart to build a temple for my Name, you did well to have this in your heart.
2CHR|6|9|Nevertheless, you are not the one to build the temple, but your son, who is your own flesh and blood-he is the one who will build the temple for my Name.'
2CHR|6|10|"The LORD has kept the promise he made. I have succeeded David my father and now I sit on the throne of Israel, just as the LORD promised, and I have built the temple for the Name of the LORD, the God of Israel.
2CHR|6|11|There I have placed the ark, in which is the covenant of the LORD that he made with the people of Israel."
2CHR|6|12|Then Solomon stood before the altar of the LORD in front of the whole assembly of Israel and spread out his hands.
2CHR|6|13|Now he had made a bronze platform, five cubits long, five cubits wide and three cubits high, and had placed it in the center of the outer court. He stood on the platform and then knelt down before the whole assembly of Israel and spread out his hands toward heaven.
2CHR|6|14|He said: "O LORD, God of Israel, there is no God like you in heaven or on earth-you who keep your covenant of love with your servants who continue wholeheartedly in your way.
2CHR|6|15|You have kept your promise to your servant David my father; with your mouth you have promised and with your hand you have fulfilled it-as it is today.
2CHR|6|16|"Now LORD, God of Israel, keep for your servant David my father the promises you made to him when you said, 'You shall never fail to have a man to sit before me on the throne of Israel, if only your sons are careful in all they do to walk before me according to my law, as you have done.'
2CHR|6|17|And now, O LORD, God of Israel, let your word that you promised your servant David come true.
2CHR|6|18|"But will God really dwell on earth with men? The heavens, even the highest heavens, cannot contain you. How much less this temple I have built!
2CHR|6|19|Yet give attention to your servant's prayer and his plea for mercy, O LORD my God. Hear the cry and the prayer that your servant is praying in your presence.
2CHR|6|20|May your eyes be open toward this temple day and night, this place of which you said you would put your Name there. May you hear the prayer your servant prays toward this place.
2CHR|6|21|Hear the supplications of your servant and of your people Israel when they pray toward this place. Hear from heaven, your dwelling place; and when you hear, forgive.
2CHR|6|22|"When a man wrongs his neighbor and is required to take an oath and he comes and swears the oath before your altar in this temple,
2CHR|6|23|then hear from heaven and act. Judge between your servants, repaying the guilty by bringing down on his own head what he has done. Declare the innocent not guilty and so establish his innocence.
2CHR|6|24|"When your people Israel have been defeated by an enemy because they have sinned against you and when they turn back and confess your name, praying and making supplication before you in this temple,
2CHR|6|25|then hear from heaven and forgive the sin of your people Israel and bring them back to the land you gave to them and their fathers.
2CHR|6|26|"When the heavens are shut up and there is no rain because your people have sinned against you, and when they pray toward this place and confess your name and turn from their sin because you have afflicted them,
2CHR|6|27|then hear from heaven and forgive the sin of your servants, your people Israel. Teach them the right way to live, and send rain on the land you gave your people for an inheritance.
2CHR|6|28|"When famine or plague comes to the land, or blight or mildew, locusts or grasshoppers, or when enemies besiege them in any of their cities, whatever disaster or disease may come,
2CHR|6|29|and when a prayer or plea is made by any of your people Israel-each one aware of his afflictions and pains, and spreading out his hands toward this temple-
2CHR|6|30|then hear from heaven, your dwelling place. Forgive, and deal with each man according to all he does, since you know his heart (for you alone know the hearts of men),
2CHR|6|31|so that they will fear you and walk in your ways all the time they live in the land you gave our fathers.
2CHR|6|32|"As for the foreigner who does not belong to your people Israel but has come from a distant land because of your great name and your mighty hand and your outstretched arm-when he comes and prays toward this temple,
2CHR|6|33|then hear from heaven, your dwelling place, and do whatever the foreigner asks of you, so that all the peoples of the earth may know your name and fear you, as do your own people Israel, and may know that this house I have built bears your Name.
2CHR|6|34|"When your people go to war against their enemies, wherever you send them, and when they pray to you toward this city you have chosen and the temple I have built for your Name,
2CHR|6|35|then hear from heaven their prayer and their plea, and uphold their cause.
2CHR|6|36|"When they sin against you-for there is no one who does not sin-and you become angry with them and give them over to the enemy, who takes them captive to a land far away or near;
2CHR|6|37|and if they have a change of heart in the land where they are held captive, and repent and plead with you in the land of their captivity and say, 'We have sinned, we have done wrong and acted wickedly';
2CHR|6|38|and if they turn back to you with all their heart and soul in the land of their captivity where they were taken, and pray toward the land you gave their fathers, toward the city you have chosen and toward the temple I have built for your Name;
2CHR|6|39|then from heaven, your dwelling place, hear their prayer and their pleas, and uphold their cause. And forgive your people, who have sinned against you.
2CHR|6|40|"Now, my God, may your eyes be open and your ears attentive to the prayers offered in this place.
2CHR|6|41|"Now arise, O LORD God, and come to your resting place, you and the ark of your might. May your priests, O LORD God, be clothed with salvation, may your saints rejoice in your goodness.
2CHR|6|42|O LORD God, do not reject your anointed one. Remember the great love promised to David your servant."
2CHR|7|1|When Solomon finished praying, fire came down from heaven and consumed the burnt offering and the sacrifices, and the glory of the LORD filled the temple.
2CHR|7|2|The priests could not enter the temple of the LORD because the glory of the LORD filled it.
2CHR|7|3|When all the Israelites saw the fire coming down and the glory of the LORD above the temple, they knelt on the pavement with their faces to the ground, and they worshiped and gave thanks to the LORD, saying, "He is good; his love endures forever."
2CHR|7|4|Then the king and all the people offered sacrifices before the LORD.
2CHR|7|5|And King Solomon offered a sacrifice of twenty-two thousand head of cattle and a hundred and twenty thousand sheep and goats. So the king and all the people dedicated the temple of God.
2CHR|7|6|The priests took their positions, as did the Levites with the LORD's musical instruments, which King David had made for praising the LORD and which were used when he gave thanks, saying, "His love endures forever." Opposite the Levites, the priests blew their trumpets, and all the Israelites were standing.
2CHR|7|7|Solomon consecrated the middle part of the courtyard in front of the temple of the LORD, and there he offered burnt offerings and the fat of the fellowship offerings, because the bronze altar he had made could not hold the burnt offerings, the grain offerings and the fat portions.
2CHR|7|8|So Solomon observed the festival at that time for seven days, and all Israel with him-a vast assembly, people from Lebo Hamath to the Wadi of Egypt.
2CHR|7|9|On the eighth day they held an assembly, for they had celebrated the dedication of the altar for seven days and the festival for seven days more.
2CHR|7|10|On the twenty-third day of the seventh month he sent the people to their homes, joyful and glad in heart for the good things the LORD had done for David and Solomon and for his people Israel.
2CHR|7|11|When Solomon had finished the temple of the LORD and the royal palace, and had succeeded in carrying out all he had in mind to do in the temple of the LORD and in his own palace,
2CHR|7|12|the LORD appeared to him at night and said: "I have heard your prayer and have chosen this place for myself as a temple for sacrifices.
2CHR|7|13|"When I shut up the heavens so that there is no rain, or command locusts to devour the land or send a plague among my people,
2CHR|7|14|if my people, who are called by my name, will humble themselves and pray and seek my face and turn from their wicked ways, then will I hear from heaven and will forgive their sin and will heal their land.
2CHR|7|15|Now my eyes will be open and my ears attentive to the prayers offered in this place.
2CHR|7|16|I have chosen and consecrated this temple so that my Name may be there forever. My eyes and my heart will always be there.
2CHR|7|17|"As for you, if you walk before me as David your father did, and do all I command, and observe my decrees and laws,
2CHR|7|18|I will establish your royal throne, as I covenanted with David your father when I said, 'You shall never fail to have a man to rule over Israel.'
2CHR|7|19|"But if you turn away and forsake the decrees and commands I have given you and go off to serve other gods and worship them,
2CHR|7|20|then I will uproot Israel from my land, which I have given them, and will reject this temple I have consecrated for my Name. I will make it a byword and an object of ridicule among all peoples.
2CHR|7|21|And though this temple is now so imposing, all who pass by will be appalled and say, 'Why has the LORD done such a thing to this land and to this temple?'
2CHR|7|22|People will answer, 'Because they have forsaken the LORD, the God of their fathers, who brought them out of Egypt, and have embraced other gods, worshiping and serving them-that is why he brought all this disaster on them.'"
2CHR|8|1|At the end of twenty years, during which Solomon built the temple of the LORD and his own palace,
2CHR|8|2|Solomon rebuilt the villages that Hiram had given him, and settled Israelites in them.
2CHR|8|3|Solomon then went to Hamath Zobah and captured it.
2CHR|8|4|He also built up Tadmor in the desert and all the store cities he had built in Hamath.
2CHR|8|5|He rebuilt Upper Beth Horon and Lower Beth Horon as fortified cities, with walls and with gates and bars,
2CHR|8|6|as well as Baalath and all his store cities, and all the cities for his chariots and for his horses -whatever he desired to build in Jerusalem, in Lebanon and throughout all the territory he ruled.
2CHR|8|7|All the people left from the Hittites, Amorites, Perizzites, Hivites and Jebusites (these peoples were not Israelites),
2CHR|8|8|that is, their descendants remaining in the land, whom the Israelites had not destroyed-these Solomon conscripted for his slave labor force, as it is to this day.
2CHR|8|9|But Solomon did not make slaves of the Israelites for his work; they were his fighting men, commanders of his captains, and commanders of his chariots and charioteers.
2CHR|8|10|They were also King Solomon's chief officials-two hundred and fifty officials supervising the men.
2CHR|8|11|Solomon brought Pharaoh's daughter up from the City of David to the palace he had built for her, for he said, "My wife must not live in the palace of David king of Israel, because the places the ark of the LORD has entered are holy."
2CHR|8|12|On the altar of the LORD that he had built in front of the portico, Solomon sacrificed burnt offerings to the LORD,
2CHR|8|13|according to the daily requirement for offerings commanded by Moses for Sabbaths, New Moons and the three annual feasts-the Feast of Unleavened Bread, the Feast of Weeks and the Feast of Tabernacles.
2CHR|8|14|In keeping with the ordinance of his father David, he appointed the divisions of the priests for their duties, and the Levites to lead the praise and to assist the priests according to each day's requirement. He also appointed the gatekeepers by divisions for the various gates, because this was what David the man of God had ordered.
2CHR|8|15|They did not deviate from the king's commands to the priests or to the Levites in any matter, including that of the treasuries.
2CHR|8|16|All Solomon's work was carried out, from the day the foundation of the temple of the LORD was laid until its completion. So the temple of the LORD was finished.
2CHR|8|17|Then Solomon went to Ezion Geber and Elath on the coast of Edom.
2CHR|8|18|And Hiram sent him ships commanded by his own officers, men who knew the sea. These, with Solomon's men, sailed to Ophir and brought back four hundred and fifty talents of gold, which they delivered to King Solomon.
2CHR|9|1|When the queen of Sheba heard of Solomon's fame, she came to Jerusalem to test him with hard questions. Arriving with a very great caravan-with camels carrying spices, large quantities of gold, and precious stones-she came to Solomon and talked with him about all she had on her mind.
2CHR|9|2|Solomon answered all her questions; nothing was too hard for him to explain to her.
2CHR|9|3|When the queen of Sheba saw the wisdom of Solomon, as well as the palace he had built,
2CHR|9|4|the food on his table, the seating of his officials, the attending servants in their robes, the cupbearers in their robes and the burnt offerings he made at the temple of the LORD, she was overwhelmed.
2CHR|9|5|She said to the king, "The report I heard in my own country about your achievements and your wisdom is true.
2CHR|9|6|But I did not believe what they said until I came and saw with my own eyes. Indeed, not even half the greatness of your wisdom was told me; you have far exceeded the report I heard.
2CHR|9|7|How happy your men must be! How happy your officials, who continually stand before you and hear your wisdom!
2CHR|9|8|Praise be to the LORD your God, who has delighted in you and placed you on his throne as king to rule for the LORD your God. Because of the love of your God for Israel and his desire to uphold them forever, he has made you king over them, to maintain justice and righteousness."
2CHR|9|9|Then she gave the king 120 talents of gold, large quantities of spices, and precious stones. There had never been such spices as those the queen of Sheba gave to King Solomon.
2CHR|9|10|(The men of Hiram and the men of Solomon brought gold from Ophir; they also brought algumwood and precious stones.
2CHR|9|11|The king used the algumwood to make steps for the temple of the LORD and for the royal palace, and to make harps and lyres for the musicians. Nothing like them had ever been seen in Judah.)
2CHR|9|12|King Solomon gave the queen of Sheba all she desired and asked for; he gave her more than she had brought to him. Then she left and returned with her retinue to her own country.
2CHR|9|13|The weight of the gold that Solomon received yearly was 666 talents,
2CHR|9|14|not including the revenues brought in by merchants and traders. Also all the kings of Arabia and the governors of the land brought gold and silver to Solomon.
2CHR|9|15|King Solomon made two hundred large shields of hammered gold; six hundred bekas of hammered gold went into each shield.
2CHR|9|16|He also made three hundred small shields of hammered gold, with three hundred bekas of gold in each shield. The king put them in the Palace of the Forest of Lebanon.
2CHR|9|17|Then the king made a great throne inlaid with ivory and overlaid with pure gold.
2CHR|9|18|The throne had six steps, and a footstool of gold was attached to it. On both sides of the seat were armrests, with a lion standing beside each of them.
2CHR|9|19|Twelve lions stood on the six steps, one at either end of each step. Nothing like it had ever been made for any other kingdom.
2CHR|9|20|All King Solomon's goblets were gold, and all the household articles in the Palace of the Forest of Lebanon were pure gold. Nothing was made of silver, because silver was considered of little value in Solomon's day.
2CHR|9|21|The king had a fleet of trading ships manned by Hiram's men. Once every three years it returned, carrying gold, silver and ivory, and apes and baboons.
2CHR|9|22|King Solomon was greater in riches and wisdom than all the other kings of the earth.
2CHR|9|23|All the kings of the earth sought audience with Solomon to hear the wisdom God had put in his heart.
2CHR|9|24|Year after year, everyone who came brought a gift-articles of silver and gold, and robes, weapons and spices, and horses and mules.
2CHR|9|25|Solomon had four thousand stalls for horses and chariots, and twelve thousand horses, which he kept in the chariot cities and also with him in Jerusalem.
2CHR|9|26|He ruled over all the kings from the River to the land of the Philistines, as far as the border of Egypt.
2CHR|9|27|The king made silver as common in Jerusalem as stones, and cedar as plentiful as sycamore-fig trees in the foothills.
2CHR|9|28|Solomon's horses were imported from Egypt and from all other countries.
2CHR|9|29|As for the other events of Solomon's reign, from beginning to end, are they not written in the records of Nathan the prophet, in the prophecy of Ahijah the Shilonite and in the visions of Iddo the seer concerning Jeroboam son of Nebat?
2CHR|9|30|Solomon reigned in Jerusalem over all Israel forty years.
2CHR|9|31|Then he rested with his fathers and was buried in the city of David his father. And Rehoboam his son succeeded him as king.
2CHR|10|1|Rehoboam went to Shechem, for all the Israelites had gone there to make him king.
2CHR|10|2|When Jeroboam son of Nebat heard this (he was in Egypt, where he had fled from King Solomon), he returned from Egypt.
2CHR|10|3|So they sent for Jeroboam, and he and all Israel went to Rehoboam and said to him:
2CHR|10|4|"Your father put a heavy yoke on us, but now lighten the harsh labor and the heavy yoke he put on us, and we will serve you."
2CHR|10|5|Rehoboam answered, "Come back to me in three days." So the people went away.
2CHR|10|6|Then King Rehoboam consulted the elders who had served his father Solomon during his lifetime. "How would you advise me to answer these people?" he asked.
2CHR|10|7|They replied, "If you will be kind to these people and please them and give them a favorable answer, they will always be your servants."
2CHR|10|8|But Rehoboam rejected the advice the elders gave him and consulted the young men who had grown up with him and were serving him.
2CHR|10|9|He asked them, "What is your advice? How should we answer these people who say to me, 'Lighten the yoke your father put on us'?"
2CHR|10|10|The young men who had grown up with him replied, "Tell the people who have said to you, 'Your father put a heavy yoke on us, but make our yoke lighter'-tell them, 'My little finger is thicker than my father's waist.
2CHR|10|11|My father laid on you a heavy yoke; I will make it even heavier. My father scourged you with whips; I will scourge you with scorpions.'"
2CHR|10|12|Three days later Jeroboam and all the people returned to Rehoboam, as the king had said, "Come back to me in three days."
2CHR|10|13|The king answered them harshly. Rejecting the advice of the elders,
2CHR|10|14|he followed the advice of the young men and said, "My father made your yoke heavy; I will make it even heavier. My father scourged you with whips; I will scourge you with scorpions."
2CHR|10|15|So the king did not listen to the people, for this turn of events was from God, to fulfill the word the LORD had spoken to Jeroboam son of Nebat through Ahijah the Shilonite.
2CHR|10|16|When all Israel saw that the king refused to listen to them, they answered the king: "What share do we have in David, what part in Jesse's son? To your tents, O Israel! Look after your own house, O David!" So all the Israelites went home.
2CHR|10|17|But as for the Israelites who were living in the towns of Judah, Rehoboam still ruled over them.
2CHR|10|18|King Rehoboam sent out Adoniram, who was in charge of forced labor, but the Israelites stoned him to death. King Rehoboam, however, managed to get into his chariot and escape to Jerusalem.
2CHR|10|19|So Israel has been in rebellion against the house of David to this day.
2CHR|11|1|When Rehoboam arrived in Jerusalem, he mustered the house of Judah and Benjamin-a hundred and eighty thousand fighting men-to make war against Israel and to regain the kingdom for Rehoboam.
2CHR|11|2|But this word of the LORD came to Shemaiah the man of God:
2CHR|11|3|"Say to Rehoboam son of Solomon king of Judah and to all the Israelites in Judah and Benjamin,
2CHR|11|4|'This is what the LORD says: Do not go up to fight against your brothers. Go home, every one of you, for this is my doing.'" So they obeyed the words of the LORD and turned back from marching against Jeroboam.
2CHR|11|5|Rehoboam lived in Jerusalem and built up towns for defense in Judah:
2CHR|11|6|Bethlehem, Etam, Tekoa,
2CHR|11|7|Beth Zur, Soco, Adullam,
2CHR|11|8|Gath, Mareshah, Ziph,
2CHR|11|9|Adoraim, Lachish, Azekah,
2CHR|11|10|Zorah, Aijalon and Hebron. These were fortified cities in Judah and Benjamin.
2CHR|11|11|He strengthened their defenses and put commanders in them, with supplies of food, olive oil and wine.
2CHR|11|12|He put shields and spears in all the cities, and made them very strong. So Judah and Benjamin were his.
2CHR|11|13|The priests and Levites from all their districts throughout Israel sided with him.
2CHR|11|14|The Levites even abandoned their pasturelands and property, and came to Judah and Jerusalem because Jeroboam and his sons had rejected them as priests of the LORD.
2CHR|11|15|And he appointed his own priests for the high places and for the goat and calf idols he had made.
2CHR|11|16|Those from every tribe of Israel who set their hearts on seeking the LORD, the God of Israel, followed the Levites to Jerusalem to offer sacrifices to the LORD, the God of their fathers.
2CHR|11|17|They strengthened the kingdom of Judah and supported Rehoboam son of Solomon three years, walking in the ways of David and Solomon during this time.
2CHR|11|18|Rehoboam married Mahalath, who was the daughter of David's son Jerimoth and of Abihail, the daughter of Jesse's son Eliab.
2CHR|11|19|She bore him sons: Jeush, Shemariah and Zaham.
2CHR|11|20|Then he married Maacah daughter of Absalom, who bore him Abijah, Attai, Ziza and Shelomith.
2CHR|11|21|Rehoboam loved Maacah daughter of Absalom more than any of his other wives and concubines. In all, he had eighteen wives and sixty concubines, twenty-eight sons and sixty daughters.
2CHR|11|22|Rehoboam appointed Abijah son of Maacah to be the chief prince among his brothers, in order to make him king.
2CHR|11|23|He acted wisely, dispersing some of his sons throughout the districts of Judah and Benjamin, and to all the fortified cities. He gave them abundant provisions and took many wives for them.
2CHR|12|1|After Rehoboam's position as king was established and he had become strong, he and all Israel with him abandoned the law of the LORD.
2CHR|12|2|Because they had been unfaithful to the LORD, Shishak king of Egypt attacked Jerusalem in the fifth year of King Rehoboam.
2CHR|12|3|With twelve hundred chariots and sixty thousand horsemen and the innumerable troops of Libyans, Sukkites and Cushites that came with him from Egypt,
2CHR|12|4|he captured the fortified cities of Judah and came as far as Jerusalem.
2CHR|12|5|Then the prophet Shemaiah came to Rehoboam and to the leaders of Judah who had assembled in Jerusalem for fear of Shishak, and he said to them, "This is what the LORD says, 'You have abandoned me; therefore, I now abandon you to Shishak.'"
2CHR|12|6|The leaders of Israel and the king humbled themselves and said, "The LORD is just."
2CHR|12|7|When the LORD saw that they humbled themselves, this word of the LORD came to Shemaiah: "Since they have humbled themselves, I will not destroy them but will soon give them deliverance. My wrath will not be poured out on Jerusalem through Shishak.
2CHR|12|8|They will, however, become subject to him, so that they may learn the difference between serving me and serving the kings of other lands."
2CHR|12|9|When Shishak king of Egypt attacked Jerusalem, he carried off the treasures of the temple of the LORD and the treasures of the royal palace. He took everything, including the gold shields Solomon had made.
2CHR|12|10|So King Rehoboam made bronze shields to replace them and assigned these to the commanders of the guard on duty at the entrance to the royal palace.
2CHR|12|11|Whenever the king went to the LORD's temple, the guards went with him, bearing the shields, and afterward they returned them to the guardroom.
2CHR|12|12|Because Rehoboam humbled himself, the LORD's anger turned from him, and he was not totally destroyed. Indeed, there was some good in Judah.
2CHR|12|13|King Rehoboam established himself firmly in Jerusalem and continued as king. He was forty-one years old when he became king, and he reigned seventeen years in Jerusalem, the city the LORD had chosen out of all the tribes of Israel in which to put his Name. His mother's name was Naamah; she was an Ammonite.
2CHR|12|14|He did evil because he had not set his heart on seeking the LORD.
2CHR|12|15|As for the events of Rehoboam's reign, from beginning to end, are they not written in the records of Shemaiah the prophet and of Iddo the seer that deal with genealogies? There was continual warfare between Rehoboam and Jeroboam.
2CHR|12|16|Rehoboam rested with his fathers and was buried in the City of David. And Abijah his son succeeded him as king.
2CHR|13|1|In the eighteenth year of the reign of Jeroboam, Abijah became king of Judah,
2CHR|13|2|and he reigned in Jerusalem three years. His mother's name was Maacah, a daughter of Uriel of Gibeah. There was war between Abijah and Jeroboam.
2CHR|13|3|Abijah went into battle with a force of four hundred thousand able fighting men, and Jeroboam drew up a battle line against him with eight hundred thousand able troops.
2CHR|13|4|Abijah stood on Mount Zemaraim, in the hill country of Ephraim, and said, "Jeroboam and all Israel, listen to me!
2CHR|13|5|Don't you know that the LORD, the God of Israel, has given the kingship of Israel to David and his descendants forever by a covenant of salt?
2CHR|13|6|Yet Jeroboam son of Nebat, an official of Solomon son of David, rebelled against his master.
2CHR|13|7|Some worthless scoundrels gathered around him and opposed Rehoboam son of Solomon when he was young and indecisive and not strong enough to resist them.
2CHR|13|8|"And now you plan to resist the kingdom of the LORD, which is in the hands of David's descendants. You are indeed a vast army and have with you the golden calves that Jeroboam made to be your gods.
2CHR|13|9|But didn't you drive out the priests of the LORD, the sons of Aaron, and the Levites, and make priests of your own as the peoples of other lands do? Whoever comes to consecrate himself with a young bull and seven rams may become a priest of what are not gods.
2CHR|13|10|"As for us, the LORD is our God, and we have not forsaken him. The priests who serve the LORD are sons of Aaron, and the Levites assist them.
2CHR|13|11|Every morning and evening they present burnt offerings and fragrant incense to the LORD. They set out the bread on the ceremonially clean table and light the lamps on the gold lampstand every evening. We are observing the requirements of the LORD our God. But you have forsaken him.
2CHR|13|12|God is with us; he is our leader. His priests with their trumpets will sound the battle cry against you. Men of Israel, do not fight against the LORD, the God of your fathers, for you will not succeed."
2CHR|13|13|Now Jeroboam had sent troops around to the rear, so that while he was in front of Judah the ambush was behind them.
2CHR|13|14|Judah turned and saw that they were being attacked at both front and rear. Then they cried out to the LORD. The priests blew their trumpets
2CHR|13|15|and the men of Judah raised the battle cry. At the sound of their battle cry, God routed Jeroboam and all Israel before Abijah and Judah.
2CHR|13|16|The Israelites fled before Judah, and God delivered them into their hands.
2CHR|13|17|Abijah and his men inflicted heavy losses on them, so that there were five hundred thousand casualties among Israel's able men.
2CHR|13|18|The men of Israel were subdued on that occasion, and the men of Judah were victorious because they relied on the LORD, the God of their fathers.
2CHR|13|19|Abijah pursued Jeroboam and took from him the towns of Bethel, Jeshanah and Ephron, with their surrounding villages.
2CHR|13|20|Jeroboam did not regain power during the time of Abijah. And the LORD struck him down and he died.
2CHR|13|21|But Abijah grew in strength. He married fourteen wives and had twenty-two sons and sixteen daughters.
2CHR|13|22|The other events of Abijah's reign, what he did and what he said, are written in the annotations of the prophet Iddo.
2CHR|14|1|And Abijah rested with his fathers and was buried in the City of David. Asa his son succeeded him as king, and in his days the country was at peace for ten years.
2CHR|14|2|Asa did what was good and right in the eyes of the LORD his God.
2CHR|14|3|He removed the foreign altars and the high places, smashed the sacred stones and cut down the Asherah poles.
2CHR|14|4|He commanded Judah to seek the LORD, the God of their fathers, and to obey his laws and commands.
2CHR|14|5|He removed the high places and incense altars in every town in Judah, and the kingdom was at peace under him.
2CHR|14|6|He built up the fortified cities of Judah, since the land was at peace. No one was at war with him during those years, for the LORD gave him rest.
2CHR|14|7|"Let us build up these towns," he said to Judah, "and put walls around them, with towers, gates and bars. The land is still ours, because we have sought the LORD our God; we sought him and he has given us rest on every side." So they built and prospered.
2CHR|14|8|Asa had an army of three hundred thousand men from Judah, equipped with large shields and with spears, and two hundred and eighty thousand from Benjamin, armed with small shields and with bows. All these were brave fighting men.
2CHR|14|9|Zerah the Cushite marched out against them with a vast army and three hundred chariots, and came as far as Mareshah.
2CHR|14|10|Asa went out to meet him, and they took up battle positions in the Valley of Zephathah near Mareshah.
2CHR|14|11|Then Asa called to the LORD his God and said, "LORD, there is no one like you to help the powerless against the mighty. Help us, O LORD our God, for we rely on you, and in your name we have come against this vast army. O LORD, you are our God; do not let man prevail against you."
2CHR|14|12|The LORD struck down the Cushites before Asa and Judah. The Cushites fled,
2CHR|14|13|and Asa and his army pursued them as far as Gerar. Such a great number of Cushites fell that they could not recover; they were crushed before the LORD and his forces. The men of Judah carried off a large amount of plunder.
2CHR|14|14|They destroyed all the villages around Gerar, for the terror of the LORD had fallen upon them. They plundered all these villages, since there was much booty there.
2CHR|14|15|They also attacked the camps of the herdsmen and carried off droves of sheep and goats and camels. Then they returned to Jerusalem.
2CHR|15|1|The Spirit of God came upon Azariah son of Oded.
2CHR|15|2|He went out to meet Asa and said to him, "Listen to me, Asa and all Judah and Benjamin. The LORD is with you when you are with him. If you seek him, he will be found by you, but if you forsake him, he will forsake you.
2CHR|15|3|For a long time Israel was without the true God, without a priest to teach and without the law.
2CHR|15|4|But in their distress they turned to the LORD, the God of Israel, and sought him, and he was found by them.
2CHR|15|5|In those days it was not safe to travel about, for all the inhabitants of the lands were in great turmoil.
2CHR|15|6|One nation was being crushed by another and one city by another, because God was troubling them with every kind of distress.
2CHR|15|7|But as for you, be strong and do not give up, for your work will be rewarded."
2CHR|15|8|When Asa heard these words and the prophecy of Azariah son of Oded the prophet, he took courage. He removed the detestable idols from the whole land of Judah and Benjamin and from the towns he had captured in the hills of Ephraim. He repaired the altar of the LORD that was in front of the portico of the LORD's temple.
2CHR|15|9|Then he assembled all Judah and Benjamin and the people from Ephraim, Manasseh and Simeon who had settled among them, for large numbers had come over to him from Israel when they saw that the LORD his God was with him.
2CHR|15|10|They assembled at Jerusalem in the third month of the fifteenth year of Asa's reign.
2CHR|15|11|At that time they sacrificed to the LORD seven hundred head of cattle and seven thousand sheep and goats from the plunder they had brought back.
2CHR|15|12|They entered into a covenant to seek the LORD, the God of their fathers, with all their heart and soul.
2CHR|15|13|All who would not seek the LORD, the God of Israel, were to be put to death, whether small or great, man or woman.
2CHR|15|14|They took an oath to the LORD with loud acclamation, with shouting and with trumpets and horns.
2CHR|15|15|All Judah rejoiced about the oath because they had sworn it wholeheartedly. They sought God eagerly, and he was found by them. So the LORD gave them rest on every side.
2CHR|15|16|King Asa also deposed his grandmother Maacah from her position as queen mother, because she had made a repulsive Asherah pole. Asa cut the pole down, broke it up and burned it in the Kidron Valley.
2CHR|15|17|Although he did not remove the high places from Israel, Asa's heart was fully committed to the LORD all his life.
2CHR|15|18|He brought into the temple of God the silver and gold and the articles that he and his father had dedicated.
2CHR|15|19|There was no more war until the thirty-fifth year of Asa's reign.
2CHR|16|1|In the thirty-sixth year of Asa's reign Baasha king of Israel went up against Judah and fortified Ramah to prevent anyone from leaving or entering the territory of Asa king of Judah.
2CHR|16|2|Asa then took the silver and gold out of the treasuries of the LORD's temple and of his own palace and sent it to Ben-Hadad king of Aram, who was ruling in Damascus.
2CHR|16|3|"Let there be a treaty between me and you," he said, "as there was between my father and your father. See, I am sending you silver and gold. Now break your treaty with Baasha king of Israel so he will withdraw from me."
2CHR|16|4|Ben-Hadad agreed with King Asa and sent the commanders of his forces against the towns of Israel. They conquered Ijon, Dan, Abel Maim and all the store cities of Naphtali.
2CHR|16|5|When Baasha heard this, he stopped building Ramah and abandoned his work.
2CHR|16|6|Then King Asa brought all the men of Judah, and they carried away from Ramah the stones and timber Baasha had been using. With them he built up Geba and Mizpah.
2CHR|16|7|At that time Hanani the seer came to Asa king of Judah and said to him: "Because you relied on the king of Aram and not on the LORD your God, the army of the king of Aram has escaped from your hand.
2CHR|16|8|Were not the Cushites and Libyans a mighty army with great numbers of chariots and horsemen? Yet when you relied on the LORD, he delivered them into your hand.
2CHR|16|9|For the eyes of the LORD range throughout the earth to strengthen those whose hearts are fully committed to him. You have done a foolish thing, and from now on you will be at war."
2CHR|16|10|Asa was angry with the seer because of this; he was so enraged that he put him in prison. At the same time Asa brutally oppressed some of the people.
2CHR|16|11|The events of Asa's reign, from beginning to end, are written in the book of the kings of Judah and Israel.
2CHR|16|12|In the thirty-ninth year of his reign Asa was afflicted with a disease in his feet. Though his disease was severe, even in his illness he did not seek help from the LORD, but only from the physicians.
2CHR|16|13|Then in the forty-first year of his reign Asa died and rested with his fathers.
2CHR|16|14|They buried him in the tomb that he had cut out for himself in the City of David. They laid him on a bier covered with spices and various blended perfumes, and they made a huge fire in his honor.
2CHR|17|1|Jehoshaphat his son succeeded him as king and strengthened himself against Israel.
2CHR|17|2|He stationed troops in all the fortified cities of Judah and put garrisons in Judah and in the towns of Ephraim that his father Asa had captured.
2CHR|17|3|The LORD was with Jehoshaphat because in his early years he walked in the ways his father David had followed. He did not consult the Baals
2CHR|17|4|but sought the God of his father and followed his commands rather than the practices of Israel.
2CHR|17|5|The LORD established the kingdom under his control; and all Judah brought gifts to Jehoshaphat, so that he had great wealth and honor.
2CHR|17|6|His heart was devoted to the ways of the LORD; furthermore, he removed the high places and the Asherah poles from Judah.
2CHR|17|7|In the third year of his reign he sent his officials Ben-Hail, Obadiah, Zechariah, Nethanel and Micaiah to teach in the towns of Judah.
2CHR|17|8|With them were certain Levites-Shemaiah, Nethaniah, Zebadiah, Asahel, Shemiramoth, Jehonathan, Adonijah, Tobijah and Tob-Adonijah-and the priests Elishama and Jehoram.
2CHR|17|9|They taught throughout Judah, taking with them the Book of the Law of the LORD; they went around to all the towns of Judah and taught the people.
2CHR|17|10|The fear of the LORD fell on all the kingdoms of the lands surrounding Judah, so that they did not make war with Jehoshaphat.
2CHR|17|11|Some Philistines brought Jehoshaphat gifts and silver as tribute, and the Arabs brought him flocks: seven thousand seven hundred rams and seven thousand seven hundred goats.
2CHR|17|12|Jehoshaphat became more and more powerful; he built forts and store cities in Judah
2CHR|17|13|and had large supplies in the towns of Judah. He also kept experienced fighting men in Jerusalem.
2CHR|17|14|Their enrollment by families was as follows: From Judah, commanders of units of 1,000: Adnah the commander, with 300,000 fighting men;
2CHR|17|15|next, Jehohanan the commander, with 280,000;
2CHR|17|16|next, Amasiah son of Zicri, who volunteered himself for the service of the LORD, with 200,000.
2CHR|17|17|From Benjamin: Eliada, a valiant soldier, with 200,000 men armed with bows and shields;
2CHR|17|18|next, Jehozabad, with 180,000 men armed for battle.
2CHR|17|19|These were the men who served the king, besides those he stationed in the fortified cities throughout Judah.
2CHR|18|1|Now Jehoshaphat had great wealth and honor, and he allied himself with Ahab by marriage.
2CHR|18|2|Some years later he went down to visit Ahab in Samaria. Ahab slaughtered many sheep and cattle for him and the people with him and urged him to attack Ramoth Gilead.
2CHR|18|3|Ahab king of Israel asked Jehoshaphat king of Judah, "Will you go with me against Ramoth Gilead?" Jehoshaphat replied, "I am as you are, and my people as your people; we will join you in the war."
2CHR|18|4|But Jehoshaphat also said to the king of Israel, "First seek the counsel of the LORD."
2CHR|18|5|So the king of Israel brought together the prophets-four hundred men-and asked them, "Shall we go to war against Ramoth Gilead, or shall I refrain?Go," they answered, "for God will give it into the king's hand."
2CHR|18|6|But Jehoshaphat asked, "Is there not a prophet of the LORD here whom we can inquire of?"
2CHR|18|7|The king of Israel answered Jehoshaphat, "There is still one man through whom we can inquire of the LORD, but I hate him because he never prophesies anything good about me, but always bad. He is Micaiah son of Imlah.The king should not say that," Jehoshaphat replied.
2CHR|18|8|So the king of Israel called one of his officials and said, "Bring Micaiah son of Imlah at once."
2CHR|18|9|Dressed in their royal robes, the king of Israel and Jehoshaphat king of Judah were sitting on their thrones at the threshing floor by the entrance to the gate of Samaria, with all the prophets prophesying before them.
2CHR|18|10|Now Zedekiah son of Kenaanah had made iron horns, and he declared, "This is what the LORD says: 'With these you will gore the Arameans until they are destroyed.'"
2CHR|18|11|All the other prophets were prophesying the same thing. "Attack Ramoth Gilead and be victorious," they said, "for the LORD will give it into the king's hand."
2CHR|18|12|The messenger who had gone to summon Micaiah said to him, "Look, as one man the other prophets are predicting success for the king. Let your word agree with theirs, and speak favorably."
2CHR|18|13|But Micaiah said, "As surely as the LORD lives, I can tell him only what my God says."
2CHR|18|14|When he arrived, the king asked him, "Micaiah, shall we go to war against Ramoth Gilead, or shall I refrain?Attack and be victorious," he answered, "for they will be given into your hand."
2CHR|18|15|The king said to him, "How many times must I make you swear to tell me nothing but the truth in the name of the LORD?"
2CHR|18|16|Then Micaiah answered, "I saw all Israel scattered on the hills like sheep without a shepherd, and the LORD said, 'These people have no master. Let each one go home in peace.'"
2CHR|18|17|The king of Israel said to Jehoshaphat, "Didn't I tell you that he never prophesies anything good about me, but only bad?"
2CHR|18|18|Micaiah continued, "Therefore hear the word of the LORD: I saw the LORD sitting on his throne with all the host of heaven standing on his right and on his left.
2CHR|18|19|And the LORD said, 'Who will entice Ahab king of Israel into attacking Ramoth Gilead and going to his death there?'"One suggested this, and another that.
2CHR|18|20|Finally, a spirit came forward, stood before the LORD and said, 'I will entice him.'"'By what means?' the LORD asked.
2CHR|18|21|"'I will go and be a lying spirit in the mouths of all his prophets,' he said. "'You will succeed in enticing him,' said the LORD. 'Go and do it.'
2CHR|18|22|"So now the LORD has put a lying spirit in the mouths of these prophets of yours. The LORD has decreed disaster for you."
2CHR|18|23|Then Zedekiah son of Kenaanah went up and slapped Micaiah in the face. "Which way did the spirit from the LORD go when he went from me to speak to you?" he asked.
2CHR|18|24|Micaiah replied, "You will find out on the day you go to hide in an inner room."
2CHR|18|25|The king of Israel then ordered, "Take Micaiah and send him back to Amon the ruler of the city and to Joash the king's son,
2CHR|18|26|and say, 'This is what the king says: Put this fellow in prison and give him nothing but bread and water until I return safely.'"
2CHR|18|27|Micaiah declared, "If you ever return safely, the LORD has not spoken through me." Then he added, "Mark my words, all you people!"
2CHR|18|28|So the king of Israel and Jehoshaphat king of Judah went up to Ramoth Gilead.
2CHR|18|29|The king of Israel said to Jehoshaphat, "I will enter the battle in disguise, but you wear your royal robes." So the king of Israel disguised himself and went into battle.
2CHR|18|30|Now the king of Aram had ordered his chariot commanders, "Do not fight with anyone, small or great, except the king of Israel."
2CHR|18|31|When the chariot commanders saw Jehoshaphat, they thought, "This is the king of Israel." So they turned to attack him, but Jehoshaphat cried out, and the LORD helped him. God drew them away from him,
2CHR|18|32|for when the chariot commanders saw that he was not the king of Israel, they stopped pursuing him.
2CHR|18|33|But someone drew his bow at random and hit the king of Israel between the sections of his armor. The king told the chariot driver, "Wheel around and get me out of the fighting. I've been wounded."
2CHR|18|34|All day long the battle raged, and the king of Israel propped himself up in his chariot facing the Arameans until evening. Then at sunset he died.
2CHR|19|1|When Jehoshaphat king of Judah returned safely to his palace in Jerusalem,
2CHR|19|2|Jehu the seer, the son of Hanani, went out to meet him and said to the king, "Should you help the wicked and love those who hate the LORD? Because of this, the wrath of the LORD is upon you.
2CHR|19|3|There is, however, some good in you, for you have rid the land of the Asherah poles and have set your heart on seeking God."
2CHR|19|4|Jehoshaphat lived in Jerusalem, and he went out again among the people from Beersheba to the hill country of Ephraim and turned them back to the LORD, the God of their fathers.
2CHR|19|5|He appointed judges in the land, in each of the fortified cities of Judah.
2CHR|19|6|He told them, "Consider carefully what you do, because you are not judging for man but for the LORD, who is with you whenever you give a verdict.
2CHR|19|7|Now let the fear of the LORD be upon you. Judge carefully, for with the LORD our God there is no injustice or partiality or bribery."
2CHR|19|8|In Jerusalem also, Jehoshaphat appointed some of the Levites, priests and heads of Israelite families to administer the law of the LORD and to settle disputes. And they lived in Jerusalem.
2CHR|19|9|He gave them these orders: "You must serve faithfully and wholeheartedly in the fear of the LORD.
2CHR|19|10|In every case that comes before you from your fellow countrymen who live in the cities-whether bloodshed or other concerns of the law, commands, decrees or ordinances-you are to warn them not to sin against the LORD; otherwise his wrath will come on you and your brothers. Do this, and you will not sin.
2CHR|19|11|"Amariah the chief priest will be over you in any matter concerning the LORD, and Zebadiah son of Ishmael, the leader of the tribe of Judah, will be over you in any matter concerning the king, and the Levites will serve as officials before you. Act with courage, and may the LORD be with those who do well."
2CHR|20|1|After this, the Moabites and Ammonites with some of the Meunites came to make war on Jehoshaphat.
2CHR|20|2|Some men came and told Jehoshaphat, "A vast army is coming against you from Edom, from the other side of the Sea. It is already in Hazazon Tamar" (that is, En Gedi).
2CHR|20|3|Alarmed, Jehoshaphat resolved to inquire of the LORD, and he proclaimed a fast for all Judah.
2CHR|20|4|The people of Judah came together to seek help from the LORD; indeed, they came from every town in Judah to seek him.
2CHR|20|5|Then Jehoshaphat stood up in the assembly of Judah and Jerusalem at the temple of the LORD in the front of the new courtyard
2CHR|20|6|and said: "O LORD, God of our fathers, are you not the God who is in heaven? You rule over all the kingdoms of the nations. Power and might are in your hand, and no one can withstand you.
2CHR|20|7|O our God, did you not drive out the inhabitants of this land before your people Israel and give it forever to the descendants of Abraham your friend?
2CHR|20|8|They have lived in it and have built in it a sanctuary for your Name, saying,
2CHR|20|9|'If calamity comes upon us, whether the sword of judgment, or plague or famine, we will stand in your presence before this temple that bears your Name and will cry out to you in our distress, and you will hear us and save us.'
2CHR|20|10|"But now here are men from Ammon, Moab and Mount Seir, whose territory you would not allow Israel to invade when they came from Egypt; so they turned away from them and did not destroy them.
2CHR|20|11|See how they are repaying us by coming to drive us out of the possession you gave us as an inheritance.
2CHR|20|12|O our God, will you not judge them? For we have no power to face this vast army that is attacking us. We do not know what to do, but our eyes are upon you."
2CHR|20|13|All the men of Judah, with their wives and children and little ones, stood there before the LORD.
2CHR|20|14|Then the Spirit of the LORD came upon Jahaziel son of Zechariah, the son of Benaiah, the son of Jeiel, the son of Mattaniah, a Levite and descendant of Asaph, as he stood in the assembly.
2CHR|20|15|He said: "Listen, King Jehoshaphat and all who live in Judah and Jerusalem! This is what the LORD says to you: 'Do not be afraid or discouraged because of this vast army. For the battle is not yours, but God's.
2CHR|20|16|Tomorrow march down against them. They will be climbing up by the Pass of Ziz, and you will find them at the end of the gorge in the Desert of Jeruel.
2CHR|20|17|You will not have to fight this battle. Take up your positions; stand firm and see the deliverance the LORD will give you, O Judah and Jerusalem. Do not be afraid; do not be discouraged. Go out to face them tomorrow, and the LORD will be with you.'"
2CHR|20|18|Jehoshaphat bowed with his face to the ground, and all the people of Judah and Jerusalem fell down in worship before the LORD.
2CHR|20|19|Then some Levites from the Kohathites and Korahites stood up and praised the LORD, the God of Israel, with very loud voice.
2CHR|20|20|Early in the morning they left for the Desert of Tekoa. As they set out, Jehoshaphat stood and said, "Listen to me, Judah and people of Jerusalem! Have faith in the LORD your God and you will be upheld; have faith in his prophets and you will be successful."
2CHR|20|21|After consulting the people, Jehoshaphat appointed men to sing to the LORD and to praise him for the splendor of his holiness as they went out at the head of the army, saying: "Give thanks to the LORD, for his love endures forever."
2CHR|20|22|As they began to sing and praise, the LORD set ambushes against the men of Ammon and Moab and Mount Seir who were invading Judah, and they were defeated.
2CHR|20|23|The men of Ammon and Moab rose up against the men from Mount Seir to destroy and annihilate them. After they finished slaughtering the men from Seir, they helped to destroy one another.
2CHR|20|24|When the men of Judah came to the place that overlooks the desert and looked toward the vast army, they saw only dead bodies lying on the ground; no one had escaped.
2CHR|20|25|So Jehoshaphat and his men went to carry off their plunder, and they found among them a great amount of equipment and clothing and also articles of value-more than they could take away. There was so much plunder that it took three days to collect it.
2CHR|20|26|On the fourth day they assembled in the Valley of Beracah, where they praised the LORD. This is why it is called the Valley of Beracah to this day.
2CHR|20|27|Then, led by Jehoshaphat, all the men of Judah and Jerusalem returned joyfully to Jerusalem, for the LORD had given them cause to rejoice over their enemies.
2CHR|20|28|They entered Jerusalem and went to the temple of the LORD with harps and lutes and trumpets.
2CHR|20|29|The fear of God came upon all the kingdoms of the countries when they heard how the LORD had fought against the enemies of Israel.
2CHR|20|30|And the kingdom of Jehoshaphat was at peace, for his God had given him rest on every side.
2CHR|20|31|So Jehoshaphat reigned over Judah. He was thirty-five years old when he became king of Judah, and he reigned in Jerusalem twenty-five years. His mother's name was Azubah daughter of Shilhi.
2CHR|20|32|He walked in the ways of his father Asa and did not stray from them; he did what was right in the eyes of the LORD.
2CHR|20|33|The high places, however, were not removed, and the people still had not set their hearts on the God of their fathers.
2CHR|20|34|The other events of Jehoshaphat's reign, from beginning to end, are written in the annals of Jehu son of Hanani, which are recorded in the book of the kings of Israel.
2CHR|20|35|Later, Jehoshaphat king of Judah made an alliance with Ahaziah king of Israel, who was guilty of wickedness.
2CHR|20|36|He agreed with him to construct a fleet of trading ships. After these were built at Ezion Geber,
2CHR|20|37|Eliezer son of Dodavahu of Mareshah prophesied against Jehoshaphat, saying, "Because you have made an alliance with Ahaziah, the LORD will destroy what you have made." The ships were wrecked and were not able to set sail to trade.
2CHR|21|1|Then Jehoshaphat rested with his fathers and was buried with them in the City of David. And Jehoram his son succeeded him as king.
2CHR|21|2|Jehoram's brothers, the sons of Jehoshaphat, were Azariah, Jehiel, Zechariah, Azariahu, Michael and Shephatiah. All these were sons of Jehoshaphat king of Israel.
2CHR|21|3|Their father had given them many gifts of silver and gold and articles of value, as well as fortified cities in Judah, but he had given the kingdom to Jehoram because he was his firstborn son.
2CHR|21|4|When Jehoram established himself firmly over his father's kingdom, he put all his brothers to the sword along with some of the princes of Israel.
2CHR|21|5|Jehoram was thirty-two years old when he became king, and he reigned in Jerusalem eight years.
2CHR|21|6|He walked in the ways of the kings of Israel, as the house of Ahab had done, for he married a daughter of Ahab. He did evil in the eyes of the LORD.
2CHR|21|7|Nevertheless, because of the covenant the LORD had made with David, the LORD was not willing to destroy the house of David. He had promised to maintain a lamp for him and his descendants forever.
2CHR|21|8|In the time of Jehoram, Edom rebelled against Judah and set up its own king.
2CHR|21|9|So Jehoram went there with his officers and all his chariots. The Edomites surrounded him and his chariot commanders, but he rose up and broke through by night.
2CHR|21|10|To this day Edom has been in rebellion against Judah. Libnah revolted at the same time, because Jehoram had forsaken the LORD, the God of his fathers.
2CHR|21|11|He had also built high places on the hills of Judah and had caused the people of Jerusalem to prostitute themselves and had led Judah astray.
2CHR|21|12|Jehoram received a letter from Elijah the prophet, which said: "This is what the LORD, the God of your father David, says: 'You have not walked in the ways of your father Jehoshaphat or of Asa king of Judah.
2CHR|21|13|But you have walked in the ways of the kings of Israel, and you have led Judah and the people of Jerusalem to prostitute themselves, just as the house of Ahab did. You have also murdered your own brothers, members of your father's house, men who were better than you.
2CHR|21|14|So now the LORD is about to strike your people, your sons, your wives and everything that is yours, with a heavy blow.
2CHR|21|15|You yourself will be very ill with a lingering disease of the bowels, until the disease causes your bowels to come out.'"
2CHR|21|16|The LORD aroused against Jehoram the hostility of the Philistines and of the Arabs who lived near the Cushites.
2CHR|21|17|They attacked Judah, invaded it and carried off all the goods found in the king's palace, together with his sons and wives. Not a son was left to him except Ahaziah, the youngest.
2CHR|21|18|After all this, the LORD afflicted Jehoram with an incurable disease of the bowels.
2CHR|21|19|In the course of time, at the end of the second year, his bowels came out because of the disease, and he died in great pain. His people made no fire in his honor, as they had for his fathers.
2CHR|21|20|Jehoram was thirty-two years old when he became king, and he reigned in Jerusalem eight years. He passed away, to no one's regret, and was buried in the City of David, but not in the tombs of the kings.
2CHR|22|1|The people of Jerusalem made Ahaziah, Jehoram's youngest son, king in his place, since the raiders, who came with the Arabs into the camp, had killed all the older sons. So Ahaziah son of Jehoram king of Judah began to reign.
2CHR|22|2|Ahaziah was twenty-two years old when he became king, and he reigned in Jerusalem one year. His mother's name was Athaliah, a granddaughter of Omri.
2CHR|22|3|He too walked in the ways of the house of Ahab, for his mother encouraged him in doing wrong.
2CHR|22|4|He did evil in the eyes of the LORD, as the house of Ahab had done, for after his father's death they became his advisers, to his undoing.
2CHR|22|5|He also followed their counsel when he went with Joram son of Ahab king of Israel to war against Hazael king of Aram at Ramoth Gilead. The Arameans wounded Joram;
2CHR|22|6|so he returned to Jezreel to recover from the wounds they had inflicted on him at Ramoth in his battle with Hazael king of Aram. Then Ahaziah son of Jehoram king of Judah went down to Jezreel to see Joram son of Ahab because he had been wounded.
2CHR|22|7|Through Ahaziah's visit to Joram, God brought about Ahaziah's downfall. When Ahaziah arrived, he went out with Joram to meet Jehu son of Nimshi, whom the LORD had anointed to destroy the house of Ahab.
2CHR|22|8|While Jehu was executing judgment on the house of Ahab, he found the princes of Judah and the sons of Ahaziah's relatives, who had been attending Ahaziah, and he killed them.
2CHR|22|9|He then went in search of Ahaziah, and his men captured him while he was hiding in Samaria. He was brought to Jehu and put to death. They buried him, for they said, "He was a son of Jehoshaphat, who sought the LORD with all his heart." So there was no one in the house of Ahaziah powerful enough to retain the kingdom.
2CHR|22|10|When Athaliah the mother of Ahaziah saw that her son was dead, she proceeded to destroy the whole royal family of the house of Judah.
2CHR|22|11|But Jehosheba, the daughter of King Jehoram, took Joash son of Ahaziah and stole him away from among the royal princes who were about to be murdered and put him and his nurse in a bedroom. Because Jehosheba, the daughter of King Jehoram and wife of the priest Jehoiada, was Ahaziah's sister, she hid the child from Athaliah so she could not kill him.
2CHR|22|12|He remained hidden with them at the temple of God for six years while Athaliah ruled the land.
2CHR|23|1|In the seventh year Jehoiada showed his strength. He made a covenant with the commanders of units of a hundred: Azariah son of Jeroham, Ishmael son of Jehohanan, Azariah son of Obed, Maaseiah son of Adaiah, and Elishaphat son of Zicri.
2CHR|23|2|They went throughout Judah and gathered the Levites and the heads of Israelite families from all the towns. When they came to Jerusalem,
2CHR|23|3|the whole assembly made a covenant with the king at the temple of God. Jehoiada said to them, "The king's son shall reign, as the LORD promised concerning the descendants of David.
2CHR|23|4|Now this is what you are to do: A third of you priests and Levites who are going on duty on the Sabbath are to keep watch at the doors,
2CHR|23|5|a third of you at the royal palace and a third at the Foundation Gate, and all the other men are to be in the courtyards of the temple of the LORD.
2CHR|23|6|No one is to enter the temple of the LORD except the priests and Levites on duty; they may enter because they are consecrated, but all the other men are to guard what the LORD has assigned to them.
2CHR|23|7|The Levites are to station themselves around the king, each man with his weapons in his hand. Anyone who enters the temple must be put to death. Stay close to the king wherever he goes."
2CHR|23|8|The Levites and all the men of Judah did just as Jehoiada the priest ordered. Each one took his men-those who were going on duty on the Sabbath and those who were going off duty-for Jehoiada the priest had not released any of the divisions.
2CHR|23|9|Then he gave the commanders of units of a hundred the spears and the large and small shields that had belonged to King David and that were in the temple of God.
2CHR|23|10|He stationed all the men, each with his weapon in his hand, around the king-near the altar and the temple, from the south side to the north side of the temple.
2CHR|23|11|Jehoiada and his sons brought out the king's son and put the crown on him; they presented him with a copy of the covenant and proclaimed him king. They anointed him and shouted, "Long live the king!"
2CHR|23|12|When Athaliah heard the noise of the people running and cheering the king, she went to them at the temple of the LORD.
2CHR|23|13|She looked, and there was the king, standing by his pillar at the entrance. The officers and the trumpeters were beside the king, and all the people of the land were rejoicing and blowing trumpets, and singers with musical instruments were leading the praises. Then Athaliah tore her robes and shouted, "Treason! Treason!"
2CHR|23|14|Jehoiada the priest sent out the commanders of units of a hundred, who were in charge of the troops, and said to them: "Bring her out between the ranks and put to the sword anyone who follows her." For the priest had said, "Do not put her to death at the temple of the LORD."
2CHR|23|15|So they seized her as she reached the entrance of the Horse Gate on the palace grounds, and there they put her to death.
2CHR|23|16|Jehoiada then made a covenant that he and the people and the king would be the LORD's people.
2CHR|23|17|All the people went to the temple of Baal and tore it down. They smashed the altars and idols and killed Mattan the priest of Baal in front of the altars.
2CHR|23|18|Then Jehoiada placed the oversight of the temple of the LORD in the hands of the priests, who were Levites, to whom David had made assignments in the temple, to present the burnt offerings of the LORD as written in the Law of Moses, with rejoicing and singing, as David had ordered.
2CHR|23|19|He also stationed doorkeepers at the gates of the LORD's temple so that no one who was in any way unclean might enter.
2CHR|23|20|He took with him the commanders of hundreds, the nobles, the rulers of the people and all the people of the land and brought the king down from the temple of the LORD. They went into the palace through the Upper Gate and seated the king on the royal throne,
2CHR|23|21|and all the people of the land rejoiced. And the city was quiet, because Athaliah had been slain with the sword.
2CHR|24|1|Joash was seven years old when he became king, and he reigned in Jerusalem forty years. His mother's name was Zibiah; she was from Beersheba.
2CHR|24|2|Joash did what was right in the eyes of the LORD all the years of Jehoiada the priest.
2CHR|24|3|Jehoiada chose two wives for him, and he had sons and daughters.
2CHR|24|4|Some time later Joash decided to restore the temple of the LORD.
2CHR|24|5|He called together the priests and Levites and said to them, "Go to the towns of Judah and collect the money due annually from all Israel, to repair the temple of your God. Do it now." But the Levites did not act at once.
2CHR|24|6|Therefore the king summoned Jehoiada the chief priest and said to him, "Why haven't you required the Levites to bring in from Judah and Jerusalem the tax imposed by Moses the servant of the LORD and by the assembly of Israel for the Tent of the Testimony?"
2CHR|24|7|Now the sons of that wicked woman Athaliah had broken into the temple of God and had used even its sacred objects for the Baals.
2CHR|24|8|At the king's command, a chest was made and placed outside, at the gate of the temple of the LORD.
2CHR|24|9|A proclamation was then issued in Judah and Jerusalem that they should bring to the LORD the tax that Moses the servant of God had required of Israel in the desert.
2CHR|24|10|All the officials and all the people brought their contributions gladly, dropping them into the chest until it was full.
2CHR|24|11|Whenever the chest was brought in by the Levites to the king's officials and they saw that there was a large amount of money, the royal secretary and the officer of the chief priest would come and empty the chest and carry it back to its place. They did this regularly and collected a great amount of money.
2CHR|24|12|The king and Jehoiada gave it to the men who carried out the work required for the temple of the LORD. They hired masons and carpenters to restore the LORD's temple, and also workers in iron and bronze to repair the temple.
2CHR|24|13|The men in charge of the work were diligent, and the repairs progressed under them. They rebuilt the temple of God according to its original design and reinforced it.
2CHR|24|14|When they had finished, they brought the rest of the money to the king and Jehoiada, and with it were made articles for the LORD's temple: articles for the service and for the burnt offerings, and also dishes and other objects of gold and silver. As long as Jehoiada lived, burnt offerings were presented continually in the temple of the LORD.
2CHR|24|15|Now Jehoiada was old and full of years, and he died at the age of a hundred and thirty.
2CHR|24|16|He was buried with the kings in the City of David, because of the good he had done in Israel for God and his temple.
2CHR|24|17|After the death of Jehoiada, the officials of Judah came and paid homage to the king, and he listened to them.
2CHR|24|18|They abandoned the temple of the LORD, the God of their fathers, and worshiped Asherah poles and idols. Because of their guilt, God's anger came upon Judah and Jerusalem.
2CHR|24|19|Although the LORD sent prophets to the people to bring them back to him, and though they testified against them, they would not listen.
2CHR|24|20|Then the Spirit of God came upon Zechariah son of Jehoiada the priest. He stood before the people and said, "This is what God says: 'Why do you disobey the LORD's commands? You will not prosper. Because you have forsaken the LORD, he has forsaken you.'"
2CHR|24|21|But they plotted against him, and by order of the king they stoned him to death in the courtyard of the LORD's temple.
2CHR|24|22|King Joash did not remember the kindness Zechariah's father Jehoiada had shown him but killed his son, who said as he lay dying, "May the LORD see this and call you to account."
2CHR|24|23|At the turn of the year, the army of Aram marched against Joash; it invaded Judah and Jerusalem and killed all the leaders of the people. They sent all the plunder to their king in Damascus.
2CHR|24|24|Although the Aramean army had come with only a few men, the LORD delivered into their hands a much larger army. Because Judah had forsaken the LORD, the God of their fathers, judgment was executed on Joash.
2CHR|24|25|When the Arameans withdrew, they left Joash severely wounded. His officials conspired against him for murdering the son of Jehoiada the priest, and they killed him in his bed. So he died and was buried in the City of David, but not in the tombs of the kings.
2CHR|24|26|Those who conspired against him were Zabad, son of Shimeath an Ammonite woman, and Jehozabad, son of Shimrith a Moabite woman.
2CHR|24|27|The account of his sons, the many prophecies about him, and the record of the restoration of the temple of God are written in the annotations on the book of the kings. And Amaziah his son succeeded him as king.
2CHR|25|1|Amaziah was twenty-five years old when he became king, and he reigned in Jerusalem twenty-nine years. His mother's name was Jehoaddin; she was from Jerusalem.
2CHR|25|2|He did what was right in the eyes of the LORD, but not wholeheartedly.
2CHR|25|3|After the kingdom was firmly in his control, he executed the officials who had murdered his father the king.
2CHR|25|4|Yet he did not put their sons to death, but acted in accordance with what is written in the Law, in the Book of Moses, where the LORD commanded: "Fathers shall not be put to death for their children, nor children put to death for their fathers; each is to die for his own sins."
2CHR|25|5|Amaziah called the people of Judah together and assigned them according to their families to commanders of thousands and commanders of hundreds for all Judah and Benjamin. He then mustered those twenty years old or more and found that there were three hundred thousand men ready for military service, able to handle the spear and shield.
2CHR|25|6|He also hired a hundred thousand fighting men from Israel for a hundred talents of silver.
2CHR|25|7|But a man of God came to him and said, "O king, these troops from Israel must not march with you, for the LORD is not with Israel-not with any of the people of Ephraim.
2CHR|25|8|Even if you go and fight courageously in battle, God will overthrow you before the enemy, for God has the power to help or to overthrow."
2CHR|25|9|Amaziah asked the man of God, "But what about the hundred talents I paid for these Israelite troops?" The man of God replied, "The LORD can give you much more than that."
2CHR|25|10|So Amaziah dismissed the troops who had come to him from Ephraim and sent them home. They were furious with Judah and left for home in a great rage.
2CHR|25|11|Amaziah then marshaled his strength and led his army to the Valley of Salt, where he killed ten thousand men of Seir.
2CHR|25|12|The army of Judah also captured ten thousand men alive, took them to the top of a cliff and threw them down so that all were dashed to pieces.
2CHR|25|13|Meanwhile the troops that Amaziah had sent back and had not allowed to take part in the war raided Judean towns from Samaria to Beth Horon. They killed three thousand people and carried off great quantities of plunder.
2CHR|25|14|When Amaziah returned from slaughtering the Edomites, he brought back the gods of the people of Seir. He set them up as his own gods, bowed down to them and burned sacrifices to them.
2CHR|25|15|The anger of the LORD burned against Amaziah, and he sent a prophet to him, who said, "Why do you consult this people's gods, which could not save their own people from your hand?"
2CHR|25|16|While he was still speaking, the king said to him, "Have we appointed you an adviser to the king? Stop! Why be struck down?" So the prophet stopped but said, "I know that God has determined to destroy you, because you have done this and have not listened to my counsel."
2CHR|25|17|After Amaziah king of Judah consulted his advisers, he sent this challenge to Jehoash son of Jehoahaz, the son of Jehu, king of Israel: "Come, meet me face to face."
2CHR|25|18|But Jehoash king of Israel replied to Amaziah king of Judah: "A thistle in Lebanon sent a message to a cedar in Lebanon, 'Give your daughter to my son in marriage.' Then a wild beast in Lebanon came along and trampled the thistle underfoot.
2CHR|25|19|You say to yourself that you have defeated Edom, and now you are arrogant and proud. But stay at home! Why ask for trouble and cause your own downfall and that of Judah also?"
2CHR|25|20|Amaziah, however, would not listen, for God so worked that he might hand them over to Jehoash, because they sought the gods of Edom.
2CHR|25|21|So Jehoash king of Israel attacked. He and Amaziah king of Judah faced each other at Beth Shemesh in Judah.
2CHR|25|22|Judah was routed by Israel, and every man fled to his home.
2CHR|25|23|Jehoash king of Israel captured Amaziah king of Judah, the son of Joash, the son of Ahaziah, at Beth Shemesh. Then Jehoash brought him to Jerusalem and broke down the wall of Jerusalem from the Ephraim Gate to the Corner Gate-a section about six hundred feet long.
2CHR|25|24|He took all the gold and silver and all the articles found in the temple of God that had been in the care of Obed-Edom, together with the palace treasures and the hostages, and returned to Samaria.
2CHR|25|25|Amaziah son of Joash king of Judah lived for fifteen years after the death of Jehoash son of Jehoahaz king of Israel.
2CHR|25|26|As for the other events of Amaziah's reign, from beginning to end, are they not written in the book of the kings of Judah and Israel?
2CHR|25|27|From the time that Amaziah turned away from following the LORD, they conspired against him in Jerusalem and he fled to Lachish, but they sent men after him to Lachish and killed him there.
2CHR|25|28|He was brought back by horse and was buried with his fathers in the City of Judah.
2CHR|26|1|Then all the people of Judah took Uzziah, who was sixteen years old, and made him king in place of his father Amaziah.
2CHR|26|2|He was the one who rebuilt Elath and restored it to Judah after Amaziah rested with his fathers.
2CHR|26|3|Uzziah was sixteen years old when he became king, and he reigned in Jerusalem fifty-two years. His mother's name was Jecoliah; she was from Jerusalem.
2CHR|26|4|He did what was right in the eyes of the LORD, just as his father Amaziah had done.
2CHR|26|5|He sought God during the days of Zechariah, who instructed him in the fear of God. As long as he sought the LORD, God gave him success.
2CHR|26|6|He went to war against the Philistines and broke down the walls of Gath, Jabneh and Ashdod. He then rebuilt towns near Ashdod and elsewhere among the Philistines.
2CHR|26|7|God helped him against the Philistines and against the Arabs who lived in Gur Baal and against the Meunites.
2CHR|26|8|The Ammonites brought tribute to Uzziah, and his fame spread as far as the border of Egypt, because he had become very powerful.
2CHR|26|9|Uzziah built towers in Jerusalem at the Corner Gate, at the Valley Gate and at the angle of the wall, and he fortified them.
2CHR|26|10|He also built towers in the desert and dug many cisterns, because he had much livestock in the foothills and in the plain. He had people working his fields and vineyards in the hills and in the fertile lands, for he loved the soil.
2CHR|26|11|Uzziah had a well-trained army, ready to go out by divisions according to their numbers as mustered by Jeiel the secretary and Maaseiah the officer under the direction of Hananiah, one of the royal officials.
2CHR|26|12|The total number of family leaders over the fighting men was 2,600.
2CHR|26|13|Under their command was an army of 307,500 men trained for war, a powerful force to support the king against his enemies.
2CHR|26|14|Uzziah provided shields, spears, helmets, coats of armor, bows and slingstones for the entire army.
2CHR|26|15|In Jerusalem he made machines designed by skillful men for use on the towers and on the corner defenses to shoot arrows and hurl large stones. His fame spread far and wide, for he was greatly helped until he became powerful.
2CHR|26|16|But after Uzziah became powerful, his pride led to his downfall. He was unfaithful to the LORD his God, and entered the temple of the LORD to burn incense on the altar of incense.
2CHR|26|17|Azariah the priest with eighty other courageous priests of the LORD followed him in.
2CHR|26|18|They confronted him and said, "It is not right for you, Uzziah, to burn incense to the LORD. That is for the priests, the descendants of Aaron, who have been consecrated to burn incense. Leave the sanctuary, for you have been unfaithful; and you will not be honored by the LORD God."
2CHR|26|19|Uzziah, who had a censer in his hand ready to burn incense, became angry. While he was raging at the priests in their presence before the incense altar in the LORD's temple, leprosy broke out on his forehead.
2CHR|26|20|When Azariah the chief priest and all the other priests looked at him, they saw that he had leprosy on his forehead, so they hurried him out. Indeed, he himself was eager to leave, because the LORD had afflicted him.
2CHR|26|21|King Uzziah had leprosy until the day he died. He lived in a separate house -leprous, and excluded from the temple of the LORD. Jotham his son had charge of the palace and governed the people of the land.
2CHR|26|22|The other events of Uzziah's reign, from beginning to end, are recorded by the prophet Isaiah son of Amoz.
2CHR|26|23|Uzziah rested with his fathers and was buried near them in a field for burial that belonged to the kings, for people said, "He had leprosy." And Jotham his son succeeded him as king.
2CHR|27|1|Jotham was twenty-five years old when he became king, and he reigned in Jerusalem sixteen years. His mother's name was Jerusha daughter of Zadok.
2CHR|27|2|He did what was right in the eyes of the LORD, just as his father Uzziah had done, but unlike him he did not enter the temple of the LORD. The people, however, continued their corrupt practices.
2CHR|27|3|Jotham rebuilt the Upper Gate of the temple of the LORD and did extensive work on the wall at the hill of Ophel.
2CHR|27|4|He built towns in the Judean hills and forts and towers in the wooded areas.
2CHR|27|5|Jotham made war on the king of the Ammonites and conquered them. That year the Ammonites paid him a hundred talents of silver, ten thousand cors of wheat and ten thousand cors of barley. The Ammonites brought him the same amount also in the second and third years.
2CHR|27|6|Jotham grew powerful because he walked steadfastly before the LORD his God.
2CHR|27|7|The other events in Jotham's reign, including all his wars and the other things he did, are written in the book of the kings of Israel and Judah.
2CHR|27|8|He was twenty-five years old when he became king, and he reigned in Jerusalem sixteen years.
2CHR|27|9|Jotham rested with his fathers and was buried in the City of David. And Ahaz his son succeeded him as king.
2CHR|28|1|Ahaz was twenty years old when he became king, and he reigned in Jerusalem sixteen years. Unlike David his father, he did not do what was right in the eyes of the LORD.
2CHR|28|2|He walked in the ways of the kings of Israel and also made cast idols for worshiping the Baals.
2CHR|28|3|He burned sacrifices in the Valley of Ben Hinnom and sacrificed his sons in the fire, following the detestable ways of the nations the LORD had driven out before the Israelites.
2CHR|28|4|He offered sacrifices and burned incense at the high places, on the hilltops and under every spreading tree.
2CHR|28|5|Therefore the LORD his God handed him over to the king of Aram. The Arameans defeated him and took many of his people as prisoners and brought them to Damascus. He was also given into the hands of the king of Israel, who inflicted heavy casualties on him.
2CHR|28|6|In one day Pekah son of Remaliah killed a hundred and twenty thousand soldiers in Judah-because Judah had forsaken the LORD, the God of their fathers.
2CHR|28|7|Zicri, an Ephraimite warrior, killed Maaseiah the king's son, Azrikam the officer in charge of the palace, and Elkanah, second to the king.
2CHR|28|8|The Israelites took captive from their kinsmen two hundred thousand wives, sons and daughters. They also took a great deal of plunder, which they carried back to Samaria.
2CHR|28|9|But a prophet of the LORD named Oded was there, and he went out to meet the army when it returned to Samaria. He said to them, "Because the LORD, the God of your fathers, was angry with Judah, he gave them into your hand. But you have slaughtered them in a rage that reaches to heaven.
2CHR|28|10|And now you intend to make the men and women of Judah and Jerusalem your slaves. But aren't you also guilty of sins against the LORD your God?
2CHR|28|11|Now listen to me! Send back your fellow countrymen you have taken as prisoners, for the LORD's fierce anger rests on you."
2CHR|28|12|Then some of the leaders in Ephraim-Azariah son of Jehohanan, Berekiah son of Meshillemoth, Jehizkiah son of Shallum, and Amasa son of Hadlai-confronted those who were arriving from the war.
2CHR|28|13|"You must not bring those prisoners here," they said, "or we will be guilty before the LORD. Do you intend to add to our sin and guilt? For our guilt is already great, and his fierce anger rests on Israel."
2CHR|28|14|So the soldiers gave up the prisoners and plunder in the presence of the officials and all the assembly.
2CHR|28|15|The men designated by name took the prisoners, and from the plunder they clothed all who were naked. They provided them with clothes and sandals, food and drink, and healing balm. All those who were weak they put on donkeys. So they took them back to their fellow countrymen at Jericho, the City of Palms, and returned to Samaria.
2CHR|28|16|At that time King Ahaz sent to the king of Assyria for help.
2CHR|28|17|The Edomites had again come and attacked Judah and carried away prisoners,
2CHR|28|18|while the Philistines had raided towns in the foothills and in the Negev of Judah. They captured and occupied Beth Shemesh, Aijalon and Gederoth, as well as Soco, Timnah and Gimzo, with their surrounding villages.
2CHR|28|19|The LORD had humbled Judah because of Ahaz king of Israel, for he had promoted wickedness in Judah and had been most unfaithful to the LORD.
2CHR|28|20|Tiglath-Pileser king of Assyria came to him, but he gave him trouble instead of help.
2CHR|28|21|Ahaz took some of the things from the temple of the LORD and from the royal palace and from the princes and presented them to the king of Assyria, but that did not help him.
2CHR|28|22|In his time of trouble King Ahaz became even more unfaithful to the LORD.
2CHR|28|23|He offered sacrifices to the gods of Damascus, who had defeated him; for he thought, "Since the gods of the kings of Aram have helped them, I will sacrifice to them so they will help me." But they were his downfall and the downfall of all Israel.
2CHR|28|24|Ahaz gathered together the furnishings from the temple of God and took them away. He shut the doors of the LORD's temple and set up altars at every street corner in Jerusalem.
2CHR|28|25|In every town in Judah he built high places to burn sacrifices to other gods and provoked the LORD, the God of his fathers, to anger.
2CHR|28|26|The other events of his reign and all his ways, from beginning to end, are written in the book of the kings of Judah and Israel.
2CHR|28|27|Ahaz rested with his fathers and was buried in the city of Jerusalem, but he was not placed in the tombs of the kings of Israel. And Hezekiah his son succeeded him as king.
2CHR|29|1|Hezekiah was twenty-five years old when he became king, and he reigned in Jerusalem twenty-nine years. His mother's name was Abijah daughter of Zechariah.
2CHR|29|2|He did what was right in the eyes of the LORD, just as his father David had done.
2CHR|29|3|In the first month of the first year of his reign, he opened the doors of the temple of the LORD and repaired them.
2CHR|29|4|He brought in the priests and the Levites, assembled them in the square on the east side
2CHR|29|5|and said: "Listen to me, Levites! Consecrate yourselves now and consecrate the temple of the LORD, the God of your fathers. Remove all defilement from the sanctuary.
2CHR|29|6|Our fathers were unfaithful; they did evil in the eyes of the LORD our God and forsook him. They turned their faces away from the LORD's dwelling place and turned their backs on him.
2CHR|29|7|They also shut the doors of the portico and put out the lamps. They did not burn incense or present any burnt offerings at the sanctuary to the God of Israel.
2CHR|29|8|Therefore, the anger of the LORD has fallen on Judah and Jerusalem; he has made them an object of dread and horror and scorn, as you can see with your own eyes.
2CHR|29|9|This is why our fathers have fallen by the sword and why our sons and daughters and our wives are in captivity.
2CHR|29|10|Now I intend to make a covenant with the LORD, the God of Israel, so that his fierce anger will turn away from us.
2CHR|29|11|My sons, do not be negligent now, for the LORD has chosen you to stand before him and serve him, to minister before him and to burn incense."
2CHR|29|12|Then these Levites set to work: from the Kohathites, Mahath son of Amasai and Joel son of Azariah; from the Merarites, Kish son of Abdi and Azariah son of Jehallelel; from the Gershonites, Joah son of Zimmah and Eden son of Joah;
2CHR|29|13|from the descendants of Elizaphan, Shimri and Jeiel; from the descendants of Asaph, Zechariah and Mattaniah;
2CHR|29|14|from the descendants of Heman, Jehiel and Shimei; from the descendants of Jeduthun, Shemaiah and Uzziel.
2CHR|29|15|When they had assembled their brothers and consecrated themselves, they went in to purify the temple of the LORD, as the king had ordered, following the word of the LORD.
2CHR|29|16|The priests went into the sanctuary of the LORD to purify it. They brought out to the courtyard of the LORD's temple everything unclean that they found in the temple of the LORD. The Levites took it and carried it out to the Kidron Valley.
2CHR|29|17|They began the consecration on the first day of the first month, and by the eighth day of the month they reached the portico of the LORD. For eight more days they consecrated the temple of the LORD itself, finishing on the sixteenth day of the first month.
2CHR|29|18|Then they went in to King Hezekiah and reported: "We have purified the entire temple of the LORD, the altar of burnt offering with all its utensils, and the table for setting out the consecrated bread, with all its articles.
2CHR|29|19|We have prepared and consecrated all the articles that King Ahaz removed in his unfaithfulness while he was king. They are now in front of the LORD's altar."
2CHR|29|20|Early the next morning King Hezekiah gathered the city officials together and went up to the temple of the LORD.
2CHR|29|21|They brought seven bulls, seven rams, seven male lambs and seven male goats as a sin offering for the kingdom, for the sanctuary and for Judah. The king commanded the priests, the descendants of Aaron, to offer these on the altar of the LORD.
2CHR|29|22|So they slaughtered the bulls, and the priests took the blood and sprinkled it on the altar; next they slaughtered the rams and sprinkled their blood on the altar; then they slaughtered the lambs and sprinkled their blood on the altar.
2CHR|29|23|The goats for the sin offering were brought before the king and the assembly, and they laid their hands on them.
2CHR|29|24|The priests then slaughtered the goats and presented their blood on the altar for a sin offering to atone for all Israel, because the king had ordered the burnt offering and the sin offering for all Israel.
2CHR|29|25|He stationed the Levites in the temple of the LORD with cymbals, harps and lyres in the way prescribed by David and Gad the king's seer and Nathan the prophet; this was commanded by the LORD through his prophets.
2CHR|29|26|So the Levites stood ready with David's instruments, and the priests with their trumpets.
2CHR|29|27|Hezekiah gave the order to sacrifice the burnt offering on the altar. As the offering began, singing to the LORD began also, accompanied by trumpets and the instruments of David king of Israel.
2CHR|29|28|The whole assembly bowed in worship, while the singers sang and the trumpeters played. All this continued until the sacrifice of the burnt offering was completed.
2CHR|29|29|When the offerings were finished, the king and everyone present with him knelt down and worshiped.
2CHR|29|30|King Hezekiah and his officials ordered the Levites to praise the LORD with the words of David and of Asaph the seer. So they sang praises with gladness and bowed their heads and worshiped.
2CHR|29|31|Then Hezekiah said, "You have now dedicated yourselves to the LORD. Come and bring sacrifices and thank offerings to the temple of the LORD." So the assembly brought sacrifices and thank offerings, and all whose hearts were willing brought burnt offerings.
2CHR|29|32|The number of burnt offerings the assembly brought was seventy bulls, a hundred rams and two hundred male lambs-all of them for burnt offerings to the LORD.
2CHR|29|33|The animals consecrated as sacrifices amounted to six hundred bulls and three thousand sheep and goats.
2CHR|29|34|The priests, however, were too few to skin all the burnt offerings; so their kinsmen the Levites helped them until the task was finished and until other priests had been consecrated, for the Levites had been more conscientious in consecrating themselves than the priests had been.
2CHR|29|35|There were burnt offerings in abundance, together with the fat of the fellowship offerings and the drink offerings that accompanied the burnt offerings. So the service of the temple of the LORD was reestablished.
2CHR|29|36|Hezekiah and all the people rejoiced at what God had brought about for his people, because it was done so quickly.
2CHR|30|1|Hezekiah sent word to all Israel and Judah and also wrote letters to Ephraim and Manasseh, inviting them to come to the temple of the LORD in Jerusalem and celebrate the Passover to the LORD, the God of Israel.
2CHR|30|2|The king and his officials and the whole assembly in Jerusalem decided to celebrate the Passover in the second month.
2CHR|30|3|They had not been able to celebrate it at the regular time because not enough priests had consecrated themselves and the people had not assembled in Jerusalem.
2CHR|30|4|The plan seemed right both to the king and to the whole assembly.
2CHR|30|5|They decided to send a proclamation throughout Israel, from Beersheba to Dan, calling the people to come to Jerusalem and celebrate the Passover to the LORD, the God of Israel. It had not been celebrated in large numbers according to what was written.
2CHR|30|6|At the king's command, couriers went throughout Israel and Judah with letters from the king and from his officials, which read: "People of Israel, return to the LORD, the God of Abraham, Isaac and Israel, that he may return to you who are left, who have escaped from the hand of the kings of Assyria.
2CHR|30|7|Do not be like your fathers and brothers, who were unfaithful to the LORD, the God of their fathers, so that he made them an object of horror, as you see.
2CHR|30|8|Do not be stiff-necked, as your fathers were; submit to the LORD. Come to the sanctuary, which he has consecrated forever. Serve the LORD your God, so that his fierce anger will turn away from you.
2CHR|30|9|If you return to the LORD, then your brothers and your children will be shown compassion by their captors and will come back to this land, for the LORD your God is gracious and compassionate. He will not turn his face from you if you return to him."
2CHR|30|10|The couriers went from town to town in Ephraim and Manasseh, as far as Zebulun, but the people scorned and ridiculed them.
2CHR|30|11|Nevertheless, some men of Asher, Manasseh and Zebulun humbled themselves and went to Jerusalem.
2CHR|30|12|Also in Judah the hand of God was on the people to give them unity of mind to carry out what the king and his officials had ordered, following the word of the LORD.
2CHR|30|13|A very large crowd of people assembled in Jerusalem to celebrate the Feast of Unleavened Bread in the second month.
2CHR|30|14|They removed the altars in Jerusalem and cleared away the incense altars and threw them into the Kidron Valley.
2CHR|30|15|They slaughtered the Passover lamb on the fourteenth day of the second month. The priests and the Levites were ashamed and consecrated themselves and brought burnt offerings to the temple of the LORD.
2CHR|30|16|Then they took up their regular positions as prescribed in the Law of Moses the man of God. The priests sprinkled the blood handed to them by the Levites.
2CHR|30|17|Since many in the crowd had not consecrated themselves, the Levites had to kill the Passover lambs for all those who were not ceremonially clean and could not consecrate their lambs to the LORD.
2CHR|30|18|Although most of the many people who came from Ephraim, Manasseh, Issachar and Zebulun had not purified themselves, yet they ate the Passover, contrary to what was written. But Hezekiah prayed for them, saying, "May the LORD, who is good, pardon everyone
2CHR|30|19|who sets his heart on seeking God-the LORD, the God of his fathers-even if he is not clean according to the rules of the sanctuary."
2CHR|30|20|And the LORD heard Hezekiah and healed the people.
2CHR|30|21|The Israelites who were present in Jerusalem celebrated the Feast of Unleavened Bread for seven days with great rejoicing, while the Levites and priests sang to the LORD every day, accompanied by the LORD's instruments of praise.
2CHR|30|22|Hezekiah spoke encouragingly to all the Levites, who showed good understanding of the service of the LORD. For the seven days they ate their assigned portion and offered fellowship offerings and praised the LORD, the God of their fathers.
2CHR|30|23|The whole assembly then agreed to celebrate the festival seven more days; so for another seven days they celebrated joyfully.
2CHR|30|24|Hezekiah king of Judah provided a thousand bulls and seven thousand sheep and goats for the assembly, and the officials provided them with a thousand bulls and ten thousand sheep and goats. A great number of priests consecrated themselves.
2CHR|30|25|The entire assembly of Judah rejoiced, along with the priests and Levites and all who had assembled from Israel, including the aliens who had come from Israel and those who lived in Judah.
2CHR|30|26|There was great joy in Jerusalem, for since the days of Solomon son of David king of Israel there had been nothing like this in Jerusalem.
2CHR|30|27|The priests and the Levites stood to bless the people, and God heard them, for their prayer reached heaven, his holy dwelling place.
2CHR|31|1|When all this had ended, the Israelites who were there went out to the towns of Judah, smashed the sacred stones and cut down the Asherah poles. They destroyed the high places and the altars throughout Judah and Benjamin and in Ephraim and Manasseh. After they had destroyed all of them, the Israelites returned to their own towns and to their own property.
2CHR|31|2|Hezekiah assigned the priests and Levites to divisions-each of them according to their duties as priests or Levites-to offer burnt offerings and fellowship offerings, to minister, to give thanks and to sing praises at the gates of the LORD's dwelling.
2CHR|31|3|The king contributed from his own possessions for the morning and evening burnt offerings and for the burnt offerings on the Sabbaths, New Moons and appointed feasts as written in the Law of the LORD.
2CHR|31|4|He ordered the people living in Jerusalem to give the portion due the priests and Levites so they could devote themselves to the Law of the LORD.
2CHR|31|5|As soon as the order went out, the Israelites generously gave the firstfruits of their grain, new wine, oil and honey and all that the fields produced. They brought a great amount, a tithe of everything.
2CHR|31|6|The men of Israel and Judah who lived in the towns of Judah also brought a tithe of their herds and flocks and a tithe of the holy things dedicated to the LORD their God, and they piled them in heaps.
2CHR|31|7|They began doing this in the third month and finished in the seventh month.
2CHR|31|8|When Hezekiah and his officials came and saw the heaps, they praised the LORD and blessed his people Israel.
2CHR|31|9|Hezekiah asked the priests and Levites about the heaps;
2CHR|31|10|and Azariah the chief priest, from the family of Zadok, answered, "Since the people began to bring their contributions to the temple of the LORD, we have had enough to eat and plenty to spare, because the LORD has blessed his people, and this great amount is left over."
2CHR|31|11|Hezekiah gave orders to prepare storerooms in the temple of the LORD, and this was done.
2CHR|31|12|Then they faithfully brought in the contributions, tithes and dedicated gifts. Conaniah, a Levite, was in charge of these things, and his brother Shimei was next in rank.
2CHR|31|13|Jehiel, Azaziah, Nahath, Asahel, Jerimoth, Jozabad, Eliel, Ismakiah, Mahath and Benaiah were supervisors under Conaniah and Shimei his brother, by appointment of King Hezekiah and Azariah the official in charge of the temple of God.
2CHR|31|14|Kore son of Imnah the Levite, keeper of the East Gate, was in charge of the freewill offerings given to God, distributing the contributions made to the LORD and also the consecrated gifts.
2CHR|31|15|Eden, Miniamin, Jeshua, Shemaiah, Amariah and Shecaniah assisted him faithfully in the towns of the priests, distributing to their fellow priests according to their divisions, old and young alike.
2CHR|31|16|In addition, they distributed to the males three years old or more whose names were in the genealogical records-all who would enter the temple of the LORD to perform the daily duties of their various tasks, according to their responsibilities and their divisions.
2CHR|31|17|And they distributed to the priests enrolled by their families in the genealogical records and likewise to the Levites twenty years old or more, according to their responsibilities and their divisions.
2CHR|31|18|They included all the little ones, the wives, and the sons and daughters of the whole community listed in these genealogical records. For they were faithful in consecrating themselves.
2CHR|31|19|As for the priests, the descendants of Aaron, who lived on the farm lands around their towns or in any other towns, men were designated by name to distribute portions to every male among them and to all who were recorded in the genealogies of the Levites.
2CHR|31|20|This is what Hezekiah did throughout Judah, doing what was good and right and faithful before the LORD his God.
2CHR|31|21|In everything that he undertook in the service of God's temple and in obedience to the law and the commands, he sought his God and worked wholeheartedly. And so he prospered.
2CHR|32|1|After all that Hezekiah had so faithfully done, Sennacherib king of Assyria came and invaded Judah. He laid siege to the fortified cities, thinking to conquer them for himself.
2CHR|32|2|When Hezekiah saw that Sennacherib had come and that he intended to make war on Jerusalem,
2CHR|32|3|he consulted with his officials and military staff about blocking off the water from the springs outside the city, and they helped him.
2CHR|32|4|A large force of men assembled, and they blocked all the springs and the stream that flowed through the land. "Why should the kings of Assyria come and find plenty of water?" they said.
2CHR|32|5|Then he worked hard repairing all the broken sections of the wall and building towers on it. He built another wall outside that one and reinforced the supporting terraces of the City of David. He also made large numbers of weapons and shields.
2CHR|32|6|He appointed military officers over the people and assembled them before him in the square at the city gate and encouraged them with these words:
2CHR|32|7|"Be strong and courageous. Do not be afraid or discouraged because of the king of Assyria and the vast army with him, for there is a greater power with us than with him.
2CHR|32|8|With him is only the arm of flesh, but with us is the LORD our God to help us and to fight our battles." And the people gained confidence from what Hezekiah the king of Judah said.
2CHR|32|9|Later, when Sennacherib king of Assyria and all his forces were laying siege to Lachish, he sent his officers to Jerusalem with this message for Hezekiah king of Judah and for all the people of Judah who were there:
2CHR|32|10|"This is what Sennacherib king of Assyria says: On what are you basing your confidence, that you remain in Jerusalem under siege?
2CHR|32|11|When Hezekiah says, 'The LORD our God will save us from the hand of the king of Assyria,' he is misleading you, to let you die of hunger and thirst.
2CHR|32|12|Did not Hezekiah himself remove this god's high places and altars, saying to Judah and Jerusalem, 'You must worship before one altar and burn sacrifices on it'?
2CHR|32|13|"Do you not know what I and my fathers have done to all the peoples of the other lands? Were the gods of those nations ever able to deliver their land from my hand?
2CHR|32|14|Who of all the gods of these nations that my fathers destroyed has been able to save his people from me? How then can your god deliver you from my hand?
2CHR|32|15|Now do not let Hezekiah deceive you and mislead you like this. Do not believe him, for no god of any nation or kingdom has been able to deliver his people from my hand or the hand of my fathers. How much less will your god deliver you from my hand!"
2CHR|32|16|Sennacherib's officers spoke further against the LORD God and against his servant Hezekiah.
2CHR|32|17|The king also wrote letters insulting the LORD, the God of Israel, and saying this against him: "Just as the gods of the peoples of the other lands did not rescue their people from my hand, so the god of Hezekiah will not rescue his people from my hand."
2CHR|32|18|Then they called out in Hebrew to the people of Jerusalem who were on the wall, to terrify them and make them afraid in order to capture the city.
2CHR|32|19|They spoke about the God of Jerusalem as they did about the gods of the other peoples of the world-the work of men's hands.
2CHR|32|20|King Hezekiah and the prophet Isaiah son of Amoz cried out in prayer to heaven about this.
2CHR|32|21|And the LORD sent an angel, who annihilated all the fighting men and the leaders and officers in the camp of the Assyrian king. So he withdrew to his own land in disgrace. And when he went into the temple of his god, some of his sons cut him down with the sword.
2CHR|32|22|So the LORD saved Hezekiah and the people of Jerusalem from the hand of Sennacherib king of Assyria and from the hand of all others. He took care of them on every side.
2CHR|32|23|Many brought offerings to Jerusalem for the LORD and valuable gifts for Hezekiah king of Judah. From then on he was highly regarded by all the nations.
2CHR|32|24|In those days Hezekiah became ill and was at the point of death. He prayed to the LORD, who answered him and gave him a miraculous sign.
2CHR|32|25|But Hezekiah's heart was proud and he did not respond to the kindness shown him; therefore the LORD's wrath was on him and on Judah and Jerusalem.
2CHR|32|26|Then Hezekiah repented of the pride of his heart, as did the people of Jerusalem; therefore the LORD's wrath did not come upon them during the days of Hezekiah.
2CHR|32|27|Hezekiah had very great riches and honor, and he made treasuries for his silver and gold and for his precious stones, spices, shields and all kinds of valuables.
2CHR|32|28|He also made buildings to store the harvest of grain, new wine and oil; and he made stalls for various kinds of cattle, and pens for the flocks.
2CHR|32|29|He built villages and acquired great numbers of flocks and herds, for God had given him very great riches.
2CHR|32|30|It was Hezekiah who blocked the upper outlet of the Gihon spring and channeled the water down to the west side of the City of David. He succeeded in everything he undertook.
2CHR|32|31|But when envoys were sent by the rulers of Babylon to ask him about the miraculous sign that had occurred in the land, God left him to test him and to know everything that was in his heart.
2CHR|32|32|The other events of Hezekiah's reign and his acts of devotion are written in the vision of the prophet Isaiah son of Amoz in the book of the kings of Judah and Israel.
2CHR|32|33|Hezekiah rested with his fathers and was buried on the hill where the tombs of David's descendants are. All Judah and the people of Jerusalem honored him when he died. And Manasseh his son succeeded him as king.
2CHR|33|1|Manasseh was twelve years old when he became king, and he reigned in Jerusalem fifty-five years.
2CHR|33|2|He did evil in the eyes of the LORD, following the detestable practices of the nations the LORD had driven out before the Israelites.
2CHR|33|3|He rebuilt the high places his father Hezekiah had demolished; he also erected altars to the Baals and made Asherah poles. He bowed down to all the starry hosts and worshiped them.
2CHR|33|4|He built altars in the temple of the LORD, of which the LORD had said, "My Name will remain in Jerusalem forever."
2CHR|33|5|In both courts of the temple of the LORD, he built altars to all the starry hosts.
2CHR|33|6|He sacrificed his sons in the fire in the Valley of Ben Hinnom, practiced sorcery, divination and witchcraft, and consulted mediums and spiritists. He did much evil in the eyes of the LORD, provoking him to anger.
2CHR|33|7|He took the carved image he had made and put it in God's temple, of which God had said to David and to his son Solomon, "In this temple and in Jerusalem, which I have chosen out of all the tribes of Israel, I will put my Name forever.
2CHR|33|8|I will not again make the feet of the Israelites leave the land I assigned to your forefathers, if only they will be careful to do everything I commanded them concerning all the laws, decrees and ordinances given through Moses."
2CHR|33|9|But Manasseh led Judah and the people of Jerusalem astray, so that they did more evil than the nations the LORD had destroyed before the Israelites.
2CHR|33|10|The LORD spoke to Manasseh and his people, but they paid no attention.
2CHR|33|11|So the LORD brought against them the army commanders of the king of Assyria, who took Manasseh prisoner, put a hook in his nose, bound him with bronze shackles and took him to Babylon.
2CHR|33|12|In his distress he sought the favor of the LORD his God and humbled himself greatly before the God of his fathers.
2CHR|33|13|And when he prayed to him, the LORD was moved by his entreaty and listened to his plea; so he brought him back to Jerusalem and to his kingdom. Then Manasseh knew that the LORD is God.
2CHR|33|14|Afterward he rebuilt the outer wall of the City of David, west of the Gihon spring in the valley, as far as the entrance of the Fish Gate and encircling the hill of Ophel; he also made it much higher. He stationed military commanders in all the fortified cities in Judah.
2CHR|33|15|He got rid of the foreign gods and removed the image from the temple of the LORD, as well as all the altars he had built on the temple hill and in Jerusalem; and he threw them out of the city.
2CHR|33|16|Then he restored the altar of the LORD and sacrificed fellowship offerings and thank offerings on it, and told Judah to serve the LORD, the God of Israel.
2CHR|33|17|The people, however, continued to sacrifice at the high places, but only to the LORD their God.
2CHR|33|18|The other events of Manasseh's reign, including his prayer to his God and the words the seers spoke to him in the name of the LORD, the God of Israel, are written in the annals of the kings of Israel.
2CHR|33|19|His prayer and how God was moved by his entreaty, as well as all his sins and unfaithfulness, and the sites where he built high places and set up Asherah poles and idols before he humbled himself-all are written in the records of the seers.
2CHR|33|20|Manasseh rested with his fathers and was buried in his palace. And Amon his son succeeded him as king.
2CHR|33|21|Amon was twenty-two years old when he became king, and he reigned in Jerusalem two years.
2CHR|33|22|He did evil in the eyes of the LORD, as his father Manasseh had done. Amon worshiped and offered sacrifices to all the idols Manasseh had made.
2CHR|33|23|But unlike his father Manasseh, he did not humble himself before the LORD; Amon increased his guilt.
2CHR|33|24|Amon's officials conspired against him and assassinated him in his palace.
2CHR|33|25|Then the people of the land killed all who had plotted against King Amon, and they made Josiah his son king in his place.
2CHR|34|1|Josiah was eight years old when he became king, and he reigned in Jerusalem thirty-one years.
2CHR|34|2|He did what was right in the eyes of the LORD and walked in the ways of his father David, not turning aside to the right or to the left.
2CHR|34|3|In the eighth year of his reign, while he was still young, he began to seek the God of his father David. In his twelfth year he began to purge Judah and Jerusalem of high places, Asherah poles, carved idols and cast images.
2CHR|34|4|Under his direction the altars of the Baals were torn down; he cut to pieces the incense altars that were above them, and smashed the Asherah poles, the idols and the images. These he broke to pieces and scattered over the graves of those who had sacrificed to them.
2CHR|34|5|He burned the bones of the priests on their altars, and so he purged Judah and Jerusalem.
2CHR|34|6|In the towns of Manasseh, Ephraim and Simeon, as far as Naphtali, and in the ruins around them,
2CHR|34|7|he tore down the altars and the Asherah poles and crushed the idols to powder and cut to pieces all the incense altars throughout Israel. Then he went back to Jerusalem.
2CHR|34|8|In the eighteenth year of Josiah's reign, to purify the land and the temple, he sent Shaphan son of Azaliah and Maaseiah the ruler of the city, with Joah son of Joahaz, the recorder, to repair the temple of the LORD his God.
2CHR|34|9|They went to Hilkiah the high priest and gave him the money that had been brought into the temple of God, which the Levites who were the doorkeepers had collected from the people of Manasseh, Ephraim and the entire remnant of Israel and from all the people of Judah and Benjamin and the inhabitants of Jerusalem.
2CHR|34|10|Then they entrusted it to the men appointed to supervise the work on the LORD's temple. These men paid the workers who repaired and restored the temple.
2CHR|34|11|They also gave money to the carpenters and builders to purchase dressed stone, and timber for joists and beams for the buildings that the kings of Judah had allowed to fall into ruin.
2CHR|34|12|The men did the work faithfully. Over them to direct them were Jahath and Obadiah, Levites descended from Merari, and Zechariah and Meshullam, descended from Kohath. The Levites-all who were skilled in playing musical instruments-
2CHR|34|13|had charge of the laborers and supervised all the workers from job to job. Some of the Levites were secretaries, scribes and doorkeepers.
2CHR|34|14|While they were bringing out the money that had been taken into the temple of the LORD, Hilkiah the priest found the Book of the Law of the LORD that had been given through Moses.
2CHR|34|15|Hilkiah said to Shaphan the secretary, "I have found the Book of the Law in the temple of the LORD." He gave it to Shaphan.
2CHR|34|16|Then Shaphan took the book to the king and reported to him: "Your officials are doing everything that has been committed to them.
2CHR|34|17|They have paid out the money that was in the temple of the LORD and have entrusted it to the supervisors and workers."
2CHR|34|18|Then Shaphan the secretary informed the king, "Hilkiah the priest has given me a book." And Shaphan read from it in the presence of the king.
2CHR|34|19|When the king heard the words of the Law, he tore his robes.
2CHR|34|20|He gave these orders to Hilkiah, Ahikam son of Shaphan, Abdon son of Micah, Shaphan the secretary and Asaiah the king's attendant:
2CHR|34|21|"Go and inquire of the LORD for me and for the remnant in Israel and Judah about what is written in this book that has been found. Great is the LORD's anger that is poured out on us because our fathers have not kept the word of the LORD; they have not acted in accordance with all that is written in this book."
2CHR|34|22|Hilkiah and those the king had sent with him went to speak to the prophetess Huldah, who was the wife of Shallum son of Tokhath, the son of Hasrah, keeper of the wardrobe. She lived in Jerusalem, in the Second District.
2CHR|34|23|She said to them, "This is what the LORD, the God of Israel, says: Tell the man who sent you to me,
2CHR|34|24|'This is what the LORD says: I am going to bring disaster on this place and its people-all the curses written in the book that has been read in the presence of the king of Judah.
2CHR|34|25|Because they have forsaken me and burned incense to other gods and provoked me to anger by all that their hands have made, my anger will be poured out on this place and will not be quenched.'
2CHR|34|26|Tell the king of Judah, who sent you to inquire of the LORD, 'This is what the LORD, the God of Israel, says concerning the words you heard:
2CHR|34|27|Because your heart was responsive and you humbled yourself before God when you heard what he spoke against this place and its people, and because you humbled yourself before me and tore your robes and wept in my presence, I have heard you, declares the LORD.
2CHR|34|28|Now I will gather you to your fathers, and you will be buried in peace. Your eyes will not see all the disaster I am going to bring on this place and on those who live here.'" So they took her answer back to the king.
2CHR|34|29|Then the king called together all the elders of Judah and Jerusalem.
2CHR|34|30|He went up to the temple of the LORD with the men of Judah, the people of Jerusalem, the priests and the Levites-all the people from the least to the greatest. He read in their hearing all the words of the Book of the Covenant, which had been found in the temple of the LORD.
2CHR|34|31|The king stood by his pillar and renewed the covenant in the presence of the LORD -to follow the LORD and keep his commands, regulations and decrees with all his heart and all his soul, and to obey the words of the covenant written in this book.
2CHR|34|32|Then he had everyone in Jerusalem and Benjamin pledge themselves to it; the people of Jerusalem did this in accordance with the covenant of God, the God of their fathers.
2CHR|34|33|Josiah removed all the detestable idols from all the territory belonging to the Israelites, and he had all who were present in Israel serve the LORD their God. As long as he lived, they did not fail to follow the LORD, the God of their fathers.
2CHR|35|1|Josiah celebrated the Passover to the LORD in Jerusalem, and the Passover lamb was slaughtered on the fourteenth day of the first month.
2CHR|35|2|He appointed the priests to their duties and encouraged them in the service of the LORD's temple.
2CHR|35|3|He said to the Levites, who instructed all Israel and who had been consecrated to the LORD: "Put the sacred ark in the temple that Solomon son of David king of Israel built. It is not to be carried about on your shoulders. Now serve the LORD your God and his people Israel.
2CHR|35|4|Prepare yourselves by families in your divisions, according to the directions written by David king of Israel and by his son Solomon.
2CHR|35|5|"Stand in the holy place with a group of Levites for each subdivision of the families of your fellow countrymen, the lay people.
2CHR|35|6|Slaughter the Passover lambs, consecrate yourselves and prepare the lambs for your fellow countrymen, doing what the LORD commanded through Moses."
2CHR|35|7|Josiah provided for all the lay people who were there a total of thirty thousand sheep and goats for the Passover offerings, and also three thousand cattle-all from the king's own possessions.
2CHR|35|8|His officials also contributed voluntarily to the people and the priests and Levites. Hilkiah, Zechariah and Jehiel, the administrators of God's temple, gave the priests twenty-six hundred Passover offerings and three hundred cattle.
2CHR|35|9|Also Conaniah along with Shemaiah and Nethanel, his brothers, and Hashabiah, Jeiel and Jozabad, the leaders of the Levites, provided five thousand Passover offerings and five hundred head of cattle for the Levites.
2CHR|35|10|The service was arranged and the priests stood in their places with the Levites in their divisions as the king had ordered.
2CHR|35|11|The Passover lambs were slaughtered, and the priests sprinkled the blood handed to them, while the Levites skinned the animals.
2CHR|35|12|They set aside the burnt offerings to give them to the subdivisions of the families of the people to offer to the LORD, as is written in the Book of Moses. They did the same with the cattle.
2CHR|35|13|They roasted the Passover animals over the fire as prescribed, and boiled the holy offerings in pots, caldrons and pans and served them quickly to all the people.
2CHR|35|14|After this, they made preparations for themselves and for the priests, because the priests, the descendants of Aaron, were sacrificing the burnt offerings and the fat portions until nightfall. So the Levites made preparations for themselves and for the Aaronic priests.
2CHR|35|15|The musicians, the descendants of Asaph, were in the places prescribed by David, Asaph, Heman and Jeduthun the king's seer. The gatekeepers at each gate did not need to leave their posts, because their fellow Levites made the preparations for them.
2CHR|35|16|So at that time the entire service of the LORD was carried out for the celebration of the Passover and the offering of burnt offerings on the altar of the LORD, as King Josiah had ordered.
2CHR|35|17|The Israelites who were present celebrated the Passover at that time and observed the Feast of Unleavened Bread for seven days.
2CHR|35|18|The Passover had not been observed like this in Israel since the days of the prophet Samuel; and none of the kings of Israel had ever celebrated such a Passover as did Josiah, with the priests, the Levites and all Judah and Israel who were there with the people of Jerusalem.
2CHR|35|19|This Passover was celebrated in the eighteenth year of Josiah's reign.
2CHR|35|20|After all this, when Josiah had set the temple in order, Neco king of Egypt went up to fight at Carchemish on the Euphrates, and Josiah marched out to meet him in battle.
2CHR|35|21|But Neco sent messengers to him, saying, "What quarrel is there between you and me, O king of Judah? It is not you I am attacking at this time, but the house with which I am at war. God has told me to hurry; so stop opposing God, who is with me, or he will destroy you."
2CHR|35|22|Josiah, however, would not turn away from him, but disguised himself to engage him in battle. He would not listen to what Neco had said at God's command but went to fight him on the plain of Megiddo.
2CHR|35|23|Archers shot King Josiah, and he told his officers, "Take me away; I am badly wounded."
2CHR|35|24|So they took him out of his chariot, put him in the other chariot he had and brought him to Jerusalem, where he died. He was buried in the tombs of his fathers, and all Judah and Jerusalem mourned for him.
2CHR|35|25|Jeremiah composed laments for Josiah, and to this day all the men and women singers commemorate Josiah in the laments. These became a tradition in Israel and are written in the Laments.
2CHR|35|26|The other events of Josiah's reign and his acts of devotion, according to what is written in the Law of the LORD -
2CHR|35|27|all the events, from beginning to end, are written in the book of the kings of Israel and Judah.
2CHR|36|1|And the people of the land took Jehoahaz son of Josiah and made him king in Jerusalem in place of his father.
2CHR|36|2|Jehoahaz was twenty-three years old when he became king, and he reigned in Jerusalem three months.
2CHR|36|3|The king of Egypt dethroned him in Jerusalem and imposed on Judah a levy of a hundred talents of silver and a talent of gold.
2CHR|36|4|The king of Egypt made Eliakim, a brother of Jehoahaz, king over Judah and Jerusalem and changed Eliakim's name to Jehoiakim. But Neco took Eliakim's brother Jehoahaz and carried him off to Egypt.
2CHR|36|5|Jehoiakim was twenty-five years old when he became king, and he reigned in Jerusalem eleven years. He did evil in the eyes of the LORD his God.
2CHR|36|6|Nebuchadnezzar king of Babylon attacked him and bound him with bronze shackles to take him to Babylon.
2CHR|36|7|Nebuchadnezzar also took to Babylon articles from the temple of the LORD and put them in his temple there.
2CHR|36|8|The other events of Jehoiakim's reign, the detestable things he did and all that was found against him, are written in the book of the kings of Israel and Judah. And Jehoiachin his son succeeded him as king.
2CHR|36|9|Jehoiachin was eighteen years old when he became king, and he reigned in Jerusalem three months and ten days. He did evil in the eyes of the LORD.
2CHR|36|10|In the spring, King Nebuchadnezzar sent for him and brought him to Babylon, together with articles of value from the temple of the LORD, and he made Jehoiachin's uncle, Zedekiah, king over Judah and Jerusalem.
2CHR|36|11|Zedekiah was twenty-one years old when he became king, and he reigned in Jerusalem eleven years.
2CHR|36|12|He did evil in the eyes of the LORD his God and did not humble himself before Jeremiah the prophet, who spoke the word of the LORD.
2CHR|36|13|He also rebelled against King Nebuchadnezzar, who had made him take an oath in God's name. He became stiff-necked and hardened his heart and would not turn to the LORD, the God of Israel.
2CHR|36|14|Furthermore, all the leaders of the priests and the people became more and more unfaithful, following all the detestable practices of the nations and defiling the temple of the LORD, which he had consecrated in Jerusalem.
2CHR|36|15|The LORD, the God of their fathers, sent word to them through his messengers again and again, because he had pity on his people and on his dwelling place.
2CHR|36|16|But they mocked God's messengers, despised his words and scoffed at his prophets until the wrath of the LORD was aroused against his people and there was no remedy.
2CHR|36|17|He brought up against them the king of the Babylonians, who killed their young men with the sword in the sanctuary, and spared neither young man nor young woman, old man or aged. God handed all of them over to Nebuchadnezzar.
2CHR|36|18|He carried to Babylon all the articles from the temple of God, both large and small, and the treasures of the LORD's temple and the treasures of the king and his officials.
2CHR|36|19|They set fire to God's temple and broke down the wall of Jerusalem; they burned all the palaces and destroyed everything of value there.
2CHR|36|20|He carried into exile to Babylon the remnant, who escaped from the sword, and they became servants to him and his sons until the kingdom of Persia came to power.
2CHR|36|21|The land enjoyed its sabbath rests; all the time of its desolation it rested, until the seventy years were completed in fulfillment of the word of the LORD spoken by Jeremiah.
2CHR|36|22|In the first year of Cyrus king of Persia, in order to fulfill the word of the LORD spoken by Jeremiah, the LORD moved the heart of Cyrus king of Persia to make a proclamation throughout his realm and to put it in writing:
2CHR|36|23|"This is what Cyrus king of Persia says: "'The LORD, the God of heaven, has given me all the kingdoms of the earth and he has appointed me to build a temple for him at Jerusalem in Judah. Anyone of his people among you-may the LORD his God be with him, and let him go up.'"
