2THESS|1|1|Павло, і Силуан, і Тимофій до Солунської Церкви в нашім Бозі Отці й Господі Ісусі Христі:
2THESS|1|2|благодать вам і мир від Бога Отця й Господа Ісуса Христа!
2THESS|1|3|Ми завжди повинні подяку складати за вас Богові, браття, як і годиться, бо сильно росте віра ваша, і примножується любов кожного з усіх вас один до одного.
2THESS|1|4|Так що ми самі хвалимось вами по Божих Церквах за ваші страждання та віру в усіх переслідуваннях ваших та в утисках, що їх переносите ви.
2THESS|1|5|А це доказ праведного Божого суду, щоб стали ви гідні Божого Царства, що за нього й страждаєте ви!
2THESS|1|6|Бо то справедливе в Бога віддати утиском тим, хто вас утискає,
2THESS|1|7|а вам, хто утиски терпить, відпочинок із нами, коли з'явиться з неба Господь Ісус з Анголами сили Своєї,
2THESS|1|8|в огні полум'яному, що даватиме помсту на тих, хто Бога не знає, і не слухає Євангелії Господа нашого Ісуса.
2THESS|1|9|Вони кару приймуть, вічну погибіль від лиця Господнього та від слави потуги Його,
2THESS|1|10|як Він прийде того дня прославитися в Своїх святих, і стати дивним у всіх віруючих, бо свідчення наше знайшло віру між вами.
2THESS|1|11|За це ми й молимось завжди за вас, щоб наш Бог учинив вас гідними покликання, і міццю наповнив усю добру волю добрости й діло віри,
2THESS|1|12|щоб прославилося Ім'я Господа нашого Ісуса в вас, а ви в Ньому, за благодаттю Бога нашого й Господа Ісуса Христа.
2THESS|2|1|Благаємо ж, браття, ми вас, щодо приходу Господа нашого Ісуса Христа й нашого згромадження до Нього,
2THESS|2|2|щоб ви не хвилювалися зараз умом та не жахались ані через духа, ані через слово, ані через листа, що він ніби від нас, ніби вже настав день Господній.
2THESS|2|3|Хай ніхто жадним способом вас не зведе! Бо той день не настане, аж перше прийде відступлення, і виявиться беззаконник, призначений на погибіль,
2THESS|2|4|що противиться та несеться над усе, зване Богом чи святощами, так що в Божому храмі він сяде, як Бог, і за Бога себе видаватиме.
2THESS|2|5|Чи ви не пам'ятаєте, як, ще в вас живши, я це вам говорив був?
2THESS|2|6|І тепер ви знаєте, що саме не допускає з'явитись йому своєчасно.
2THESS|2|7|Бо вже діється таємниця беззаконня; тільки той, хто тримає тепер, буде тримати, аж поки не буде усунений він із середини.
2THESS|2|8|І тоді то з'явиться той беззаконник, що його Господь Ісус заб'є Духом уст Своїх і знищить з'явленням приходу Свого.
2THESS|2|9|Його прихід за чином сатани буде з усякою силою й знаками та з неправдивими чудами,
2THESS|2|10|і з усякою обманою неправди між тими, хто гине, бо любови правди вони не прийняли, щоб їм спастися.
2THESS|2|11|І за це Бог пошле їм дію обмани, щоб у неправду повірили,
2THESS|2|12|щоб стали засуджені всі, хто не вірив у правду, але полюбив неправду.
2THESS|2|13|А ми завжди повинні дякувати Богові за вас, улюблені Господом браття, що Бог вибрав вас спочатку на спасіння освяченням Духа та вірою в правду,
2THESS|2|14|до чого покликав Він вас через нашу Євангелію, щоб отримати славу Господа нашого Ісуса Христа.
2THESS|2|15|Отже, браття, стійте й тримайтеся передань, яких ви навчились чи то словом, чи нашим посланням.
2THESS|2|16|Сам же Господь наш Ісус Христос і Бог Отець наш, що нас полюбив і дав у благодаті вічну потіху та добру надію,
2THESS|2|17|нехай ваші серця Він потішить, і нехай Він зміцнить вас у всякому доброму ділі та в слові!
2THESS|3|1|Наостанку, моліться, браття, за нас, щоб ширилось Слово Господнє та славилось, як і в вас,
2THESS|3|2|і щоб ми визволилися від злих та лукавих людей, бо віра не в усіх.
2THESS|3|3|І вірний Господь, що зміцнить вас і збереже від лукавого.
2THESS|3|4|А про вас покладаємо надію на Господа, що й чините ви, і чинити будете те, що наказуємо вам.
2THESS|3|5|Господь же нехай серця ваші спрямує на Божу любов та терпеливість Христову!
2THESS|3|6|А ми вам наказуємо, браття, Ім'ям Господа Ісуса Христа, щоб ви цуралися кожного брата, що живе по-ледачому, а не за переданням, яке прийняли ви від нас.
2THESS|3|7|Самі бо ви знаєте, як належить наслідувати нас. Бо ми поміж вами не сидні справляли,
2THESS|3|8|і хліба не їли ні в кого даремно, але в перевтомі й напруженні день і ніч працювали, щоб не бути нікому із вас тягарем,
2THESS|3|9|не тому, щоб ми влади не мали, але щоб себе за взірця дати вам, щоб нас ви наслідували.
2THESS|3|10|Бо коли ми в вас перебували, то це вам наказували, що як хто працювати не хоче, нехай той не їсть!
2THESS|3|11|Бо ми чуємо, що дехто між вами живуть по-ледачому, нічого не роблять, а тільки вдають, ніби роблять.
2THESS|3|12|Таким ми наказуємо та благаємо Господом нашим Ісусом Христом, щоб мовчки вони працювали та власний хліб їли.
2THESS|3|13|А ви, браття, не втомлюйтеся, коли чините добре.
2THESS|3|14|Коли ж хто не послухає нашого слова через цього листа, зауважте того, і не майте з ним зносин, щоб він був посоромлений.
2THESS|3|15|Та не майте його за неприятеля, а навчайте, як брата.
2THESS|3|16|А Сам Господь миру нехай завжди дасть вам мир усяким способом. Господь з вами всіма!
2THESS|3|17|Привіт вам моєю рукою Павловою, це править за знака в усякім листі. Так пишу я.
2THESS|3|18|Благодать Господа нашого Ісуса Христа нехай буде з вами всіма! Амінь.
