2PET|1|1|Simon Peter, a servant and apostle of Jesus Christ, To those who through the righteousness of our God and Savior Jesus Christ have received a faith as precious as ours:
2PET|1|2|Grace and peace be yours in abundance through the knowledge of God and of Jesus our Lord.
2PET|1|3|His divine power has given us everything we need for life and godliness through our knowledge of him who called us by his own glory and goodness.
2PET|1|4|Through these he has given us his very great and precious promises, so that through them you may participate in the divine nature and escape the corruption in the world caused by evil desires.
2PET|1|5|For this very reason, make every effort to add to your faith goodness; and to goodness, knowledge;
2PET|1|6|and to knowledge, self-control; and to self-control, perseverance; and to perseverance, godliness;
2PET|1|7|and to godliness, brotherly kindness; and to brotherly kindness, love.
2PET|1|8|For if you possess these qualities in increasing measure, they will keep you from being ineffective and unproductive in your knowledge of our Lord Jesus Christ.
2PET|1|9|But if anyone does not have them, he is nearsighted and blind, and has forgotten that he has been cleansed from his past sins.
2PET|1|10|Therefore, my brothers, be all the more eager to make your calling and election sure. For if you do these things, you will never fall,
2PET|1|11|and you will receive a rich welcome into the eternal kingdom of our Lord and Savior Jesus Christ.
2PET|1|12|So I will always remind you of these things, even though you know them and are firmly established in the truth you now have.
2PET|1|13|I think it is right to refresh your memory as long as I live in the tent of this body,
2PET|1|14|because I know that I will soon put it aside, as our Lord Jesus Christ has made clear to me.
2PET|1|15|And I will make every effort to see that after my departure you will always be able to remember these things.
2PET|1|16|We did not follow cleverly invented stories when we told you about the power and coming of our Lord Jesus Christ, but we were eyewitnesses of his majesty.
2PET|1|17|For he received honor and glory from God the Father when the voice came to him from the Majestic Glory, saying, "This is my Son, whom I love; with him I am well pleased."
2PET|1|18|We ourselves heard this voice that came from heaven when we were with him on the sacred mountain.
2PET|1|19|And we have the word of the prophets made more certain, and you will do well to pay attention to it, as to a light shining in a dark place, until the day dawns and the morning star rises in your hearts.
2PET|1|20|Above all, you must understand that no prophecy of Scripture came about by the prophet's own interpretation.
2PET|1|21|For prophecy never had its origin in the will of man, but men spoke from God as they were carried along by the Holy Spirit.
2PET|2|1|But there were also false prophets among the people, just as there will be false teachers among you. They will secretly introduce destructive heresies, even denying the sovereign Lord who bought them--bringing swift destruction on themselves.
2PET|2|2|Many will follow their shameful ways and will bring the way of truth into disrepute.
2PET|2|3|In their greed these teachers will exploit you with stories they have made up. Their condemnation has long been hanging over them, and their destruction has not been sleeping.
2PET|2|4|For if God did not spare angels when they sinned, but sent them to hell, putting them into gloomy dungeons to be held for judgment;
2PET|2|5|if he did not spare the ancient world when he brought the flood on its ungodly people, but protected Noah, a preacher of righteousness, and seven others;
2PET|2|6|if he condemned the cities of Sodom and Gomorrah by burning them to ashes, and made them an example of what is going to happen to the ungodly;
2PET|2|7|and if he rescued Lot, a righteous man, who was distressed by the filthy lives of lawless men
2PET|2|8|(for that righteous man, living among them day after day, was tormented in his righteous soul by the lawless deeds he saw and heard)--
2PET|2|9|if this is so, then the Lord knows how to rescue godly men from trials and to hold the unrighteous for the day of judgment, while continuing their punishment.
2PET|2|10|This is especially true of those who follow the corrupt desire of the sinful nature and despise authority.
2PET|2|11|Bold and arrogant, these men are not afraid to slander celestial beings; yet even angels, although they are stronger and more powerful, do not bring slanderous accusations against such beings in the presence of the Lord.
2PET|2|12|But these men blaspheme in matters they do not understand. They are like brute beasts, creatures of instinct, born only to be caught and destroyed, and like beasts they too will perish.
2PET|2|13|They will be paid back with harm for the harm they have done. Their idea of pleasure is to carouse in broad daylight. They are blots and blemishes, reveling in their pleasures while they feast with you.
2PET|2|14|With eyes full of adultery, they never stop sinning; they seduce the unstable; they are experts in greed--an accursed brood!
2PET|2|15|They have left the straight way and wandered off to follow the way of Balaam son of Beor, who loved the wages of wickedness.
2PET|2|16|But he was rebuked for his wrongdoing by a donkey--a beast without speech--who spoke with a man's voice and restrained the prophet's madness.
2PET|2|17|These men are springs without water and mists driven by a storm. Blackest darkness is reserved for them.
2PET|2|18|For they mouth empty, boastful words and, by appealing to the lustful desires of sinful human nature, they entice people who are just escaping from those who live in error.
2PET|2|19|They promise them freedom, while they themselves are slaves of depravity--for a man is a slave to whatever has mastered him.
2PET|2|20|If they have escaped the corruption of the world by knowing our Lord and Savior Jesus Christ and are again entangled in it and overcome, they are worse off at the end than they were at the beginning.
2PET|2|21|It would have been better for them not to have known the way of righteousness, than to have known it and then to turn their backs on the sacred command that was passed on to them.
2PET|2|22|Of them the proverbs are true: "A dog returns to its vomit," and, "A sow that is washed goes back to her wallowing in the mud."
2PET|3|1|Dear friends, this is now my second letter to you. I have written both of them as reminders to stimulate you to wholesome thinking.
2PET|3|2|I want you to recall the words spoken in the past by the holy prophets and the command given by our Lord and Savior through your apostles.
2PET|3|3|First of all, you must understand that in the last days scoffers will come, scoffing and following their own evil desires.
2PET|3|4|They will say, "Where is this 'coming' he promised? Ever since our fathers died, everything goes on as it has since the beginning of creation."
2PET|3|5|But they deliberately forget that long ago by God's word the heavens existed and the earth was formed out of water and by water.
2PET|3|6|By these waters also the world of that time was deluged and destroyed.
2PET|3|7|By the same word the present heavens and earth are reserved for fire, being kept for the day of judgment and destruction of ungodly men.
2PET|3|8|But do not forget this one thing, dear friends: With the Lord a day is like a thousand years, and a thousand years are like a day.
2PET|3|9|The Lord is not slow in keeping his promise, as some understand slowness. He is patient with you, not wanting anyone to perish, but everyone to come to repentance.
2PET|3|10|But the day of the Lord will come like a thief. The heavens will disappear with a roar; the elements will be destroyed by fire, and the earth and everything in it will be laid bare.
2PET|3|11|Since everything will be destroyed in this way, what kind of people ought you to be? You ought to live holy and godly lives
2PET|3|12|as you look forward to the day of God and speed its coming. That day will bring about the destruction of the heavens by fire, and the elements will melt in the heat.
2PET|3|13|But in keeping with his promise we are looking forward to a new heaven and a new earth, the home of righteousness.
2PET|3|14|So then, dear friends, since you are looking forward to this, make every effort to be found spotless, blameless and at peace with him.
2PET|3|15|Bear in mind that our Lord's patience means salvation, just as our dear brother Paul also wrote you with the wisdom that God gave him.
2PET|3|16|He writes the same way in all his letters, speaking in them of these matters. His letters contain some things that are hard to understand, which ignorant and unstable people distort, as they do the other Scriptures, to their own destruction.
2PET|3|17|Therefore, dear friends, since you already know this, be on your guard so that you may not be carried away by the error of lawless men and fall from your secure position.
2PET|3|18|But grow in the grace and knowledge of our Lord and Savior Jesus Christ. To him be glory both now and forever! Amen.
