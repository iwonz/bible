MATT|1|1|亚伯拉罕 的后裔、 大卫 的子孙 耶稣基督的家谱：
MATT|1|2|亚伯拉罕 生 以撒 ， 以撒 生 雅各 ， 雅各 生 犹大 和他的兄弟，
MATT|1|3|犹大 从 她玛 氏生 法勒斯 和 谢拉 ， 法勒斯 生 希斯仑 ， 希斯仑 生 亚兰 ，
MATT|1|4|亚兰 生 亚米拿达 ， 亚米拿达 生 拿顺 ， 拿顺 生 撒门 ，
MATT|1|5|撒门 从 喇合 氏生 波阿斯 ， 波阿斯 从 路得 氏生 俄备得 ， 俄备得 生 耶西 ，
MATT|1|6|耶西 生 大卫 王。 大卫 从 乌利亚 的妻子生 所罗门 ，
MATT|1|7|所罗门 生 罗波安 ， 罗波安 生 亚比雅 ， 亚比雅 生 亚撒 ，
MATT|1|8|亚撒 生 约沙法 ， 约沙法 生 约兰 ， 约兰 生 乌西雅 ，
MATT|1|9|乌西雅 生 约坦 ， 约坦 生 亚哈斯 ， 亚哈斯 生 希西家 ，
MATT|1|10|希西家 生 玛拿西 ， 玛拿西 生 亚们 ， 亚们 生 约西亚 ，
MATT|1|11|百姓被迁到 巴比伦 的时候， 约西亚 生 耶哥尼雅 和他的兄弟。
MATT|1|12|迁到 巴比伦 之后， 耶哥尼雅 生 撒拉铁 ， 撒拉铁 生 所罗巴伯 ，
MATT|1|13|所罗巴伯 生 亚比玉 ， 亚比玉 生 以利亚敬 ， 以利亚敬 生 亚所 ，
MATT|1|14|亚所 生 撒督 ， 撒督 生 亚金 ， 亚金 生 以律 ，
MATT|1|15|以律 生 以利亚撒 ， 以利亚撒 生 马但 ， 马但 生 雅各 ，
MATT|1|16|雅各 生 约瑟 ，就是 马利亚 的丈夫；那称为基督的耶稣是从 马利亚 生的。
MATT|1|17|这样，从 亚伯拉罕 到 大卫 共有十四代，从 大卫 到迁至 巴比伦 的时候也有十四代，从迁至 巴比伦 的时候到基督又有十四代。
MATT|1|18|耶稣基督降生的事记在下面：他母亲 马利亚 已经许配给 约瑟 ，还没有迎娶， 马利亚 就从圣灵怀了孕。
MATT|1|19|她丈夫 约瑟 是个义人，不愿意当众羞辱她，想要暗地里把她休了。
MATT|1|20|正考虑这些事的时候，忽然主的使者在 约瑟 梦中向他显现，说：“ 大卫 的子孙 约瑟 ，不要怕，把你的妻子 马利亚 娶过来，因她所怀的孕是从圣灵来的。
MATT|1|21|她将要生一个儿子，你要给他起名叫耶稣，因他要将自己的百姓从罪恶里救出来。”
MATT|1|22|这整件事的发生，是要应验主藉先知所说的话：
MATT|1|23|“必有童女怀孕生子； 人要称他的名为 以马内利 。” （ 以马内利 翻出来就是“上帝与我们同在”。）
MATT|1|24|约瑟 醒来，就遵照主的使者的吩咐把妻子娶过来；
MATT|1|25|但是没有和她同房，直到她生了儿子 ，就给他起名叫耶稣。
MATT|2|1|在 希律 作王的时候，耶稣生在 犹太 的 伯利恒 。有几个博学之士 从东方来到 耶路撒冷 ，说：
MATT|2|2|“那生下来作 犹太 人之王的在哪里？我们在东方看见他的星，特来拜他。”
MATT|2|3|希律 王听见了，就心里不安； 耶路撒冷 全城的人也都不安。
MATT|2|4|他就召集了祭司长和民间的文士，问他们：“基督该生在哪里？”
MATT|2|5|他们说：“在 犹太 的 伯利恒 。因为有先知记着：
MATT|2|6|‘ 犹大 地的 伯利恒 啊， 你在 犹大 诸城中并不是最小的； 因为将来有一位统治者要从你那里出来， 牧养我 以色列 民。’”
MATT|2|7|于是， 希律 暗地里召了博学之士来，查问那星是什么时候出现的，
MATT|2|8|就派他们往 伯利恒 去，说：“你们去仔细寻访那小孩子，找到了就来报信，我也好去拜他。”
MATT|2|9|他们听了王的话就去了。忽然，在东方所看到的那颗星在前面引领他们，一直行到小孩子所在地方的上方就停住了。
MATT|2|10|他们看见那星，就非常欢喜；
MATT|2|11|进了房子，看见小孩子和他母亲 马利亚 ，就俯伏拜那小孩子，揭开宝盒，拿出黄金、乳香、没药，作为礼物献给他。
MATT|2|12|因为在梦中得到主的指示，不要回去见 希律 ，他们就从别的路回自己的家乡去了。
MATT|2|13|他们走后，忽然主的使者在 约瑟 梦中向他显现，说：“起来！带着小孩子和他母亲逃往 埃及 ，住在那里，等我的指示；因为 希律 要搜寻那小孩子来杀害他。”
MATT|2|14|约瑟 就起来，连夜带着小孩子和他母亲往 埃及 去，
MATT|2|15|住在那里，直到 希律 死了。这是要应验主藉先知所说的话：“我从 埃及 召我的儿子出来。”
MATT|2|16|希律 见自己被博学之士愚弄，极其愤怒，差人将 伯利恒 城里和四境所有的男孩，根据他向博学之士仔细查问到的时间，凡两岁以内的，都杀尽了。
MATT|2|17|这就应验了 耶利米 先知所说的话：
MATT|2|18|“在 拉玛 听见号啕大哭的声音， 是 拉结 哭她儿女； 她不肯受安慰， 因为他们都不在了。”
MATT|2|19|希律 死了以后，在 埃及 ，忽然主的使者在 约瑟 梦中向他显现，
MATT|2|20|说：“起来，带着小孩子和他母亲回 以色列 地去！因为要杀害这小孩子的人已经死了。”
MATT|2|21|约瑟 就起来，带着小孩子和他母亲进入 以色列 地去。
MATT|2|22|但是他因听见 亚基老 继承他父亲 希律 作了 犹太 王，怕到那里去；又在梦中得到主的指示，就往 加利利 境内去了。
MATT|2|23|他们到了一座城，名叫 拿撒勒 ，就住在那里。这是要应验先知所说的话：“他将称为 拿撒勒 人。”
MATT|3|1|在那些日子，施洗的 约翰 出来，在 犹太 的旷野宣讲：
MATT|3|2|“你们要悔改！因为天国近了。”
MATT|3|3|这人就是 以赛亚 先知所说的： “在旷野有声音呼喊着： 预备主的道， 修直他的路。”
MATT|3|4|这 约翰 身穿骆驼毛的衣服，腰束皮带，吃的是蝗虫和野蜜。
MATT|3|5|那时， 耶路撒冷 、全 犹太 和全 约旦河 地区的人，都到 约翰 那里去，
MATT|3|6|承认他们的罪，在 约旦河 里受他的洗。
MATT|3|7|约翰 看见许多法利赛人和撒都该人也来受洗，就对他们说：“毒蛇的孽种啊，谁指示你们逃避那将要来的愤怒呢？
MATT|3|8|你们要结出果子来，和悔改的心相称。
MATT|3|9|不要自己心里说：‘我们有 亚伯拉罕 为祖宗。’我告诉你们，上帝能从这些石头中给 亚伯拉罕 兴起子孙来。
MATT|3|10|现在斧子已经放在树根上，凡不结好果子的树就砍下来，丢在火里。
MATT|3|11|我是用水给你们施洗，叫你们悔改；但那在我以后来的，能力比我更大，我就是给他提鞋子也不配，他要用圣灵与火给你们施洗。
MATT|3|12|他手里拿着簸箕，要扬净他的谷物，把麦子收在仓里，把糠用不灭的火烧尽。”
MATT|3|13|当时，耶稣从 加利利 来到 约旦河 ，到了 约翰 那里，请 约翰 为他施洗。
MATT|3|14|约翰 想要阻止他，说：“我应该受你的洗，你怎么到我这里来呢？”
MATT|3|15|耶稣回答他：“暂且这样做吧，因为我们理当这样履行全部的义 。”于是 约翰 就依了他。
MATT|3|16|耶稣受了洗，随即从水里上来。天忽然为他 开了，他看见上帝的灵降下，仿佛鸽子落在他身上。
MATT|3|17|这时，天上有声音说：“这是我的爱子，我所喜爱的。”
MATT|4|1|当时，耶稣被圣灵引到旷野，受魔鬼的试探。
MATT|4|2|他禁食四十昼夜，后来就饿了。
MATT|4|3|那试探者进前来对他说：“你若是上帝的儿子，叫这些石头变成食物吧。”
MATT|4|4|耶稣却回答说：“经上记着： ‘人活着，不是单靠食物， 乃是靠上帝口里所出的一切话。’”
MATT|4|5|魔鬼就带他进了圣城，叫他站在圣殿顶上，
MATT|4|6|对他说：“你若是上帝的儿子，就跳下去！因为经上记着： ‘主要为你命令他的使者， 用手托住你， 免得你的脚碰在石头上。’”
MATT|4|7|耶稣对他说：“经上又记着：‘不可试探主—你的上帝。’”
MATT|4|8|魔鬼又带他上了一座很高的山，将世上的万国和万国的荣华都指给他看，
MATT|4|9|对他说：“你若俯伏拜我，我就把这一切赐给你。”
MATT|4|10|耶稣说：“撒但 ，退去！因为经上记着： ‘要拜主—你的上帝， 惟独事奉他。’”
MATT|4|11|于是，魔鬼离开了耶稣，立刻有天使来伺候他。
MATT|4|12|耶稣听见 约翰 下了监，就退到 加利利 去；
MATT|4|13|后来离开 拿撒勒 ，往 迦百农 去，住在那里。那地方靠海，在 西布伦 和 拿弗他利 地区。
MATT|4|14|这是要应验 以赛亚 先知所说的话：
MATT|4|15|“ 西布伦 ， 拿弗他利 ， 沿海的路， 约旦河 的东边， 外邦人的 加利利 —
MATT|4|16|那坐在黑暗里的百姓 看见了大光； 坐在死荫之地的人 有光照耀他们。”
MATT|4|17|从那时候，耶稣开始宣讲，说：“你们要悔改！因为天国近了。”
MATT|4|18|耶稣沿着 加利利 海边行走，看见两兄弟，就是那叫 彼得 的 西门 和他弟弟 安得烈 ，正往海里撒网；他们本是打鱼的。
MATT|4|19|耶稣对他们说：“来跟从我，我要叫你们得人如得鱼一样。”
MATT|4|20|他们立刻舍了网，跟从他。
MATT|4|21|耶稣从那里往前走，看见另外两兄弟，就是 西庇太 的儿子 雅各 和他弟弟 约翰 ，同他们的父亲 西庇太 在船上补网，耶稣就呼召他们。
MATT|4|22|他们立刻舍了船，辞别父亲，跟从了耶稣。
MATT|4|23|耶稣走遍 加利利 ，在各会堂里教导人，宣讲天国的福音，医治百姓各样的疾病。
MATT|4|24|他的名声传遍了 叙利亚 。那里的人把一切病人，就是有各样疾病和疼痛的、被鬼附的、癫痫的、瘫痪的，都带了来，耶稣就治好了他们。
MATT|4|25|当时，有一大群人从 加利利 、 低加坡里 、 耶路撒冷 、 犹太 、 约旦河 的东边，来跟从他。
MATT|5|1|耶稣看见这一群人，就上了山，坐下后，门徒到他跟前来，
MATT|5|2|他开口教导他们说：
MATT|5|3|“心灵贫穷的人有福了！ 因为天国是他们的。
MATT|5|4|哀恸的人有福了！ 因为他们必得安慰。
MATT|5|5|谦和的人有福了！ 因为他们必承受土地。
MATT|5|6|饥渴慕义的人有福了！ 因为他们必得饱足。
MATT|5|7|怜悯人的人有福了！ 因为他们必蒙怜悯。
MATT|5|8|清心的人有福了！ 因为他们必得见上帝。
MATT|5|9|缔造和平的人有福了！ 因为他们必称为上帝的儿子。
MATT|5|10|为义受迫害的人有福了！ 因为天国是他们的。
MATT|5|11|“人若因我辱骂你们，迫害你们，捏造各样坏话毁谤你们 ，你们就有福了！
MATT|5|12|要欢喜快乐，因为你们在天上的赏赐是很多的。在你们以前的先知，人也是这样迫害他们。”
MATT|5|13|“你们是地上的盐。盐若失了味，怎能叫它再咸呢？它不再有用，只好被丢在外面，任人践踏。
MATT|5|14|你们是世上的光。城造在山上是不能隐藏的。
MATT|5|15|人点灯，不放在斗底下，而是放在灯台上，就照亮一家的人。
MATT|5|16|你们的光也要这样照在人前，叫他们看见你们的好行为，把荣耀归给你们在天上的父。”
MATT|5|17|“不要以为我来是要废掉律法和先知。我来不是要废掉，而是要成全。
MATT|5|18|我实在告诉你们，就是到天地都废去，律法的一点一画也不能废去，直到一切都实现。
MATT|5|19|所以，无论谁废掉这诫命中最小的一条，又教导人也这样做，他在天国里要称为最小的。但无论谁遵行并如此教导人的，他在天国里要称为大。
MATT|5|20|我告诉你们，你们的义若不胜过文士和法利赛人的义，绝不能进天国。”
MATT|5|21|“你们听过有对古人说：‘不可杀人’；‘凡杀人的，必须受审判。’
MATT|5|22|但是我告诉你们：凡向弟兄动怒的，必须受审判；凡骂弟兄是废物的，必须受议会的审判；凡骂弟兄是白痴的，必须遭受地狱的火。
MATT|5|23|所以，你在祭坛上献祭物的时候，若想起有弟兄对你怀恨，
MATT|5|24|就要把祭物留在坛前，先去跟弟兄和好，然后来献祭物。
MATT|5|25|你同告你的冤家还在路上，就要赶快与他讲和，免得他把你送交给法官，法官交给警卫，你就下在监里了。
MATT|5|26|我实在告诉你，就是有一个大文钱 还没有还清，你也绝不能从那里出来。”
MATT|5|27|“你们听过有话说：‘不可奸淫。’
MATT|5|28|但是我告诉你们：凡看见妇女就动淫念的，这人心里已经与她犯奸淫了。
MATT|5|29|若是你的右眼使你跌倒，就把它挖出来，丢掉。宁可失去身体中的一部分，也不让整个身体被扔进地狱。
MATT|5|30|若是你的右手使你跌倒，就把它砍下来，丢掉。宁可失去身体中的一部分，也不让整个身体下地狱。”
MATT|5|31|“又有话说：‘无论谁休妻，都要给她休书。’
MATT|5|32|但是我告诉你们：凡休妻的，除非是因不贞的缘故，否则就是使她犯奸淫了；人若娶被休的妇人，也是犯奸淫了。”
MATT|5|33|“你们又听过有对古人说：‘不可背誓，所起的誓总要向主谨守。’
MATT|5|34|但是我告诉你们：什么誓都不可起。不可指着天起誓，因为天是上帝的宝座。
MATT|5|35|不可指着地起誓，因为地是他的脚凳；也不可指着 耶路撒冷 起誓，因为 耶路撒冷 是大君王的京城。
MATT|5|36|又不可指着你的头起誓，因为你不能使一根头发变黑变白。
MATT|5|37|你们的话，是，就说是；不是，就说不是。若再多说，就是出于那恶者。”
MATT|5|38|“你们听过有话说：‘以眼还眼，以牙还牙。’
MATT|5|39|但是我告诉你们：不要与恶人作对。有人打你的右脸，连另一边也转过去由他打。
MATT|5|40|有人想要告你，要拿你的里衣，连外衣也由他拿去。
MATT|5|41|有人强迫你走一里 路，你就跟他走二里。
MATT|5|42|有求你的，就给他；有向你借贷的，不可推辞。”
MATT|5|43|“你们听过有话说：‘要爱你的邻舍，恨你的仇敌。’
MATT|5|44|但是我告诉你们：要爱你们的仇敌，为那迫害你们的祷告。
MATT|5|45|这样，你们就可以作天父的儿女了。因为他叫太阳照好人，也照坏人；降雨给义人，也给不义的人。
MATT|5|46|你们若只爱那爱你们的人，有什么赏赐呢？就是税吏不也是这样做吗？
MATT|5|47|你们若只请你弟兄的安，有什么比别人强呢？就是外邦人不也是这样做吗？
MATT|5|48|所以，你们要完全，如同你们的天父是完全的。”
MATT|6|1|“你们要谨慎，不可故意在人面前表现虔诚，叫他们看见，若是这样，就不能得你们天父的赏赐了。
MATT|6|2|“所以，你施舍的时候，不可叫人在你前面吹号，像那假冒为善的人在会堂里和街道上所做的，故意要得人的称赞。我实在告诉你们，他们已经得了他们的赏赐。
MATT|6|3|你施舍的时候，不要让左手知道右手所做的，
MATT|6|4|好使你隐秘地施舍；你父在隐秘中察看，必然赏赐你。”
MATT|6|5|“你们祷告的时候，不可像那假冒为善的人，爱站在会堂里和十字路口祷告，故意让人看见。我实在告诉你们，他们已经得了他们的赏赐。
MATT|6|6|你祷告的时候，要进入内室，关上门，向那在隐秘中的父祷告；你父在隐秘中察看，必将赏赐你。
MATT|6|7|你们祷告，不可像外邦人那样重复一些空话，他们以为话多了必蒙垂听。
MATT|6|8|你们不可效法他们。因为在你们祈求以前，你们所需要的，你们的父早已知道了。”
MATT|6|9|“所以，你们要这样祷告： ‘我们在天上的父： 愿人都尊你的名为圣。
MATT|6|10|愿你的国降临； 愿你的旨意行在地上， 如同行在天上。
MATT|6|11|我们日用的饮食，今日赐给我们。
MATT|6|12|免我们的债， 如同我们免了人的债。
MATT|6|13|不叫我们陷入试探； 救我们脱离那恶者。 因为国度、权柄、荣耀，全是你的， 直到永远。阿们！ ’
MATT|6|14|“你们若饶恕人的过犯，你们的天父也必饶恕你们；
MATT|6|15|你们若不饶恕人 ，你们的天父也必不饶恕你们的过犯。”
MATT|6|16|“你们禁食的时候，不可像那假冒为善的人，脸上带着愁容；因为他们蓬头垢面，故意让人看出他们在禁食。我实在告诉你们，他们已经得了他们的赏赐。
MATT|6|17|你禁食的时候，要梳头洗脸，
MATT|6|18|不要让人看出你在禁食，只让你隐秘中的父看见；你父在隐秘中察看，必然赏赐你。”
MATT|6|19|“不要为自己在地上积蓄财宝；地上有虫子咬，能锈坏，也有贼挖洞来偷。
MATT|6|20|要在天上积蓄财宝；天上没有虫子咬，不会锈坏，也没有贼挖洞来偷。
MATT|6|21|因为你的财宝在哪里，你的心也在哪里。”
MATT|6|22|“眼睛是身体的灯。你的眼睛若明亮，全身就光明；
MATT|6|23|你的眼睛若昏花，全身就黑暗。你里面的光若黑暗了，那黑暗是何等大呢！”
MATT|6|24|“一个人不能服侍两个主；他不是恨这个爱那个，就是重这个轻那个。你们不能又服侍上帝，又服侍 玛门 。”
MATT|6|25|“所以，我告诉你们，不要为你们的生命忧虑吃什么喝什么 ，或为你们的身体忧虑穿什么。生命不胜于饮食吗？身体不胜于衣裳吗？
MATT|6|26|你们看一看那天上的飞鸟，也不种也不收，也不在仓里存粮，你们的天父尚且养活它们。你们不比飞鸟贵重得多吗？
MATT|6|27|你们哪一个能藉着忧虑使寿数多加一刻呢 ？
MATT|6|28|何必为衣裳忧虑呢？你们想一想野地里的百合花是怎么长起来的：它也不劳动也不纺线。
MATT|6|29|然而我告诉你们，就是 所罗门 极荣华的时候，他所穿戴的还不如这些花的一朵呢！
MATT|6|30|你们这小信的人哪！野地里的草今天还在，明天就丢在炉里，上帝还给它这样的妆饰，何况你们呢？
MATT|6|31|所以，不要忧虑，说：‘我们吃什么？喝什么？穿什么？’
MATT|6|32|这都是外邦人所求的。你们需要这一切东西，你们的天父都知道。
MATT|6|33|你们要先求上帝的国和他的义，这些东西都要加给你们了。
MATT|6|34|所以，不要为明天忧虑，因为明天自有明天的忧虑；一天的难处一天当就够了。”
MATT|7|1|“你们不要评断别人，免得你们被审判。
MATT|7|2|因为你们怎样评断别人，也必怎样被审判；你们用什么量器量给人，也必用什么量器量给你们。
MATT|7|3|为什么看见你弟兄眼中有刺，却不想自己眼中有梁木呢？
MATT|7|4|你自己眼中有梁木，怎能对你弟兄说‘让我去掉你眼中的刺’呢？
MATT|7|5|你这假冒为善的人！先去掉自己眼中的梁木，然后才能看得清楚，好去掉你弟兄眼中的刺。
MATT|7|6|不要把圣物给狗，也不要把你们的珍珠丢在猪面前，恐怕它们践踏了珍珠，转过来咬你们。”
MATT|7|7|“你们祈求，就给你们；寻找，就找到；叩门，就给你们开门。
MATT|7|8|因为凡祈求的，就得着；寻找的，就找到；叩门的，就给他开门。
MATT|7|9|你们中间谁有儿子求饼，反给他石头呢？
MATT|7|10|求鱼，反给他蛇呢？
MATT|7|11|你们虽然不好，尚且知道拿好东西给儿女，何况你们在天上的父，他岂不更要把好东西赐给求他的人吗？
MATT|7|12|所以，无论何事，你们想要人怎样待你们，你们也要怎样待人，因为这就是律法和先知的道理。”
MATT|7|13|“你们要进窄门。因为通往灭亡的门是宽的，路是大的，进去的人也多；
MATT|7|14|通往生命的门是窄的，路是小的，找到的人也少。”
MATT|7|15|“你们要防备假先知。他们到你们这里来，外面披着羊皮，里面却是残暴的狼。
MATT|7|16|岂能在荆棘上摘葡萄呢？岂能在蒺藜里摘无花果呢？凭着他们的果子，就可以认出他们来。
MATT|7|17|这样，凡好树都结好果子，而坏树结坏果子。
MATT|7|18|好树不能结坏果子，坏树也不能结好果子。
MATT|7|19|凡不结好果子的树就砍下来，丢在火里。
MATT|7|20|所以，凭着他们的果子就可以认出他们来。”
MATT|7|21|“不是每一个称呼我‘主啊，主啊’的人都能进天国；惟有遵行我天父旨意的人才能进去。
MATT|7|22|在那日必有许多人对我说：‘主啊，主啊，我们不是奉你的名传道，奉你的名赶鬼，奉你的名行许多异能吗？’
MATT|7|23|我要向他们宣告：‘我从来不认识你们，你们这些作恶的人，给我走开！’”
MATT|7|24|“所以，凡听了我这些话又去做的，好比一个聪明人把房子盖在磐石上。
MATT|7|25|风吹，雨打，水冲，撞击那房子，房子总不倒塌，因为根基立在磐石上。
MATT|7|26|凡听了我这些话而不去做的，好比一个无知的人把房子盖在沙土上。
MATT|7|27|风吹，雨打，水冲，撞击那房子，房子就倒塌了，并且倒塌得很厉害。”
MATT|7|28|耶稣讲完了这些话，众人对他的教导都感到惊奇，
MATT|7|29|因为他教导他们正像有权柄的人，不像他们的文士。
MATT|8|1|耶稣下了山，有一大群人跟着他。
MATT|8|2|这时，一个痲疯病人前来拜他，说：“主啊，你若肯，你能使我洁净。”
MATT|8|3|耶稣伸手摸他，说：“我肯，你洁净了吧！”他的痲疯病立刻就洁净了。
MATT|8|4|耶稣对他说：“你要注意，不可告诉任何人，只要去，让祭司为你检查，并献上 摩西 所吩咐的祭物，作为证据给众人看。”
MATT|8|5|耶稣进了 迦百农 ，有一个百夫长进前来，求他，
MATT|8|6|说：“主啊，我的僮仆瘫痪了，躺在家里，非常痛苦。”
MATT|8|7|耶稣说：“我去医治他。”
MATT|8|8|百夫长回答：“主啊，你到舍下来，我不敢当；只要你说一句话，我的僮仆就会痊愈。
MATT|8|9|因为我在人的权下，也有兵在我以下。我对这个说：‘去！’他就去；对那个说：‘来！’他就来；对我的仆人说：‘做这事！’他就去做。”
MATT|8|10|耶稣听了就很惊讶，对跟从的人说：“我实在告诉你们，这么大的信心，就是在 以色列 ，我也没有见过。
MATT|8|11|我又告诉你们，从东从西，将有许多人来，在天国里与 亚伯拉罕 、 以撒 、 雅各 一同坐席；
MATT|8|12|本国的子民反而被赶到外边黑暗里去，在那里要哀哭切齿了。”
MATT|8|13|耶稣对百夫长说：“你回去吧！照你的信心成全你了。”就在那时，他的僮仆好了。
MATT|8|14|耶稣到了 彼得 家里，见 彼得 的岳母正发烧躺着。
MATT|8|15|耶稣一摸她的手，烧就退了，于是她起来服事耶稣。
MATT|8|16|傍晚的时候，有人带着许多被鬼附的来到耶稣跟前，他只用一句话就把邪灵都赶出去，并且治好了一切有病的人。
MATT|8|17|这是要应验 以赛亚 先知所说的话： “他代替了我们的软弱， 担当了我们的疾病。”
MATT|8|18|耶稣见许多人围着他，就吩咐渡到对岸去。
MATT|8|19|有一个文士进前来对他说：“老师，你无论往哪里去，我都要跟从你。”
MATT|8|20|耶稣说：“狐狸有洞，天空的飞鸟有窝，人子却没有枕头的地方。”
MATT|8|21|又有一个门徒对耶稣说：“主啊，容许我先回去埋葬我的父亲。”
MATT|8|22|耶稣说：“让死人埋葬他们的死人。你跟从我吧！”
MATT|8|23|耶稣上了船，门徒跟着他。
MATT|8|24|海里忽然起了猛烈的风暴，以致船几乎被波浪淹没，耶稣却睡着了。
MATT|8|25|门徒去叫醒他，说：“主啊，救命啊，我们快没命啦！”
MATT|8|26|耶稣说：“你们这些小信的人哪，为什么胆怯呢？”于是他起来，斥责风和海，风和海就大大平静了。
MATT|8|27|众人惊讶地说：“这是怎样的一个人？连风和海都听从他。”
MATT|8|28|耶稣渡到对岸去，到 加大拉 人 的地区，有两个被鬼附的人从坟墓迎着他走来。他们极其凶猛，甚至没有人敢从那条路经过。
MATT|8|29|他们喊着说：“上帝的儿子，你为什么干扰我们？时候还没有到，你就上这里来叫我们受苦吗？”
MATT|8|30|离他们很远，有一大群猪正在吃食。
MATT|8|31|鬼就央求耶稣，说：“若要把我们赶出去，就打发我们进入猪群吧！”
MATT|8|32|耶稣对他们说：“去吧！”鬼就出来，进入猪群。一转眼，整群猪都闯下山崖，投进海里，淹死了。
MATT|8|33|放猪的就逃进城去，把这一切事和被鬼附的人所遭遇的都告诉众人。
MATT|8|34|全城的人都出来迎见耶稣，见了他以后，就央求他离开他们的地区。
MATT|9|1|耶稣上了船，渡过海，来到自己的城里。
MATT|9|2|有人用褥子抬着一个瘫子到耶稣跟前来。耶稣见他们的信心，就对瘫子说：“孩子，放心吧，你的罪赦了。”
MATT|9|3|这时，有几个文士心里说：“这个人说亵渎的话了。”
MATT|9|4|耶稣知道他们的心思，就说：“你们心里为什么怀着恶念呢？
MATT|9|5|说‘你的罪赦了’，或说‘你起来行走’，哪一样容易呢？
MATT|9|6|但要让你们知道，人子在地上有赦罪的权柄”，于是对瘫子说：“起来！拿你的褥子回家去吧。”
MATT|9|7|那人就起来，回家去了。
MATT|9|8|众人看见都畏惧，归荣耀给上帝，因为他把这样的权柄赐给人。
MATT|9|9|耶稣从那里往前走，看见一个人名叫 马太 ，在税关坐着，就对他说：“来跟从我！”他就起来跟从耶稣。
MATT|9|10|耶稣在屋里坐席的时候，有好些税吏和罪人来，与耶稣和他的门徒一同坐席。
MATT|9|11|法利赛人看见，就对耶稣的门徒说：“你们的老师为什么与税吏和罪人一同吃饭呢？”
MATT|9|12|耶稣听见，就说：“健康的人用不着医生；有病的人才用得着。
MATT|9|13|经上说：‘我喜爱怜悯，不喜爱祭祀。’这句话的意思，你们去揣摩。我不是来召义人，而是召罪人。”
MATT|9|14|那时， 约翰 的门徒来见耶稣，说：“我们和法利赛人常常 禁食，你的门徒却不禁食，这是为什么呢？”
MATT|9|15|耶稣对他们说：“新郎和宾客在一起的时候，宾客怎么能哀恸呢？但日子将到，新郎要被带走，那时候他们就要禁食了。
MATT|9|16|没有人把新布补在旧衣服上；因为所补上的会撕破那衣服，裂口就更大了。
MATT|9|17|也没有人把新酒装在旧皮袋里，若是这样，皮袋会胀破，酒就漏出来，皮袋也糟蹋了。相反地，把新酒装在新皮袋里，两样就都保全了。”
MATT|9|18|耶稣说这些话的时候，有一个会堂主管来，向他下跪，说：“我女儿刚死了，求你去按手在她身上，她就会活过来。”
MATT|9|19|耶稣就起来跟他去；门徒也跟了去。
MATT|9|20|这时，有一个女人，患了经血不止的病有十二年，来到耶稣背后，摸他的衣裳繸子；
MATT|9|21|因为她心里说：“我只要摸他的衣裳，就会痊愈。”
MATT|9|22|耶稣转过来，看见她，就说：“女儿，放心！你的信救了你。”从那时起，这女人就痊愈了。
MATT|9|23|耶稣到了会堂主管的家里，看见吹鼓手和乱哄哄的一群人，
MATT|9|24|就说：“退去吧！这女孩不是死了，而是睡着了。”他们就嘲笑他。
MATT|9|25|众人被赶出后，耶稣就进去，拉着女孩的手，女孩就起来了。
MATT|9|26|于是这消息传遍了那地方。
MATT|9|27|耶稣从那里往前走，有两个盲人跟着他，喊叫说：“ 大卫 之子，可怜我们吧！”
MATT|9|28|耶稣进了屋子，盲人就来到他跟前。耶稣说：“你们信我能做这事吗？”他们说：“主啊，我们信。”
MATT|9|29|耶稣就摸他们的眼睛，说：“照着你们的信心成全你们吧。”
MATT|9|30|他们的眼睛就开了。耶稣严严地叮嘱他们说：“要小心，不可让人知道。”
MATT|9|31|他们出去，竟把他的名声传遍了那地方。
MATT|9|32|他们出去的时候，有人把一个被鬼附的哑巴带到耶稣跟前来。
MATT|9|33|鬼被赶出去，哑巴就说出话来。众人都很惊讶，说：“在 以色列 ，从来没有见过这样的事。”
MATT|9|34|法利赛人却说：“他是靠着鬼王赶鬼的。”
MATT|9|35|耶稣走遍各城各乡，在他们的会堂里教导人，宣讲天国的福音，又医治各样的病症。
MATT|9|36|他看见一大群人，就怜悯他们；因为他们困苦无助，如同羊没有牧人一样。
MATT|9|37|于是他对门徒说：“要收的庄稼多，做工的人少。
MATT|9|38|所以，你们要求庄稼的主差遣做工的人出去收他的庄稼。”
MATT|10|1|耶稣叫了十二个门徒来，给他们权柄，能驱赶污灵和医治各样的疾病。
MATT|10|2|这十二使徒的名字如下：头一个叫 西门 （又称 彼得 ），还有他弟弟 安得烈 ， 西庇太 的儿子 雅各 和 雅各 的弟弟 约翰 ，
MATT|10|3|腓力 和 巴多罗买 ， 多马 和税吏 马太 ， 亚勒腓 的儿子 雅各 ，和 达太 ，
MATT|10|4|激进党的 西门 ，还有出卖耶稣的 加略 人 犹大 。
MATT|10|5|耶稣差遣这十二个人出去，吩咐他们说：“外邦人的路，你们不要走； 撒玛利亚 人的城，你们不要进；
MATT|10|6|宁可往 以色列 家迷失的羊那里去。
MATT|10|7|要边走边传，说‘天国近了’。
MATT|10|8|要医治病人，使死人复活，使痲疯病人洁净，把鬼赶出去。你们白白地得来，也要白白地给人。
MATT|10|9|腰袋里不要带金银铜钱；
MATT|10|10|途中不要带行囊，不要带两件内衣，也不要带鞋子和手杖，因为工人得饮食是应当的。
MATT|10|11|你们无论进哪一城、哪一村，要打听那里谁是合适的人，就住在他家，直住到离开的时候。
MATT|10|12|进他家时，要向那家请安。
MATT|10|13|那家若配得平安，你们所求的平安就临到那家；若不配得，你们所求的平安仍归你们。
MATT|10|14|凡不接待你们，不听你们话的人，你们离开那家，或是那城的时候，要跺掉你们脚上的尘土。
MATT|10|15|我实在告诉你们，在审判的日子， 所多玛 和 蛾摩拉 地方所受的，比那城还容易受呢！”
MATT|10|16|“看哪！我差你们出去，如同羊进入狼群，所以你们要机警如蛇，纯真如鸽。
MATT|10|17|你们要防备那些人，因为他们要把你们交给议会，也要在会堂里鞭打你们。
MATT|10|18|你们要为我的缘故被送到统治者和君王面前，对他们和外邦人作见证。
MATT|10|19|当人把你们交出时，不要担心怎样说话，或说什么话。到那时候，必赐给你们该说的话，
MATT|10|20|因为不是你们自己说的，而是你们父的灵在你们里面说的。
MATT|10|21|兄弟要把兄弟、父亲要把儿女置于死地；儿女要起来与父母为敌，害死他们。
MATT|10|22|而且你们要为我的名被众人憎恨。但坚忍到底的终必得救。
MATT|10|23|有人在这城迫害你们，就逃到另一城去。 我实在告诉你们， 以色列 的城镇，你们还没有走遍，人子就要来临。
MATT|10|24|“学生不高过老师，仆人不高过主人。
MATT|10|25|学生所遭遇的与老师一样，仆人所遭遇的与主人一样，也就够了。既然有人骂一家的主人是‘ 别西卜 ’ ，更何况他的家人呢？”
MATT|10|26|“所以，不要怕他们，因为掩盖的事没有不显露出来的，隐藏的事也没有不被知道的。
MATT|10|27|我在暗中告诉你们的，你们要在明处说出来；你们耳中所听的，要在屋顶上宣扬出来。
MATT|10|28|那杀人身体但不能灭人灵魂的，不要怕他们；惟有那能在地狱里毁灭身体和灵魂的，才要怕他。
MATT|10|29|两只麻雀不是卖一铜钱 吗？你们的父若不许，一只也不会掉在地上。
MATT|10|30|就是你们的头发也都数过了。
MATT|10|31|所以，不要惧怕，你们比许多的麻雀还贵重！”
MATT|10|32|“所以，凡在人面前认我的，我在我天上的父面前也必认他；
MATT|10|33|凡在人面前不认我的，我在我天上的父面前也必不认他。”
MATT|10|34|“你们不要以为我来是带给地上和平，我来并不是带来和平，而是刀剑。
MATT|10|35|因为我来是要叫 ‘人与父亲对立， 女儿与母亲对立， 媳妇与婆婆对立。
MATT|10|36|人的仇敌就是自己家里的人。’
MATT|10|37|爱父母胜过爱我的，不配作我的门徒；爱儿女胜过爱我的，不配作我的门徒。
MATT|10|38|不背自己的十字架跟从我的，不配作我的门徒。
MATT|10|39|得着性命的，要丧失性命；为我丧失性命的，要得着性命。”
MATT|10|40|“接纳你们的就是接纳我；接纳我的就是接纳差遣我来的那位。
MATT|10|41|把先知当作先知接纳的，必得先知的赏赐；把义人当作义人接纳的，必得义人的赏赐。
MATT|10|42|无论谁，只因门徒的名，就算把一杯凉水给这些小子中的一个喝，我实在告诉你们，他一定会得到赏赐。”
MATT|11|1|耶稣吩咐完了十二个门徒，就离开那里，往各城去传道，教导人。
MATT|11|2|约翰 在监狱里听见基督所做的事，就派他的门徒去，
MATT|11|3|问耶稣：“将要来的那位就是你吗？还是我们要等候另一位呢？”
MATT|11|4|耶稣回答他们：“你们去，把所听见、所看见的告诉 约翰 ：
MATT|11|5|就是盲人看见，瘸子行走，痲疯病人得洁净，聋子听见，死人复活，穷人听到福音。
MATT|11|6|凡不因我跌倒的有福了！”
MATT|11|7|他们一走，耶稣就对众人谈到 约翰 ，说：“你们从前到旷野去，是要看什么呢？看风吹动的芦苇吗？
MATT|11|8|你们出去到底是要看什么？看穿细软衣服的人吗？那穿细软衣服的人是在王宫里。
MATT|11|9|你们出去究竟是要看什么？是先知吗？是的，我告诉你们，他比先知大多了。
MATT|11|10|这个人就是经上所说的： ‘看哪，我要差遣我的使者在你面前， 他要在你前面为你预备道路。’
MATT|11|11|我实在告诉你们，凡女子所生的，没有一个比施洗 约翰 大；但在天国里，最小的比他还大。
MATT|11|12|从施洗 约翰 的日子到今天，天国受到强烈的攻击，强者夺取它 。
MATT|11|13|众先知和律法，直到 约翰 为止，都说了预言。
MATT|11|14|如果你们愿意接受，这人就是那要来的 以利亚 。
MATT|11|15|有耳的，就应当听！
MATT|11|16|“我该用什么来比这世代呢？这正像孩童坐在街市上向同伴呼喊：
MATT|11|17|‘我们为你们吹笛，你们不跳舞； 我们唱哀歌，你们不捶胸。’
MATT|11|18|约翰 来了，既不吃也不喝，人们就说他是被鬼附的；
MATT|11|19|人子来了，也吃也喝，他们又说这人贪食好酒，是税吏和罪人的朋友。而智慧是由它的果子来证实的 。”
MATT|11|20|那时，耶稣在一些城行了许多异能。因为城里的人不肯悔改，他就责备那些城说：
MATT|11|21|“ 哥拉汛 哪，你有祸了！ 伯赛大 啊，你有祸了！因为在你们中间所行的异能若行在 推罗 、 西顿 ，他们早已披麻蒙灰悔改了。
MATT|11|22|但我告诉你们，在审判的日子， 推罗 和 西顿 所受的，比你们还容易受呢！
MATT|11|23|迦百农 啊， 你以为要被举到天上吗？ 你要被推下阴间！ 因为在你那里所行的异能，若行在 所多玛 ，它还可以存留到今日。
MATT|11|24|但我告诉你们，在审判的日子， 所多玛 地方所受的，比你们还容易受呢！”
MATT|11|25|那时，耶稣说：“父啊，天地的主，我感谢你！因为你把这些事向聪明智慧的人隐藏起来，而向婴孩启示出来。
MATT|11|26|父啊，是的，因为你的美意本是如此。
MATT|11|27|一切都是我父交给我的；除了父，没有人知道子；除了子和子所愿意启示的人，没有人知道父。
MATT|11|28|凡劳苦担重担的人都到我这里来，我要使你们得安息。
MATT|11|29|我心里柔和谦卑，你们当负我的轭，向我学习；这样，你们的心灵就必得安息。
MATT|11|30|因为我的轭是容易的，我的担子是轻省的。”
MATT|12|1|那时，耶稣在安息日从麦田经过。他的门徒饿了，就摘麦穗来吃。
MATT|12|2|法利赛人看见，对耶稣说：“看哪，你的门徒在安息日做不合法的事了。”
MATT|12|3|耶稣对他们说：“ 大卫 和跟从他的人饥饿时所做的事，你们没有念过吗？
MATT|12|4|他怎么进了上帝的居所，吃了供饼呢？这饼是他和跟从他的人不可以吃的，惟独祭司才可以吃。
MATT|12|5|再者，律法上所记的，在安息日，祭司在圣殿里犯了安息日也不算有罪，你们没有念过吗？
MATT|12|6|但我告诉你们，比圣殿更大的在这里。
MATT|12|7|‘我喜爱怜悯，不喜爱祭祀。’你们若明白这话的意思，就不将无罪的当作有罪了。
MATT|12|8|因为人子是安息日的主。”
MATT|12|9|耶稣离开那地方，进了 犹太 人的会堂；
MATT|12|10|那里有个一只手萎缩了的人。有人为了要控告耶稣，就问他：“安息日治病合不合法？”
MATT|12|11|耶稣对他们说：“你们中间谁有一只羊在安息日掉在坑里，不抓住它，把它拉上来呢？
MATT|12|12|人比羊贵重得多了！所以，在安息日做善事是合法的。”
MATT|12|13|于是对那人说：“伸出手来！”他把手一伸，手就复原了，和另一只一样。
MATT|12|14|法利赛人出去，商议怎样除掉耶稣。
MATT|12|15|耶稣知道了，就离开那里，有一大群人跟着他。他把所有的病人都治好了，
MATT|12|16|又嘱咐他们不要把他宣扬出去。
MATT|12|17|这是要应验 以赛亚 先知所说的话：
MATT|12|18|“看哪，我所拣选的仆人， 我所亲爱，心所喜悦的； 我要将我的灵赐给他， 他必将公理传给外邦。
MATT|12|19|他不争吵，不喧嚷， 街上也没有人听见他的声音。
MATT|12|20|压伤的芦苇，他不折断， 将残的灯火，他不吹灭， 直到他使公理得胜。
MATT|12|21|外邦人都要仰望他的名。”
MATT|12|22|当时，有人把一个被鬼附，又盲又哑的人带到耶稣那里，耶稣医治他，那哑巴就能说话，又能看见。
MATT|12|23|众人都惊奇，说：“这不是 大卫 之子吗？”
MATT|12|24|但法利赛人听见，就说：“这个人赶鬼，无非是靠着鬼王 别西卜 罢了。”
MATT|12|25|耶稣知道他们的心思，就对他们说：“一国自相纷争，必定荒芜；一城一家自相纷争，必立不住。
MATT|12|26|若撒但赶出撒但，就是自相纷争，他的国怎能立得住呢？
MATT|12|27|我若靠着 别西卜 赶鬼，你们的子弟赶鬼又靠着谁呢？这样，他们要作你们的判官。
MATT|12|28|我若靠着上帝的灵赶鬼，那么，上帝的国就已临到你们了。
MATT|12|29|人怎能进壮士家里抢夺他的东西呢？除非先绑住那壮士，否则无法抢夺他的家。
MATT|12|30|不跟我一起的，就是反对我；不与我一起收聚的，就是在拆散。
MATT|12|31|所以我告诉你们，人一切的罪和亵渎的话都可得赦免，但是亵渎圣灵，总不得赦免。
MATT|12|32|凡说话干犯人子的，还可得赦免；但是说话干犯圣灵的，今世来世总不得赦免。”
MATT|12|33|“你们知道树好，果子也好；又知道树坏，果子也坏；因为看果子就可以知道树。
MATT|12|34|毒蛇的孽种啊，你们既是恶人，怎能说出好话来呢？因为心里所充满的，口里就说出来。
MATT|12|35|善人从他所存的善发出善来；恶人从他所存的恶发出恶来。
MATT|12|36|我告诉你们，凡是人所说的闲话，在审判的日子，要句句供出来；
MATT|12|37|因为要凭你的话定你为义，也要凭你的话定你有罪。”
MATT|12|38|当时，有几个文士和法利赛人对耶稣说：“老师，我们想请你显个神迹给我们看看。”
MATT|12|39|耶稣回答他们：“邪恶淫乱的世代求看神迹，除了先知 约拿 的神迹以外，再没有神迹给他们看了。
MATT|12|40|约拿 三日三夜在大鱼肚腹中，同样，人子也要三日三夜在地里面。
MATT|12|41|在审判的时候， 尼尼微 人要起来定这世代的罪，因为 尼尼微 人听了 约拿 所传的就悔改了。看哪，比 约拿 更大的在这里！
MATT|12|42|在审判的时候，南方的女王要起来定这世代的罪，因为她从地极而来，要听 所罗门 智慧的话。看哪，比 所罗门 更大的在这里！”
MATT|12|43|“污灵离了人身，走遍无水之地寻找安歇之处，却找不到。
MATT|12|44|于是他说：‘我要回到我原来的屋里去。’他到了，看见里面空着，打扫干净，修饰好了，
MATT|12|45|就去另带了七个比自己更恶的灵来，都进去住在那里。那人后来的景况比先前更坏了。这邪恶的世代也要如此。”
MATT|12|46|耶稣还在对众人说话的时候，不料，他母亲和他兄弟站在外边想要跟他说话。
MATT|12|47|有人告诉他：“看哪！你母亲和你兄弟站在外边，想要跟你说话。”
MATT|12|48|他却回答那对他说话的人，说：“谁是我的母亲？谁是我的兄弟？”
MATT|12|49|于是他伸手指着门徒，说：“看哪，我的母亲，我的兄弟！
MATT|12|50|凡遵行我天父旨意的人就是我的兄弟、姊妹和母亲。”
MATT|13|1|就在那天，耶稣从房子里出来，坐在海边。
MATT|13|2|有一大群人到他那里聚集，他只好上船坐下，众人都站在岸上。
MATT|13|3|他用比喻对他们讲了许多话。他说：“有一个撒种的出去撒种。
MATT|13|4|他撒的时候，有的落在路旁，飞鸟来把它们吃掉了。
MATT|13|5|有的落在土浅的石头地上，因为土不深，很快就长出苗来，
MATT|13|6|太阳出来一晒，因为没有根就枯干了。
MATT|13|7|有的落在荆棘里，荆棘长起来，把它挤住了。
MATT|13|8|又有的落在好土里，就结出果实，有一百倍的，有六十倍的，有三十倍的。
MATT|13|9|有耳的，就应当听！”
MATT|13|10|门徒进前来问耶稣：“对众人讲话，为什么用比喻呢？”
MATT|13|11|耶稣回答他们说：“因为天国的奥秘只让你们知道，不让他们知道。
MATT|13|12|凡有的，还要给他，让他有余；凡没有的，连他所有的也要夺去。
MATT|13|13|我之所以用比喻对他们讲，是因为 他们看却看不清， 听却听不见，也不明白。
MATT|13|14|在他们身上，正应验了 以赛亚 的预言： ‘你们听了又听，却不明白， 看了又看，却看不清。
MATT|13|15|因为这百姓的心麻木， 耳朵发沉， 眼睛闭着， 免得眼睛看见， 耳朵听见， 心里明白，回转过来， 我会医治他们。’
MATT|13|16|但你们的眼睛是有福的，因为看得见；你们的耳朵也是有福的，因为听得见。
MATT|13|17|我实在告诉你们，从前有许多先知和义人要看你们所看的，却没有看见；要听你们所听的，却没有听见。”
MATT|13|18|“所以，你们要听这撒种的比喻。
MATT|13|19|凡听见天国的道而不明白的，那恶者就来，把撒在他心里的夺了去；这就是撒在路旁的了。
MATT|13|20|撒在石头地上的，就是人听了道，立刻欢喜领受，
MATT|13|21|只因心里没有根，不过是暂时的，一旦为道遭受患难或迫害，立刻就跌倒。
MATT|13|22|撒在荆棘里的，就是人听了道，后来有世上的忧虑、钱财的迷惑把道挤住了，结不出果实。
MATT|13|23|撒在好土里的，就是人听了道，明白了，后来结了果实，有一百倍的，有六十倍的，有三十倍的。”
MATT|13|24|耶稣又设个比喻对他们说：“天国好比人撒好种在田里，
MATT|13|25|在人睡觉的时候，他的仇敌来，把杂草撒在麦子里就走了。
MATT|13|26|到长苗吐穗的时候，杂草也显出来。
MATT|13|27|地主的仆人进前来对他说：‘主人，你不是撒好种在田里吗？哪里来的杂草呢？’
MATT|13|28|主人回答他们：‘这是仇敌做的。’仆人对他说：‘你要我们去拔掉吗？’
MATT|13|29|主人说：‘不必，恐怕拔杂草，也把麦子连根拔出来。
MATT|13|30|让这两样一起长，等到收割。当收割的时候，我会对收割的人说，先把杂草拔出来，捆成捆，留着烧，把麦子收在我的仓里。’”
MATT|13|31|他又设个比喻对他们说：“天国好比一粒芥菜种，有人拿去种在田里。
MATT|13|32|它原比所有的种子都小，等到长起来，却比各样的菜都大，且成了树，以致天上的飞鸟来在它的枝上筑巢。”
MATT|13|33|他又对他们讲另一个比喻：“天国好比面酵，有妇人拿来放进三斗面里，直到全团都发起来。”
MATT|13|34|这都是耶稣用比喻对众人说的话，不用比喻，他就不对他们说什么。
MATT|13|35|这是要应验先知 所说的话： “我要开口说比喻， 说出从创世以来所隐藏的事。”
MATT|13|36|当时，耶稣离开众人，进了屋子。他的门徒进前来，说：“请把田间杂草的比喻讲给我们听。”
MATT|13|37|他回答：“那撒好种的就是人子，
MATT|13|38|田地就是世界，好种就是天国之子，杂草就是那恶者之子，
MATT|13|39|撒杂草的仇敌就是魔鬼，收割的时候就是世代的终结，收割的人就是天使。
MATT|13|40|正如把杂草拔出来用火焚烧，世代的终结也要如此。
MATT|13|41|人子要差遣他的使者，把一切使人跌倒的和作恶的从他国里挑出来，
MATT|13|42|丢在火炉里，在那里要哀哭切齿了。
MATT|13|43|那时，义人要在他们父的国里发出光来，像太阳一样。有耳的，就应当听！”
MATT|13|44|“天国好比宝贝藏在地里，人发现了就把它藏起来，欢欢喜喜地去变卖一切所有的，买这块地。
MATT|13|45|“天国又好比商人寻找好的珍珠，
MATT|13|46|发现一颗贵重的珍珠，就去变卖他一切所有的，买下这颗珍珠。”
MATT|13|47|“天国又好比网撒在海里，聚拢各种鱼类，
MATT|13|48|网一满，人们就把它拉上岸，坐下来，拣好的收在桶里，不好的丢掉。
MATT|13|49|世代的终结也要这样：天使要出来，把恶人从义人中分别出来，
MATT|13|50|丢在火炉里，在那里要哀哭切齿了。”
MATT|13|51|耶稣说：“这一切的话你们都明白了吗？”他们对他说：“明白了。”
MATT|13|52|他对他们说：“凡文士学习作天国的门徒，就像一个家的主人从他库里拿出新的和旧的东西来。”
MATT|13|53|耶稣说完了这些比喻，就离开那里，
MATT|13|54|来到自己的家乡，在会堂里教导人，以致他们都很惊奇，说：“这人哪来这样的智慧和异能呢？
MATT|13|55|这不是那木匠的儿子吗？他母亲不是叫 马利亚 吗？他兄弟们不是叫 雅各 、 约瑟 、 西门 、 犹大 吗？
MATT|13|56|他姊妹们不是都在我们这里吗？他这一切是从哪里来的呢？”
MATT|13|57|他们就厌弃他。耶稣对他们说：“先知除了在本乡和自己的家之外，没有不被尊敬的。”
MATT|13|58|耶稣因为他们不信，没有在那里行很多异能。
MATT|14|1|那时， 希律 分封王听见耶稣的名声，
MATT|14|2|就对臣仆说：“这是施洗的 约翰 从死人中复活，因此才有这些异能在他里面运行。”
MATT|14|3|原来， 希律 为他兄弟 腓力 的妻子 希罗底 的缘故，把 约翰 抓住绑了，关进监狱，
MATT|14|4|因为 约翰 曾对他说：“你占有这妇人是不合法的。”
MATT|14|5|希律 就想要杀他，可是怕民众，因为他们认为 约翰 是先知。
MATT|14|6|到了 希律 的生日， 希罗底 的女儿在众人面前跳舞，使 希律 欢喜，
MATT|14|7|于是 希律 发誓许诺随她所求的给她。
MATT|14|8|女儿被母亲指使，就说：“请把施洗 约翰 的头放在盘子里，拿来给我。”
MATT|14|9|王就忧愁，然而因他所发的誓，又因同席的人，就下令给她；
MATT|14|10|于是打发人去，在监狱里斩了 约翰 ，
MATT|14|11|把头放在盘子里，拿来给那女孩，她拿去给她母亲。
MATT|14|12|约翰 的门徒来，把尸体领去埋葬了，又去告诉耶稣。
MATT|14|13|耶稣听到了，就从那里上船，私下退到荒野的地方去。众人听到后，从各城来，步行跟随他。
MATT|14|14|耶稣出来，见有一大群人，就怜悯他们，治好了他们的病人。
MATT|14|15|傍晚的时候，门徒进前来，说：“这地方偏僻，而且时候已经晚了，请叫众人散去，他们好进村子，自己买些食物。”
MATT|14|16|耶稣对他们说：“不用他们去，你们给他们吃吧！”
MATT|14|17|门徒说：“我们这里只有五个饼、两条鱼。”
MATT|14|18|耶稣说：“拿过来给我。”
MATT|14|19|于是他吩咐众人坐在草地上，就拿着这五个饼和两条鱼，望着天祝福，擘开饼，递给门徒，门徒又递给众人。
MATT|14|20|他们都吃，并且吃饱了。门徒把剩下的碎屑收拾起来，装满了十二个篮子。
MATT|14|21|吃的人中，男的约有五千，还不算妇女和孩子。
MATT|14|22|耶稣随即催门徒上船，先渡到对岸，等他叫众人散去。
MATT|14|23|疏散了众人以后，他独自上山去祷告。到了晚上，只有他一人在那里。
MATT|14|24|那时船已离岸好几里 ，因风不顺，被浪颠簸。
MATT|14|25|天快亮的时候，耶稣在海面上走，往门徒那里去。
MATT|14|26|但门徒看见他在海面上走，就惊慌了，说：“是个鬼怪！”他们害怕得喊叫起来。
MATT|14|27|耶稣连忙对他们说：“放心！是我，不要怕！”
MATT|14|28|彼得 回答他说：“主啊，如果是你，请叫我从水面上走到你那里去。”
MATT|14|29|耶稣说：“你来吧！” 彼得 就从船上下去，在水面上走，往耶稣那里去；
MATT|14|30|只因见风很强 ，害怕起来，将要沉下去，就喊着说：“主啊，救我！”
MATT|14|31|耶稣立刻伸手拉住他，说：“你这小信的人哪，为什么疑惑呢？”
MATT|14|32|他们一上船，风就停了。
MATT|14|33|在船上的人都拜他，说：“你真是上帝的儿子。”
MATT|14|34|他们渡过了海，在 革尼撒勒 上岸。
MATT|14|35|那里的人认出耶稣，就打发人到整个周围地区去，把所有的病人带到他那里，
MATT|14|36|求耶稣让他们只摸一摸他的衣裳繸子，摸着的人就都好了。
MATT|15|1|那时，有法利赛人和文士从 耶路撒冷 来见耶稣，说：
MATT|15|2|“你的门徒为什么违反古人的传统？因为他们吃饭的时候不洗手。”
MATT|15|3|耶稣回答他们：“你们为什么因你们的传统而违反上帝的诫命呢？
MATT|15|4|上帝说：‘当孝敬父母’；又说：‘咒骂父母的，必须处死。’
MATT|15|5|你们倒说：‘无论谁对父母说：我所当供奉你的已经作了奉献，
MATT|15|6|就可以不孝敬他的父亲 。’这就是你们藉着传统，废了上帝的话。
MATT|15|7|假冒为善的人哪！ 以赛亚 指着你们所预言的说得好：
MATT|15|8|‘这百姓用嘴唇尊敬我， 他们的心却远离我。
MATT|15|9|他们把人的规条当作教义教导人； 他们拜我也是枉然。’”
MATT|15|10|耶稣叫了众人来，对他们说：“你们要听，也要明白。
MATT|15|11|从口里进去的不玷污人，从口里出来的才玷污人。”
MATT|15|12|当时，门徒进前来对他说：“法利赛人听见这话很反感，你知道吗？”
MATT|15|13|耶稣回答：“一切植物，若不是我天父栽植的，都要连根拔出来。
MATT|15|14|由他们吧！他们是瞎子作瞎子的向导 ；若是瞎子领瞎子，两个人都要掉在坑里。”
MATT|15|15|彼得 回应他说：“请将这比喻讲解给我们听。”
MATT|15|16|耶稣说：“连你们也还不明白吗？
MATT|15|17|难道你们不了解，凡进到口里的，是经过肚子，又排入厕所吗？
MATT|15|18|然而口里出来的是出于心里，这才玷污人。
MATT|15|19|因为出于心里的有种种恶念，如凶杀、奸淫、淫乱、偷盗、伪证、毁谤。
MATT|15|20|这些才玷污人。至于不洗手吃饭，那并不玷污人。”
MATT|15|21|耶稣离开那里，退到 推罗 、 西顿 境内。
MATT|15|22|有一个 迦南 妇人从那地方出来，喊着说：“主啊， 大卫 之子，可怜我！我女儿被鬼缠得很苦。”
MATT|15|23|耶稣却一言不答。门徒进前来，求他说：“这妇人在我们后头喊叫，请打发她走吧。”
MATT|15|24|耶稣回答：“我奉差遣只到 以色列 家迷失的羊那里去。”
MATT|15|25|那妇人来拜他，说：“主啊，帮帮我！”
MATT|15|26|他回答：“拿孩子的饼丢给小狗吃是不妥的。”
MATT|15|27|妇人说：“主啊，不错，可是小狗也吃它主人桌上掉下来的碎屑。”
MATT|15|28|于是耶稣回答她说：“妇人，你的信心很大！照你所要的成全你吧。”从那时起，她的女儿就好了。
MATT|15|29|耶稣离开那地方，来到靠近 加利利 的海边，就上山坐下。
MATT|15|30|有一大群人到他那里，带着瘸子、盲人、肢残的、聋哑的，和好些别的病人，都放在他脚前，他就治好了他们。
MATT|15|31|于是众人都惊讶，因为看见聋哑的说话，肢残的痊愈，瘸子行走，盲人看见，他们就归荣耀给 以色列 的上帝。
MATT|15|32|耶稣叫门徒来，说：“我怜悯这群人，因为他们同我在这里已经三天，没有吃的东西了。我不愿意叫他们饿着回去，恐怕他们在路上饿昏了。”
MATT|15|33|门徒说：“我们在这野地，哪里有这么多的饼让这许多人吃饱呢？”
MATT|15|34|耶稣对他们说：“你们有多少饼？”他们说：“有七个，还有几条小鱼。”
MATT|15|35|他就吩咐众人坐在地上，
MATT|15|36|拿着这七个饼和几条鱼，祝谢了，擘开，递给门徒；门徒又递给众人。
MATT|15|37|他们都吃，并且吃饱了，收拾剩下的碎屑，装满了七个筐子。
MATT|15|38|吃的人中，男的有四千，还不算妇女和孩子。
MATT|15|39|耶稣叫众人散去，就上船，来到 马加丹 境内。
MATT|16|1|法利赛人和撒都该人来试探耶稣，请他显个来自天上的神迹给他们看。
MATT|16|2|耶稣回答他们：“傍晚天发红，你们就说：‘明日天晴。’
MATT|16|3|早晨天色又红又暗，你们就说：‘今日有风雨。’你们知道分辨天上的气象，倒不能分辨这个时代的神迹 。
MATT|16|4|邪恶淫乱的世代求看神迹，除了 约拿 的神迹以外，再没有神迹给他们看了。”于是耶稣离开他们走了。
MATT|16|5|门徒渡到对岸，忘了带饼。
MATT|16|6|耶稣对他们说：“你们要谨慎，要防备法利赛人和撒都该人的酵。”
MATT|16|7|门徒彼此议论说：“这是因为我们没有带饼吧。”
MATT|16|8|耶稣知道了，就说：“你们这小信的人，为什么因为没有饼就彼此议论呢？
MATT|16|9|你们还不明白吗？不记得那五个饼分给五千人，你们收拾了多少篮子的碎屑吗？
MATT|16|10|也不记得那七个饼分给四千人，你们又收拾了多少筐子的碎屑吗？
MATT|16|11|我对你们说‘要防备法利赛人和撒都该人的酵’，这话不是指着饼说的，你们怎么不明白呢？”
MATT|16|12|门徒这才明白他所说的不是要他们防备饼的酵 ，而是要防备法利赛人和撒都该人的教训。
MATT|16|13|耶稣到了 凯撒利亚．腓立比 的境内，就问门徒：“人们说人子是谁？”
MATT|16|14|他们说：“有人说是施洗的 约翰 ；有人说是 以利亚 ；又有人说是 耶利米 或是先知中的一位。”
MATT|16|15|耶稣问他们：“你们说我是谁？”
MATT|16|16|西门．彼得 回答说：“你是基督，是永生上帝的儿子。”
MATT|16|17|耶稣回答他说：“ 约拿 的儿子 西门 ，你是有福的！因为这不是属血肉的启示你的，而是我在天上的父启示的。
MATT|16|18|我还告诉你，你是 彼得 ，我要把我的教会建造在这磐石上，阴间的权柄不能胜过它。
MATT|16|19|我要把天国的钥匙给你，凡你在地上所捆绑的，在天上也要捆绑；凡你在地上所释放的，在天上也要释放。”
MATT|16|20|当时，耶稣嘱咐门徒不可对任何人说他是基督。
MATT|16|21|从那时起，耶稣才向门徒明说，他必须上 耶路撒冷 去，受长老、祭司长和文士许多的苦，并且被杀，第三天复活。
MATT|16|22|彼得 就拉着他，责备他说：“主啊，千万不可如此！这事绝不可临到你身上。”
MATT|16|23|耶稣转过来，对 彼得 说：“撒但，退到我后边去！你是我的绊脚石，因为你不体会上帝的心意，而是体会人的意思。”
MATT|16|24|于是耶稣对门徒说：“若有人要跟从我，就当舍己，背起自己的十字架来跟从我。
MATT|16|25|因为凡要救自己生命的，要丧失生命；凡为我丧失生命的，要得着生命。
MATT|16|26|人若赚得全世界，赔上自己的生命，有什么益处呢？人还能拿什么换生命呢？
MATT|16|27|人子要在他父的荣耀里与他的众使者一起来临，那时候，他要照各人的行为报应各人。
MATT|16|28|我实在告诉你们，站在这里的，有人在没经历死亡以前，必定看见人子来到他的国里。”
MATT|17|1|过了六天，耶稣带着 彼得 、 雅各 和 雅各 的弟弟 约翰 ，领他们悄悄地上了高山。
MATT|17|2|他在他们面前变了形像，他的脸明亮如太阳，衣裳洁白如光。
MATT|17|3|忽然，有 摩西 和 以利亚 向他们显现，与耶稣说话。
MATT|17|4|彼得 回应，对耶稣说：“主啊，我们在这里真好！你若愿意，我就在这里搭三座棚，一座为你，一座为 摩西 ，一座为 以利亚 。”
MATT|17|5|说话之间，忽然有一朵明亮的云彩遮盖他们，又有声音从云彩里出来，说：“这是我的爱子，我所喜爱的。你们要听从他！”
MATT|17|6|门徒听见，就俯伏在地，极其害怕。
MATT|17|7|耶稣进前来，拍拍他们，说：“起来，不要害怕！”
MATT|17|8|他们举目，不见一人，只见耶稣独自一人。
MATT|17|9|下山的时候，耶稣嘱咐他们说：“人子还没有从死人中复活，你们不要把所看到的告诉人。”
MATT|17|10|门徒问耶稣：“那么，文士为什么说 以利亚 必须先来？”
MATT|17|11|耶稣回答：“ 以利亚 的确要来，并要复兴万事；
MATT|17|12|可是我告诉你们， 以利亚 已经来了，人不认识他，反倒任意待他。人子也将这样受他们的苦。”
MATT|17|13|门徒这才明白耶稣所说的是指施洗的 约翰 。
MATT|17|14|耶稣和门徒到了众人那里，有一个人来见耶稣，跪下，
MATT|17|15|说：“主啊，可怜我的儿子。他害癫痫病很苦，屡次跌进火里，屡次跌进水里。
MATT|17|16|我带他到你门徒那里，他们却不能医治他。”
MATT|17|17|耶稣回答：“唉！这又不信又悖谬的世代啊，我和你们在一起要到几时呢？我忍耐你们要到几时呢？把他带到我这里来！”
MATT|17|18|耶稣斥责那鬼，鬼就出来；从那时起，孩子就痊愈了。
MATT|17|19|门徒私下进前来问耶稣：“我们为什么不能赶出那鬼呢？”
MATT|17|20|耶稣对他们说：“是因你们的信心小。我实在告诉你们，你们若有信心像一粒芥菜种，就是对这座山说：‘你从这边移到那边’，它也会移过去，并且你们没有一件不能做的事了。 ”
MATT|17|21|
MATT|17|22|他们聚集在 加利利 的时候，耶稣对门徒说：“人子将要被交在人手里。
MATT|17|23|他们要杀害他，第三天他要复活。”门徒就非常忧愁。
MATT|17|24|他们到了 迦百农 ，收圣殿税 的人来见 彼得 ，说：“你们的老师不纳圣殿税吗？”
MATT|17|25|彼得 说：“纳。”他进了屋子，耶稣先对他说：“ 西门 ，你的意见如何？世上的君王向谁征收关税或丁税？是向自己的儿子呢？还是向外人呢？”
MATT|17|26|彼得 说：“是向外人。”耶稣对他说：“既然如此，儿子就可以免了。
MATT|17|27|但恐怕触犯他们，你往海边去钓鱼，把先钓上来的鱼拿起来，开了它的口，会发现一个司塔特 ，可以拿去给他们，作你我的税钱。”
MATT|18|1|当时，门徒前来问耶稣：“天国里谁是最大的？”
MATT|18|2|耶稣叫一个小孩子来，让他站在他们当中，
MATT|18|3|说：“我实在告诉你们，你们若不回转，变成像小孩子一样，绝不能进天国。
MATT|18|4|所以，凡自己谦卑像这小孩子的，他在天国里就是最大的。
MATT|18|5|凡为我的名接纳一个像这小孩子的，就是接纳我。”
MATT|18|6|“凡使这些信我的小子中的一个跌倒的，倒不如把大磨石拴在这人的颈项上，沉在深海里。
MATT|18|7|这世界有祸了，因为它使人跌倒；绊倒人的事是免不了的，但那绊倒人的有祸了！
MATT|18|8|如果你一只手或是一只脚使你跌倒，就把它砍下来扔掉。你缺一只手或是一只脚进入永生，比有两手两脚被扔进永火里还好。
MATT|18|9|如果你一只眼使你跌倒，就把它挖出来扔掉。你只有一只眼进入永生，比有两只眼被扔进地狱的火里还好。”
MATT|18|10|“你们要小心，不可轻看这些小子中的一个；我告诉你们，他们的天使在天上，常见我天父的面。
MATT|18|11|
MATT|18|12|“一个人若有一百只羊，其中一只走迷了路，你们的意见如何？他岂不留下这九十九只在山上，去找那只迷路的羊吗？
MATT|18|13|若是找到了，我实在告诉你们，他为这一只羊欢喜，比为那没有迷路的九十九只欢喜还大呢！
MATT|18|14|你们 在天上的父也是这样，不愿意失去这些小子中的一个。”
MATT|18|15|“若是你的弟兄得罪你 ，你要去，趁着只有他和你在一起的时候，指出他的错来。他若听你，你就赢得了你的弟兄；
MATT|18|16|他若不听，你就另外带一个或两个人同去，因为‘任何指控都要凭两个或三个证人的口述才能成立’。
MATT|18|17|他若是不听他们，就去告诉教会；若是不听教会，就把他看作外邦人和税吏。
MATT|18|18|“我实在告诉你们，凡你们在地上所捆绑的，在天上也要捆绑；凡你们在地上所释放的，在天上也要释放。
MATT|18|19|我又实在 告诉你们，若是你们中间有两个人在地上同心合意地求什么事，我在天上的父必为他们成全。
MATT|18|20|因为，哪里有两三个人奉我的名聚会，哪里就有我在他们中间。”
MATT|18|21|那时， 彼得 进前来，对耶稣说：“主啊，我弟兄得罪我，我当饶恕他几次呢？到七次够吗？”
MATT|18|22|耶稣说：“我告诉你，不是到七次，而是到七十个七次。
MATT|18|23|因为天国好像一个王要和他仆人算账。
MATT|18|24|他开始算的时候，有人带了一个欠一万他连得的仆人来。
MATT|18|25|因为他没有什么偿还之物，主人下令把他和他妻子儿女，以及一切所有的都卖了来偿还。
MATT|18|26|那仆人就俯伏向他叩头，说：‘宽容我吧，我都会还你的。’
MATT|18|27|那仆人的主人就动了慈心，把他释放了，并且免了他的债。
MATT|18|28|那仆人出来，遇见一个欠他一百个银币的同伴，就揪着他，扼住他的喉咙，说：‘把你所欠的还我！’
MATT|18|29|他的同伴就俯伏央求他，说：‘宽容我吧，我会还你的。’
MATT|18|30|他不肯，却把他下在监里，直到他还了所欠的债。
MATT|18|31|同伴们看见他所做的事就很悲愤，把这一切的事都告诉了主人。
MATT|18|32|于是主人叫了他来，对他说：‘你这恶奴才！你央求我，我就把你所欠的都免了；
MATT|18|33|你不应该怜悯你的同伴，像我怜悯你吗？’
MATT|18|34|主人就大怒，把他交给司刑的，直到他还清了所欠的债。
MATT|18|35|你们各人若不从心里饶恕你的弟兄，我天父也要这样待你们。”
MATT|19|1|耶稣说完了这些话，就离开 加利利 ，来到 犹太 的境内、 约旦河 的东边。
MATT|19|2|有一大群人跟着他，他就在那里治好了他们。
MATT|19|3|有些法利赛人来试探耶稣说：“无论什么缘故，人休妻都合法吗？”
MATT|19|4|耶稣回答：“那起初造人的，是造男造女，并且说：‘因此，人要离开父母，与妻子结合，二人成为一体。’这经文你们没有念过吗？
MATT|19|5|
MATT|19|6|既然如此，夫妻不再是两个人，而是一体的了。所以，上帝配合的，人不可分开。”
MATT|19|7|法利赛人说：“这样， 摩西 为什么吩咐给妻子休书就可以休她呢？”
MATT|19|8|耶稣说：“ 摩西 因为你们的心硬，所以准许你们休妻，但起初并不是这样。
MATT|19|9|我告诉你们，凡休妻另娶的，若不是为不贞的缘故，就是犯奸淫了。 ”
MATT|19|10|门徒对耶稣说：“丈夫和妻子的关系既是这样，倒不如不娶。”
MATT|19|11|耶稣对他们说：“这话不是人人都能领受的，惟独赐给谁，谁才能领受。
MATT|19|12|因为有人从母腹里就是不宜结婚的，也有因人为的缘故不宜结婚的，并有为天国的缘故自己不结婚的 。这话谁能领受，就领受吧。”
MATT|19|13|那时，有人带着小孩子来见耶稣，要他给他们按手祷告，门徒就责备那些人。
MATT|19|14|耶稣说：“让小孩子到我这里来，不要阻止他们，因为在天国的正是这样的人。”
MATT|19|15|耶稣给他们按手，然后离开那地方。
MATT|19|16|有一个人进前来问耶稣：“老师，我该做什么善事才能得永生？”
MATT|19|17|耶稣对他说：“你为什么问我关于善的事呢？只有一位是善良的。你若要进入永生，就该遵守诫命。”
MATT|19|18|他说：“哪些诫命？”耶稣说：“就是不可杀人；不可奸淫；不可偷盗；不可作假见证；
MATT|19|19|当孝敬父母；又当爱邻 如己。”
MATT|19|20|那青年说：“这一切我都遵守了，还缺少什么呢？”
MATT|19|21|耶稣说：“你若愿意作完全人，去变卖你所拥有的，分给穷人，就必有财宝在天上；然后来跟从我。”
MATT|19|22|那青年听见这话，就忧忧愁愁地走了，因为他的产业很多。
MATT|19|23|耶稣对门徒说：“我实在告诉你们，财主进天国是难的。
MATT|19|24|我再告诉你们，骆驼穿过针眼比财主进上帝的国还容易呢！”
MATT|19|25|门徒听见这话，就非常惊奇，说：“这样，谁能得救呢？”
MATT|19|26|耶稣看着他们，说：“在人这是不能，在上帝凡事都能。”
MATT|19|27|于是 彼得 回应，对他说：“看哪，我们已经撇下一切跟从你了，我们会得到什么呢？”
MATT|19|28|耶稣对他们说：“我实在告诉你们，你们这些跟从我的人，到了万物更新、人子坐在他荣耀宝座上的时候，你们也要坐在十二个宝座上，审判 以色列 十二个支派。
MATT|19|29|凡为我的名撇下房屋，或是兄弟、姊妹、父亲、母亲、 儿女、田地的，将得着百倍，并且承受永生。
MATT|19|30|然而，有许多在前的，将要在后；在后的，将要在前。”
MATT|20|1|“因为天国好比一家的主人清早去雇人进他的葡萄园做工。
MATT|20|2|他和工人讲定一天一个银币 ，就打发他们进葡萄园去。
MATT|20|3|约在上午九点钟出去，看见市场上还有闲站的人，
MATT|20|4|就对那些人说：‘你们也进葡萄园去，我会给你们合理的工钱。’
MATT|20|5|他们也进去了。约在正午和下午三点钟又出去，他也是这么做。
MATT|20|6|约在下午五点钟出去，他看见还有人站在那里，就问他们：‘你们为什么整天在这里闲站呢？’
MATT|20|7|他们说：‘因为没有人雇我们。’他说：‘你们也进葡萄园去。’
MATT|20|8|到了晚上，园主对工头说：‘叫工人都来，给他们工钱，从后来的起，到先来的为止。’
MATT|20|9|约在下午五点钟雇的人来了，各人领了一个银币。
MATT|20|10|那些最先雇的来了，以为可以多领，谁知也是各领一个银币。
MATT|20|11|他们领了工钱，就埋怨那家的主人说：
MATT|20|12|‘我们整天劳苦受热，那些后来的只做了一小时，你竟待他们和我们一样吗？’
MATT|20|13|主人回答其中的一人说：‘朋友，我没亏待你，你与我讲定的不是一个银币吗？
MATT|20|14|拿你的钱走吧！我乐意给那后来的和给你的一样，
MATT|20|15|难道我的东西不可随我的意思用吗？因为我作好人，你就眼红了吗？’
MATT|20|16|这样，那在后的，将要在前；在前的，将要在后了。”
MATT|20|17|耶稣上 耶路撒冷 去的时候，在路上把十二个门徒带到一边，对他们说：
MATT|20|18|“看哪，我们上 耶路撒冷 去，人子将被交给祭司长和文士；他们要定他死罪，
MATT|20|19|把他交给外邦人戏弄，鞭打，钉在十字架上；第三天他要复活。”
MATT|20|20|那时， 西庇太 儿子的母亲和她两个儿子上前来，向耶稣叩头，求他一件事。
MATT|20|21|耶稣问她：“你要什么呢？”她对耶稣说：“在你的国里，请让我这两个儿子一个坐在你右边，一个坐在你左边。”
MATT|20|22|耶稣回答：“你们不知道所求的是什么。我将要喝的杯，你们能喝吗？”他们对他说：“我们能。”
MATT|20|23|耶稣说：“我所喝的杯，你们要喝。可是坐在我的左右，不是我可以赐的，而是我父为谁预备就赐给谁。”
MATT|20|24|其余十个门徒听见，就对他们兄弟二人很生气。
MATT|20|25|耶稣叫了他们来，说：“你们知道，外邦人有君王作主治理他们，有大臣操权管辖他们。
MATT|20|26|但是在你们中间，不可这样。你们中间谁愿为大，就要作你们的用人；
MATT|20|27|谁愿为首，就要作你们的仆人。
MATT|20|28|正如人子来，不是要受人的服事，乃是要服事人，并且要舍命，作多人的赎价。”
MATT|20|29|他们出 耶利哥 的时候，有一大群人跟随耶稣。
MATT|20|30|有两个盲人坐在路旁，听说是耶稣经过，就喊着说：“主啊 ， 大卫 之子，可怜我们吧！”
MATT|20|31|众人责备他们，不许他们作声，他们却越发喊着说：“主啊 ， 大卫 之子，可怜我们吧！”
MATT|20|32|耶稣就站住，叫他们来，说：“你们要我为你们做什么？”
MATT|20|33|他们说：“主啊，让我们的眼睛能看见。”
MATT|20|34|耶稣动了慈心，摸了他们的眼睛，他们立刻看得见，就跟从耶稣。
MATT|21|1|耶稣和门徒快到 耶路撒冷 ，进了 橄榄山 的 伯法其 时，打发两个门徒，
MATT|21|2|对他们说：“你们往对面村子里去，会立刻看见一匹驴拴在那里，还有驴驹同在一处，解开它们，牵到我这里来。
MATT|21|3|若有人对你们说什么，你们就说：‘主要用它们。’那人会立刻让你们牵来。”
MATT|21|4|这事发生是要应验先知所说的话：
MATT|21|5|“要对 锡安 的儿女 说： 看哪，你的王来到你这里， 谦和地骑着驴， 骑着小驴—驴的驹子。”
MATT|21|6|门徒就照耶稣所吩咐的去做，
MATT|21|7|牵了驴和驴驹来，把他们的衣服搭在上面，耶稣就骑上。
MATT|21|8|许许多多的人把自己的衣服铺在路上，还有人砍下树枝来铺在路上。
MATT|21|9|前呼后拥的人群喊着说： “和散那 归于 大卫 之子！ 奉主名来的是应当称颂的！ 至高无上的，和散那！”
MATT|21|10|耶稣进了 耶路撒冷 ，全城都惊动了，说：“这是谁？”
MATT|21|11|众人说：“这是从 加利利 的 拿撒勒 来的先知耶稣。”
MATT|21|12|耶稣进了圣殿 ，赶出圣殿里所有在做买卖的人，推倒兑换银钱之人的桌子和卖鸽子之人的凳子，
MATT|21|13|对他们说：“经上记着： ‘我的殿要称为祷告的殿， 你们倒使它成为贼窝了。’”
MATT|21|14|在圣殿里有盲人和瘸子到耶稣跟前，他就治好了他们。
MATT|21|15|祭司长和文士看见耶稣所行的奇事，又见小孩子在圣殿里喊着说：“和散那归于 大卫 之子！”就很生气，
MATT|21|16|对他说：“这些人所喊的，你听到了吗？”耶稣对他们说：“听到了。经上说：‘你藉孩童和吃奶的口发出完全的赞美’，你们没有念过吗？”
MATT|21|17|于是他离开他们，出城到 伯大尼 去，在那里过夜。
MATT|21|18|早晨回城的时候，他饿了，
MATT|21|19|看见路旁有一棵无花果树，就走到跟前，在树上找不到什么，只有叶子，就对树说：“从今以后，你永不结果子！”那无花果树立刻枯干了。
MATT|21|20|门徒看见了，惊讶地说：“无花果树怎么立刻枯干了呢？”
MATT|21|21|耶稣回答他们：“我实在告诉你们，你们若有信心，不疑惑，不但能行我对无花果树所行的事，就是对这座山说：‘离开此地，投在海里！’也会实现。
MATT|21|22|你们祷告，无论求什么，只要信，就必得着。”
MATT|21|23|耶稣进了圣殿，正教导人的时候，祭司长和百姓的长老来问他：“你仗着什么权柄做这些事？给你这权柄的是谁呢？”
MATT|21|24|耶稣回答他们说：“我也要问你们一句话，你们若告诉我，我就告诉你们我仗着什么权柄做这些事。
MATT|21|25|约翰 的洗礼是从哪里来的？是从天上来的，还是从人间来的呢？”他们彼此商议说：“我们若说‘从天上来的’，他会对我们说：‘这样，你们为什么不信他呢？’
MATT|21|26|若说‘从人间来的’，我们又怕众人，因为大家都认为 约翰 是先知。”
MATT|21|27|于是他们回答耶稣：“我们不知道。”耶稣也对他们说：“我也不告诉你们，我仗着什么权柄做这些事。”
MATT|21|28|“有一件事，你们的意见如何？一个人有两个儿子。他来对大儿子说：‘孩子，今天到葡萄园里做工去。’
MATT|21|29|他回答：‘我不去’，以后自己懊悔，就去了。
MATT|21|30|他来对小儿子也是这样说。他回答：‘父亲大人，我去’，却不去。
MATT|21|31|这两个儿子是哪一个照着父亲的意愿做了呢？”他们说：“大儿子。”耶稣说：“我实在告诉你们，税吏和娼妓倒比你们先进上帝的国。
MATT|21|32|因为 约翰 到你们这里来指引你们走义路，你们却不信他，税吏和娼妓倒信了他。你们看见了以后，还是不悔悟去信他。”
MATT|21|33|“你们再听一个比喻：有一个家的主人开垦了一个葡萄园，四周围上篱笆，里面挖了一个榨酒池，盖了一座守望楼，租给园户，就出外远行去了。
MATT|21|34|收果子的时候快到了，他打发仆人到园户那里去收果子。
MATT|21|35|园户拿住仆人，打了一个，杀了一个，用石头打死了一个。
MATT|21|36|主人又打发别的仆人去，比先前更多；园户还是照样对待他们。
MATT|21|37|最后他打发自己的儿子到他们那里去，说：‘他们会尊敬我的儿子。’
MATT|21|38|可是，园户看见他儿子，彼此说：‘这是承受产业的。来，我们杀了他，占他的产业！’
MATT|21|39|于是他们拿住他，把他扔出葡萄园外，杀了。
MATT|21|40|葡萄园的主人来的时候，要怎样处置那些园户呢？”
MATT|21|41|他们说：“要狠狠地除灭那些恶人，将葡萄园转租给那些按时候交果子的园户。”
MATT|21|42|耶稣对他们说： “‘匠人所丢弃的石头 已作了房角的头块石头。 这是主所做的， 在我们眼中看为奇妙。’ 这段经文你们从来没有念过吗？
MATT|21|43|所以我告诉你们，上帝的国必从你们夺去，赐给那能结果子的民。
MATT|21|44|谁跌在这石头上，一定会跌得粉碎；这石头掉在谁的身上，就要把谁压得稀烂。 ”
MATT|21|45|祭司长和法利赛人听见他的比喻，就看出他是指着他们说的。
MATT|21|46|他们想要捉拿他，但是惧怕众人，因为众人认为他是先知。
MATT|22|1|耶稣又用比喻对他们说：
MATT|22|2|“天国好比一个王为他儿子摆设娶亲的宴席。
MATT|22|3|他打发仆人去，请那些被邀的人来赴宴，他们却不肯来。
MATT|22|4|王又打发别的仆人，说：‘你们去告诉那被邀的人，我的宴席已经预备好了，牛和肥畜已经宰了，各样都齐备，请你们来赴宴。’
MATT|22|5|那些人不理就走了，一个到自己田里去，一个做买卖去。
MATT|22|6|其余的抓住仆人，凌辱他们，把他们杀了。
MATT|22|7|王就大怒，发兵除灭那些凶手，烧毁他们的城。
MATT|22|8|于是王对仆人说：‘喜宴已经齐备，只是所邀的人不配。
MATT|22|9|所以你们要往岔路口上去，凡遇见的，都邀来赴宴。’
MATT|22|10|那些仆人就出去，到大路上，凡遇见的，不论善恶都招聚了来，宴席上就坐满了客人。
MATT|22|11|王进来见宾客，看到那里有一个没有穿礼服的，
MATT|22|12|就对他说：‘朋友，你到这里来怎么不穿礼服呢？’那人无言可答。
MATT|22|13|于是王对侍从说：‘捆起他的手脚，把他扔在外边的黑暗里；在那里他要哀哭切齿了。’
MATT|22|14|因为被召的人多，选上的人少。”
MATT|22|15|于是，法利赛人出去商议，怎样找话柄来陷害耶稣，
MATT|22|16|就打发他们的门徒同 希律 党人去见耶稣，说：“老师，我们知道你是诚实的，并且诚诚实实传上帝的道，无论谁你都一视同仁，因为你不看人的面子。
MATT|22|17|请告诉我们，你的意见如何？纳税给凯撒合不合法？”
MATT|22|18|耶稣看出他们的恶意，就说：“假冒为善的人哪，为什么试探我？
MATT|22|19|拿一个纳税的钱给我看！”他们就拿一个银币来给他。
MATT|22|20|耶稣问他们：“这像和这名号是谁的？”
MATT|22|21|他们说：“是凯撒的。”于是耶稣说：“这样，凯撒的归凯撒；上帝的归上帝。”
MATT|22|22|他们听了十分惊讶，就离开他走了。
MATT|22|23|那天，撒都该人来见耶稣。他们说没有复活这回事，于是问耶稣：
MATT|22|24|“老师， 摩西 说：‘某人若死了，没有孩子，他弟弟该娶他的妻子，为哥哥生子立后。’
MATT|22|25|从前，在我们这里有兄弟七人，第一个娶了妻，死了，没有孩子，撇下妻子给弟弟。
MATT|22|26|第二、第三，直到第七个，都是如此。
MATT|22|27|后来，那妇人也死了。
MATT|22|28|那么，在复活的时候，她是七个人中哪一个的妻子呢？因为他们都娶过她。”
MATT|22|29|耶稣回答他们说：“你们错了，因为不明白圣经，也不知道上帝的大能。
MATT|22|30|在复活的时候，人也不娶也不嫁，而是像天上的天使一样。
MATT|22|31|论到死人复活，上帝向你们所说的话，你们没有念过吗？
MATT|22|32|他说：‘我是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。’上帝不是死人的上帝，而是活人的上帝。”
MATT|22|33|众人听见这话，对他的教导非常惊讶。
MATT|22|34|法利赛人听见耶稣堵住了撒都该人的口，他们就聚集在一起。
MATT|22|35|其中有一个人是律法师 ，要试探耶稣，就问他：
MATT|22|36|“老师，律法上的诫命哪一条是最大的呢？”
MATT|22|37|耶稣对他说：“你要尽心、尽性、尽意爱主—你的上帝。
MATT|22|38|这是最大的，且是第一条诫命。
MATT|22|39|第二条也如此，就是要爱邻 如己。
MATT|22|40|这两条诫命是一切律法和先知书的总纲。”
MATT|22|41|法利赛人聚集的时候，耶稣问他们：
MATT|22|42|“论到基督，你们的意见如何？他是谁的后裔呢？”他们说：“是 大卫 的。”
MATT|22|43|耶稣说：“这样， 大卫 被圣灵感动，怎么还称他为主，说：
MATT|22|44|‘主对我主说： 你坐在我的右边， 等我把你的仇敌放在你脚下？’
MATT|22|45|大卫 既称他为主，他怎么又是 大卫 的后裔呢？”
MATT|22|46|没有一个人能回答一句话，从那日以后没有人敢再问他什么。
MATT|23|1|那时，耶稣对众人和门徒讲论，
MATT|23|2|说：“文士和法利赛人坐在 摩西 的位上，
MATT|23|3|所以凡他们所吩咐你们的，你们都要谨守遵行。但不要效法他们的行为，因为他们能说不能行。
MATT|23|4|他们把难挑的 重担捆起来，搁在人的肩上，但自己一个指头也不肯动。
MATT|23|5|他们所做的一切事都是要让人看见，所以把佩戴的经匣 加宽了，衣裳的繸子加长了，
MATT|23|6|喜爱宴席上的首座、会堂里的高位，
MATT|23|7|又喜欢人们在街市上向他们问安，称呼他们拉比 。
MATT|23|8|但你们不要接受拉比的称呼，因为只有一位是你们的老师；你们都是弟兄。
MATT|23|9|也不要称呼地上的人为父，因为只有一位是你们的父，就是在天上的父。
MATT|23|10|不要接受师傅的称呼，因为只有一位是你们的师傅，就是基督。
MATT|23|11|你们中间谁为大，谁就要作你们的用人。
MATT|23|12|凡自高的，必降为卑；自甘卑微的，必升为高。
MATT|23|13|“你们这假冒为善的文士和法利赛人有祸了！因为你们当着人的面把天国的门关了，自己不进去，要进去的人，你们也不容他们进去。
MATT|23|14|
MATT|23|15|“你们这假冒为善的文士和法利赛人有祸了！因为你们走遍海洋陆地，说服一个人入教，既入了教，却使他成为比你们加倍坏的地狱之子。
MATT|23|16|“你们这瞎眼的向导有祸了！你们说：‘凡指着圣所起誓的算不得什么；但是凡指着圣所中的金子起誓的，他就该谨守。’
MATT|23|17|你们这无知的瞎子啊，哪个更大呢？是金子，还是使金子成圣的圣所呢？
MATT|23|18|你们又说：‘凡指着祭坛起誓的算不得什么；但是凡指着坛上祭物起誓的，他就该谨守。’
MATT|23|19|你们这些瞎子啊，哪个更大呢？是祭物，还是使祭物成圣的坛呢？
MATT|23|20|所以，人指着祭坛起誓，就是指着坛和坛上一切所有的起誓；
MATT|23|21|人指着圣所起誓，就是指着圣所和那住在圣所里的起誓；
MATT|23|22|人指着天起誓，就是指着上帝的宝座和那坐在上面的起誓。
MATT|23|23|“你们这假冒为善的文士和法利赛人有祸了！因为你们将薄荷、大茴香、小茴香献上十分之一，那律法上更重要的事，就是公义、怜悯、信实，你们反倒不做；这原是你们该做的－至于那些奉献也不可废弃。
MATT|23|24|你们这瞎眼的向导，蠓虫你们就滤出来，骆驼你们倒吞下去。
MATT|23|25|“你们这假冒为善的文士和法利赛人有祸了！因为你们洗净杯盘的外面，里面却满了贪婪和放荡。
MATT|23|26|你这瞎眼的法利赛人，先洗净杯子 的里面，好使外面也干净了。
MATT|23|27|“你们这假冒为善的文士和法利赛人有祸了！因为你们好像粉饰了的坟墓，外面好看，里面却满了死人的骨头和一切的污秽。
MATT|23|28|你们也是如此，外面对人显出公义，里面却满了虚伪和不法的事。
MATT|23|29|“你们这假冒为善的文士和法利赛人有祸了！因为你们建造先知的坟，装修义人的墓，
MATT|23|30|说：‘若是我们在先祖的时代，必不和他们一同流先知的血。’
MATT|23|31|这样，你们就证明自己是杀害先知的人的子孙了。
MATT|23|32|你们去充满你们祖宗的恶贯吧！
MATT|23|33|你们这些蛇啊，毒蛇的孽种啊，怎能逃脱地狱的惩罚呢？
MATT|23|34|所以，我差遣先知、智慧人和文士到你们这里来，有的你们要杀害，要钉十字架；有的你们要在会堂里鞭打，从这城追逼到那城，
MATT|23|35|如此，地上所有义人流的血都归到你们身上，从义人 亚伯 的血起，直到你们在圣所和祭坛中间所杀的 巴拉加 的儿子 撒迦利亚 的血为止。
MATT|23|36|我实在告诉你们，这一切的罪都要归到这世代了。”
MATT|23|37|“ 耶路撒冷 啊， 耶路撒冷 啊，你常杀害先知，又用石头打死那奉差遣到你这里来的人。我多少次想聚集你的儿女，好像母鸡把小鸡聚集在翅膀底下，但是你们不愿意。
MATT|23|38|看吧，你们的家要被废弃成为荒芜。
MATT|23|39|我告诉你们，从今以后，你们绝不会再见到我，直到你们说：‘奉主名来的是应当称颂的！’”
MATT|24|1|耶稣出了圣殿，正离开的时候，门徒前来，把圣殿的建筑指给他看。
MATT|24|2|耶稣回应他们说：“你们不是看见这一切吗？我实在告诉你们，这里将没有一块石头会留在另一块石头上，而不被拆毁的。”
MATT|24|3|耶稣在 橄榄山 上坐着，门徒私下进前来问他：“请告诉我们，什么时候有这些事呢？你来临和世代的终结有什么预兆呢？”
MATT|24|4|耶稣回答他们：“你们要谨慎，免得有人迷惑你们。
MATT|24|5|因为将有好些人冒我的名来，说‘我是基督’，并且要迷惑许多人。
MATT|24|6|你们也将听见打仗和打仗的风声。注意，不要惊慌！因为这些事必须发生，但这还不是终结。
MATT|24|7|民要攻打民，国要攻打国，多处必有饥荒、地震。
MATT|24|8|这都是灾难 的起头。
MATT|24|9|那时，人要使你们陷在患难里，也要杀害你们；你们又要为我的名被万民憎恨。
MATT|24|10|那时，会有许多人跌倒，也会彼此陷害，彼此憎恨；
MATT|24|11|且有好些假先知起来，迷惑许多人。
MATT|24|12|因为不法的事增多，许多人的爱心渐渐冷淡了。
MATT|24|13|但坚忍到底的终必得救。
MATT|24|14|这天国的福音要传遍天下，对万民作见证，然后终结才来到。”
MATT|24|15|“当你们看见先知 但以理 所说的那‘施行毁灭的亵渎者’站在圣地（读这经的人要会意），
MATT|24|16|那时，在 犹太 的，应当逃到山上；
MATT|24|17|在屋顶上的，不要下来拿家里的东西；
MATT|24|18|在田里的，不要回去取衣裳。
MATT|24|19|在那些日子，怀孕的和奶孩子的就苦了。
MATT|24|20|你们要祈求，好让你们逃走的时候，不遇见冬天或安息日。
MATT|24|21|因为那时必有大灾难，自从世界的起头直到如今，从没有这样的灾难，将来也不会有。
MATT|24|22|若不减少那些日子，凡血肉之躯的，就没有一个能得救；可是为了选民，那些日子将减少。
MATT|24|23|那时，若有人对你们说：‘看哪，基督在这里！’或‘在那里！’你们不要信。
MATT|24|24|因为假基督和假先知将要起来，显大神迹、大奇事，如果可能，要把选民也迷惑了。
MATT|24|25|看哪，我已经预先告诉你们了。
MATT|24|26|若有人对你们说：‘看哪，基督在旷野里！’你们不要出去；或说：‘看哪，基督在内室中！’你们不要信。
MATT|24|27|好像闪电从东边发出，直照到西边，人子来临也要这样。
MATT|24|28|尸首在哪里，鹰也会聚在哪里。”
MATT|24|29|“那些日子的灾难一过去， 太阳要变黑， 月亮也不放光， 众星要从天上坠落， 天上的万象都要震动。
MATT|24|30|那时，人子的预兆要显在天上，地上的万族都要哀哭。他们要看见人子带着能力和大荣耀，驾着天上的云来临。
MATT|24|31|他要差遣天使，用大声的号筒，从四方，从天这边直到天那边，召集他的选民。”
MATT|24|32|“你们要从无花果树学习功课：当树枝发芽长叶的时候，你们就知道夏天近了。
MATT|24|33|同样，当你们看见这一切，就知道那时候近了，就在门口了。
MATT|24|34|我实在告诉你们，这世代还没有过去，这一切都要发生。
MATT|24|35|天地要废去，我的话却绝不废去。”
MATT|24|36|“但那日子，那时辰，没有人知道，连天上的天使也不知道，子也不知道，惟有父知道。
MATT|24|37|挪亚 的日子怎样，人子来临也要怎样。
MATT|24|38|在洪水以前的那些日子，人照常吃喝嫁娶，直到 挪亚 进方舟的那日，
MATT|24|39|不知不觉洪水来了，把他们全都冲去。人子来临也要这样。
MATT|24|40|那时，两个人在田里，一个被接去，一个被撇下。
MATT|24|41|两个女人推磨，一个被接去，一个被撇下。
MATT|24|42|所以，你们要警醒，因为不知道你们的主哪一天来到。
MATT|24|43|你们要知道，一家的主人若知道晚上什么时候有贼来，就必警醒，不让贼挖穿房屋。
MATT|24|44|所以，你们也要预备，因为在你们想不到的时候，人子就来了。”
MATT|24|45|“那么，谁是那忠心又精明的仆人，主人派他管理自己的家仆、按时分粮给他们的呢？
MATT|24|46|主人来到，看见仆人这样做，那仆人就有福了。
MATT|24|47|我实在告诉你们，主人要派他管理所有的财产。
MATT|24|48|如果那恶仆心里说：‘我的主人会来得迟’，
MATT|24|49|就动手打他的同伴，又和醉酒的人一同吃喝，
MATT|24|50|在想不到的日子，不知道的时候，那仆人的主人要来，
MATT|24|51|重重地惩罚他 ，定他和假冒为善的人同罪，在那里他要哀哭切齿了。”
MATT|25|1|“那时，天国好比十个童女拿着灯出去迎接新郎。
MATT|25|2|其中有五个是愚拙的，五个是聪明的。
MATT|25|3|愚拙的拿着灯，却没有带油；
MATT|25|4|聪明的拿着灯，又盛了油在器皿里。
MATT|25|5|新郎迟延的时候，她们都打盹，睡着了。
MATT|25|6|半夜有人喊：‘看，新郎来了，你们出来迎接他。’
MATT|25|7|那些童女就都起来挑亮她们的灯。
MATT|25|8|愚拙的对聪明的说：‘请分点油给我们，因为我们的灯要灭了。’
MATT|25|9|聪明的回答：‘恐怕不够你我用的；你们还是自己到卖油的那里去买吧。’
MATT|25|10|她们去买的时候，新郎到了。那预备好了的，与他进去共赴婚宴，门就关了。
MATT|25|11|其余的童女随后也来了，说：‘主啊，主啊，给我们开门！’
MATT|25|12|他却回答：‘我实在告诉你们，我不认识你们。’
MATT|25|13|所以，你们要警醒，因为那日子，那时辰，你们不知道。”
MATT|25|14|“天国又好比一个人要出外远行，就叫了仆人来，把他的家业交给他们。
MATT|25|15|他按着各人的才干，给他们银子：一个给了五千 ，一个给了二千 ，一个给了一千 ，就出外远行去了。
MATT|25|16|那领五千的立刻拿去做买卖，另外赚了五千。
MATT|25|17|那领二千的也照样另赚了二千。
MATT|25|18|但那领一千的去掘开地，把主人的银子埋藏了。
MATT|25|19|过了许久，那些仆人的主人来了，和他们算账。
MATT|25|20|那领五千的又带着另外的五千来，说：‘主啊，你交给我五千。请看，我又赚了五千。’
MATT|25|21|主人说：‘好，你这又善良又忠心的仆人，你在少许的事上忠心，我要派你管理许多的事，进来享受你主人的快乐吧！’
MATT|25|22|那领二千的也进前来，说：‘主啊，你交给我二千。请看，我又赚了二千。’
MATT|25|23|主人说：‘好，你这又善良又忠心的仆人，你在少许的事上忠心，我要派你管理许多的事，进来享受你主人的快乐吧！’
MATT|25|24|那领一千的也进前来，说：‘主啊，我知道你，你是个严厉的人：没有种的地方也要收割，没有播的地方也要收获，
MATT|25|25|我就害怕，去把你的一千银子埋藏在地里。请看，你的银子在这里。’
MATT|25|26|他的主人回答他说：‘你这又恶又懒的仆人，你既知道我没有种的地方也要收割，没有播的地方也要收获，
MATT|25|27|就该把我的银子放给兑换银钱的人，到我来的时候可以连本带利收回。
MATT|25|28|把他这一千夺过来，给那有一万 的。
MATT|25|29|因为凡有的，还要加给他，叫他有余；没有的，连他所有的也要夺过来。
MATT|25|30|把这无用的仆人丢在外面黑暗里，在那里他要哀哭切齿了。’”
MATT|25|31|“当人子在他荣耀里，同着众天使来临的时候，要坐在他荣耀的宝座上。
MATT|25|32|万民都要聚集在他面前。他要把他们分别出来，好像牧人分别绵羊、山羊一般，
MATT|25|33|把绵羊安置在右边，山羊在左边。
MATT|25|34|于是王要向他右边的说：‘你们这蒙我父赐福的，可来承受那创世以来为你们所预备的国。
MATT|25|35|因为我饿了，你们给我吃；渴了，你们给我喝；我流浪在外，你们留我住；
MATT|25|36|我赤身露体，你们给我穿；我病了，你们看顾我；我在监狱里，你们来看我。’
MATT|25|37|义人就回答：‘主啊，我们什么时候见你饿了，给你吃；渴了，给你喝？
MATT|25|38|什么时候见你流浪在外，留你住；或是赤身露体，给你穿？
MATT|25|39|又什么时候见你病了，或是在监狱里，来看你呢？’
MATT|25|40|王回答他们说：‘我实在告诉你们，这些事你们做在我弟兄中一个最小的身上，就是做在我身上了。’
MATT|25|41|“王又要向那左边的说：‘你们这被诅咒的人，离开我！进入那为魔鬼和他的使者所预备的永火里去！
MATT|25|42|因为我饿了，你们没有给我吃；渴了，你们没有给我喝；
MATT|25|43|我流浪在外，你们没有留我住；我赤身露体，你们没有给我穿；我病了，我在监狱里，你们没有来看顾我。’
MATT|25|44|他们也要回答：‘主啊，我们什么时候见你饿了，或渴了，或流浪在外，或赤身露体，或病了，或在监狱里，没有伺候你呢？’
MATT|25|45|王要回答：‘我实在告诉你们，这些事你们没有做在任何一个最小的弟兄身上，就是没有做在我身上了。’
MATT|25|46|这些人要往永刑里去；那些义人要往永生里去。”
MATT|26|1|耶稣说完了这一切的话，就对门徒说：
MATT|26|2|“你们知道，过两天是逾越节，人子将要被出卖，钉在十字架上。”
MATT|26|3|那时，祭司长和百姓的长老聚集在那称为 该亚法 的大祭司的院里。
MATT|26|4|大家商议要设计捉拿耶稣，把他杀掉。
MATT|26|5|可是他们说：“不可在过节的日子，恐怕百姓生乱。”
MATT|26|6|耶稣在 伯大尼 的痲疯病人 西门 家里，
MATT|26|7|有一个女人拿着一玉瓶极贵的香膏来，趁耶稣坐席的时候，浇在他的头上。
MATT|26|8|门徒看见就很不高兴，说：“何必这样浪费呢！
MATT|26|9|这香膏可以卖许多钱，周济穷人。”
MATT|26|10|耶稣看出他们的意思，就说：“为什么难为这女人呢？她在我身上做的是一件美事。
MATT|26|11|因为常有穷人和你们在一起，但是你们不常有我。
MATT|26|12|她把这香膏浇在我身上是为我安葬作准备的。
MATT|26|13|我实在告诉你们，普天之下，无论在什么地方传这福音，都要述说这女人所做的，来记念她。”
MATT|26|14|当时，十二使徒中有一个叫 加略 人 犹大 的，去见祭司长，
MATT|26|15|说：“我把他交给你们，你们愿意给我多少钱？”他们给了他三十块银钱。
MATT|26|16|从那时候起，他就找机会要把耶稣交给他们。
MATT|26|17|除酵节的第一天，门徒来问耶稣：“你要我们在哪里给你预备吃逾越节的宴席呢？”
MATT|26|18|耶稣说：“你们进城去，到某人那里，对他说：‘老师说：我的时候快到了，我要和我的门徒在你家里守逾越节。’”
MATT|26|19|门徒遵照耶稣所吩咐的去预备了逾越节的宴席。
MATT|26|20|到了晚上，耶稣和十二使徒坐席。
MATT|26|21|他们吃的时候，耶稣说：“我实在告诉你们，你们中间有一个人要出卖我。”
MATT|26|22|他们就非常忧愁，一个一个地问他：“主，该不是我吧？”
MATT|26|23|耶稣回答说：“同我蘸手在盘子里的，就是要出卖我的。
MATT|26|24|人子要去了，正如经上所写有关他的；但出卖人子的人有祸了！那人没有出生倒好。”
MATT|26|25|出卖耶稣的 犹大 回答他说：“拉比，该不是我吧？”耶稣说：“你自己说了。”
MATT|26|26|他们吃的时候，耶稣拿起饼来，祝福了，就擘开，递给门徒，说：“你们拿去，吃吧。这是我的身体。”
MATT|26|27|他又拿起杯来，祝谢了，递给他们，说：“你们都喝这个，
MATT|26|28|因为这是我立约的血，为许多人流出来，使罪得赦。
MATT|26|29|但我告诉你们，从今以后，我不再喝这葡萄汁，直到我在我父的国里与你们同喝新的那日子。”
MATT|26|30|他们唱了诗，就出来往 橄榄山 去。
MATT|26|31|那时，耶稣对他们说：“今夜，你们为我的缘故都要跌倒。因为经上记着： ‘我要击打牧人， 羊就分散了。’
MATT|26|32|但我复活以后，要在你们之前往 加利利 去。”
MATT|26|33|彼得 回答他说：“即使众人为你的缘故跌倒，我也绝不跌倒。”
MATT|26|34|耶稣说：“我实在告诉你，今夜鸡叫以前，你要三次不认我。”
MATT|26|35|彼得 说：“我就是必须和你同死，也绝不会不认你。”所有的门徒都是这样说。
MATT|26|36|耶稣和门徒来到一个地方，名叫 客西马尼 。他对他们说：“你们坐在这里，我到那边去祷告。”
MATT|26|37|于是他带着 彼得 和 西庇太 的两个儿子同去。他忧愁起来，极其难过，
MATT|26|38|就对他们说：“我心里非常忧伤，几乎要死；你们留在这里，和我一同警醒。”
MATT|26|39|他就稍往前走，俯伏在地，祷告说：“我父啊，如果可能，求你使这杯离开我。然而，不是照我所愿的，而是照你所愿的。”
MATT|26|40|他回到门徒那里，见他们睡着了，就对 彼得 说：“怎么样？你们不能同我警醒一小时吗？
MATT|26|41|总要警醒祷告，免得陷入试探。你们心灵固然愿意，肉体却软弱了。”
MATT|26|42|他第二次又去祷告说：“我父啊，这杯若不能离开我，必须我喝，就愿你的旨意成全。”
MATT|26|43|他又来，见他们睡着了，因为他们的眼睛困倦。
MATT|26|44|耶稣又离开他们，第三次去祷告，说的话跟先前一样。
MATT|26|45|然后他来到门徒那里，对他们说：“现在你们仍在睡觉安歇吗？看哪，时候到了，人子被出卖在罪人手里了。
MATT|26|46|起来，我们走吧！看哪，那出卖我的人快来了。”
MATT|26|47|耶稣还在说话的时候，十二使徒之一的 犹大 来了，还有一大群人带着刀棒，从祭司长和百姓的长老那里跟他同来。
MATT|26|48|那出卖耶稣的给了他们一个暗号，说：“我亲谁，谁就是。你们把他抓住。”
MATT|26|49|犹大 立刻进前来对耶稣说：“拉比，你好！”就跟他亲吻。
MATT|26|50|耶稣对他说：“朋友，你来要做的事，就做吧。 ”于是那些人上前，下手抓住耶稣。
MATT|26|51|忽然，有一个和耶稣一起的人伸手拔出刀来，把大祭司的仆人砍了一刀，削掉了他一只耳朵。
MATT|26|52|耶稣对他说：“收刀入鞘吧！凡动刀的，必死在刀下。
MATT|26|53|你想我不能求我父，现在为我差遣比十二营还多的天使来吗？
MATT|26|54|若是这样，经上所说事情必须如此发生的话怎么应验呢？”
MATT|26|55|就在那时，耶稣对众人说：“你们带着刀棒出来抓我，如同拿强盗吗？我天天坐在圣殿里教导人，你们并没有抓我。
MATT|26|56|但这整件事的发生，是要应验先知书上的话。”那时，门徒都离开他，逃走了。
MATT|26|57|抓耶稣的人把他带到大祭司 该亚法 那里去，文士和长老已经在那里聚集。
MATT|26|58|彼得 远远地跟着耶稣，直到大祭司的院子，进到里面，就和警卫同坐，要看结局怎样。
MATT|26|59|祭司长和全议会寻找假见证控告耶稣，要处死他。
MATT|26|60|虽然有好些人来作假见证，总找不到实据。最后有两个人前来，
MATT|26|61|说：“这个人曾说：‘我能拆毁上帝的殿，三日内又建造起来。’”
MATT|26|62|大祭司就站起来，对耶稣说：“这些人作证告你的事，你什么都不回答吗？”
MATT|26|63|耶稣却不言语。大祭司对他说：“我指着永生上帝命令你起誓告诉我们，你是不是基督—上帝的儿子？”
MATT|26|64|耶稣对他说：“你自己说了。然而，我告诉你们， 此后你们要看见人子 坐在权能者的右边， 驾着天上的云来临。”
MATT|26|65|大祭司就撕裂衣服，说：“他说了亵渎的话，我们何必再要证人呢？现在你们已经听见他这亵渎的话了。
MATT|26|66|你们的意见如何？”他们回答：“他该处死。”
MATT|26|67|他们就吐唾沫在他脸上，用拳头打他，也有打他耳光的，
MATT|26|68|说：“基督啊，向我们说预言吧！打你的是谁？”
MATT|26|69|彼得 在外面院子里坐着，有一个使女进前来，说：“你素来也是同那 加利利 人耶稣一起的。”
MATT|26|70|彼得 在众人面前却不承认，说：“我不知道你说的是什么！”
MATT|26|71|他出去，到了门口，又有一个使女看见他，就对那里的人说：“这个人是同 拿撒勒 人耶稣一起的。”
MATT|26|72|彼得 又不承认，起誓说：“我不认得那个人。”
MATT|26|73|过了不久，旁边站着的人前来，对 彼得 说：“你的确是他们一伙的，你的口音把你显露出来了。”
MATT|26|74|彼得 就赌咒发誓说：“我不认得那个人。”立刻鸡就叫了。
MATT|26|75|彼得 想起耶稣所说的话：“鸡叫以前，你要三次不认我。”他就出去痛哭。
MATT|27|1|到了早晨，众祭司长和百姓的长老商议要处死耶稣，
MATT|27|2|就把他绑着，解去，交给 彼拉多 总督。
MATT|27|3|这时，出卖耶稣的 犹大 看见耶稣已经定了罪，就后悔，把那三十块银钱拿回来给祭司长和长老，
MATT|27|4|说：“我出卖了无辜人的血有罪了。”他们说：“那跟我们有什么相干？你自己承当吧！”
MATT|27|5|犹大 就把那银钱丢在殿里，出去吊死了。
MATT|27|6|祭司长拾起银钱来，说：“这是血价，不可放在圣殿的银库里。”
MATT|27|7|他们商议，就用那银钱买了窑户的一块田，用来埋葬外乡人。
MATT|27|8|所以，那块田直到今日还叫做“血田”。
MATT|27|9|这就应验了先知 耶利米 所说的话：“他们用那三十块银钱，就是 以色列 人给那被估定的人所估定的价钱，
MATT|27|10|买了窑户的一块田；这是照着主所吩咐我的。”
MATT|27|11|耶稣站在总督面前，总督问他：“你是 犹太 人的王吗？”耶稣说：“是你说的。”
MATT|27|12|他被祭司长和长老控告的时候，什么都不回答。
MATT|27|13|彼拉多 就对他说：“他们作证告你这么多的事，你没有听见吗？”
MATT|27|14|耶稣仍不回答，连一句话也不说，以致总督觉得非常惊讶。
MATT|27|15|总督有一个常例，每逢这节期，随众人的意愿释放一个囚犯给他们。
MATT|27|16|当时有一个出名的囚犯叫 巴拉巴 。
MATT|27|17|众人聚集的时候， 彼拉多 就对他们说：“你们要我释放哪一个给你们？是 巴拉巴 呢？是称为基督的耶稣呢？”
MATT|27|18|总督原知道他们是因为嫉妒才把他解了来。
MATT|27|19|正坐堂的时候，他的夫人打发人来说：“这义人的事，你一点不可管，因为我今天在梦中因他受了许多的苦。”
MATT|27|20|祭司长和长老挑唆众人，要求释放 巴拉巴 ，除掉耶稣。
MATT|27|21|总督回答他们说：“这两个人，你们要我释放哪一个给你们呢？”他们说：“ 巴拉巴 。”
MATT|27|22|彼拉多 说：“这样，那称为基督的耶稣我怎么办他呢？”他们都说：“把他钉十字架！”
MATT|27|23|总督说：“为什么？他做了什么恶事呢？”他们更加喊着说：“把他钉十字架！”
MATT|27|24|彼拉多 见说也无济于事，反要生乱，就拿水在众人面前洗手，说：“流这人 的血，罪不在我，你们承当吧。”
MATT|27|25|众人都回答：“他的血归到我们和我们的子孙身上！”
MATT|27|26|于是 彼拉多 释放 巴拉巴 给他们，把耶稣鞭打后交给人钉十字架。
MATT|27|27|总督的兵把耶稣带进总督府，把全营的兵都聚集在耶稣那里。
MATT|27|28|他们脱了他的衣服，穿上一件朱红色的袍子，
MATT|27|29|用荆棘编了冠冕，戴在他头上，拿一根芦苇秆放在他右手里，跪在他面前，戏弄他，说：“万岁， 犹太 人的王！”
MATT|27|30|他们又向他吐唾沫，拿芦苇秆打他的头。
MATT|27|31|他们戏弄完了，就给他脱了袍子，又穿上他自己的衣服，带他出去，要钉十字架。
MATT|27|32|他们出去的时候，遇见一个 古利奈 人，名叫 西门 ，就强迫他同去，好背耶稣的十字架。
MATT|27|33|他们到了一个地方，名叫 各各他 ，就是“髑髅地”。
MATT|27|34|士兵拿苦胆调和的酒给耶稣喝。他尝了，不肯喝。
MATT|27|35|他们把他钉在十字架上，然后抽签分了他的衣服，
MATT|27|36|又坐在那里看守他。
MATT|27|37|他们在他头上方安了一个罪状牌，写着：“这是 犹太 人的王耶稣。”
MATT|27|38|当时，有两个强盗和他同钉十字架，一个在右边，一个在左边。
MATT|27|39|从那里经过的人讥笑他，摇着头，
MATT|27|40|说：“你这拆毁殿、三日又建造起来的，救救你自己吧！如果你是上帝的儿子，就从十字架上下来呀！”
MATT|27|41|众祭司长、文士和长老也同样嘲笑他，说：
MATT|27|42|“他救了别人，不能救自己。他是 以色列 的王，现在从十字架上下来，我们就信他。
MATT|27|43|他倚靠上帝，上帝若愿意，现在就来救他，因为他曾说‘我是上帝的儿子’。”
MATT|27|44|和他同钉的强盗也这样讥讽他。
MATT|27|45|从正午到下午三点钟，遍地都黑暗了。
MATT|27|46|约在下午三点钟，耶稣大声高呼，说：“以利！以利！拉马撒巴各大尼？”就是说：“我的上帝！我的上帝！为什么离弃我？”
MATT|27|47|站在那里的人，有的听见就说：“这个人呼叫 以利亚 呢！”
MATT|27|48|其中有一个人立刻跑去，拿海绵蘸满了醋，绑在芦苇秆上，送给他喝。
MATT|27|49|其余的人说：“且等着，看 以利亚 来不来救他。”
MATT|27|50|耶稣又大喊一声，气就断了。
MATT|27|51|忽然，殿的幔子从上到下裂为两半，地震动，磐石崩裂，
MATT|27|52|坟墓也开了，有许多已睡了的圣徒的身体也复活了。
MATT|27|53|耶稣复活以后，他们从坟墓里出来，进了圣城，向许多人显现。
MATT|27|54|百夫长和跟他一同看守耶稣的人看见地震和所经历的事，非常害怕，说：“他真是上帝的儿子！”
MATT|27|55|有好些妇女在那里，远远地观看，她们是从 加利利 跟随耶稣，来服事他的；
MATT|27|56|其中有 抹大拉 的 马利亚 ，又有 雅各 和 约瑟 的母亲 马利亚 ，并有 西庇太 两个儿子的母亲。
MATT|27|57|到了晚上，有一个财主，名叫 约瑟 ，是 亚利马太 来的，他也是耶稣的门徒。
MATT|27|58|这人去见 彼拉多 ，请求要耶稣的身体， 彼拉多 就吩咐给他。
MATT|27|59|约瑟 取了身体，用干净的细麻布裹好，
MATT|27|60|然后把他安放在自己的新墓穴里，就是他凿在岩石里的。他又把大石头滚到墓门口，然后离开。
MATT|27|61|有 抹大拉 的 马利亚 和另一个 马利亚 在那里，对着坟墓坐着。
MATT|27|62|次日，就是预备日的第二天，祭司长和法利赛人聚集来见 彼拉多 ，
MATT|27|63|说：“大人，我们记得那迷惑人的还活着的时候曾说：‘三天后我要复活。’
MATT|27|64|因此，请吩咐人将坟墓把守妥当，直到第三天，恐怕他的门徒来把他偷了去，就告诉百姓说：‘他从死人中复活了。’这样的话，那后来的迷惑就比先前的更厉害了。”
MATT|27|65|彼拉多 说：“你们有看守的兵，去吧！尽你们所能的把守妥当。”
MATT|27|66|他们就带着看守的兵同去，封了石头，将坟墓把守妥当。
MATT|28|1|安息日过后，七日的第一日，天快亮的时候， 抹大拉 的 马利亚 和另一个 马利亚 来看坟墓。
MATT|28|2|忽然，地大震动；因为有主的一个使者从天上下来，把石头滚开，坐在上面。
MATT|28|3|他的相貌如同闪电，衣服洁白如雪。
MATT|28|4|看守的人吓得浑身颤抖，甚至和死人一样。
MATT|28|5|天使回应妇女说：“不要害怕！我知道你们是寻找那钉十字架的耶稣。
MATT|28|6|他不在这里，照他所说的，他已经复活了。你们来！看看安放他的地方。
MATT|28|7|快去告诉他的门徒，说他已从死人中复活了，并且要比你们先到 加利利 去，在那里你们会看见他。看哪！我已经告诉你们了。”
MATT|28|8|妇女们急忙离开坟墓，又害怕，又大为欢喜，跑去告诉他的门徒。
MATT|28|9|忽然，耶稣迎上她们，说：“平安！”她们就上前抱住他的脚拜他。
MATT|28|10|耶稣对她们说：“不要害怕！你们去告诉我的弟兄，叫他们往 加利利 去，在那里会见到我。”
MATT|28|11|她们去的时候，看守的兵有几个进城去，把所发生的事都报告祭司长。
MATT|28|12|祭司长和长老聚集商议，就拿许多银钱给士兵，
MATT|28|13|说：“你们要这样说：‘夜间我们睡觉的时候，他的门徒来把他偷去了。’
MATT|28|14|若是这话被总督听见，有我们劝他，保你们无事。”
MATT|28|15|士兵收了银钱，就照所嘱咐他们的去做。这话就在 犹太 人中间流传，直到今日。
MATT|28|16|十一个门徒往 加利利 去，到了耶稣指定他们去的山上。
MATT|28|17|他们见了耶稣就拜他，然而还有人疑惑。
MATT|28|18|耶稣进前来，对他们说：“天上地下所有的权柄都赐给我了。
MATT|28|19|所以，你们要去，使万民作我的门徒，奉父、子、圣灵的名给他们施洗 ，
MATT|28|20|凡我所吩咐你们的，都教导他们遵守。看哪，我天天与你们同在，直到世代的终结。”
