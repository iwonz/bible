JOB|1|1|In the land of Uz there lived a man whose name was Job. This man was blameless and upright; he feared God and shunned evil.
JOB|1|2|He had seven sons and three daughters,
JOB|1|3|and he owned seven thousand sheep, three thousand camels, five hundred yoke of oxen and five hundred donkeys, and had a large number of servants. He was the greatest man among all the people of the East.
JOB|1|4|His sons used to take turns holding feasts in their homes, and they would invite their three sisters to eat and drink with them.
JOB|1|5|When a period of feasting had run its course, Job would send and have them purified. Early in the morning he would sacrifice a burnt offering for each of them, thinking, "Perhaps my children have sinned and cursed God in their hearts." This was Job's regular custom.
JOB|1|6|One day the angels came to present themselves before the LORD, and Satan also came with them.
JOB|1|7|The LORD said to Satan, "Where have you come from?" Satan answered the LORD, "From roaming through the earth and going back and forth in it."
JOB|1|8|Then the LORD said to Satan, "Have you considered my servant Job? There is no one on earth like him; he is blameless and upright, a man who fears God and shuns evil."
JOB|1|9|"Does Job fear God for nothing?" Satan replied.
JOB|1|10|"Have you not put a hedge around him and his household and everything he has? You have blessed the work of his hands, so that his flocks and herds are spread throughout the land.
JOB|1|11|But stretch out your hand and strike everything he has, and he will surely curse you to your face."
JOB|1|12|The LORD said to Satan, "Very well, then, everything he has is in your hands, but on the man himself do not lay a finger." Then Satan went out from the presence of the LORD.
JOB|1|13|One day when Job's sons and daughters were feasting and drinking wine at the oldest brother's house,
JOB|1|14|a messenger came to Job and said, "The oxen were plowing and the donkeys were grazing nearby,
JOB|1|15|and the Sabeans attacked and carried them off. They put the servants to the sword, and I am the only one who has escaped to tell you!"
JOB|1|16|While he was still speaking, another messenger came and said, "The fire of God fell from the sky and burned up the sheep and the servants, and I am the only one who has escaped to tell you!"
JOB|1|17|While he was still speaking, another messenger came and said, "The Chaldeans formed three raiding parties and swept down on your camels and carried them off. They put the servants to the sword, and I am the only one who has escaped to tell you!"
JOB|1|18|While he was still speaking, yet another messenger came and said, "Your sons and daughters were feasting and drinking wine at the oldest brother's house,
JOB|1|19|when suddenly a mighty wind swept in from the desert and struck the four corners of the house. It collapsed on them and they are dead, and I am the only one who has escaped to tell you!"
JOB|1|20|At this, Job got up and tore his robe and shaved his head. Then he fell to the ground in worship
JOB|1|21|and said: "Naked I came from my mother's womb, and naked I will depart. The LORD gave and the LORD has taken away; may the name of the LORD be praised."
JOB|1|22|In all this, Job did not sin by charging God with wrongdoing.
JOB|2|1|On another day the angels came to present themselves before the LORD, and Satan also came with them to present himself before him.
JOB|2|2|And the LORD said to Satan, "Where have you come from?" Satan answered the LORD, "From roaming through the earth and going back and forth in it."
JOB|2|3|Then the LORD said to Satan, "Have you considered my servant Job? There is no one on earth like him; he is blameless and upright, a man who fears God and shuns evil. And he still maintains his integrity, though you incited me against him to ruin him without any reason."
JOB|2|4|"Skin for skin!" Satan replied. "A man will give all he has for his own life.
JOB|2|5|But stretch out your hand and strike his flesh and bones, and he will surely curse you to your face."
JOB|2|6|The LORD said to Satan, "Very well, then, he is in your hands; but you must spare his life."
JOB|2|7|So Satan went out from the presence of the LORD and afflicted Job with painful sores from the soles of his feet to the top of his head.
JOB|2|8|Then Job took a piece of broken pottery and scraped himself with it as he sat among the ashes.
JOB|2|9|His wife said to him, "Are you still holding on to your integrity? Curse God and die!"
JOB|2|10|He replied, "You are talking like a foolish woman. Shall we accept good from God, and not trouble?" In all this, Job did not sin in what he said.
JOB|2|11|When Job's three friends, Eliphaz the Temanite, Bildad the Shuhite and Zophar the Naamathite, heard about all the troubles that had come upon him, they set out from their homes and met together by agreement to go and sympathize with him and comfort him.
JOB|2|12|When they saw him from a distance, they could hardly recognize him; they began to weep aloud, and they tore their robes and sprinkled dust on their heads.
JOB|2|13|Then they sat on the ground with him for seven days and seven nights. No one said a word to him, because they saw how great his suffering was.
JOB|3|1|After this, Job opened his mouth and cursed the day of his birth.
JOB|3|2|He said:
JOB|3|3|"May the day of my birth perish, and the night it was said, 'A boy is born!'
JOB|3|4|That day-may it turn to darkness; may God above not care about it; may no light shine upon it.
JOB|3|5|May darkness and deep shadow claim it once more; may a cloud settle over it; may blackness overwhelm its light.
JOB|3|6|That night-may thick darkness seize it; may it not be included among the days of the year nor be entered in any of the months.
JOB|3|7|May that night be barren; may no shout of joy be heard in it.
JOB|3|8|May those who curse days curse that day, those who are ready to rouse Leviathan.
JOB|3|9|May its morning stars become dark; may it wait for daylight in vain and not see the first rays of dawn,
JOB|3|10|for it did not shut the doors of the womb on me to hide trouble from my eyes.
JOB|3|11|"Why did I not perish at birth, and die as I came from the womb?
JOB|3|12|Why were there knees to receive me and breasts that I might be nursed?
JOB|3|13|For now I would be lying down in peace; I would be asleep and at rest
JOB|3|14|with kings and counselors of the earth, who built for themselves places now lying in ruins,
JOB|3|15|with rulers who had gold, who filled their houses with silver.
JOB|3|16|Or why was I not hidden in the ground like a stillborn child, like an infant who never saw the light of day?
JOB|3|17|There the wicked cease from turmoil, and there the weary are at rest.
JOB|3|18|Captives also enjoy their ease; they no longer hear the slave driver's shout.
JOB|3|19|The small and the great are there, and the slave is freed from his master.
JOB|3|20|"Why is light given to those in misery, and life to the bitter of soul,
JOB|3|21|to those who long for death that does not come, who search for it more than for hidden treasure,
JOB|3|22|who are filled with gladness and rejoice when they reach the grave?
JOB|3|23|Why is life given to a man whose way is hidden, whom God has hedged in?
JOB|3|24|For sighing comes to me instead of food; my groans pour out like water.
JOB|3|25|What I feared has come upon me; what I dreaded has happened to me.
JOB|3|26|I have no peace, no quietness; I have no rest, but only turmoil."
JOB|4|1|Then Eliphaz the Temanite replied:
JOB|4|2|"If someone ventures a word with you, will you be impatient? But who can keep from speaking?
JOB|4|3|Think how you have instructed many, how you have strengthened feeble hands.
JOB|4|4|Your words have supported those who stumbled; you have strengthened faltering knees.
JOB|4|5|But now trouble comes to you, and you are discouraged; it strikes you, and you are dismayed.
JOB|4|6|Should not your piety be your confidence and your blameless ways your hope?
JOB|4|7|"Consider now: Who, being innocent, has ever perished? Where were the upright ever destroyed?
JOB|4|8|As I have observed, those who plow evil and those who sow trouble reap it.
JOB|4|9|At the breath of God they are destroyed; at the blast of his anger they perish.
JOB|4|10|The lions may roar and growl, yet the teeth of the great lions are broken.
JOB|4|11|The lion perishes for lack of prey, and the cubs of the lioness are scattered.
JOB|4|12|"A word was secretly brought to me, my ears caught a whisper of it.
JOB|4|13|Amid disquieting dreams in the night, when deep sleep falls on men,
JOB|4|14|fear and trembling seized me and made all my bones shake.
JOB|4|15|A spirit glided past my face, and the hair on my body stood on end.
JOB|4|16|It stopped, but I could not tell what it was. A form stood before my eyes, and I heard a hushed voice:
JOB|4|17|'Can a mortal be more righteous than God? Can a man be more pure than his Maker?
JOB|4|18|If God places no trust in his servants, if he charges his angels with error,
JOB|4|19|how much more those who live in houses of clay, whose foundations are in the dust, who are crushed more readily than a moth!
JOB|4|20|Between dawn and dusk they are broken to pieces; unnoticed, they perish forever.
JOB|4|21|Are not the cords of their tent pulled up, so that they die without wisdom?'
JOB|5|1|"Call if you will, but who will answer you? To which of the holy ones will you turn?
JOB|5|2|Resentment kills a fool, and envy slays the simple.
JOB|5|3|I myself have seen a fool taking root, but suddenly his house was cursed.
JOB|5|4|His children are far from safety, crushed in court without a defender.
JOB|5|5|The hungry consume his harvest, taking it even from among thorns, and the thirsty pant after his wealth.
JOB|5|6|For hardship does not spring from the soil, nor does trouble sprout from the ground.
JOB|5|7|Yet man is born to trouble as surely as sparks fly upward.
JOB|5|8|"But if it were I, I would appeal to God; I would lay my cause before him.
JOB|5|9|He performs wonders that cannot be fathomed, miracles that cannot be counted.
JOB|5|10|He bestows rain on the earth; he sends water upon the countryside.
JOB|5|11|The lowly he sets on high, and those who mourn are lifted to safety.
JOB|5|12|He thwarts the plans of the crafty, so that their hands achieve no success.
JOB|5|13|He catches the wise in their craftiness, and the schemes of the wily are swept away.
JOB|5|14|Darkness comes upon them in the daytime; at noon they grope as in the night.
JOB|5|15|He saves the needy from the sword in their mouth; he saves them from the clutches of the powerful.
JOB|5|16|So the poor have hope, and injustice shuts its mouth.
JOB|5|17|"Blessed is the man whom God corrects; so do not despise the discipline of the Almighty.
JOB|5|18|For he wounds, but he also binds up; he injures, but his hands also heal.
JOB|5|19|From six calamities he will rescue you; in seven no harm will befall you.
JOB|5|20|In famine he will ransom you from death, and in battle from the stroke of the sword.
JOB|5|21|You will be protected from the lash of the tongue, and need not fear when destruction comes.
JOB|5|22|You will laugh at destruction and famine, and need not fear the beasts of the earth.
JOB|5|23|For you will have a covenant with the stones of the field, and the wild animals will be at peace with you.
JOB|5|24|You will know that your tent is secure; you will take stock of your property and find nothing missing.
JOB|5|25|You will know that your children will be many, and your descendants like the grass of the earth.
JOB|5|26|You will come to the grave in full vigor, like sheaves gathered in season.
JOB|5|27|"We have examined this, and it is true. So hear it and apply it to yourself."
JOB|6|1|Then Job replied:
JOB|6|2|"If only my anguish could be weighed and all my misery be placed on the scales!
JOB|6|3|It would surely outweigh the sand of the seas- no wonder my words have been impetuous.
JOB|6|4|The arrows of the Almighty are in me, my spirit drinks in their poison; God's terrors are marshaled against me.
JOB|6|5|Does a wild donkey bray when it has grass, or an ox bellow when it has fodder?
JOB|6|6|Is tasteless food eaten without salt, or is there flavor in the white of an egg?
JOB|6|7|I refuse to touch it; such food makes me ill.
JOB|6|8|"Oh, that I might have my request, that God would grant what I hope for,
JOB|6|9|that God would be willing to crush me, to let loose his hand and cut me off!
JOB|6|10|Then I would still have this consolation- my joy in unrelenting pain- that I had not denied the words of the Holy One.
JOB|6|11|"What strength do I have, that I should still hope? What prospects, that I should be patient?
JOB|6|12|Do I have the strength of stone? Is my flesh bronze?
JOB|6|13|Do I have any power to help myself, now that success has been driven from me?
JOB|6|14|"A despairing man should have the devotion of his friends, even though he forsakes the fear of the Almighty.
JOB|6|15|But my brothers are as undependable as intermittent streams, as the streams that overflow
JOB|6|16|when darkened by thawing ice and swollen with melting snow,
JOB|6|17|but that cease to flow in the dry season, and in the heat vanish from their channels.
JOB|6|18|Caravans turn aside from their routes; they go up into the wasteland and perish.
JOB|6|19|The caravans of Tema look for water, the traveling merchants of Sheba look in hope.
JOB|6|20|They are distressed, because they had been confident; they arrive there, only to be disappointed.
JOB|6|21|Now you too have proved to be of no help; you see something dreadful and are afraid.
JOB|6|22|Have I ever said, 'Give something on my behalf, pay a ransom for me from your wealth,
JOB|6|23|deliver me from the hand of the enemy, ransom me from the clutches of the ruthless'?
JOB|6|24|"Teach me, and I will be quiet; show me where I have been wrong.
JOB|6|25|How painful are honest words! But what do your arguments prove?
JOB|6|26|Do you mean to correct what I say, and treat the words of a despairing man as wind?
JOB|6|27|You would even cast lots for the fatherless and barter away your friend.
JOB|6|28|"But now be so kind as to look at me. Would I lie to your face?
JOB|6|29|Relent, do not be unjust; reconsider, for my integrity is at stake.
JOB|6|30|Is there any wickedness on my lips? Can my mouth not discern malice?
JOB|7|1|"Does not man have hard service on earth? Are not his days like those of a hired man?
JOB|7|2|Like a slave longing for the evening shadows, or a hired man waiting eagerly for his wages,
JOB|7|3|so I have been allotted months of futility, and nights of misery have been assigned to me.
JOB|7|4|When I lie down I think, 'How long before I get up?' The night drags on, and I toss till dawn.
JOB|7|5|My body is clothed with worms and scabs, my skin is broken and festering.
JOB|7|6|"My days are swifter than a weaver's shuttle, and they come to an end without hope.
JOB|7|7|Remember, O God, that my life is but a breath; my eyes will never see happiness again.
JOB|7|8|The eye that now sees me will see me no longer; you will look for me, but I will be no more.
JOB|7|9|As a cloud vanishes and is gone, so he who goes down to the grave does not return.
JOB|7|10|He will never come to his house again; his place will know him no more.
JOB|7|11|"Therefore I will not keep silent; I will speak out in the anguish of my spirit, I will complain in the bitterness of my soul.
JOB|7|12|Am I the sea, or the monster of the deep, that you put me under guard?
JOB|7|13|When I think my bed will comfort me and my couch will ease my complaint,
JOB|7|14|even then you frighten me with dreams and terrify me with visions,
JOB|7|15|so that I prefer strangling and death, rather than this body of mine.
JOB|7|16|I despise my life; I would not live forever. Let me alone; my days have no meaning.
JOB|7|17|"What is man that you make so much of him, that you give him so much attention,
JOB|7|18|that you examine him every morning and test him every moment?
JOB|7|19|Will you never look away from me, or let me alone even for an instant?
JOB|7|20|If I have sinned, what have I done to you, O watcher of men? Why have you made me your target? Have I become a burden to you?
JOB|7|21|Why do you not pardon my offenses and forgive my sins? For I will soon lie down in the dust; you will search for me, but I will be no more."
JOB|8|1|Then Bildad the Shuhite replied:
JOB|8|2|"How long will you say such things? Your words are a blustering wind.
JOB|8|3|Does God pervert justice? Does the Almighty pervert what is right?
JOB|8|4|When your children sinned against him, he gave them over to the penalty of their sin.
JOB|8|5|But if you will look to God and plead with the Almighty,
JOB|8|6|if you are pure and upright, even now he will rouse himself on your behalf and restore you to your rightful place.
JOB|8|7|Your beginnings will seem humble, so prosperous will your future be.
JOB|8|8|"Ask the former generations and find out what their fathers learned,
JOB|8|9|for we were born only yesterday and know nothing, and our days on earth are but a shadow.
JOB|8|10|Will they not instruct you and tell you? Will they not bring forth words from their understanding?
JOB|8|11|Can papyrus grow tall where there is no marsh? Can reeds thrive without water?
JOB|8|12|While still growing and uncut, they wither more quickly than grass.
JOB|8|13|Such is the destiny of all who forget God; so perishes the hope of the godless.
JOB|8|14|What he trusts in is fragile; what he relies on is a spider's web.
JOB|8|15|He leans on his web, but it gives way; he clings to it, but it does not hold.
JOB|8|16|He is like a well-watered plant in the sunshine, spreading its shoots over the garden;
JOB|8|17|it entwines its roots around a pile of rocks and looks for a place among the stones.
JOB|8|18|But when it is torn from its spot, that place disowns it and says, 'I never saw you.'
JOB|8|19|Surely its life withers away, and from the soil other plants grow.
JOB|8|20|"Surely God does not reject a blameless man or strengthen the hands of evildoers.
JOB|8|21|He will yet fill your mouth with laughter and your lips with shouts of joy.
JOB|8|22|Your enemies will be clothed in shame, and the tents of the wicked will be no more."
JOB|9|1|Then Job replied:
JOB|9|2|"Indeed, I know that this is true. But how can a mortal be righteous before God?
JOB|9|3|Though one wished to dispute with him, he could not answer him one time out of a thousand.
JOB|9|4|His wisdom is profound, his power is vast. Who has resisted him and come out unscathed?
JOB|9|5|He moves mountains without their knowing it and overturns them in his anger.
JOB|9|6|He shakes the earth from its place and makes its pillars tremble.
JOB|9|7|He speaks to the sun and it does not shine; he seals off the light of the stars.
JOB|9|8|He alone stretches out the heavens and treads on the waves of the sea.
JOB|9|9|He is the Maker of the Bear and Orion, the Pleiades and the constellations of the south.
JOB|9|10|He performs wonders that cannot be fathomed, miracles that cannot be counted.
JOB|9|11|When he passes me, I cannot see him; when he goes by, I cannot perceive him.
JOB|9|12|If he snatches away, who can stop him? Who can say to him, 'What are you doing?'
JOB|9|13|God does not restrain his anger; even the cohorts of Rahab cowered at his feet.
JOB|9|14|"How then can I dispute with him? How can I find words to argue with him?
JOB|9|15|Though I were innocent, I could not answer him; I could only plead with my Judge for mercy.
JOB|9|16|Even if I summoned him and he responded, I do not believe he would give me a hearing.
JOB|9|17|He would crush me with a storm and multiply my wounds for no reason.
JOB|9|18|He would not let me regain my breath but would overwhelm me with misery.
JOB|9|19|If it is a matter of strength, he is mighty! And if it is a matter of justice, who will summon him?
JOB|9|20|Even if I were innocent, my mouth would condemn me; if I were blameless, it would pronounce me guilty.
JOB|9|21|"Although I am blameless, I have no concern for myself; I despise my own life.
JOB|9|22|It is all the same; that is why I say, 'He destroys both the blameless and the wicked.'
JOB|9|23|When a scourge brings sudden death, he mocks the despair of the innocent.
JOB|9|24|When a land falls into the hands of the wicked, he blindfolds its judges. If it is not he, then who is it?
JOB|9|25|"My days are swifter than a runner; they fly away without a glimpse of joy.
JOB|9|26|They skim past like boats of papyrus, like eagles swooping down on their prey.
JOB|9|27|If I say, 'I will forget my complaint, I will change my expression, and smile,'
JOB|9|28|I still dread all my sufferings, for I know you will not hold me innocent.
JOB|9|29|Since I am already found guilty, why should I struggle in vain?
JOB|9|30|Even if I washed myself with soap and my hands with washing soda,
JOB|9|31|you would plunge me into a slime pit so that even my clothes would detest me.
JOB|9|32|"He is not a man like me that I might answer him, that we might confront each other in court.
JOB|9|33|If only there were someone to arbitrate between us, to lay his hand upon us both,
JOB|9|34|someone to remove God's rod from me, so that his terror would frighten me no more.
JOB|9|35|Then I would speak up without fear of him, but as it now stands with me, I cannot.
JOB|10|1|"I loathe my very life; therefore I will give free rein to my complaint and speak out in the bitterness of my soul.
JOB|10|2|I will say to God: Do not condemn me, but tell me what charges you have against me.
JOB|10|3|Does it please you to oppress me, to spurn the work of your hands, while you smile on the schemes of the wicked?
JOB|10|4|Do you have eyes of flesh? Do you see as a mortal sees?
JOB|10|5|Are your days like those of a mortal or your years like those of a man,
JOB|10|6|that you must search out my faults and probe after my sin-
JOB|10|7|though you know that I am not guilty and that no one can rescue me from your hand?
JOB|10|8|"Your hands shaped me and made me. Will you now turn and destroy me?
JOB|10|9|Remember that you molded me like clay. Will you now turn me to dust again?
JOB|10|10|Did you not pour me out like milk and curdle me like cheese,
JOB|10|11|clothe me with skin and flesh and knit me together with bones and sinews?
JOB|10|12|You gave me life and showed me kindness, and in your providence watched over my spirit.
JOB|10|13|"But this is what you concealed in your heart, and I know that this was in your mind:
JOB|10|14|If I sinned, you would be watching me and would not let my offense go unpunished.
JOB|10|15|If I am guilty-woe to me! Even if I am innocent, I cannot lift my head, for I am full of shame and drowned in my affliction.
JOB|10|16|If I hold my head high, you stalk me like a lion and again display your awesome power against me.
JOB|10|17|You bring new witnesses against me and increase your anger toward me; your forces come against me wave upon wave.
JOB|10|18|"Why then did you bring me out of the womb? I wish I had died before any eye saw me.
JOB|10|19|If only I had never come into being, or had been carried straight from the womb to the grave!
JOB|10|20|Are not my few days almost over? Turn away from me so I can have a moment's joy
JOB|10|21|before I go to the place of no return, to the land of gloom and deep shadow,
JOB|10|22|to the land of deepest night, of deep shadow and disorder, where even the light is like darkness."
JOB|11|1|Then Zophar the Naamathite replied:
JOB|11|2|"Are all these words to go unanswered? Is this talker to be vindicated?
JOB|11|3|Will your idle talk reduce men to silence? Will no one rebuke you when you mock?
JOB|11|4|You say to God, 'My beliefs are flawless and I am pure in your sight.'
JOB|11|5|Oh, how I wish that God would speak, that he would open his lips against you
JOB|11|6|and disclose to you the secrets of wisdom, for true wisdom has two sides. Know this: God has even forgotten some of your sin.
JOB|11|7|"Can you fathom the mysteries of God? Can you probe the limits of the Almighty?
JOB|11|8|They are higher than the heavens-what can you do? They are deeper than the depths of the grave -what can you know?
JOB|11|9|Their measure is longer than the earth and wider than the sea.
JOB|11|10|"If he comes along and confines you in prison and convenes a court, who can oppose him?
JOB|11|11|Surely he recognizes deceitful men; and when he sees evil, does he not take note?
JOB|11|12|But a witless man can no more become wise than a wild donkey's colt can be born a man.
JOB|11|13|"Yet if you devote your heart to him and stretch out your hands to him,
JOB|11|14|if you put away the sin that is in your hand and allow no evil to dwell in your tent,
JOB|11|15|then you will lift up your face without shame; you will stand firm and without fear.
JOB|11|16|You will surely forget your trouble, recalling it only as waters gone by.
JOB|11|17|Life will be brighter than noonday, and darkness will become like morning.
JOB|11|18|You will be secure, because there is hope; you will look about you and take your rest in safety.
JOB|11|19|You will lie down, with no one to make you afraid, and many will court your favor.
JOB|11|20|But the eyes of the wicked will fail, and escape will elude them; their hope will become a dying gasp."
JOB|12|1|Then Job replied:
JOB|12|2|"Doubtless you are the people, and wisdom will die with you!
JOB|12|3|But I have a mind as well as you; I am not inferior to you. Who does not know all these things?
JOB|12|4|"I have become a laughingstock to my friends, though I called upon God and he answered- a mere laughingstock, though righteous and blameless!
JOB|12|5|Men at ease have contempt for misfortune as the fate of those whose feet are slipping.
JOB|12|6|The tents of marauders are undisturbed, and those who provoke God are secure- those who carry their god in their hands.
JOB|12|7|"But ask the animals, and they will teach you, or the birds of the air, and they will tell you;
JOB|12|8|or speak to the earth, and it will teach you, or let the fish of the sea inform you.
JOB|12|9|Which of all these does not know that the hand of the LORD has done this?
JOB|12|10|In his hand is the life of every creature and the breath of all mankind.
JOB|12|11|Does not the ear test words as the tongue tastes food?
JOB|12|12|Is not wisdom found among the aged? Does not long life bring understanding?
JOB|12|13|"To God belong wisdom and power; counsel and understanding are his.
JOB|12|14|What he tears down cannot be rebuilt; the man he imprisons cannot be released.
JOB|12|15|If he holds back the waters, there is drought; if he lets them loose, they devastate the land.
JOB|12|16|To him belong strength and victory; both deceived and deceiver are his.
JOB|12|17|He leads counselors away stripped and makes fools of judges.
JOB|12|18|He takes off the shackles put on by kings and ties a loincloth around their waist.
JOB|12|19|He leads priests away stripped and overthrows men long established.
JOB|12|20|He silences the lips of trusted advisers and takes away the discernment of elders.
JOB|12|21|He pours contempt on nobles and disarms the mighty.
JOB|12|22|He reveals the deep things of darkness and brings deep shadows into the light.
JOB|12|23|He makes nations great, and destroys them; he enlarges nations, and disperses them.
JOB|12|24|He deprives the leaders of the earth of their reason; he sends them wandering through a trackless waste.
JOB|12|25|They grope in darkness with no light; he makes them stagger like drunkards.
JOB|13|1|"My eyes have seen all this, my ears have heard and understood it.
JOB|13|2|What you know, I also know; I am not inferior to you.
JOB|13|3|But I desire to speak to the Almighty and to argue my case with God.
JOB|13|4|You, however, smear me with lies; you are worthless physicians, all of you!
JOB|13|5|If only you would be altogether silent! For you, that would be wisdom.
JOB|13|6|Hear now my argument; listen to the plea of my lips.
JOB|13|7|Will you speak wickedly on God's behalf? Will you speak deceitfully for him?
JOB|13|8|Will you show him partiality? Will you argue the case for God?
JOB|13|9|Would it turn out well if he examined you? Could you deceive him as you might deceive men?
JOB|13|10|He would surely rebuke you if you secretly showed partiality.
JOB|13|11|Would not his splendor terrify you? Would not the dread of him fall on you?
JOB|13|12|Your maxims are proverbs of ashes; your defenses are defenses of clay.
JOB|13|13|"Keep silent and let me speak; then let come to me what may.
JOB|13|14|Why do I put myself in jeopardy and take my life in my hands?
JOB|13|15|Though he slay me, yet will I hope in him; I will surely defend my ways to his face.
JOB|13|16|Indeed, this will turn out for my deliverance, for no godless man would dare come before him!
JOB|13|17|Listen carefully to my words; let your ears take in what I say.
JOB|13|18|Now that I have prepared my case, I know I will be vindicated.
JOB|13|19|Can anyone bring charges against me? If so, I will be silent and die.
JOB|13|20|"Only grant me these two things, O God, and then I will not hide from you:
JOB|13|21|Withdraw your hand far from me, and stop frightening me with your terrors.
JOB|13|22|Then summon me and I will answer, or let me speak, and you reply.
JOB|13|23|How many wrongs and sins have I committed? Show me my offense and my sin.
JOB|13|24|Why do you hide your face and consider me your enemy?
JOB|13|25|Will you torment a windblown leaf? Will you chase after dry chaff?
JOB|13|26|For you write down bitter things against me and make me inherit the sins of my youth.
JOB|13|27|You fasten my feet in shackles; you keep close watch on all my paths by putting marks on the soles of my feet.
JOB|13|28|"So man wastes away like something rotten, like a garment eaten by moths.
JOB|14|1|"Man born of woman is of few days and full of trouble.
JOB|14|2|He springs up like a flower and withers away; like a fleeting shadow, he does not endure.
JOB|14|3|Do you fix your eye on such a one? Will you bring him before you for judgment?
JOB|14|4|Who can bring what is pure from the impure? No one!
JOB|14|5|Man's days are determined; you have decreed the number of his months and have set limits he cannot exceed.
JOB|14|6|So look away from him and let him alone, till he has put in his time like a hired man.
JOB|14|7|"At least there is hope for a tree: If it is cut down, it will sprout again, and its new shoots will not fail.
JOB|14|8|Its roots may grow old in the ground and its stump die in the soil,
JOB|14|9|yet at the scent of water it will bud and put forth shoots like a plant.
JOB|14|10|But man dies and is laid low; he breathes his last and is no more.
JOB|14|11|As water disappears from the sea or a riverbed becomes parched and dry,
JOB|14|12|so man lies down and does not rise; till the heavens are no more, men will not awake or be roused from their sleep.
JOB|14|13|"If only you would hide me in the grave and conceal me till your anger has passed! If only you would set me a time and then remember me!
JOB|14|14|If a man dies, will he live again? All the days of my hard service I will wait for my renewal to come.
JOB|14|15|You will call and I will answer you; you will long for the creature your hands have made.
JOB|14|16|Surely then you will count my steps but not keep track of my sin.
JOB|14|17|My offenses will be sealed up in a bag; you will cover over my sin.
JOB|14|18|"But as a mountain erodes and crumbles and as a rock is moved from its place,
JOB|14|19|as water wears away stones and torrents wash away the soil, so you destroy man's hope.
JOB|14|20|You overpower him once for all, and he is gone; you change his countenance and send him away.
JOB|14|21|If his sons are honored, he does not know it; if they are brought low, he does not see it.
JOB|14|22|He feels but the pain of his own body and mourns only for himself."
JOB|15|1|Then Eliphaz the Temanite replied:
JOB|15|2|"Would a wise man answer with empty notions or fill his belly with the hot east wind?
JOB|15|3|Would he argue with useless words, with speeches that have no value?
JOB|15|4|But you even undermine piety and hinder devotion to God.
JOB|15|5|Your sin prompts your mouth; you adopt the tongue of the crafty.
JOB|15|6|Your own mouth condemns you, not mine; your own lips testify against you.
JOB|15|7|"Are you the first man ever born? Were you brought forth before the hills?
JOB|15|8|Do you listen in on God's council? Do you limit wisdom to yourself?
JOB|15|9|What do you know that we do not know? What insights do you have that we do not have?
JOB|15|10|The gray-haired and the aged are on our side, men even older than your father.
JOB|15|11|Are God's consolations not enough for you, words spoken gently to you?
JOB|15|12|Why has your heart carried you away, and why do your eyes flash,
JOB|15|13|so that you vent your rage against God and pour out such words from your mouth?
JOB|15|14|"What is man, that he could be pure, or one born of woman, that he could be righteous?
JOB|15|15|If God places no trust in his holy ones, if even the heavens are not pure in his eyes,
JOB|15|16|how much less man, who is vile and corrupt, who drinks up evil like water!
JOB|15|17|"Listen to me and I will explain to you; let me tell you what I have seen,
JOB|15|18|what wise men have declared, hiding nothing received from their fathers
JOB|15|19|(to whom alone the land was given when no alien passed among them):
JOB|15|20|All his days the wicked man suffers torment, the ruthless through all the years stored up for him.
JOB|15|21|Terrifying sounds fill his ears; when all seems well, marauders attack him.
JOB|15|22|He despairs of escaping the darkness; he is marked for the sword.
JOB|15|23|He wanders about-food for vultures; he knows the day of darkness is at hand.
JOB|15|24|Distress and anguish fill him with terror; they overwhelm him, like a king poised to attack,
JOB|15|25|because he shakes his fist at God and vaunts himself against the Almighty,
JOB|15|26|defiantly charging against him with a thick, strong shield.
JOB|15|27|"Though his face is covered with fat and his waist bulges with flesh,
JOB|15|28|he will inhabit ruined towns and houses where no one lives, houses crumbling to rubble.
JOB|15|29|He will no longer be rich and his wealth will not endure, nor will his possessions spread over the land.
JOB|15|30|He will not escape the darkness; a flame will wither his shoots, and the breath of God's mouth will carry him away.
JOB|15|31|Let him not deceive himself by trusting what is worthless, for he will get nothing in return.
JOB|15|32|Before his time he will be paid in full, and his branches will not flourish.
JOB|15|33|He will be like a vine stripped of its unripe grapes, like an olive tree shedding its blossoms.
JOB|15|34|For the company of the godless will be barren, and fire will consume the tents of those who love bribes.
JOB|15|35|They conceive trouble and give birth to evil; their womb fashions deceit."
JOB|16|1|Then Job replied:
JOB|16|2|"I have heard many things like these; miserable comforters are you all!
JOB|16|3|Will your long-winded speeches never end? What ails you that you keep on arguing?
JOB|16|4|I also could speak like you, if you were in my place; I could make fine speeches against you and shake my head at you.
JOB|16|5|But my mouth would encourage you; comfort from my lips would bring you relief.
JOB|16|6|"Yet if I speak, my pain is not relieved; and if I refrain, it does not go away.
JOB|16|7|Surely, O God, you have worn me out; you have devastated my entire household.
JOB|16|8|You have bound me-and it has become a witness; my gauntness rises up and testifies against me.
JOB|16|9|God assails me and tears me in his anger and gnashes his teeth at me; my opponent fastens on me his piercing eyes.
JOB|16|10|Men open their mouths to jeer at me; they strike my cheek in scorn and unite together against me.
JOB|16|11|God has turned me over to evil men and thrown me into the clutches of the wicked.
JOB|16|12|All was well with me, but he shattered me; he seized me by the neck and crushed me. He has made me his target;
JOB|16|13|his archers surround me. Without pity, he pierces my kidneys and spills my gall on the ground.
JOB|16|14|Again and again he bursts upon me; he rushes at me like a warrior.
JOB|16|15|"I have sewed sackcloth over my skin and buried my brow in the dust.
JOB|16|16|My face is red with weeping, deep shadows ring my eyes;
JOB|16|17|yet my hands have been free of violence and my prayer is pure.
JOB|16|18|"O earth, do not cover my blood; may my cry never be laid to rest!
JOB|16|19|Even now my witness is in heaven; my advocate is on high.
JOB|16|20|My intercessor is my friend as my eyes pour out tears to God;
JOB|16|21|on behalf of a man he pleads with God as a man pleads for his friend.
JOB|16|22|"Only a few years will pass before I go on the journey of no return.
JOB|17|1|My spirit is broken, my days are cut short, the grave awaits me.
JOB|17|2|Surely mockers surround me; my eyes must dwell on their hostility.
JOB|17|3|"Give me, O God, the pledge you demand. Who else will put up security for me?
JOB|17|4|You have closed their minds to understanding; therefore you will not let them triumph.
JOB|17|5|If a man denounces his friends for reward, the eyes of his children will fail.
JOB|17|6|"God has made me a byword to everyone, a man in whose face people spit.
JOB|17|7|My eyes have grown dim with grief; my whole frame is but a shadow.
JOB|17|8|Upright men are appalled at this; the innocent are aroused against the ungodly.
JOB|17|9|Nevertheless, the righteous will hold to their ways, and those with clean hands will grow stronger.
JOB|17|10|"But come on, all of you, try again! I will not find a wise man among you.
JOB|17|11|My days have passed, my plans are shattered, and so are the desires of my heart.
JOB|17|12|These men turn night into day; in the face of darkness they say, 'Light is near.'
JOB|17|13|If the only home I hope for is the grave, if I spread out my bed in darkness,
JOB|17|14|if I say to corruption, 'You are my father,' and to the worm, 'My mother' or 'My sister,'
JOB|17|15|where then is my hope? Who can see any hope for me?
JOB|17|16|Will it go down to the gates of death? Will we descend together into the dust?"
JOB|18|1|Then Bildad the Shuhite replied:
JOB|18|2|"When will you end these speeches? Be sensible, and then we can talk.
JOB|18|3|Why are we regarded as cattle and considered stupid in your sight?
JOB|18|4|You who tear yourself to pieces in your anger, is the earth to be abandoned for your sake? Or must the rocks be moved from their place?
JOB|18|5|"The lamp of the wicked is snuffed out; the flame of his fire stops burning.
JOB|18|6|The light in his tent becomes dark; the lamp beside him goes out.
JOB|18|7|The vigor of his step is weakened; his own schemes throw him down.
JOB|18|8|His feet thrust him into a net and he wanders into its mesh.
JOB|18|9|A trap seizes him by the heel; a snare holds him fast.
JOB|18|10|A noose is hidden for him on the ground; a trap lies in his path.
JOB|18|11|Terrors startle him on every side and dog his every step.
JOB|18|12|Calamity is hungry for him; disaster is ready for him when he falls.
JOB|18|13|It eats away parts of his skin; death's firstborn devours his limbs.
JOB|18|14|He is torn from the security of his tent and marched off to the king of terrors.
JOB|18|15|Fire resides in his tent; burning sulfur is scattered over his dwelling.
JOB|18|16|His roots dry up below and his branches wither above.
JOB|18|17|The memory of him perishes from the earth; he has no name in the land.
JOB|18|18|He is driven from light into darkness and is banished from the world.
JOB|18|19|He has no offspring or descendants among his people, no survivor where once he lived.
JOB|18|20|Men of the west are appalled at his fate; men of the east are seized with horror.
JOB|18|21|Surely such is the dwelling of an evil man; such is the place of one who knows not God."
JOB|19|1|Then Job replied:
JOB|19|2|"How long will you torment me and crush me with words?
JOB|19|3|Ten times now you have reproached me; shamelessly you attack me.
JOB|19|4|If it is true that I have gone astray, my error remains my concern alone.
JOB|19|5|If indeed you would exalt yourselves above me and use my humiliation against me,
JOB|19|6|then know that God has wronged me and drawn his net around me.
JOB|19|7|"Though I cry, 'I've been wronged!' I get no response; though I call for help, there is no justice.
JOB|19|8|He has blocked my way so I cannot pass; he has shrouded my paths in darkness.
JOB|19|9|He has stripped me of my honor and removed the crown from my head.
JOB|19|10|He tears me down on every side till I am gone; he uproots my hope like a tree.
JOB|19|11|His anger burns against me; he counts me among his enemies.
JOB|19|12|His troops advance in force; they build a siege ramp against me and encamp around my tent.
JOB|19|13|"He has alienated my brothers from me; my acquaintances are completely estranged from me.
JOB|19|14|My kinsmen have gone away; my friends have forgotten me.
JOB|19|15|My guests and my maidservants count me a stranger; they look upon me as an alien.
JOB|19|16|I summon my servant, but he does not answer, though I beg him with my own mouth.
JOB|19|17|My breath is offensive to my wife; I am loathsome to my own brothers.
JOB|19|18|Even the little boys scorn me; when I appear, they ridicule me.
JOB|19|19|All my intimate friends detest me; those I love have turned against me.
JOB|19|20|I am nothing but skin and bones; I have escaped with only the skin of my teeth.
JOB|19|21|"Have pity on me, my friends, have pity, for the hand of God has struck me.
JOB|19|22|Why do you pursue me as God does? Will you never get enough of my flesh?
JOB|19|23|"Oh, that my words were recorded, that they were written on a scroll,
JOB|19|24|that they were inscribed with an iron tool on lead, or engraved in rock forever!
JOB|19|25|I know that my Redeemer lives, and that in the end he will stand upon the earth.
JOB|19|26|And after my skin has been destroyed, yet in my flesh I will see God;
JOB|19|27|I myself will see him with my own eyes-I, and not another. How my heart yearns within me!
JOB|19|28|"If you say, 'How we will hound him, since the root of the trouble lies in him, '
JOB|19|29|you should fear the sword yourselves; for wrath will bring punishment by the sword, and then you will know that there is judgment. "
JOB|20|1|Then Zophar the Naamathite replied:
JOB|20|2|"My troubled thoughts prompt me to answer because I am greatly disturbed.
JOB|20|3|I hear a rebuke that dishonors me, and my understanding inspires me to reply.
JOB|20|4|"Surely you know how it has been from of old, ever since man was placed on the earth,
JOB|20|5|that the mirth of the wicked is brief, the joy of the godless lasts but a moment.
JOB|20|6|Though his pride reaches to the heavens and his head touches the clouds,
JOB|20|7|he will perish forever, like his own dung; those who have seen him will say, 'Where is he?'
JOB|20|8|Like a dream he flies away, no more to be found, banished like a vision of the night.
JOB|20|9|The eye that saw him will not see him again; his place will look on him no more.
JOB|20|10|His children must make amends to the poor; his own hands must give back his wealth.
JOB|20|11|The youthful vigor that fills his bones will lie with him in the dust.
JOB|20|12|"Though evil is sweet in his mouth and he hides it under his tongue,
JOB|20|13|though he cannot bear to let it go and keeps it in his mouth,
JOB|20|14|yet his food will turn sour in his stomach; it will become the venom of serpents within him.
JOB|20|15|He will spit out the riches he swallowed; God will make his stomach vomit them up.
JOB|20|16|He will suck the poison of serpents; the fangs of an adder will kill him.
JOB|20|17|He will not enjoy the streams, the rivers flowing with honey and cream.
JOB|20|18|What he toiled for he must give back uneaten; he will not enjoy the profit from his trading.
JOB|20|19|For he has oppressed the poor and left them destitute; he has seized houses he did not build.
JOB|20|20|"Surely he will have no respite from his craving; he cannot save himself by his treasure.
JOB|20|21|Nothing is left for him to devour; his prosperity will not endure.
JOB|20|22|In the midst of his plenty, distress will overtake him; the full force of misery will come upon him.
JOB|20|23|When he has filled his belly, God will vent his burning anger against him and rain down his blows upon him.
JOB|20|24|Though he flees from an iron weapon, a bronze-tipped arrow pierces him.
JOB|20|25|He pulls it out of his back, the gleaming point out of his liver. Terrors will come over him;
JOB|20|26|total darkness lies in wait for his treasures. A fire unfanned will consume him and devour what is left in his tent.
JOB|20|27|The heavens will expose his guilt; the earth will rise up against him.
JOB|20|28|A flood will carry off his house, rushing waters on the day of God's wrath.
JOB|20|29|Such is the fate God allots the wicked, the heritage appointed for them by God."
JOB|21|1|Then Job replied:
JOB|21|2|"Listen carefully to my words; let this be the consolation you give me.
JOB|21|3|Bear with me while I speak, and after I have spoken, mock on.
JOB|21|4|"Is my complaint directed to man? Why should I not be impatient?
JOB|21|5|Look at me and be astonished; clap your hand over your mouth.
JOB|21|6|When I think about this, I am terrified; trembling seizes my body.
JOB|21|7|Why do the wicked live on, growing old and increasing in power?
JOB|21|8|They see their children established around them, their offspring before their eyes.
JOB|21|9|Their homes are safe and free from fear; the rod of God is not upon them.
JOB|21|10|Their bulls never fail to breed; their cows calve and do not miscarry.
JOB|21|11|They send forth their children as a flock; their little ones dance about.
JOB|21|12|They sing to the music of tambourine and harp; they make merry to the sound of the flute.
JOB|21|13|They spend their years in prosperity and go down to the grave in peace.
JOB|21|14|Yet they say to God, 'Leave us alone! We have no desire to know your ways.
JOB|21|15|Who is the Almighty, that we should serve him? What would we gain by praying to him?'
JOB|21|16|But their prosperity is not in their own hands, so I stand aloof from the counsel of the wicked.
JOB|21|17|"Yet how often is the lamp of the wicked snuffed out? How often does calamity come upon them, the fate God allots in his anger?
JOB|21|18|How often are they like straw before the wind, like chaff swept away by a gale?
JOB|21|19|It is said, 'God stores up a man's punishment for his sons.' Let him repay the man himself, so that he will know it!
JOB|21|20|Let his own eyes see his destruction; let him drink of the wrath of the Almighty.
JOB|21|21|For what does he care about the family he leaves behind when his allotted months come to an end?
JOB|21|22|"Can anyone teach knowledge to God, since he judges even the highest?
JOB|21|23|One man dies in full vigor, completely secure and at ease,
JOB|21|24|his body well nourished, his bones rich with marrow.
JOB|21|25|Another man dies in bitterness of soul, never having enjoyed anything good.
JOB|21|26|Side by side they lie in the dust, and worms cover them both.
JOB|21|27|"I know full well what you are thinking, the schemes by which you would wrong me.
JOB|21|28|You say, 'Where now is the great man's house, the tents where wicked men lived?'
JOB|21|29|Have you never questioned those who travel? Have you paid no regard to their accounts-
JOB|21|30|that the evil man is spared from the day of calamity, that he is delivered from the day of wrath?
JOB|21|31|Who denounces his conduct to his face? Who repays him for what he has done?
JOB|21|32|He is carried to the grave, and watch is kept over his tomb.
JOB|21|33|The soil in the valley is sweet to him; all men follow after him, and a countless throng goes before him.
JOB|21|34|"So how can you console me with your nonsense? Nothing is left of your answers but falsehood!"
JOB|22|1|Then Eliphaz the Temanite replied:
JOB|22|2|"Can a man be of benefit to God? Can even a wise man benefit him?
JOB|22|3|What pleasure would it give the Almighty if you were righteous? What would he gain if your ways were blameless?
JOB|22|4|"Is it for your piety that he rebukes you and brings charges against you?
JOB|22|5|Is not your wickedness great? Are not your sins endless?
JOB|22|6|You demanded security from your brothers for no reason; you stripped men of their clothing, leaving them naked.
JOB|22|7|You gave no water to the weary and you withheld food from the hungry,
JOB|22|8|though you were a powerful man, owning land- an honored man, living on it.
JOB|22|9|And you sent widows away empty-handed and broke the strength of the fatherless.
JOB|22|10|That is why snares are all around you, why sudden peril terrifies you,
JOB|22|11|why it is so dark you cannot see, and why a flood of water covers you.
JOB|22|12|"Is not God in the heights of heaven? And see how lofty are the highest stars!
JOB|22|13|Yet you say, 'What does God know? Does he judge through such darkness?
JOB|22|14|Thick clouds veil him, so he does not see us as he goes about in the vaulted heavens.'
JOB|22|15|Will you keep to the old path that evil men have trod?
JOB|22|16|They were carried off before their time, their foundations washed away by a flood.
JOB|22|17|They said to God, 'Leave us alone! What can the Almighty do to us?'
JOB|22|18|Yet it was he who filled their houses with good things, so I stand aloof from the counsel of the wicked.
JOB|22|19|"The righteous see their ruin and rejoice; the innocent mock them, saying,
JOB|22|20|'Surely our foes are destroyed, and fire devours their wealth.'
JOB|22|21|"Submit to God and be at peace with him; in this way prosperity will come to you.
JOB|22|22|Accept instruction from his mouth and lay up his words in your heart.
JOB|22|23|If you return to the Almighty, you will be restored: If you remove wickedness far from your tent
JOB|22|24|and assign your nuggets to the dust, your gold of Ophir to the rocks in the ravines,
JOB|22|25|then the Almighty will be your gold, the choicest silver for you.
JOB|22|26|Surely then you will find delight in the Almighty and will lift up your face to God.
JOB|22|27|You will pray to him, and he will hear you, and you will fulfill your vows.
JOB|22|28|What you decide on will be done, and light will shine on your ways.
JOB|22|29|When men are brought low and you say, 'Lift them up!' then he will save the downcast.
JOB|22|30|He will deliver even one who is not innocent, who will be delivered through the cleanness of your hands."
JOB|23|1|Then Job replied:
JOB|23|2|"Even today my complaint is bitter; his hand is heavy in spite of my groaning.
JOB|23|3|If only I knew where to find him; if only I could go to his dwelling!
JOB|23|4|I would state my case before him and fill my mouth with arguments.
JOB|23|5|I would find out what he would answer me, and consider what he would say.
JOB|23|6|Would he oppose me with great power? No, he would not press charges against me.
JOB|23|7|There an upright man could present his case before him, and I would be delivered forever from my judge.
JOB|23|8|"But if I go to the east, he is not there; if I go to the west, I do not find him.
JOB|23|9|When he is at work in the north, I do not see him; when he turns to the south, I catch no glimpse of him.
JOB|23|10|But he knows the way that I take; when he has tested me, I will come forth as gold.
JOB|23|11|My feet have closely followed his steps; I have kept to his way without turning aside.
JOB|23|12|I have not departed from the commands of his lips; I have treasured the words of his mouth more than my daily bread.
JOB|23|13|"But he stands alone, and who can oppose him? He does whatever he pleases.
JOB|23|14|He carries out his decree against me, and many such plans he still has in store.
JOB|23|15|That is why I am terrified before him; when I think of all this, I fear him.
JOB|23|16|God has made my heart faint; the Almighty has terrified me.
JOB|23|17|Yet I am not silenced by the darkness, by the thick darkness that covers my face.
JOB|24|1|"Why does the Almighty not set times for judgment? Why must those who know him look in vain for such days?
JOB|24|2|Men move boundary stones; they pasture flocks they have stolen.
JOB|24|3|They drive away the orphan's donkey and take the widow's ox in pledge.
JOB|24|4|They thrust the needy from the path and force all the poor of the land into hiding.
JOB|24|5|Like wild donkeys in the desert, the poor go about their labor of foraging food; the wasteland provides food for their children.
JOB|24|6|They gather fodder in the fields and glean in the vineyards of the wicked.
JOB|24|7|Lacking clothes, they spend the night naked; they have nothing to cover themselves in the cold.
JOB|24|8|They are drenched by mountain rains and hug the rocks for lack of shelter.
JOB|24|9|The fatherless child is snatched from the breast; the infant of the poor is seized for a debt.
JOB|24|10|Lacking clothes, they go about naked; they carry the sheaves, but still go hungry.
JOB|24|11|They crush olives among the terraces; they tread the winepresses, yet suffer thirst.
JOB|24|12|The groans of the dying rise from the city, and the souls of the wounded cry out for help. But God charges no one with wrongdoing.
JOB|24|13|"There are those who rebel against the light, who do not know its ways or stay in its paths.
JOB|24|14|When daylight is gone, the murderer rises up and kills the poor and needy; in the night he steals forth like a thief.
JOB|24|15|The eye of the adulterer watches for dusk; he thinks, 'No eye will see me,' and he keeps his face concealed.
JOB|24|16|In the dark, men break into houses, but by day they shut themselves in; they want nothing to do with the light.
JOB|24|17|For all of them, deep darkness is their morning; they make friends with the terrors of darkness.
JOB|24|18|"Yet they are foam on the surface of the water; their portion of the land is cursed, so that no one goes to the vineyards.
JOB|24|19|As heat and drought snatch away the melted snow, so the grave snatches away those who have sinned.
JOB|24|20|The womb forgets them, the worm feasts on them; evil men are no longer remembered but are broken like a tree.
JOB|24|21|They prey on the barren and childless woman, and to the widow show no kindness.
JOB|24|22|But God drags away the mighty by his power; though they become established, they have no assurance of life.
JOB|24|23|He may let them rest in a feeling of security, but his eyes are on their ways.
JOB|24|24|For a little while they are exalted, and then they are gone; they are brought low and gathered up like all others; they are cut off like heads of grain.
JOB|24|25|"If this is not so, who can prove me false and reduce my words to nothing?"
JOB|25|1|Then Bildad the Shuhite replied:
JOB|25|2|"Dominion and awe belong to God; he establishes order in the heights of heaven.
JOB|25|3|Can his forces be numbered? Upon whom does his light not rise?
JOB|25|4|How then can a man be righteous before God? How can one born of woman be pure?
JOB|25|5|If even the moon is not bright and the stars are not pure in his eyes,
JOB|25|6|how much less man, who is but a maggot- a son of man, who is only a worm!"
JOB|26|1|Then Job replied:
JOB|26|2|"How you have helped the powerless! How you have saved the arm that is feeble!
JOB|26|3|What advice you have offered to one without wisdom! And what great insight you have displayed!
JOB|26|4|Who has helped you utter these words? And whose spirit spoke from your mouth?
JOB|26|5|"The dead are in deep anguish, those beneath the waters and all that live in them.
JOB|26|6|Death is naked before God; Destruction lies uncovered.
JOB|26|7|He spreads out the northern skies over empty space; he suspends the earth over nothing.
JOB|26|8|He wraps up the waters in his clouds, yet the clouds do not burst under their weight.
JOB|26|9|He covers the face of the full moon, spreading his clouds over it.
JOB|26|10|He marks out the horizon on the face of the waters for a boundary between light and darkness.
JOB|26|11|The pillars of the heavens quake, aghast at his rebuke.
JOB|26|12|By his power he churned up the sea; by his wisdom he cut Rahab to pieces.
JOB|26|13|By his breath the skies became fair; his hand pierced the gliding serpent.
JOB|26|14|And these are but the outer fringe of his works; how faint the whisper we hear of him! Who then can understand the thunder of his power?"
JOB|27|1|And Job continued his discourse:
JOB|27|2|"As surely as God lives, who has denied me justice, the Almighty, who has made me taste bitterness of soul,
JOB|27|3|as long as I have life within me, the breath of God in my nostrils,
JOB|27|4|my lips will not speak wickedness, and my tongue will utter no deceit.
JOB|27|5|I will never admit you are in the right; till I die, I will not deny my integrity.
JOB|27|6|I will maintain my righteousness and never let go of it; my conscience will not reproach me as long as I live.
JOB|27|7|"May my enemies be like the wicked, my adversaries like the unjust!
JOB|27|8|For what hope has the godless when he is cut off, when God takes away his life?
JOB|27|9|Does God listen to his cry when distress comes upon him?
JOB|27|10|Will he find delight in the Almighty? Will he call upon God at all times?
JOB|27|11|"I will teach you about the power of God; the ways of the Almighty I will not conceal.
JOB|27|12|You have all seen this yourselves. Why then this meaningless talk?
JOB|27|13|"Here is the fate God allots to the wicked, the heritage a ruthless man receives from the Almighty:
JOB|27|14|However many his children, their fate is the sword; his offspring will never have enough to eat.
JOB|27|15|The plague will bury those who survive him, and their widows will not weep for them.
JOB|27|16|Though he heaps up silver like dust and clothes like piles of clay,
JOB|27|17|what he lays up the righteous will wear, and the innocent will divide his silver.
JOB|27|18|The house he builds is like a moth's cocoon, like a hut made by a watchman.
JOB|27|19|He lies down wealthy, but will do so no more; when he opens his eyes, all is gone.
JOB|27|20|Terrors overtake him like a flood; a tempest snatches him away in the night.
JOB|27|21|The east wind carries him off, and he is gone; it sweeps him out of his place.
JOB|27|22|It hurls itself against him without mercy as he flees headlong from its power.
JOB|27|23|It claps its hands in derision and hisses him out of his place.
JOB|28|1|"There is a mine for silver and a place where gold is refined.
JOB|28|2|Iron is taken from the earth, and copper is smelted from ore.
JOB|28|3|Man puts an end to the darkness; he searches the farthest recesses for ore in the blackest darkness.
JOB|28|4|Far from where people dwell he cuts a shaft, in places forgotten by the foot of man; far from men he dangles and sways.
JOB|28|5|The earth, from which food comes, is transformed below as by fire;
JOB|28|6|sapphires come from its rocks, and its dust contains nuggets of gold.
JOB|28|7|No bird of prey knows that hidden path, no falcon's eye has seen it.
JOB|28|8|Proud beasts do not set foot on it, and no lion prowls there.
JOB|28|9|Man's hand assaults the flinty rock and lays bare the roots of the mountains.
JOB|28|10|He tunnels through the rock; his eyes see all its treasures.
JOB|28|11|He searches the sources of the rivers and brings hidden things to light.
JOB|28|12|"But where can wisdom be found? Where does understanding dwell?
JOB|28|13|Man does not comprehend its worth; it cannot be found in the land of the living.
JOB|28|14|The deep says, 'It is not in me'; the sea says, 'It is not with me.'
JOB|28|15|It cannot be bought with the finest gold, nor can its price be weighed in silver.
JOB|28|16|It cannot be bought with the gold of Ophir, with precious onyx or sapphires.
JOB|28|17|Neither gold nor crystal can compare with it, nor can it be had for jewels of gold.
JOB|28|18|Coral and jasper are not worthy of mention; the price of wisdom is beyond rubies.
JOB|28|19|The topaz of Cush cannot compare with it; it cannot be bought with pure gold.
JOB|28|20|"Where then does wisdom come from? Where does understanding dwell?
JOB|28|21|It is hidden from the eyes of every living thing, concealed even from the birds of the air.
JOB|28|22|Destruction and Death say, 'Only a rumor of it has reached our ears.'
JOB|28|23|God understands the way to it and he alone knows where it dwells,
JOB|28|24|for he views the ends of the earth and sees everything under the heavens.
JOB|28|25|When he established the force of the wind and measured out the waters,
JOB|28|26|when he made a decree for the rain and a path for the thunderstorm,
JOB|28|27|then he looked at wisdom and appraised it; he confirmed it and tested it.
JOB|28|28|And he said to man, 'The fear of the Lord-that is wisdom, and to shun evil is understanding.'"
JOB|29|1|Job continued his discourse:
JOB|29|2|"How I long for the months gone by, for the days when God watched over me,
JOB|29|3|when his lamp shone upon my head and by his light I walked through darkness!
JOB|29|4|Oh, for the days when I was in my prime, when God's intimate friendship blessed my house,
JOB|29|5|when the Almighty was still with me and my children were around me,
JOB|29|6|when my path was drenched with cream and the rock poured out for me streams of olive oil.
JOB|29|7|"When I went to the gate of the city and took my seat in the public square,
JOB|29|8|the young men saw me and stepped aside and the old men rose to their feet;
JOB|29|9|the chief men refrained from speaking and covered their mouths with their hands;
JOB|29|10|the voices of the nobles were hushed, and their tongues stuck to the roof of their mouths.
JOB|29|11|Whoever heard me spoke well of me, and those who saw me commended me,
JOB|29|12|because I rescued the poor who cried for help, and the fatherless who had none to assist him.
JOB|29|13|The man who was dying blessed me; I made the widow's heart sing.
JOB|29|14|I put on righteousness as my clothing; justice was my robe and my turban.
JOB|29|15|I was eyes to the blind and feet to the lame.
JOB|29|16|I was a father to the needy; I took up the case of the stranger.
JOB|29|17|I broke the fangs of the wicked and snatched the victims from their teeth.
JOB|29|18|"I thought, 'I will die in my own house, my days as numerous as the grains of sand.
JOB|29|19|My roots will reach to the water, and the dew will lie all night on my branches.
JOB|29|20|My glory will remain fresh in me, the bow ever new in my hand.'
JOB|29|21|"Men listened to me expectantly, waiting in silence for my counsel.
JOB|29|22|After I had spoken, they spoke no more; my words fell gently on their ears.
JOB|29|23|They waited for me as for showers and drank in my words as the spring rain.
JOB|29|24|When I smiled at them, they scarcely believed it; the light of my face was precious to them.
JOB|29|25|I chose the way for them and sat as their chief; I dwelt as a king among his troops; I was like one who comforts mourners.
JOB|30|1|"But now they mock me, men younger than I, whose fathers I would have disdained to put with my sheep dogs.
JOB|30|2|Of what use was the strength of their hands to me, since their vigor had gone from them?
JOB|30|3|Haggard from want and hunger, they roamed the parched land in desolate wastelands at night.
JOB|30|4|In the brush they gathered salt herbs, and their food was the root of the broom tree.
JOB|30|5|They were banished from their fellow men, shouted at as if they were thieves.
JOB|30|6|They were forced to live in the dry stream beds, among the rocks and in holes in the ground.
JOB|30|7|They brayed among the bushes and huddled in the undergrowth.
JOB|30|8|A base and nameless brood, they were driven out of the land.
JOB|30|9|"And now their sons mock me in song; I have become a byword among them.
JOB|30|10|They detest me and keep their distance; they do not hesitate to spit in my face.
JOB|30|11|Now that God has unstrung my bow and afflicted me, they throw off restraint in my presence.
JOB|30|12|On my right the tribe attacks; they lay snares for my feet, they build their siege ramps against me.
JOB|30|13|They break up my road; they succeed in destroying me- without anyone's helping them.
JOB|30|14|They advance as through a gaping breach; amid the ruins they come rolling in.
JOB|30|15|Terrors overwhelm me; my dignity is driven away as by the wind, my safety vanishes like a cloud.
JOB|30|16|"And now my life ebbs away; days of suffering grip me.
JOB|30|17|Night pierces my bones; my gnawing pains never rest.
JOB|30|18|In his great power God becomes like clothing to me; he binds me like the neck of my garment.
JOB|30|19|He throws me into the mud, and I am reduced to dust and ashes.
JOB|30|20|"I cry out to you, O God, but you do not answer; I stand up, but you merely look at me.
JOB|30|21|You turn on me ruthlessly; with the might of your hand you attack me.
JOB|30|22|You snatch me up and drive me before the wind; you toss me about in the storm.
JOB|30|23|I know you will bring me down to death, to the place appointed for all the living.
JOB|30|24|"Surely no one lays a hand on a broken man when he cries for help in his distress.
JOB|30|25|Have I not wept for those in trouble? Has not my soul grieved for the poor?
JOB|30|26|Yet when I hoped for good, evil came; when I looked for light, then came darkness.
JOB|30|27|The churning inside me never stops; days of suffering confront me.
JOB|30|28|I go about blackened, but not by the sun; I stand up in the assembly and cry for help.
JOB|30|29|I have become a brother of jackals, a companion of owls.
JOB|30|30|My skin grows black and peels; my body burns with fever.
JOB|30|31|My harp is tuned to mourning, and my flute to the sound of wailing.
JOB|31|1|"I made a covenant with my eyes not to look lustfully at a girl.
JOB|31|2|For what is man's lot from God above, his heritage from the Almighty on high?
JOB|31|3|Is it not ruin for the wicked, disaster for those who do wrong?
JOB|31|4|Does he not see my ways and count my every step?
JOB|31|5|"If I have walked in falsehood or my foot has hurried after deceit-
JOB|31|6|let God weigh me in honest scales and he will know that I am blameless-
JOB|31|7|if my steps have turned from the path, if my heart has been led by my eyes, or if my hands have been defiled,
JOB|31|8|then may others eat what I have sown, and may my crops be uprooted.
JOB|31|9|"If my heart has been enticed by a woman, or if I have lurked at my neighbor's door,
JOB|31|10|then may my wife grind another man's grain, and may other men sleep with her.
JOB|31|11|For that would have been shameful, a sin to be judged.
JOB|31|12|It is a fire that burns to Destruction; it would have uprooted my harvest.
JOB|31|13|"If I have denied justice to my menservants and maidservants when they had a grievance against me,
JOB|31|14|what will I do when God confronts me? What will I answer when called to account?
JOB|31|15|Did not he who made me in the womb make them? Did not the same one form us both within our mothers?
JOB|31|16|"If I have denied the desires of the poor or let the eyes of the widow grow weary,
JOB|31|17|if I have kept my bread to myself, not sharing it with the fatherless-
JOB|31|18|but from my youth I reared him as would a father, and from my birth I guided the widow-
JOB|31|19|if I have seen anyone perishing for lack of clothing, or a needy man without a garment,
JOB|31|20|and his heart did not bless me for warming him with the fleece from my sheep,
JOB|31|21|if I have raised my hand against the fatherless, knowing that I had influence in court,
JOB|31|22|then let my arm fall from the shoulder, let it be broken off at the joint.
JOB|31|23|For I dreaded destruction from God, and for fear of his splendor I could not do such things.
JOB|31|24|"If I have put my trust in gold or said to pure gold, 'You are my security,'
JOB|31|25|if I have rejoiced over my great wealth, the fortune my hands had gained,
JOB|31|26|if I have regarded the sun in its radiance or the moon moving in splendor,
JOB|31|27|so that my heart was secretly enticed and my hand offered them a kiss of homage,
JOB|31|28|then these also would be sins to be judged, for I would have been unfaithful to God on high.
JOB|31|29|"If I have rejoiced at my enemy's misfortune or gloated over the trouble that came to him-
JOB|31|30|I have not allowed my mouth to sin by invoking a curse against his life-
JOB|31|31|if the men of my household have never said, 'Who has not had his fill of Job's meat?'-
JOB|31|32|but no stranger had to spend the night in the street, for my door was always open to the traveler-
JOB|31|33|if I have concealed my sin as men do, by hiding my guilt in my heart
JOB|31|34|because I so feared the crowd and so dreaded the contempt of the clans that I kept silent and would not go outside
JOB|31|35|("Oh, that I had someone to hear me! I sign now my defense-let the Almighty answer me; let my accuser put his indictment in writing.
JOB|31|36|Surely I would wear it on my shoulder, I would put it on like a crown.
JOB|31|37|I would give him an account of my every step; like a prince I would approach him.)-
JOB|31|38|"if my land cries out against me and all its furrows are wet with tears,
JOB|31|39|if I have devoured its yield without payment or broken the spirit of its tenants,
JOB|31|40|then let briers come up instead of wheat and weeds instead of barley." The words of Job are ended.
JOB|32|1|So these three men stopped answering Job, because he was righteous in his own eyes.
JOB|32|2|But Elihu son of Barakel the Buzite, of the family of Ram, became very angry with Job for justifying himself rather than God.
JOB|32|3|He was also angry with the three friends, because they had found no way to refute Job, and yet had condemned him.
JOB|32|4|Now Elihu had waited before speaking to Job because they were older than he.
JOB|32|5|But when he saw that the three men had nothing more to say, his anger was aroused.
JOB|32|6|So Elihu son of Barakel the Buzite said: "I am young in years, and you are old; that is why I was fearful, not daring to tell you what I know.
JOB|32|7|I thought, 'Age should speak; advanced years should teach wisdom.'
JOB|32|8|But it is the spirit in a man, the breath of the Almighty, that gives him understanding.
JOB|32|9|It is not only the old who are wise, not only the aged who understand what is right.
JOB|32|10|"Therefore I say: Listen to me; I too will tell you what I know.
JOB|32|11|I waited while you spoke, I listened to your reasoning; while you were searching for words,
JOB|32|12|I gave you my full attention. But not one of you has proved Job wrong; none of you has answered his arguments.
JOB|32|13|Do not say, 'We have found wisdom; let God refute him, not man.'
JOB|32|14|But Job has not marshaled his words against me, and I will not answer him with your arguments.
JOB|32|15|"They are dismayed and have no more to say; words have failed them.
JOB|32|16|Must I wait, now that they are silent, now that they stand there with no reply?
JOB|32|17|I too will have my say; I too will tell what I know.
JOB|32|18|For I am full of words, and the spirit within me compels me;
JOB|32|19|inside I am like bottled-up wine, like new wineskins ready to burst.
JOB|32|20|I must speak and find relief; I must open my lips and reply.
JOB|32|21|I will show partiality to no one, nor will I flatter any man;
JOB|32|22|for if I were skilled in flattery, my Maker would soon take me away.
JOB|33|1|"But now, Job, listen to my words; pay attention to everything I say.
JOB|33|2|I am about to open my mouth; my words are on the tip of my tongue.
JOB|33|3|My words come from an upright heart; my lips sincerely speak what I know.
JOB|33|4|The Spirit of God has made me; the breath of the Almighty gives me life.
JOB|33|5|Answer me then, if you can; prepare yourself and confront me.
JOB|33|6|I am just like you before God; I too have been taken from clay.
JOB|33|7|No fear of me should alarm you, nor should my hand be heavy upon you.
JOB|33|8|"But you have said in my hearing- I heard the very words-
JOB|33|9|'I am pure and without sin; I am clean and free from guilt.
JOB|33|10|Yet God has found fault with me; he considers me his enemy.
JOB|33|11|He fastens my feet in shackles; he keeps close watch on all my paths.'
JOB|33|12|"But I tell you, in this you are not right, for God is greater than man.
JOB|33|13|Why do you complain to him that he answers none of man's words?
JOB|33|14|For God does speak-now one way, now another- though man may not perceive it.
JOB|33|15|In a dream, in a vision of the night, when deep sleep falls on men as they slumber in their beds,
JOB|33|16|he may speak in their ears and terrify them with warnings,
JOB|33|17|to turn man from wrongdoing and keep him from pride,
JOB|33|18|to preserve his soul from the pit, his life from perishing by the sword.
JOB|33|19|Or a man may be chastened on a bed of pain with constant distress in his bones,
JOB|33|20|so that his very being finds food repulsive and his soul loathes the choicest meal.
JOB|33|21|His flesh wastes away to nothing, and his bones, once hidden, now stick out.
JOB|33|22|His soul draws near to the pit, and his life to the messengers of death.
JOB|33|23|"Yet if there is an angel on his side as a mediator, one out of a thousand, to tell a man what is right for him,
JOB|33|24|to be gracious to him and say, 'Spare him from going down to the pit; I have found a ransom for him'-
JOB|33|25|then his flesh is renewed like a child's; it is restored as in the days of his youth.
JOB|33|26|He prays to God and finds favor with him, he sees God's face and shouts for joy; he is restored by God to his righteous state.
JOB|33|27|Then he comes to men and says, 'I sinned, and perverted what was right, but I did not get what I deserved.
JOB|33|28|He redeemed my soul from going down to the pit, and I will live to enjoy the light.'
JOB|33|29|"God does all these things to a man- twice, even three times-
JOB|33|30|to turn back his soul from the pit, that the light of life may shine on him.
JOB|33|31|"Pay attention, Job, and listen to me; be silent, and I will speak.
JOB|33|32|If you have anything to say, answer me; speak up, for I want you to be cleared.
JOB|33|33|But if not, then listen to me; be silent, and I will teach you wisdom."
JOB|34|1|Then Elihu said:
JOB|34|2|"Hear my words, you wise men; listen to me, you men of learning.
JOB|34|3|For the ear tests words as the tongue tastes food.
JOB|34|4|Let us discern for ourselves what is right; let us learn together what is good.
JOB|34|5|"Job says, 'I am innocent, but God denies me justice.
JOB|34|6|Although I am right, I am considered a liar; although I am guiltless, his arrow inflicts an incurable wound.'
JOB|34|7|What man is like Job, who drinks scorn like water?
JOB|34|8|He keeps company with evildoers; he associates with wicked men.
JOB|34|9|For he says, 'It profits a man nothing when he tries to please God.'
JOB|34|10|"So listen to me, you men of understanding. Far be it from God to do evil, from the Almighty to do wrong.
JOB|34|11|He repays a man for what he has done; he brings upon him what his conduct deserves.
JOB|34|12|It is unthinkable that God would do wrong, that the Almighty would pervert justice.
JOB|34|13|Who appointed him over the earth? Who put him in charge of the whole world?
JOB|34|14|If it were his intention and he withdrew his spirit and breath,
JOB|34|15|all mankind would perish together and man would return to the dust.
JOB|34|16|"If you have understanding, hear this; listen to what I say.
JOB|34|17|Can he who hates justice govern? Will you condemn the just and mighty One?
JOB|34|18|Is he not the One who says to kings, 'You are worthless,' and to nobles, 'You are wicked,'
JOB|34|19|who shows no partiality to princes and does not favor the rich over the poor, for they are all the work of his hands?
JOB|34|20|They die in an instant, in the middle of the night; the people are shaken and they pass away; the mighty are removed without human hand.
JOB|34|21|"His eyes are on the ways of men; he sees their every step.
JOB|34|22|There is no dark place, no deep shadow, where evildoers can hide.
JOB|34|23|God has no need to examine men further, that they should come before him for judgment.
JOB|34|24|Without inquiry he shatters the mighty and sets up others in their place.
JOB|34|25|Because he takes note of their deeds, he overthrows them in the night and they are crushed.
JOB|34|26|He punishes them for their wickedness where everyone can see them,
JOB|34|27|because they turned from following him and had no regard for any of his ways.
JOB|34|28|They caused the cry of the poor to come before him, so that he heard the cry of the needy.
JOB|34|29|But if he remains silent, who can condemn him? If he hides his face, who can see him? Yet he is over man and nation alike,
JOB|34|30|to keep a godless man from ruling, from laying snares for the people.
JOB|34|31|"Suppose a man says to God, 'I am guilty but will offend no more.
JOB|34|32|Teach me what I cannot see; if I have done wrong, I will not do so again.'
JOB|34|33|Should God then reward you on your terms, when you refuse to repent? You must decide, not I; so tell me what you know.
JOB|34|34|"Men of understanding declare, wise men who hear me say to me,
JOB|34|35|'Job speaks without knowledge; his words lack insight.'
JOB|34|36|Oh, that Job might be tested to the utmost for answering like a wicked man!
JOB|34|37|To his sin he adds rebellion; scornfully he claps his hands among us and multiplies his words against God."
JOB|35|1|Then Elihu said:
JOB|35|2|"Do you think this is just? You say, 'I will be cleared by God. '
JOB|35|3|Yet you ask him, 'What profit is it to me, and what do I gain by not sinning?'
JOB|35|4|"I would like to reply to you and to your friends with you.
JOB|35|5|Look up at the heavens and see; gaze at the clouds so high above you.
JOB|35|6|If you sin, how does that affect him? If your sins are many, what does that do to him?
JOB|35|7|If you are righteous, what do you give to him, or what does he receive from your hand?
JOB|35|8|Your wickedness affects only a man like yourself, and your righteousness only the sons of men.
JOB|35|9|"Men cry out under a load of oppression; they plead for relief from the arm of the powerful.
JOB|35|10|But no one says, 'Where is God my Maker, who gives songs in the night,
JOB|35|11|who teaches more to us than to the beasts of the earth and makes us wiser than the birds of the air?'
JOB|35|12|He does not answer when men cry out because of the arrogance of the wicked.
JOB|35|13|Indeed, God does not listen to their empty plea; the Almighty pays no attention to it.
JOB|35|14|How much less, then, will he listen when you say that you do not see him, that your case is before him and you must wait for him,
JOB|35|15|and further, that his anger never punishes and he does not take the least notice of wickedness.
JOB|35|16|So Job opens his mouth with empty talk; without knowledge he multiplies words."
JOB|36|1|Elihu continued:
JOB|36|2|"Bear with me a little longer and I will show you that there is more to be said in God's behalf.
JOB|36|3|I get my knowledge from afar; I will ascribe justice to my Maker.
JOB|36|4|Be assured that my words are not false; one perfect in knowledge is with you.
JOB|36|5|"God is mighty, but does not despise men; he is mighty, and firm in his purpose.
JOB|36|6|He does not keep the wicked alive but gives the afflicted their rights.
JOB|36|7|He does not take his eyes off the righteous; he enthrones them with kings and exalts them forever.
JOB|36|8|But if men are bound in chains, held fast by cords of affliction,
JOB|36|9|he tells them what they have done- that they have sinned arrogantly.
JOB|36|10|He makes them listen to correction and commands them to repent of their evil.
JOB|36|11|If they obey and serve him, they will spend the rest of their days in prosperity and their years in contentment.
JOB|36|12|But if they do not listen, they will perish by the sword and die without knowledge.
JOB|36|13|"The godless in heart harbor resentment; even when he fetters them, they do not cry for help.
JOB|36|14|They die in their youth, among male prostitutes of the shrines.
JOB|36|15|But those who suffer he delivers in their suffering; he speaks to them in their affliction.
JOB|36|16|"He is wooing you from the jaws of distress to a spacious place free from restriction, to the comfort of your table laden with choice food.
JOB|36|17|But now you are laden with the judgment due the wicked; judgment and justice have taken hold of you.
JOB|36|18|Be careful that no one entices you by riches; do not let a large bribe turn you aside.
JOB|36|19|Would your wealth or even all your mighty efforts sustain you so you would not be in distress?
JOB|36|20|Do not long for the night, to drag people away from their homes.
JOB|36|21|Beware of turning to evil, which you seem to prefer to affliction.
JOB|36|22|"God is exalted in his power. Who is a teacher like him?
JOB|36|23|Who has prescribed his ways for him, or said to him, 'You have done wrong'?
JOB|36|24|Remember to extol his work, which men have praised in song.
JOB|36|25|All mankind has seen it; men gaze on it from afar.
JOB|36|26|How great is God-beyond our understanding! The number of his years is past finding out.
JOB|36|27|"He draws up the drops of water, which distill as rain to the streams;
JOB|36|28|the clouds pour down their moisture and abundant showers fall on mankind.
JOB|36|29|Who can understand how he spreads out the clouds, how he thunders from his pavilion?
JOB|36|30|See how he scatters his lightning about him, bathing the depths of the sea.
JOB|36|31|This is the way he governs the nations and provides food in abundance.
JOB|36|32|He fills his hands with lightning and commands it to strike its mark.
JOB|36|33|His thunder announces the coming storm; even the cattle make known its approach.
JOB|37|1|"At this my heart pounds and leaps from its place.
JOB|37|2|Listen! Listen to the roar of his voice, to the rumbling that comes from his mouth.
JOB|37|3|He unleashes his lightning beneath the whole heaven and sends it to the ends of the earth.
JOB|37|4|After that comes the sound of his roar; he thunders with his majestic voice. When his voice resounds, he holds nothing back.
JOB|37|5|God's voice thunders in marvelous ways; he does great things beyond our understanding.
JOB|37|6|He says to the snow, 'Fall on the earth,' and to the rain shower, 'Be a mighty downpour.'
JOB|37|7|So that all men he has made may know his work, he stops every man from his labor.
JOB|37|8|The animals take cover; they remain in their dens.
JOB|37|9|The tempest comes out from its chamber, the cold from the driving winds.
JOB|37|10|The breath of God produces ice, and the broad waters become frozen.
JOB|37|11|He loads the clouds with moisture; he scatters his lightning through them.
JOB|37|12|At his direction they swirl around over the face of the whole earth to do whatever he commands them.
JOB|37|13|He brings the clouds to punish men, or to water his earth and show his love.
JOB|37|14|"Listen to this, Job; stop and consider God's wonders.
JOB|37|15|Do you know how God controls the clouds and makes his lightning flash?
JOB|37|16|Do you know how the clouds hang poised, those wonders of him who is perfect in knowledge?
JOB|37|17|You who swelter in your clothes when the land lies hushed under the south wind,
JOB|37|18|can you join him in spreading out the skies, hard as a mirror of cast bronze?
JOB|37|19|"Tell us what we should say to him; we cannot draw up our case because of our darkness.
JOB|37|20|Should he be told that I want to speak? Would any man ask to be swallowed up?
JOB|37|21|Now no one can look at the sun, bright as it is in the skies after the wind has swept them clean.
JOB|37|22|Out of the north he comes in golden splendor; God comes in awesome majesty.
JOB|37|23|The Almighty is beyond our reach and exalted in power; in his justice and great righteousness, he does not oppress.
JOB|37|24|Therefore, men revere him, for does he not have regard for all the wise in heart? "
JOB|38|1|Then the LORD answered Job out of the storm. He said:
JOB|38|2|"Who is this that darkens my counsel with words without knowledge?
JOB|38|3|Brace yourself like a man; I will question you, and you shall answer me.
JOB|38|4|"Where were you when I laid the earth's foundation? Tell me, if you understand.
JOB|38|5|Who marked off its dimensions? Surely you know! Who stretched a measuring line across it?
JOB|38|6|On what were its footings set, or who laid its cornerstone-
JOB|38|7|while the morning stars sang together and all the angels shouted for joy?
JOB|38|8|"Who shut up the sea behind doors when it burst forth from the womb,
JOB|38|9|when I made the clouds its garment and wrapped it in thick darkness,
JOB|38|10|when I fixed limits for it and set its doors and bars in place,
JOB|38|11|when I said, 'This far you may come and no farther; here is where your proud waves halt'?
JOB|38|12|"Have you ever given orders to the morning, or shown the dawn its place,
JOB|38|13|that it might take the earth by the edges and shake the wicked out of it?
JOB|38|14|The earth takes shape like clay under a seal; its features stand out like those of a garment.
JOB|38|15|The wicked are denied their light, and their upraised arm is broken.
JOB|38|16|"Have you journeyed to the springs of the sea or walked in the recesses of the deep?
JOB|38|17|Have the gates of death been shown to you? Have you seen the gates of the shadow of death?
JOB|38|18|Have you comprehended the vast expanses of the earth? Tell me, if you know all this.
JOB|38|19|"What is the way to the abode of light? And where does darkness reside?
JOB|38|20|Can you take them to their places? Do you know the paths to their dwellings?
JOB|38|21|Surely you know, for you were already born! You have lived so many years!
JOB|38|22|"Have you entered the storehouses of the snow or seen the storehouses of the hail,
JOB|38|23|which I reserve for times of trouble, for days of war and battle?
JOB|38|24|What is the way to the place where the lightning is dispersed, or the place where the east winds are scattered over the earth?
JOB|38|25|Who cuts a channel for the torrents of rain, and a path for the thunderstorm,
JOB|38|26|to water a land where no man lives, a desert with no one in it,
JOB|38|27|to satisfy a desolate wasteland and make it sprout with grass?
JOB|38|28|Does the rain have a father? Who fathers the drops of dew?
JOB|38|29|From whose womb comes the ice? Who gives birth to the frost from the heavens
JOB|38|30|when the waters become hard as stone, when the surface of the deep is frozen?
JOB|38|31|"Can you bind the beautiful Pleiades? Can you loose the cords of Orion?
JOB|38|32|Can you bring forth the constellations in their seasons or lead out the Bear with its cubs?
JOB|38|33|Do you know the laws of the heavens? Can you set up God's dominion over the earth?
JOB|38|34|"Can you raise your voice to the clouds and cover yourself with a flood of water?
JOB|38|35|Do you send the lightning bolts on their way? Do they report to you, 'Here we are'?
JOB|38|36|Who endowed the heart with wisdom or gave understanding to the mind?
JOB|38|37|Who has the wisdom to count the clouds? Who can tip over the water jars of the heavens
JOB|38|38|when the dust becomes hard and the clods of earth stick together?
JOB|38|39|"Do you hunt the prey for the lioness and satisfy the hunger of the lions
JOB|38|40|when they crouch in their dens or lie in wait in a thicket?
JOB|38|41|Who provides food for the raven when its young cry out to God and wander about for lack of food?
JOB|39|1|"Do you know when the mountain goats give birth? Do you watch when the doe bears her fawn?
JOB|39|2|Do you count the months till they bear? Do you know the time they give birth?
JOB|39|3|They crouch down and bring forth their young; their labor pains are ended.
JOB|39|4|Their young thrive and grow strong in the wilds; they leave and do not return.
JOB|39|5|"Who let the wild donkey go free? Who untied his ropes?
JOB|39|6|I gave him the wasteland as his home, the salt flats as his habitat.
JOB|39|7|He laughs at the commotion in the town; he does not hear a driver's shout.
JOB|39|8|He ranges the hills for his pasture and searches for any green thing.
JOB|39|9|"Will the wild ox consent to serve you? Will he stay by your manger at night?
JOB|39|10|Can you hold him to the furrow with a harness? Will he till the valleys behind you?
JOB|39|11|Will you rely on him for his great strength? Will you leave your heavy work to him?
JOB|39|12|Can you trust him to bring in your grain and gather it to your threshing floor?
JOB|39|13|"The wings of the ostrich flap joyfully, but they cannot compare with the pinions and feathers of the stork.
JOB|39|14|She lays her eggs on the ground and lets them warm in the sand,
JOB|39|15|unmindful that a foot may crush them, that some wild animal may trample them.
JOB|39|16|She treats her young harshly, as if they were not hers; she cares not that her labor was in vain,
JOB|39|17|for God did not endow her with wisdom or give her a share of good sense.
JOB|39|18|Yet when she spreads her feathers to run, she laughs at horse and rider.
JOB|39|19|"Do you give the horse his strength or clothe his neck with a flowing mane?
JOB|39|20|Do you make him leap like a locust, striking terror with his proud snorting?
JOB|39|21|He paws fiercely, rejoicing in his strength, and charges into the fray.
JOB|39|22|He laughs at fear, afraid of nothing; he does not shy away from the sword.
JOB|39|23|The quiver rattles against his side, along with the flashing spear and lance.
JOB|39|24|In frenzied excitement he eats up the ground; he cannot stand still when the trumpet sounds.
JOB|39|25|At the blast of the trumpet he snorts, 'Aha!' He catches the scent of battle from afar, the shout of commanders and the battle cry.
JOB|39|26|"Does the hawk take flight by your wisdom and spread his wings toward the south?
JOB|39|27|Does the eagle soar at your command and build his nest on high?
JOB|39|28|He dwells on a cliff and stays there at night; a rocky crag is his stronghold.
JOB|39|29|From there he seeks out his food; his eyes detect it from afar.
JOB|39|30|His young ones feast on blood, and where the slain are, there is he."
JOB|40|1|The LORD said to Job:
JOB|40|2|"Will the one who contends with the Almighty correct him? Let him who accuses God answer him!"
JOB|40|3|Then Job answered the LORD:
JOB|40|4|"I am unworthy-how can I reply to you? I put my hand over my mouth.
JOB|40|5|I spoke once, but I have no answer- twice, but I will say no more."
JOB|40|6|Then the LORD spoke to Job out of the storm:
JOB|40|7|"Brace yourself like a man; I will question you, and you shall answer me.
JOB|40|8|"Would you discredit my justice? Would you condemn me to justify yourself?
JOB|40|9|Do you have an arm like God's, and can your voice thunder like his?
JOB|40|10|Then adorn yourself with glory and splendor, and clothe yourself in honor and majesty.
JOB|40|11|Unleash the fury of your wrath, look at every proud man and bring him low,
JOB|40|12|look at every proud man and humble him, crush the wicked where they stand.
JOB|40|13|Bury them all in the dust together; shroud their faces in the grave.
JOB|40|14|Then I myself will admit to you that your own right hand can save you.
JOB|40|15|"Look at the behemoth, which I made along with you and which feeds on grass like an ox.
JOB|40|16|What strength he has in his loins, what power in the muscles of his belly!
JOB|40|17|His tail sways like a cedar; the sinews of his thighs are close-knit.
JOB|40|18|His bones are tubes of bronze, his limbs like rods of iron.
JOB|40|19|He ranks first among the works of God, yet his Maker can approach him with his sword.
JOB|40|20|The hills bring him their produce, and all the wild animals play nearby.
JOB|40|21|Under the lotus plants he lies, hidden among the reeds in the marsh.
JOB|40|22|The lotuses conceal him in their shadow; the poplars by the stream surround him.
JOB|40|23|When the river rages, he is not alarmed; he is secure, though the Jordan should surge against his mouth.
JOB|40|24|Can anyone capture him by the eyes, or trap him and pierce his nose?
JOB|41|1|"Can you pull in the leviathan with a fishhook or tie down his tongue with a rope?
JOB|41|2|Can you put a cord through his nose or pierce his jaw with a hook?
JOB|41|3|Will he keep begging you for mercy? Will he speak to you with gentle words?
JOB|41|4|Will he make an agreement with you for you to take him as your slave for life?
JOB|41|5|Can you make a pet of him like a bird or put him on a leash for your girls?
JOB|41|6|Will traders barter for him? Will they divide him up among the merchants?
JOB|41|7|Can you fill his hide with harpoons or his head with fishing spears?
JOB|41|8|If you lay a hand on him, you will remember the struggle and never do it again!
JOB|41|9|Any hope of subduing him is false; the mere sight of him is overpowering.
JOB|41|10|No one is fierce enough to rouse him. Who then is able to stand against me?
JOB|41|11|Who has a claim against me that I must pay? Everything under heaven belongs to me.
JOB|41|12|"I will not fail to speak of his limbs, his strength and his graceful form.
JOB|41|13|Who can strip off his outer coat? Who would approach him with a bridle?
JOB|41|14|Who dares open the doors of his mouth, ringed about with his fearsome teeth?
JOB|41|15|His back has rows of shields tightly sealed together;
JOB|41|16|each is so close to the next that no air can pass between.
JOB|41|17|They are joined fast to one another; they cling together and cannot be parted.
JOB|41|18|His snorting throws out flashes of light; his eyes are like the rays of dawn.
JOB|41|19|Firebrands stream from his mouth; sparks of fire shoot out.
JOB|41|20|Smoke pours from his nostrils as from a boiling pot over a fire of reeds.
JOB|41|21|His breath sets coals ablaze, and flames dart from his mouth.
JOB|41|22|Strength resides in his neck; dismay goes before him.
JOB|41|23|The folds of his flesh are tightly joined; they are firm and immovable.
JOB|41|24|His chest is hard as rock, hard as a lower millstone.
JOB|41|25|When he rises up, the mighty are terrified; they retreat before his thrashing.
JOB|41|26|The sword that reaches him has no effect, nor does the spear or the dart or the javelin.
JOB|41|27|Iron he treats like straw and bronze like rotten wood.
JOB|41|28|Arrows do not make him flee; slingstones are like chaff to him.
JOB|41|29|A club seems to him but a piece of straw; he laughs at the rattling of the lance.
JOB|41|30|His undersides are jagged potsherds, leaving a trail in the mud like a threshing sledge.
JOB|41|31|He makes the depths churn like a boiling caldron and stirs up the sea like a pot of ointment.
JOB|41|32|Behind him he leaves a glistening wake; one would think the deep had white hair.
JOB|41|33|Nothing on earth is his equal- a creature without fear.
JOB|41|34|He looks down on all that are haughty; he is king over all that are proud."
JOB|42|1|Then Job replied to the LORD:
JOB|42|2|"I know that you can do all things; no plan of yours can be thwarted.
JOB|42|3|You asked, 'Who is this that obscures my counsel without knowledge?' Surely I spoke of things I did not understand, things too wonderful for me to know.
JOB|42|4|"You said, 'Listen now, and I will speak; I will question you, and you shall answer me.'
JOB|42|5|My ears had heard of you but now my eyes have seen you.
JOB|42|6|Therefore I despise myself and repent in dust and ashes."
JOB|42|7|After the LORD had said these things to Job, he said to Eliphaz the Temanite, "I am angry with you and your two friends, because you have not spoken of me what is right, as my servant Job has.
JOB|42|8|So now take seven bulls and seven rams and go to my servant Job and sacrifice a burnt offering for yourselves. My servant Job will pray for you, and I will accept his prayer and not deal with you according to your folly. You have not spoken of me what is right, as my servant Job has."
JOB|42|9|So Eliphaz the Temanite, Bildad the Shuhite and Zophar the Naamathite did what the LORD told them; and the LORD accepted Job's prayer.
JOB|42|10|After Job had prayed for his friends, the LORD made him prosperous again and gave him twice as much as he had before.
JOB|42|11|All his brothers and sisters and everyone who had known him before came and ate with him in his house. They comforted and consoled him over all the trouble the LORD had brought upon him, and each one gave him a piece of silver and a gold ring.
JOB|42|12|The LORD blessed the latter part of Job's life more than the first. He had fourteen thousand sheep, six thousand camels, a thousand yoke of oxen and a thousand donkeys.
JOB|42|13|And he also had seven sons and three daughters.
JOB|42|14|The first daughter he named Jemimah, the second Keziah and the third Keren-Happuch.
JOB|42|15|Nowhere in all the land were there found women as beautiful as Job's daughters, and their father granted them an inheritance along with their brothers.
JOB|42|16|After this, Job lived a hundred and forty years; he saw his children and their children to the fourth generation.
JOB|42|17|And so he died, old and full of years.
