SONG|1|1|The Song of Songs, which is Solomon's.
SONG|1|2|Let him kiss me with the kisses of his mouth! For your love is better than wine;
SONG|1|3|your anointing oils are fragrant; your name is oil poured out; therefore virgins love you.
SONG|1|4|Draw me after you; let us run. The king has brought me into his chambers. We will exult and rejoice in you; we will extol your love more than wine; rightly do they love you.
SONG|1|5|I am very dark, but lovely, O daughters of Jerusalem, like the tents of Kedar, like the curtains of Solomon.
SONG|1|6|Do not gaze at me because I am dark, because the sun has looked upon me. My mother's sons were angry with me; they made me keeper of the vineyards, but my own vineyard I have not kept!
SONG|1|7|Tell me, you whom my soul loves, where you pasture your flock, where you make it lie down at noon; for why should I be like one who veils herself beside the flocks of your companions?
SONG|1|8|If you do not know, O most beautiful among women, follow in the tracks of the flock, and pasture your young goats beside the shepherds' tents.
SONG|1|9|I compare you, my love, to a mare among Pharaoh's chariots.
SONG|1|10|Your cheeks are lovely with ornaments, your neck with strings of jewels.
SONG|1|11|We will make for you ornaments of gold, studded with silver.
SONG|1|12|While the king was on his couch, my nard gave forth its fragrance.
SONG|1|13|My beloved is to me a sachet of myrrh that lies between my breasts.
SONG|1|14|My beloved is to me a cluster of henna blossoms in the vineyards of Engedi.
SONG|1|15|Behold, you are beautiful, my love; behold, you are beautiful; your eyes are doves.
SONG|1|16|Behold, you are beautiful, my beloved, truly delightful. Our couch is green;
SONG|1|17|the beams of our house are cedar; our rafters are pine.
SONG|2|1|I am a rose of Sharon, a lily of the valleys.
SONG|2|2|As a lily among brambles, so is my love among the young women.
SONG|2|3|As an apple tree among the trees of the forest, so is my beloved among the young men. With great delight I sat in his shadow, and his fruit was sweet to my taste,
SONG|2|4|He brought me to the banqueting house, and his banner over me was love.
SONG|2|5|Sustain me with raisins; refresh me with apples, for I am sick with love.
SONG|2|6|His left hand is under my head, and his right hand embraces me!
SONG|2|7|I adjure you, O daughters of Jerusalem, by the gazelles or the does of the field, that you not stir up or awaken love until it pleases.
SONG|2|8|The voice of my beloved! Behold, he comes, leaping over the mountains, bounding over the hills.
SONG|2|9|My beloved is like a gazelle or a young stag. Behold, there he stands behind our wall, gazing through the windows, looking through the lattice.
SONG|2|10|My beloved speaks and says to me: "Arise, my love, my beautiful one, and come away,
SONG|2|11|for behold, the winter is past; the rain is over and gone.
SONG|2|12|The flowers appear on the earth, the time of singing has come, and the voice of the turtledove is heard in our land.
SONG|2|13|The fig tree ripens its figs, and the vines are in blossom; they give forth fragrance. Arise, my love, my beautiful one, and come away.
SONG|2|14|O my dove, in the clefts of the rock, in the crannies of the cliff, let me see your face, let me hear your voice, for your voice is sweet, and your face is lovely.
SONG|2|15|Catch the foxes for us, the little foxes that spoil the vineyards, for our vineyards are in blossom."
SONG|2|16|My beloved is mine, and I am his; he grazes among the lilies.
SONG|2|17|Until the day breathes and the shadows flee, turn, my beloved, be like a gazelle or a young stag on cleft mountains.
SONG|3|1|On my bed by nightI sought him whom my soul loves; I sought him, but found him not.
SONG|3|2|I will rise now and go about the city, in the streets and in the squares; I will seek him whom my soul loves. I sought him, but found him not.
SONG|3|3|The watchmen found me as they went about in the city. "Have you seen him whom my soul loves?"
SONG|3|4|Scarcely had I passed them when I found him whom my soul loves. I held him, and would not let him go until I had brought him into my mother's house, and into the chamber of her who conceived me.
SONG|3|5|I adjure you, O daughters of Jerusalem, by the gazelles or the does of the field, that you not stir up or awaken love until it pleases.
SONG|3|6|What is that coming up from the wilderness like columns of smoke, perfumed with myrrh and frankincense, with all the fragrant powders of a merchant?
SONG|3|7|Behold, it is the litter of Solomon! Around it are sixty mighty men, some of the mighty men of Israel,
SONG|3|8|all of them wearing swords and expert in war, each with his sword at his thigh, against terror by night.
SONG|3|9|King Solomon made himself a carriage from the wood of Lebanon.
SONG|3|10|He made its posts of silver, its back of gold, its seat of purple; its interior was inlaid with love by the daughters of Jerusalem.
SONG|3|11|Go out, O daughters of Zion, and look upon King Solomon, with the crown with which his mother crowned him on the day of his wedding, on the day of the gladness of his heart.
SONG|4|1|Behold, you are beautiful, my love, behold, you are beautiful! Your eyes are doves behind your veil. Your hair is like a flock of goats leaping down the slopes of Gilead.
SONG|4|2|Your teeth are like a flock of shorn ewes that have come up from the washing, all of which bear twins, and not one among them has lost its young.
SONG|4|3|Your lips are like a scarlet thread, and your mouth is lovely. Your cheeks are like halves of a pomegranate behind your veil.
SONG|4|4|Your neck is like the tower of David, built in rows of stone; on it hang a thousand shields, all of them shields of warriors.
SONG|4|5|Your two breasts are like two fawns, twins of a gazelle, that graze among the lilies.
SONG|4|6|Until the day breathes and the shadows flee, I will go away to the mountain of myrrh and the hill of frankincense.
SONG|4|7|You are altogether beautiful, my love; there is no flaw in you.
SONG|4|8|Come with me from Lebanon, my bride; come with me from Lebanon. Depart from the peak of Amana, from the peak of Senir and Hermon, from the dens of lions, from the mountains of leopards.
SONG|4|9|You have captivated my heart, my sister, my bride; you have captivated my heart with one glance of your eyes, with one jewel of your necklace.
SONG|4|10|How beautiful is your love, my sister, my bride! How much better is your love than wine, and the fragrance of your oils than any spice!
SONG|4|11|Your lips drip nectar, my bride; honey and milk are under your tongue; the fragrance of your garments is like the fragrance of Lebanon.
SONG|4|12|A garden locked is my sister, my bride, a spring locked, a fountain sealed.
SONG|4|13|Your shoots are an orchard of pomegranates with all choicest fruits, henna with nard,
SONG|4|14|nard and saffron, calamus and cinnamon, with all trees of frankincense, myrrh and aloes, with all chief spices-
SONG|4|15|a garden fountain, a well of living water, and flowing streams from Lebanon.
SONG|4|16|Awake, O north wind, and come, O south wind! Blow upon my garden, let its spices flow. Let my beloved come to his garden, and eat its choicest fruits.
SONG|5|1|I came to my garden, my sister, my bride, I gathered my myrrh with my spice, I ate my honeycomb with my honey, I drank my wine with my milk. Eat, friends, drink, and be drunk with love!
SONG|5|2|I slept, but my heart was awake. A sound! My beloved is knocking. "Open to me, my sister, my love, my dove, my perfect one, for my head is wet with dew, my locks with the drops of the night."
SONG|5|3|I had put off my garment; how could I put it on? I had bathed my feet; how could I soil them?
SONG|5|4|My beloved put his hand to the latch, and my heart was thrilled within me.
SONG|5|5|I arose to open to my beloved, and my hands dripped with myrrh, my fingers with liquid myrrh, on the handles of the bolt.
SONG|5|6|I opened to my beloved, but my beloved had turned and gone. My soul failed me when he spoke. I sought him, but found him not; I called him, but he gave no answer.
SONG|5|7|The watchmen found me as they went about in the city; they beat me, they bruised me, they took away my veil, those watchmen of the walls.
SONG|5|8|I adjure you, O daughters of Jerusalem, if you find my beloved, that you tell him I am sick with love.
SONG|5|9|What is your beloved more than another beloved, O most beautiful among women? What is your beloved more than another beloved, that you thus adjure us?
SONG|5|10|My beloved is radiant and ruddy, distinguished among ten thousand.
SONG|5|11|His head is the finest gold; his locks are wavy, black as a raven.
SONG|5|12|His eyes are like doves beside streams of water, bathed in milk, sitting beside a full pool.
SONG|5|13|His cheeks are like beds of spices, mounds of sweet-smelling herbs. His lips are lilies, dripping liquid myrrh.
SONG|5|14|His arms are rods of gold, set with jewels. His body is polished ivory, bedecked with sapphires.
SONG|5|15|His legs are alabaster columns, set on bases of gold. His appearance is like Lebanon, choice as the cedars.
SONG|5|16|His mouth is most sweet, and he is altogether desirable. This is my beloved and this is my friend, O daughters of Jerusalem.
SONG|6|1|Where has your beloved gone, O most beautiful among women? Where has your beloved turned, that we may seek him with you?
SONG|6|2|My beloved has gone down to his garden to the beds of spices, to graze in the gardens and to gather lilies.
SONG|6|3|I am my beloved's and my beloved is mine; he grazes among the lilies.
SONG|6|4|You are beautiful as Tirzah, my love, lovely as Jerusalem, awesome as an army with banners.
SONG|6|5|Turn away your eyes from me, for they overwhelm me- Your hair is like a flock of goats leaping down the slopes of Gilead.
SONG|6|6|Your teeth are like a flock of ewes that have come up from the washing; all of them bear twins; not one among them has lost its young.
SONG|6|7|Your cheeks are like halves of a pomegranate behind your veil.
SONG|6|8|There are sixty queens and eighty concubines, and virgins without number.
SONG|6|9|My dove, my perfect one, is the only one, the only one of her mother, pure to her who bore her. The young women saw her and called her blessed; the queens and concubines also, and they praised her.
SONG|6|10|"Who is this who looks down like the dawn, beautiful as the moon, bright as the sun, awesome as an army with banners?"
SONG|6|11|I went down to the nut orchard to look at the blossoms of the valley, to see whether the vines had budded, whether the pomegranates were in bloom.
SONG|6|12|Before I was aware, my desire set me among the chariots of my kinsman, a prince.
SONG|6|13|Return, return, O Shulammite, return, return, that we may look upon you. Why should you look upon the Shulammite, as upon a dance before two armies?
SONG|7|1|How beautiful are your feet in sandals, O noble daughter! Your rounded thighs are like jewels, the work of a master hand.
SONG|7|2|Your navel is a rounded bowl that never lacks mixed wine. Your belly is a heap of wheat, encircled with lilies.
SONG|7|3|Your two breasts are like two fawns, twins of a gazelle.
SONG|7|4|Your neck is like an ivory tower. Your eyes are pools in Heshbon, by the gate of Bath-rabbim. Your nose is like a tower of Lebanon, which looks toward Damascus.
SONG|7|5|Your head crowns you like Carmel, and your flowing locks are like purple; a king is held captive in the tresses.
SONG|7|6|How beautiful and pleasant you are, O loved one, with all your delights!
SONG|7|7|Your stature is like a palm tree, and your breasts are like its clusters.
SONG|7|8|I say I will climb the palm tree and lay hold of its fruit. Oh may your breasts be like clusters of the vine, and the scent of your breath like apples,
SONG|7|9|and your mouth like the best wine. It goes down smoothly for my beloved, gliding over lips and teeth.
SONG|7|10|I am my beloved's, and his desire is for me.
SONG|7|11|Come, my beloved, let us go out into the fields and lodge in the villages;
SONG|7|12|let us go out early to the vineyards and see whether the vines have budded, whether the grape blossoms have opened and the pomegranates are in bloom. There I will give you my love.
SONG|7|13|The mandrakes give forth fragrance, and beside our doors are all choice fruits, new as well as old, which I have laid up for you, O my beloved.
SONG|8|1|Oh that you were like a brother to me who nursed at my mother's breasts! If I found you outside, I would kiss you, and none would despise me.
SONG|8|2|I would lead you and bring you into the house of my mother- she who used to teach me. I would give you spiced wine to drink, the juice of my pomegranate.
SONG|8|3|His left hand is under my head, and his right hand embraces me!
SONG|8|4|I adjure you, O daughters of Jerusalem, that you not stir up or awaken love until it pleases.
SONG|8|5|Who is that coming up from the wilderness, leaning on her beloved? Under the apple tree I awakened you. There your mother was in labor with you; there she who bore you was in labor.
SONG|8|6|Set me as a seal upon your heart, as a seal upon your arm, for love is strong as death, jealousy is fierce as the grave. Its flashes are flashes of fire, the very flame of the LORD.
SONG|8|7|Many waters cannot quench love, neither can floods drown it. If a man offered for love all the wealth of his house, he would be utterly despised.
SONG|8|8|We have a little sister, and she has no breasts. What shall we do for our sister on the day when she is spoken for?
SONG|8|9|If she is a wall, we will build on her a battlement of silver, but if she is a door, we will enclose her with boards of cedar.
SONG|8|10|I was a wall, and my breasts were like towers; then I was in his eyes as one who finds peace.
SONG|8|11|Solomon had a vineyard at Baal-hamon; he let out the vineyard to keepers; each one was to bring for its fruit a thousand pieces of silver.
SONG|8|12|My vineyard, my very own, is before me; you, O Solomon, may have the thousand, and the keepers of the fruit two hundred.
SONG|8|13|O you who dwell in the gardens, with companions listening for your voice; let me hear it.
SONG|8|14|Make haste, my beloved, and be like a gazelle or a young stag on the mountains of spices.
