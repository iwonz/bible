2JOHN|1|1|Старец – избранной госпоже и детям ее, которых я люблю по истине, и не только я, но и все, познавшие истину,
2JOHN|1|2|ради истины, которая пребывает в нас и будет с нами вовек.
2JOHN|1|3|Да будет с вами благодать, милость, мир от Бога Отца и от Господа Иисуса Христа, Сына Отчего, в истине и любви.
2JOHN|1|4|Я весьма обрадовался, что нашел из детей твоих, ходящих в истине, как мы получили заповедь от Отца.
2JOHN|1|5|И ныне прошу тебя, госпожа, не как новую заповедь предписывая тебе, но ту, которую имеем от начала, чтобы мы любили друг друга.
2JOHN|1|6|Любовь же состоит в том, чтобы мы поступали по заповедям Его. Это та заповедь, которую вы слышали от начала, чтобы поступали по ней.
2JOHN|1|7|Ибо многие обольстители вошли в мир, не исповедующие Иисуса Христа, пришедшего во плоти: такой [человек] есть обольститель и антихрист.
2JOHN|1|8|Наблюдайте за собою, чтобы нам не потерять того, над чем мы трудились, но чтобы получить полную награду.
2JOHN|1|9|Всякий, преступающий учение Христово и не пребывающий в нем, не имеет Бога; пребывающий в учении Христовом имеет и Отца и Сына.
2JOHN|1|10|Кто приходит к вам и не приносит сего учения, того не принимайте в дом и не приветствуйте его.
2JOHN|1|11|Ибо приветствующий его участвует в злых делах его.
2JOHN|1|12|Многое имею писать вам, но не хочу на бумаге чернилами, а надеюсь придти к вам и говорить устами к устам, чтобы радость ваша была полна.
2JOHN|1|13|Приветствуют тебя дети сестры твоей избранной. Аминь.
