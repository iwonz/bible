AMOS|1|1|The words of Amos, one of the shepherds of Tekoa-what he saw concerning Israel two years before the earthquake, when Uzziah was king of Judah and Jeroboam son of Jehoash was king of Israel.
AMOS|1|2|He said: "The LORD roars from Zion and thunders from Jerusalem; the pastures of the shepherds dry up, and the top of Carmel withers."
AMOS|1|3|This is what the LORD says: "For three sins of Damascus, even for four, I will not turn back my wrath. Because she threshed Gilead with sledges having iron teeth,
AMOS|1|4|I will send fire upon the house of Hazael that will consume the fortresses of Ben-Hadad.
AMOS|1|5|I will break down the gate of Damascus; I will destroy the king who is in the Valley of Aven and the one who holds the scepter in Beth Eden. The people of Aram will go into exile to Kir," says the LORD.
AMOS|1|6|This is what the LORD says: "For three sins of Gaza, even for four, I will not turn back my wrath. Because she took captive whole communities and sold them to Edom,
AMOS|1|7|I will send fire upon the walls of Gaza that will consume her fortresses.
AMOS|1|8|I will destroy the king of Ashdod and the one who holds the scepter in Ashkelon. I will turn my hand against Ekron, till the last of the Philistines is dead," says the Sovereign LORD.
AMOS|1|9|This is what the LORD says: "For three sins of Tyre, even for four, I will not turn back my wrath. Because she sold whole communities of captives to Edom, disregarding a treaty of brotherhood,
AMOS|1|10|I will send fire upon the walls of Tyre that will consume her fortresses."
AMOS|1|11|This is what the LORD says: "For three sins of Edom, even for four, I will not turn back my wrath. Because he pursued his brother with a sword, stifling all compassion, because his anger raged continually and his fury flamed unchecked,
AMOS|1|12|I will send fire upon Teman that will consume the fortresses of Bozrah."
AMOS|1|13|This is what the LORD says: "For three sins of Ammon, even for four, I will not turn back {my wrath}. Because he ripped open the pregnant women of Gilead in order to extend his borders,
AMOS|1|14|I will set fire to the walls of Rabbah that will consume her fortresses amid war cries on the day of battle, amid violent winds on a stormy day.
AMOS|1|15|Her king will go into exile, he and his officials together," says the LORD.
AMOS|2|1|This is what the LORD says: "For three sins of Moab, even for four, I will not turn back {my wrath}. Because he burned, as if to lime, the bones of Edom's king,
AMOS|2|2|I will send fire upon Moab that will consume the fortresses of Kerioth. Moab will go down in great tumult amid war cries and the blast of the trumpet.
AMOS|2|3|I will destroy her ruler and kill all her officials with him," says the LORD.
AMOS|2|4|This is what the LORD says: "For three sins of Judah, even for four, I will not turn back {my wrath}. Because they have rejected the law of the LORD and have not kept his decrees, because they have been led astray by false gods, the gods their ancestors followed,
AMOS|2|5|I will send fire upon Judah that will consume the fortresses of Jerusalem."
AMOS|2|6|This is what the LORD says: "For three sins of Israel, even for four, I will not turn back {my wrath}. They sell the righteous for silver, and the needy for a pair of sandals.
AMOS|2|7|They trample on the heads of the poor as upon the dust of the ground and deny justice to the oppressed. Father and son use the same girl and so profane my holy name.
AMOS|2|8|They lie down beside every altar on garments taken in pledge. In the house of their god they drink wine taken as fines.
AMOS|2|9|"I destroyed the Amorite before them, though he was tall as the cedars and strong as the oaks. I destroyed his fruit above and his roots below.
AMOS|2|10|"I brought you up out of Egypt, and I led you forty years in the desert to give you the land of the Amorites.
AMOS|2|11|I also raised up prophets from among your sons and Nazirites from among your young men. Is this not true, people of Israel?" declares the LORD.
AMOS|2|12|"But you made the Nazirites drink wine and commanded the prophets not to prophesy.
AMOS|2|13|"Now then, I will crush you as a cart crushes when loaded with grain.
AMOS|2|14|The swift will not escape, the strong will not muster their strength, and the warrior will not save his life.
AMOS|2|15|The archer will not stand his ground, the fleet-footed soldier will not get away, and the horseman will not save his life.
AMOS|2|16|Even the bravest warriors will flee naked on that day," declares the LORD.
AMOS|3|1|Hear this word the LORD has spoken against you, O people of Israel-against the whole family I brought up out of Egypt:
AMOS|3|2|"You only have I chosen of all the families of the earth; therefore I will punish you for all your sins."
AMOS|3|3|Do two walk together unless they have agreed to do so?
AMOS|3|4|Does a lion roar in the thicket when he has no prey? Does he growl in his den when he has caught nothing?
AMOS|3|5|Does a bird fall into a trap on the ground where no snare has been set? Does a trap spring up from the earth when there is nothing to catch?
AMOS|3|6|When a trumpet sounds in a city, do not the people tremble? When disaster comes to a city, has not the LORD caused it?
AMOS|3|7|Surely the Sovereign LORD does nothing without revealing his plan to his servants the prophets.
AMOS|3|8|The lion has roared- who will not fear? The Sovereign LORD has spoken- who can but prophesy?
AMOS|3|9|Proclaim to the fortresses of Ashdod and to the fortresses of Egypt: "Assemble yourselves on the mountains of Samaria; see the great unrest within her and the oppression among her people."
AMOS|3|10|"They do not know how to do right," declares the LORD, "who hoard plunder and loot in their fortresses."
AMOS|3|11|Therefore this is what the Sovereign LORD says: "An enemy will overrun the land; he will pull down your strongholds and plunder your fortresses."
AMOS|3|12|This is what the LORD says: "As a shepherd saves from the lion's mouth only two leg bones or a piece of an ear, so will the Israelites be saved, those who sit in Samaria on the edge of their beds and in Damascus on their couches. "
AMOS|3|13|"Hear this and testify against the house of Jacob," declares the Lord, the LORD God Almighty.
AMOS|3|14|"On the day I punish Israel for her sins, I will destroy the altars of Bethel; the horns of the altar will be cut off and fall to the ground.
AMOS|3|15|I will tear down the winter house along with the summer house; the houses adorned with ivory will be destroyed and the mansions will be demolished," declares the LORD.
AMOS|4|1|Hear this word, you cows of Bashan on Mount Samaria, you women who oppress the poor and crush the needy and say to your husbands, "Bring us some drinks!"
AMOS|4|2|The Sovereign LORD has sworn by his holiness: "The time will surely come when you will be taken away with hooks, the last of you with fishhooks.
AMOS|4|3|You will each go straight out through breaks in the wall, and you will be cast out toward Harmon, "declares the LORD.
AMOS|4|4|"Go to Bethel and sin; go to Gilgal and sin yet more. Bring your sacrifices every morning, your tithes every three years.
AMOS|4|5|Burn leavened bread as a thank offering and brag about your freewill offerings- boast about them, you Israelites, for this is what you love to do," declares the Sovereign LORD.
AMOS|4|6|"I gave you empty stomachs in every city and lack of bread in every town, yet you have not returned to me," declares the LORD.
AMOS|4|7|"I also withheld rain from you when the harvest was still three months away. I sent rain on one town, but withheld it from another. One field had rain; another had none and dried up.
AMOS|4|8|People staggered from town to town for water but did not get enough to drink, yet you have not returned to me," declares the LORD.
AMOS|4|9|"Many times I struck your gardens and vineyards, I struck them with blight and mildew. Locusts devoured your fig and olive trees, yet you have not returned to me," declares the LORD.
AMOS|4|10|"I sent plagues among you as I did to Egypt. I killed your young men with the sword, along with your captured horses. I filled your nostrils with the stench of your camps, yet you have not returned to me," declares the LORD.
AMOS|4|11|"I overthrew some of you as I overthrew Sodom and Gomorrah. You were like a burning stick snatched from the fire, yet you have not returned to me," declares the LORD.
AMOS|4|12|"Therefore this is what I will do to you, Israel, and because I will do this to you, prepare to meet your God, O Israel."
AMOS|4|13|He who forms the mountains, creates the wind, and reveals his thoughts to man, he who turns dawn to darkness, and treads the high places of the earth- the LORD God Almighty is his name.
AMOS|5|1|Hear this word, O house of Israel, this lament I take up concerning you:
AMOS|5|2|"Fallen is Virgin Israel, never to rise again, deserted in her own land, with no one to lift her up."
AMOS|5|3|This is what the Sovereign LORD says: "The city that marches out a thousand strong for Israel will have only a hundred left; the town that marches out a hundred strong will have only ten left."
AMOS|5|4|This is what the LORD says to the house of Israel: "Seek me and live;
AMOS|5|5|do not seek Bethel, do not go to Gilgal, do not journey to Beersheba. For Gilgal will surely go into exile, and Bethel will be reduced to nothing. "
AMOS|5|6|Seek the LORD and live, or he will sweep through the house of Joseph like a fire; it will devour, and Bethel will have no one to quench it.
AMOS|5|7|You who turn justice into bitterness and cast righteousness to the ground
AMOS|5|8|(he who made the Pleiades and Orion, who turns blackness into dawn and darkens day into night, who calls for the waters of the sea and pours them out over the face of the land- the LORD is his name-
AMOS|5|9|he flashes destruction on the stronghold and brings the fortified city to ruin),
AMOS|5|10|you hate the one who reproves in court and despise him who tells the truth.
AMOS|5|11|You trample on the poor and force him to give you grain. Therefore, though you have built stone mansions, you will not live in them; though you have planted lush vineyards, you will not drink their wine.
AMOS|5|12|For I know how many are your offenses and how great your sins. You oppress the righteous and take bribes and you deprive the poor of justice in the courts.
AMOS|5|13|Therefore the prudent man keeps quiet in such times, for the times are evil.
AMOS|5|14|Seek good, not evil, that you may live. Then the LORD God Almighty will be with you, just as you say he is.
AMOS|5|15|Hate evil, love good; maintain justice in the courts. Perhaps the LORD God Almighty will have mercy on the remnant of Joseph.
AMOS|5|16|Therefore this is what the Lord, the LORD God Almighty, says: "There will be wailing in all the streets and cries of anguish in every public square. The farmers will be summoned to weep and the mourners to wail.
AMOS|5|17|There will be wailing in all the vineyards, for I will pass through your midst," says the LORD.
AMOS|5|18|Woe to you who long for the day of the LORD! Why do you long for the day of the LORD? That day will be darkness, not light.
AMOS|5|19|It will be as though a man fled from a lion only to meet a bear, as though he entered his house and rested his hand on the wall only to have a snake bite him.
AMOS|5|20|Will not the day of the LORD be darkness, not light- pitch-dark, without a ray of brightness?
AMOS|5|21|"I hate, I despise your religious feasts; I cannot stand your assemblies.
AMOS|5|22|Even though you bring me burnt offerings and grain offerings, I will not accept them. Though you bring choice fellowship offerings, I will have no regard for them.
AMOS|5|23|Away with the noise of your songs! I will not listen to the music of your harps.
AMOS|5|24|But let justice roll on like a river, righteousness like a never-failing stream!
AMOS|5|25|"Did you bring me sacrifices and offerings forty years in the desert, O house of Israel?
AMOS|5|26|You have lifted up the shrine of your king, the pedestal of your idols, the star of your god - which you made for yourselves.
AMOS|5|27|Therefore I will send you into exile beyond Damascus," says the LORD, whose name is God Almighty.
AMOS|6|1|Woe to you who are complacent in Zion, and to you who feel secure on Mount Samaria, you notable men of the foremost nation, to whom the people of Israel come!
AMOS|6|2|Go to Calneh and look at it; go from there to great Hamath, and then go down to Gath in Philistia. Are they better off than your two kingdoms? Is their land larger than yours?
AMOS|6|3|You put off the evil day and bring near a reign of terror.
AMOS|6|4|You lie on beds inlaid with ivory and lounge on your couches. You dine on choice lambs and fattened calves.
AMOS|6|5|You strum away on your harps like David and improvise on musical instruments.
AMOS|6|6|You drink wine by the bowlful and use the finest lotions, but you do not grieve over the ruin of Joseph.
AMOS|6|7|Therefore you will be among the first to go into exile; your feasting and lounging will end.
AMOS|6|8|The Sovereign LORD has sworn by himself-the LORD God Almighty declares: "I abhor the pride of Jacob and detest his fortresses; I will deliver up the city and everything in it."
AMOS|6|9|If ten men are left in one house, they too will die.
AMOS|6|10|And if a relative who is to burn the bodies comes to carry them out of the house and asks anyone still hiding there, "Is anyone with you?" and he says, "No," then he will say, "Hush! We must not mention the name of the LORD."
AMOS|6|11|For the LORD has given the command, and he will smash the great house into pieces and the small house into bits.
AMOS|6|12|Do horses run on the rocky crags? Does one plow there with oxen? But you have turned justice into poison and the fruit of righteousness into bitterness-
AMOS|6|13|you who rejoice in the conquest of Lo Debar and say, "Did we not take Karnaim by our own strength?"
AMOS|6|14|For the LORD God Almighty declares, "I will stir up a nation against you, O house of Israel, that will oppress you all the way from Lebo Hamath to the valley of the Arabah."
AMOS|7|1|This is what the Sovereign LORD showed me: He was preparing swarms of locusts after the king's share had been harvested and just as the second crop was coming up.
AMOS|7|2|When they had stripped the land clean, I cried out, "Sovereign LORD, forgive! How can Jacob survive? He is so small!"
AMOS|7|3|So the LORD relented. "This will not happen," the LORD said.
AMOS|7|4|This is what the Sovereign LORD showed me: The Sovereign LORD was calling for judgment by fire; it dried up the great deep and devoured the land.
AMOS|7|5|Then I cried out, "Sovereign LORD, I beg you, stop! How can Jacob survive? He is so small!"
AMOS|7|6|So the LORD relented. "This will not happen either," the Sovereign LORD said.
AMOS|7|7|This is what he showed me: The Lord was standing by a wall that had been built true to plumb, with a plumb line in his hand.
AMOS|7|8|And the LORD asked me, "What do you see, Amos?A plumb line," I replied. Then the Lord said, "Look, I am setting a plumb line among my people Israel; I will spare them no longer.
AMOS|7|9|"The high places of Isaac will be destroyed and the sanctuaries of Israel will be ruined; with my sword I will rise against the house of Jeroboam."
AMOS|7|10|Then Amaziah the priest of Bethel sent a message to Jeroboam king of Israel: "Amos is raising a conspiracy against you in the very heart of Israel. The land cannot bear all his words.
AMOS|7|11|For this is what Amos is saying: "'Jeroboam will die by the sword, and Israel will surely go into exile, away from their native land.'"
AMOS|7|12|Then Amaziah said to Amos, "Get out, you seer! Go back to the land of Judah. Earn your bread there and do your prophesying there.
AMOS|7|13|Don't prophesy anymore at Bethel, because this is the king's sanctuary and the temple of the kingdom."
AMOS|7|14|Amos answered Amaziah, "I was neither a prophet nor a prophet's son, but I was a shepherd, and I also took care of sycamore-fig trees.
AMOS|7|15|But the LORD took me from tending the flock and said to me, 'Go, prophesy to my people Israel.'
AMOS|7|16|Now then, hear the word of the LORD. You say, "'Do not prophesy against Israel, and stop preaching against the house of Isaac.'
AMOS|7|17|"Therefore this is what the LORD says: "'Your wife will become a prostitute in the city, and your sons and daughters will fall by the sword. Your land will be measured and divided up, and you yourself will die in a pagan country. And Israel will certainly go into exile, away from their native land.'"
AMOS|8|1|This is what the Sovereign LORD showed me: a basket of ripe fruit.
AMOS|8|2|"What do you see, Amos?" he asked. "A basket of ripe fruit," I answered. Then the LORD said to me, "The time is ripe for my people Israel; I will spare them no longer.
AMOS|8|3|"In that day," declares the Sovereign LORD, "the songs in the temple will turn to wailing. Many, many bodies-flung everywhere! Silence!"
AMOS|8|4|Hear this, you who trample the needy and do away with the poor of the land,
AMOS|8|5|saying, "When will the New Moon be over that we may sell grain, and the Sabbath be ended that we may market wheat?"- skimping the measure, boosting the price and cheating with dishonest scales,
AMOS|8|6|buying the poor with silver and the needy for a pair of sandals, selling even the sweepings with the wheat.
AMOS|8|7|The LORD has sworn by the Pride of Jacob: "I will never forget anything they have done.
AMOS|8|8|"Will not the land tremble for this, and all who live in it mourn? The whole land will rise like the Nile; it will be stirred up and then sink like the river of Egypt.
AMOS|8|9|"In that day," declares the Sovereign LORD, "I will make the sun go down at noon and darken the earth in broad daylight.
AMOS|8|10|I will turn your religious feasts into mourning and all your singing into weeping. I will make all of you wear sackcloth and shave your heads. I will make that time like mourning for an only son and the end of it like a bitter day.
AMOS|8|11|"The days are coming," declares the Sovereign LORD, "when I will send a famine through the land- not a famine of food or a thirst for water, but a famine of hearing the words of the LORD.
AMOS|8|12|Men will stagger from sea to sea and wander from north to east, searching for the word of the LORD, but they will not find it.
AMOS|8|13|"In that day "the lovely young women and strong young men will faint because of thirst.
AMOS|8|14|They who swear by the shame of Samaria, or say, 'As surely as your god lives, O Dan,' or, 'As surely as the god of Beersheba lives'- they will fall, never to rise again."
AMOS|9|1|I saw the Lord standing by the altar, and he said: "Strike the tops of the pillars so that the thresholds shake. Bring them down on the heads of all the people; those who are left I will kill with the sword. Not one will get away, none will escape.
AMOS|9|2|Though they dig down to the depths of the grave, from there my hand will take them. Though they climb up to the heavens, from there I will bring them down.
AMOS|9|3|Though they hide themselves on the top of Carmel, there I will hunt them down and seize them. Though they hide from me at the bottom of the sea, there I will command the serpent to bite them.
AMOS|9|4|Though they are driven into exile by their enemies, there I will command the sword to slay them. I will fix my eyes upon them for evil and not for good."
AMOS|9|5|The Lord, the LORD Almighty, he who touches the earth and it melts, and all who live in it mourn- the whole land rises like the Nile, then sinks like the river of Egypt-
AMOS|9|6|he who builds his lofty palace in the heavens and sets its foundation on the earth, who calls for the waters of the sea and pours them out over the face of the land- the LORD is his name.
AMOS|9|7|"Are not you Israelites the same to me as the Cushites?" declares the LORD. "Did I not bring Israel up from Egypt, the Philistines from Caphtor and the Arameans from Kir?
AMOS|9|8|"Surely the eyes of the Sovereign LORD are on the sinful kingdom. I will destroy it from the face of the earth- yet I will not totally destroy the house of Jacob," declares the LORD.
AMOS|9|9|"For I will give the command, and I will shake the house of Israel among all the nations as grain is shaken in a sieve, and not a pebble will reach the ground.
AMOS|9|10|All the sinners among my people will die by the sword, all those who say, 'Disaster will not overtake or meet us.'
AMOS|9|11|"In that day I will restore David's fallen tent. I will repair its broken places, restore its ruins, and build it as it used to be,
AMOS|9|12|so that they may possess the remnant of Edom and all the nations that bear my name, "declares the LORD, who will do these things.
AMOS|9|13|"The days are coming," declares the LORD, "when the reaper will be overtaken by the plowman and the planter by the one treading grapes. New wine will drip from the mountains and flow from all the hills.
AMOS|9|14|I will bring back my exiled people Israel; they will rebuild the ruined cities and live in them. They will plant vineyards and drink their wine; they will make gardens and eat their fruit.
AMOS|9|15|I will plant Israel in their own land, never again to be uprooted from the land I have given them," says the LORD your God.
