1THESS|1|1|保羅 、 西拉 、 提摩太 寫信給 帖撒羅尼迦 在父上帝和主耶穌基督裏的教會。願恩惠、平安 歸給你們！
1THESS|1|2|我們為你們眾人常常感謝上帝，禱告的時候提到你們，
1THESS|1|3|在我們的父上帝面前，不住地記念你們因信心所做的工作，因愛心所受的勞苦，因盼望我們主耶穌基督所存的堅忍。
1THESS|1|4|上帝所愛的弟兄啊，我知道你們是蒙揀選的；
1THESS|1|5|因為我們的福音傳到你們那裏，不僅在言語，也在能力，也在聖靈和充足的確信。你們知道，我們在你們那裏，為你們的緣故是怎樣為人。
1THESS|1|6|你們成為效法我們，更效法主的人，因聖靈所激發的喜樂，在大患難中領受了真道，
1THESS|1|7|從此你們作了 馬其頓 和 亞該亞 所有信主的人的榜樣。
1THESS|1|8|因為主的道已經從你們那裏傳播出去，你們向上帝的信心不只在 馬其頓 和 亞該亞 ，就是在各處也都傳開了，所以不用我們說甚麼話。
1THESS|1|9|因為他們自己已經傳講我們是怎樣進到你們那裏，你們是怎樣離棄偶像，歸向上帝來服侍那又真又活的上帝，
1THESS|1|10|等候他兒子從天降臨，就是上帝使他從死人中復活的那位救我們脫離將來憤怒的耶穌。
1THESS|2|1|弟兄們，你們自己知道我們來到你們那裏並不是徒然的。
1THESS|2|2|我們從前在 腓立比 蒙難受辱，這是你們知道的，可是我們還是靠著上帝給我們的勇氣，在強烈反對中把上帝的福音傳給你們。
1THESS|2|3|我們的勸勉不是出於錯誤，也不是出於污穢，也不是用詭詐。
1THESS|2|4|但上帝既然認定我們經得起考驗，把福音託付我們，我們就照著傳講，不是要討人喜歡，而是要討那考驗我們的心的上帝喜歡。
1THESS|2|5|因為我們從來沒有用過諂媚的話，這是你們知道的，也沒有藏著貪心，這是上帝可以作證的。
1THESS|2|6|我們作為基督的使徒，雖然可以受人尊重，卻沒有向你們或向別人求榮耀，反而在你們當中心存溫柔，如同母親哺乳自己的孩子。
1THESS|2|7|
1THESS|2|8|既然我們這樣愛你們，不但樂意將上帝的福音給你們，連自己的性命也樂意給你們，因為你們是我們所疼愛的。
1THESS|2|9|弟兄們，你們記念我們的辛苦勞碌，晝夜做工，傳上帝的福音給你們，免得你們任何人受累。
1THESS|2|10|我們對你們信主的人是何等聖潔、正直、無可指責，這有你們作證，也有上帝作證。
1THESS|2|11|正如你們知道，我們待你們好像父親待自己的兒女一樣。
1THESS|2|12|我們勸勉你們，安慰你們，囑咐你們，使你們行事對得起那召你們進他自己的國、得他榮耀的上帝。
1THESS|2|13|為此，我們也不斷地感謝上帝，因為你們聽見我們所傳上帝的道的時候，你們領受了，不以為這是人的道，而以為這確實是上帝的道，而且在你們信主的人當中運行著。
1THESS|2|14|弟兄們，你們與 猶太 地區上帝的各教會，就是在基督耶穌裏的各教會，有同樣的遭遇，因為你們也受了同胞的迫害，像他們受了 猶太 人的迫害一樣。
1THESS|2|15|這些 猶太 人不但殺了主耶穌和先知們，又把我們趕出去。他們令上帝不悅，且與眾人為敵，
1THESS|2|16|阻撓我們傳道給外邦人，使他們得救，以致常常惡貫滿盈，但上帝的憤怒終於臨到他們身上。
1THESS|2|17|弟兄們，我們被迫暫時與你們分離，身體離開，心卻沒有；我們極力想法子，渴望見你們的面。
1THESS|2|18|所以我們很想到你們那裏去。我－ 保羅 有一兩次要去，只是撒但阻擋了我們。
1THESS|2|19|當我們的主耶穌再來，我們站在他面前的時候，我們的盼望、喜樂和所誇的冠冕是甚麼呢？不正是你們嗎？
1THESS|2|20|你們就是我們的榮耀和喜樂！
1THESS|3|1|既然我們不能再忍，就決定獨自留在 雅典 ，
1THESS|3|2|於是差派我們在基督福音上作上帝同工的弟兄 提摩太 前去，在你們所信的道上堅固你們，勸勉你們，
1THESS|3|3|免得有人被這些患難動搖。因為你們自己知道，我們受患難原是命定的。
1THESS|3|4|我們在你們那裏的時候，曾預先告訴你們，我們必受患難；你們知道，這果然發生了。
1THESS|3|5|為此，既然我不能再忍，就差派人去，要知道你們的信心如何，恐怕那誘惑人的果真誘惑了你們，以致我們的勞苦歸於徒然。
1THESS|3|6|但是， 提摩太 剛從你們那裏回來，將你們信心和愛心的好消息報給我們，又說你們常常記念我們，切切想見我們，如同我們想見你們一樣。
1THESS|3|7|所以，弟兄們，我們在一切困苦患難中，因著你們的信心得到鼓勵。
1THESS|3|8|如今你們若靠主站立得穩，我們就得生了。
1THESS|3|9|我們在上帝面前，因著你們滿有喜樂。為這一切喜樂，我們能用怎樣的感謝為你們報答上帝呢？
1THESS|3|10|我們晝夜切切祈求要見你們的面，來補足你們信心的不足。
1THESS|3|11|願我們的父上帝自己和我們的主耶穌，為我們開路到你們那裏去。
1THESS|3|12|又願主使你們彼此相愛的心，和愛眾人的心，都能增長，充足，如同我們愛你們一樣，
1THESS|3|13|好堅固你們的心，使你們在我們的主耶穌同他眾聖徒來臨的時候，在我們父上帝面前，成為聖潔，無可指責。阿們！
1THESS|4|1|末了，弟兄們，我們靠著主耶穌求你們，勸你們，既然你們領受了我們的教導，知道該怎樣行事為人，討上帝的喜悅，其實你們也正這樣行，我勸你們要更加努力。
1THESS|4|2|你們原知道，我們憑主耶穌傳給你們甚麼命令。
1THESS|4|3|上帝的旨意就是要你們成為聖潔，遠避淫行；
1THESS|4|4|要你們各人知道怎樣用聖潔、尊貴控制自己的身體 ，
1THESS|4|5|不放縱私慾的邪情，像不認識上帝的外邦人。
1THESS|4|6|不准有人在這事上越軌，佔他弟兄的便宜；因為這一類的事，主必報應，正如我預先對你們說過，又切切警告過你們的。
1THESS|4|7|上帝召我們本不是要我們沾染污穢，而是要我們聖潔。
1THESS|4|8|所以，那棄絕這教導的不是棄絕人，而是棄絕那把自己的聖靈賜給你們的上帝。
1THESS|4|9|有關弟兄間的手足之情，不用人寫信給你們，因為你們自己蒙了上帝的教導要彼此相愛。
1THESS|4|10|你們向全 馬其頓 的眾弟兄固然是這樣行，但我勸弟兄們要更加努力。
1THESS|4|11|要立志過安靜的生活，管自己的事，親手 做工，正如我們從前吩咐你們的，
1THESS|4|12|好使你們的行為能得外人的尊敬，同時也不依賴任何人。
1THESS|4|13|弟兄們，至於已睡了的人，我們不願意你們不知道，恐怕你們憂傷，像那些沒有指望的人一樣。
1THESS|4|14|既然我們信耶穌死了，復活了，那些已經在耶穌裏睡了的人，上帝也必將他們與耶穌一同帶來。
1THESS|4|15|我們照主的話告訴你們一件事：我們這活著還存留到主來臨的人，絕不會在那已經睡了的人之先。
1THESS|4|16|因為，召集令一發，天使長的呼聲一叫，上帝的號角一吹，主必親自從天降臨；那在基督裏死了的人必先復活，
1THESS|4|17|然後我們這些活著還存留的人必和他們一同被提到雲裏，在空中與主相會。這樣，我們就要和主永遠同在。
1THESS|4|18|所以，你們當用這些話彼此勸勉。
1THESS|5|1|弟兄們，關於那時候和日期，不用人寫信給你們，
1THESS|5|2|因為你們自己明明知道，主的日子來到會像賊在夜間突然來到一樣。
1THESS|5|3|人正說平安穩定的時候，災禍忽然臨到他們，如同陣痛臨到懷胎的婦人一樣，他們絕逃脫不了。
1THESS|5|4|弟兄們，你們並不在黑暗裏，那日子不會像賊一樣臨到你們。
1THESS|5|5|你們都是光明之子，都是白晝之子；我們不屬黑夜，也不屬幽暗。
1THESS|5|6|所以，我們不要沉睡，像別人一樣，總要警醒謹慎。
1THESS|5|7|因為睡了的人是在夜間睡，醉了的人是在夜間醉。
1THESS|5|8|但既然我們屬於白晝，就應當謹慎，把信和愛當作護心鏡遮胸，把得救的盼望當作頭盔戴上。
1THESS|5|9|因為上帝不是預定我們受懲罰，而是預定我們藉著我們的主耶穌基督得救。
1THESS|5|10|他替我們死，讓我們無論醒著、睡著，都與他同活。
1THESS|5|11|所以，你們該彼此勸勉，互相造就，正如你們素常做的。
1THESS|5|12|弟兄們，我們勸你們要敬重那些在你們中間勞苦的，就是在主裏面督導你們、勸戒你們的人。
1THESS|5|13|又因他們所做的工作，要以愛心格外尊重他們。你們也要彼此和睦。
1THESS|5|14|弟兄們，我們勸你們，要警戒不守規矩的人，勉勵灰心的人，扶助軟弱的人，對眾人要有耐心。
1THESS|5|15|你們要謹慎，無論是誰都不要以惡報惡，彼此間和對眾人都要追求做好事。
1THESS|5|16|要常常喜樂，
1THESS|5|17|不住地禱告，
1THESS|5|18|凡事謝恩，因為這是上帝在基督耶穌裏向你們所定的旨意。
1THESS|5|19|不要熄滅聖靈；
1THESS|5|20|不要藐視先知的講論。
1THESS|5|21|但凡事要察驗：美善的事要持守，
1THESS|5|22|各樣惡事要禁戒。
1THESS|5|23|願賜平安 的上帝親自使你們完全成聖！願你們的靈、魂、體得蒙保守，在我們的主耶穌基督來臨的時候，完全無可指責。
1THESS|5|24|那召你們的本是信實的，他必成就這事。
1THESS|5|25|弟兄們，請也為 我們禱告。
1THESS|5|26|用聖潔的吻向眾弟兄問安。
1THESS|5|27|我指著主囑咐你們，要把這信宣讀給眾弟兄聽。
1THESS|5|28|願我們的主耶穌基督的恩惠與你們同在！
