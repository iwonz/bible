2SAM|1|1|І сталося по Сауловій смерті, коли Давид вернувся, розбивши Амалика, то він сидів у Ціклаґу два дні.
2SAM|1|2|І сталося третього дня, аж ось прийшов чоловік із табору від Саула, а одежа його роздерта, і порох на його голові. І сталося, як прийшов він до Давида, то впав на землю й поклонився.
2SAM|1|3|І сказав йому Давид: Звідки це ти приходиш? А той відказав: Я втік з Ізраїлевого табору.
2SAM|1|4|І сказав до нього Давид: Що це сталося, розкажи но мені! А той відказав: Народ утік із бою, а також багато з народу попадало й повмирало, і теж Саул та син його Йонатан померли.
2SAM|1|5|А Давид сказав юнакові, що розповідав йому: Як ти пізнав, що помер Саул та син його Йонатан?
2SAM|1|6|І сказав той юнак, що розповідав йому: Припадком натрапив я на горі Ґілбоа, аж ось Саул, настромлений на списа свого, а колесниці та їздці доганяють його.
2SAM|1|7|І він обернувся до мене, і побачив мене, та й покликав мене. А я відповів: Ось я!
2SAM|1|8|І сказав він до мене: Хто ти? А я відказав йому: Я амаликитянин.
2SAM|1|9|І сказав він до мене: Стань надо мною, та й убий мене, бо схопив мене корч, а вся душа ще в мені!...
2SAM|1|10|І став я при ньому, та й убив його, бо я знав, що він не буде живий по упадку своїм. І взяв я вінця, що на голові його, та наплечника, що на плечі його, і приніс сюди до пана свого.
2SAM|1|11|І схопився Давид за одежі свої, та й роздер їх, і теж усі люди, що були з ним.
2SAM|1|12|І голосили вони й плакали, та постили аж до вечора за Саулом та за сином його Йонатаном, і за народом Господнім та за Ізраїлевим домом, що попадали від меча.
2SAM|1|13|І сказав Давид юнакові, що розповідав йому: Звідки ти? А той відказав: Я син одного приходька, амаликитянина.
2SAM|1|14|І сказав йому Давид: Як ти не побоявся простягти руку свою, щоб убити Господнього помазанця?
2SAM|1|15|І покликав Давид одного з слуг своїх і сказав: Підійди, убий його! І той ударив його, і він помер.
2SAM|1|16|І сказав до нього Давид: Кров твоя на голові твоїй, бо уста твої посвідчили проти тебе, говорячи: Я вбив Господнього помазанця.
2SAM|1|17|І Давид заголосив за Саулом та за його сином Йонатаном такою жалобною піснею,
2SAM|1|18|та й сказав навчити Юдиних синів пісні про лука. Ось вона написана в книзі Праведного:
2SAM|1|19|О пишното Ізраїлева, побита із лука на згір'ях своїх, ой попадали лицарі!
2SAM|1|20|Не розказуйте в Ґаті про це, не сповіщайте на вулицях Ашкалону, щоб не тішилися филистимлянські дочки, щоб не раділи дочки необрізаних!
2SAM|1|21|Ґілбоавські гори, щоб на вас не було ні роси, ні дощу, ані поля для жертви принесення! Бо сплямлений там щит хоробрих, щит Саулів, як ніби оливою він не помазаний!
2SAM|1|22|Від крови забитих, від лою хоробрих не відривався був лук Йонатанів, і не вертався меч Саулів напорожньо!
2SAM|1|23|Саул та Йонатан, ці улюблені й милі за свойого життя, і в смерті своїй нерозлучні, прудкіші були від орлів та сильніші від левів!
2SAM|1|24|Дочки Ізраїлеві, за Саулом заплачте, що вас зодягав у багряницю з прикрасами, що оздоблював золотом вашу одежу!
2SAM|1|25|Ой, попадали лицарі посеред бою!... Йонатан на пагірках твоїх ось забитий!
2SAM|1|26|Скорблю по тобі, Йонатане, мій брате! Ти для мене був вельми улюблений, кохання твоє розкішніше для мене було від кохання жіночого!
2SAM|1|27|Ой, попадали лицарі, і загинула зброя військова!...
2SAM|2|1|І сталося потому, і запитався Давид Господа, говорячи: Чи йти мені в одне з Юдиних міст? А Господь відказав йому: Іди! І сказав Давид: Куди я піду? А Він відказав: У Хеврон!
2SAM|2|2|І ввійшов туди Давид, а також дві жінки його: їзреелітка Ахіноам та Авіґаїл, колишня жінка кармелянина Навала.
2SAM|2|3|І людей своїх, що були з ним, привів Давид кожного та дім його, і вони осілися по хевронських містах.
2SAM|2|4|І посходилися Юдині мужі, і помазали там Давида царем над Юдиним домом. А Давидові розповіли, кажучи: Люди ґілеадського Явешу поховали Саула.
2SAM|2|5|І послав Давид людей до ґілеадського Явешу, і сказав до них: Благословенні ви для Господа, що зробили цю милість із своїм паном, із Саулом, та поховали його!
2SAM|2|6|А тепер нехай Господь зробить вам милість та правду, і я теж зроблю вам те добро за те, що ви зробили цю річ.
2SAM|2|7|А тепер нехай зміцняться ваші руки, і будьте мужні, бо помер пан ваш Саул, а також Юдин дім помазав мене царем над собою.
2SAM|2|8|А Авнер, Нерів син, провідник Саулового війська, узяв Іш-Бошета, Саулового сина, та й привів його до Маханаїму.
2SAM|2|9|І він настановив його царем над Ґілеадом, і над Ашуреянином, і над Їзреелем, і над Єфремом, і над Веніямином, і над усім Ізраїлем.
2SAM|2|10|Іш-Бошет, Саулів син, був віку сорока літ, коли зацарював над Ізраїлем, і царював два роки, тільки дім Юди був за Давидом.
2SAM|2|11|А число днів, що Давид був царем у Хевроні над Юдиним домом, сім літ і шість місяців.
2SAM|2|12|І вийшов Авнер, Нерів син, та слуги Іш-Бошета, Саулового сина, з Маханаїму до Ґів'ону.
2SAM|2|13|А Йоав, син Церуї, та Давидові слуги вийшли й зустріли їх разом при ґів'онському ставі. І засіли вони ті з того боку ставу, а ті з цього боку ставу.
2SAM|2|14|І сказав Авнер до Йоава: Нехай встануть ці юнаки, і побавляться перед нами! І сказав Йоав: Нехай встануть.
2SAM|2|15|І встали, і перейшли в числі дванадцяти для Веніямина та для Іш-Бошета, Саулового сина, та дванадцять із Давидових слуг.
2SAM|2|16|І схопили один одного за голову, та й всадили свого меча до боку один одного, і попадали разом. І назвали ім'я тому місцю: Хелкат-Гаццурім, що в Ґів'оні.
2SAM|2|17|І знявся того дня дуже жорстокий бій, і був побитий Авнер та Ізраїлеві люди Давидовими слугами.
2SAM|2|18|І були там три сини Церуї: Йоав, і Авішай, і Асаїл. А Асаїл був легкий в ногах своїх, як польова та газеля.
2SAM|2|19|І гнався Асаїл за Авнером, і не збочував, ані праворуч, ані ліворуч із погоні за Авнером.
2SAM|2|20|І обернувся Авнер позад себе й сказав: Чи це ти, Асаїле? А той відказав: Я.
2SAM|2|21|І сказав йому Авнер: Збоч собі на правицю свою чи на лівицю свою, і схопи собі одного із слуг, і візьми собі зброю його. Та не хотів Асаїл спинити погоні за ним.
2SAM|2|22|А Авнер знов говорив до Асаїла: Спинися в гонитві за мною! Нащо я вб'ю тебе? І як зведу я обличчя своє до брата твого Йоава?
2SAM|2|23|А той відмовився спинитися. І вдарив його Авнер заднім кінцем списа в живіт, і спис вийшов іззаду його! І впав він там, і помер на місці... І сталося, кожен, хто приходив до того місця, де впав Асаїл та помер, то спинявся.
2SAM|2|24|І гналися Йоав та Авішай за Авнером. І сонце зайшло, а вони прийшли до згір'я Амма, що навпроти Ґіаху, на дорозі до Ґів'онської пустині.
2SAM|2|25|І зібралися Веніяминові сини при Авнері, і склали один відділ, та й спинилися на верхів'ї одного взгір'я.
2SAM|2|26|І кликнув Авнер до Йоава й сказав: Чи завжди меч буде жерти? Чи ти не знаєш, що гіркота буде наостанку? І аж доки ти не скажеш народові спинитися в гонитві за своїми братами?
2SAM|2|27|А Йоав відказав: Як живий Бог, коли б ти не сказав був іншого, то ще від ранку народ був би перестав гнатися за братом своїм.
2SAM|2|28|І засурмив Йоав у сурму, і спинився ввесь народ, і не гналися вже за Ізраїлем, і більше вже не воювали.
2SAM|2|29|А Авнер та люди його йшли степом усю ту ніч, і перейшли Йордан, і пройшли ввесь Бітрон, і прийшли до Маханаїму.
2SAM|2|30|І Йоав вернувся з погоні за Авнером, і зібрав увесь народ, і забракло з Давидових слуг дев'ятнадцяти чоловіка та Асаїла.
2SAM|2|31|А Давидові слуги побили з Веніямина та з людей Авнера, три сотні й шістдесят чоловіка, що померли.
2SAM|2|32|І винесли Асаїла, і поховали його в гробі батька його, що в Віфлеємі. І йшли цілу ніч Йоав та люди його, а розсвіло їм у Хевроні.
2SAM|3|1|І була довга та війна між домом Сауловим та між домом Давидовим. А Давид усе зміцнювався, а Саулів дім усе слабнув.
2SAM|3|2|І в Хевроні народилися Давидові сини, і був його первісток Амнон, від їзреелітки Ахіноам;
2SAM|3|3|а другий син його Кіл'ав від Авіґаїл, колишньої жінки кармелянина Навала; а третій Авесалом, син Маахи, дочки Талмая, царя ґешурського;
2SAM|3|4|а четвертий Адонійя, син Хаґґіт, а п'ятий Шефатія, син Авітал,
2SAM|3|5|а шостий Їтреам, від Еґли, Давидової жінки, оці народилися Давидові в Хевроні.
2SAM|3|6|І сталося, коли була війна між домом Сауловим та домом Давидовим, то Авнер тримався Саулового дому.
2SAM|3|7|І мав Саул наложницю, а ім'я їй Ріцпа, дочка Айї. І сказав Іш-Бошет до Авнера: Чого ти прийшов до наложниці батька мого?
2SAM|3|8|І дуже запалився Авнерові гнів на слова Іш-Бошетові, і він сказав: Чи я псяча юдська голова? Сьогодні я роблю ласку домові твого батька Саула, його братам та його приятелям, і не віддав тебе в Давидову руку, а ти сьогодні згадав на мені гріх цієї жінки?
2SAM|3|9|Нехай так зробить Бог Авнерові, і нехай ще додасть йому, якщо я не зроблю Давидові так, як Господь присягнув був йому,
2SAM|3|10|щоб перенести царство від Саулового дому, і щоб поставити Давидів трон над Ізраїлем та над Юдою від Дану й аж до Беер-Шеви.
2SAM|3|11|І той не міг уже відповідати Авнерові ані слова, бо боявся його.
2SAM|3|12|І послав Авнер замість себе послів до Давида сказати: Чия це земля? І ще сказати: Склади ж свою умову зо мною, і ось рука моя буде з тобою, щоб привернути до тебе всього Ізраїля.
2SAM|3|13|А Давид відказав: Добре, я складу з тобою умову! Тільки однієї речі я жадаю від тебе, а саме: ти не побачиш обличчя мого, якщо ти не приведеш Мелхи, Саулової дочки, коли ти прийдеш побачити мене.
2SAM|3|14|І послав Давид послів до Іш-Бошета, Саулового сина, говорячи: Віддай жінку мою Мелху, яку я заручив був собі за сотню крайніх плотів филистимських.
2SAM|3|15|І послав Іш-Бошет, і взяв її від її чоловіка, від Палтіїла, сина Лаїша.
2SAM|3|16|І пішов з нею чоловік її, і все плакав за нею аж до Бахуріму. І сказав до нього Авнер: Іди, вернися! І той вернувся.
2SAM|3|17|А Авнерове слово з Ізраїлевими старшими було таке: Ви вже давно бажаєте мати Давида царем над собою.
2SAM|3|18|А тепер зробіть це, бо Господь сказав був до Давида, говорячи: Рукою Мого раба Давида Я спасу народ Мій, Ізраїля, від руки филистимлян та від руки всіх ворогів його.
2SAM|3|19|І говорив Авнер також до ушей Веніяминових. І також пішов Авнер говорити до ушей Давидових у Хевроні, усе, що добре в очах Ізраїля та в очах усього дому Веніяминового.
2SAM|3|20|І прийшов Авнер до Давида до Хеврону, а з ним двадцятеро люда. І Давид зробив прийняття Авнерові та людям, що з ним.
2SAM|3|21|І сказав Авнер до Давида: Нехай я встану й піду, і приведу до пана, царя мого, усього Ізраїля, а вони складуть із тобою умову, і ти будеш царювати над усім, чого буде жадати душа твоя. І відпустив Давид Авнера, і він пішов із миром.
2SAM|3|22|Аж ось прийшли слуги Давидові та Йоав із походу, і принесли з собою велику здобич. А Авнера не було з Давидом у Хевроні, бо він відпустив його, і той пішов із миром.
2SAM|3|23|А Йоав та все військо, що було з ним, прийшли. І розповіли Йоаву, говорячи: Приходив Авнер, син Нерів, до царя, а він відпустив його, і той пішов із миром.
2SAM|3|24|І прийшов Йоав до царя та й сказав: Що ти зробив? Ось приходив до тебе Авнер, нащо ти відпустив його, і він відійшов?
2SAM|3|25|Ти знаєш Авнера, Нерового сина, він приходив, щоб намовити тебе та щоб вивідати твій вихід та вхід твій, і щоб вивідати все, що ти робиш.
2SAM|3|26|І вийшов Йоав від Давида, і послав посланців за Авнером, і вони завернули його з Бор-Гассіри, а Давид про те не знав.
2SAM|3|27|І вернувся Авнер до Хеврону, а Йоав відвів його в середину брами, щоб поговорити з ним таємно, та й ударив його там у живіт, і той помер за кров брата його Асаїла.
2SAM|3|28|А потім почув про це Давид і сказав: Невинний я та царство моє перед Господом аж навіки в крові Авнера, Нерового сина.
2SAM|3|29|Нехай вона спаде на голову Йоава та на ввесь дім його батька! І нехай не перестає в Йоавовому домі течивий, і прокажений, і той, хто опирається на кия, і хто падає від меча, і хто не має хліба!
2SAM|3|30|А Йоав та брат його Авішай убили Авнера за те, що він забив їхнього брата Асаїла в Ґів'оні в бою.
2SAM|3|31|І сказав Давид до Йоава та до всього народу, що був з ним: Роздеріть вашу одежу, і опережіться веретищем, та й голосіть за Авнером! А цар Давид ішов за марами.
2SAM|3|32|І поховали Авнера в Хевроні, а цар підніс свій голос та й плакав над Авнеровим гробом, і плакав увесь народ.
2SAM|3|33|І заспівав цар жалобну пісню над Авнером та й сказав: Чи Авнер мав загинути смертю негідного?
2SAM|3|34|Твої руки були не пов'язані, не забиті були твої ноги в кайдани, ти впав, як від неправедних падають! І ввесь народ ще більше плакав над ним.
2SAM|3|35|І прийшов увесь народ, щоб намовити Давида покріпитися хлібом ще того дня, та присягнув Давид, говорячи: Нехай так зробить мені Бог, і нехай ще додасть, якщо я перед заходом сонця скуштую хліба або чогобудь!
2SAM|3|36|А ввесь народ довідався про це, і це було добре в їхніх очах, як і все, що робив цар, було добре в очах усього народу.
2SAM|3|37|І того дня довідалися ввесь народ та ввесь Ізраїль, що то не було від царя, щоб забити Авнера, сина Нерового.
2SAM|3|38|І сказав цар своїм слугам: Ото ж знайте, що вождь та великий муж упав цього дня!
2SAM|3|39|А я сьогодні слабий, хоч помазаний цар, а ті люди, сини Церуї, сильніші від мене. Нехай відплатить Господь злочинцеві за його зло!
2SAM|4|1|І почув Саулів син, що помер Авнер у Хевроні, і опустилися руки його, а ввесь Ізраїль збентежився.
2SAM|4|2|А Саулів син мав двох мужів, керівників відділів, ім'я одному Баана, а ім'я другому Рехав, сини бееротянина Ріммона, а Веніяминових синів, бо й Беерот залічений був на Веніямина.
2SAM|4|3|Та повтікали бееротяни до Ґіттаїму, і мешкали там приходьками, і так є аж до цього дня.
2SAM|4|4|А Йонатан, Саулів син, мав кульгавого сина; він був віку п'яти літ, коли прийшла звістка про Саула та Йонатана з Їзреелу. А нянька його несла його й утікала; і сталося, коли вона поспішно втікала, то він упав й окривів. А ім'я його Мефівошет.
2SAM|4|5|І пішли сини бееротянина Ріммона, Рехав та Баана, і ввійшли, як була денна спекота, до Іш-Бошетового дому, а він лежав у південному спочинку.
2SAM|4|6|І ото ввійшли вони аж до середини дому, ніби взяти пшениці, та й ударили його в живіт. І Рехав та брат його Баана втекли.
2SAM|4|7|Отож, увійшли вони до дому, а він лежить на ліжку своїм у своїй спальні, і вони вдарили його, і вбили його, і зняли йому голову. І взяли вони його голову, і йшли степовою дорогою всю ніч.
2SAM|4|8|І принесли вони Іш-Бошетову голову до Давида в Хеврон, та й сказали цареві: Оце голова Іш-Бошета, Саулового сина, твого ворога, що шукав був твоєї душі. І дав Господь цього дня панові моєму, цареві, пімсту над Саулом та над насінням його.
2SAM|4|9|І відповів Давид Рехавові та братові його Баані, синам бееротеянина Ріммона, і сказав їм: Як живий Господь, що визволив душу мою від усякого утиску,
2SAM|4|10|коли того, хто розповів мені, кажучи: Ось помер Саул, а він був в очах своїх, як приємний вісник, я схопив його, і вбив його в Ціклаґу, замість дати йому нагороду за звістку,
2SAM|4|11|тим більше, коли люди несправедливі вбили справедливого чоловіка в домі його на постелі його! А тепер чи я не пошукаю його крови з вашої руки, і не вигублю вас із Краю?
2SAM|4|12|І Давид наказав слугам, і вони вбили їх, і відрубали їхні руки та їхні ноги, та й повісили над ставом у Хевроні. А Іш-Бошетову голову взяли й поховали в Авнеровім гробі в Хевроні.
2SAM|5|1|І посходилися всі Ізраїлеві племена до Давида в Хеврон та й сказали йому: Оце ми кість твоя та тіло твоє ми!
2SAM|5|2|І давніш, коли Саул був царем над нами, ти водив Ізраїля на війну і приводив назад. І Господь тобі сказав: Ти будеш пасти народа Мого, Ізраїля, і ти будеш володарем над Ізраїлем.
2SAM|5|3|І прийшли всі Ізраїлеві старші в Хеврон, а цар Давид склав із ними умову в Хевроні перед Господнім лицем. І помазали вони Давида царем над Ізраїлем.
2SAM|5|4|Давид був віку тридцяти літ, коли став царювати, і сорок літ царював він.
2SAM|5|5|У Хевроні царював він над Юдою сім літ і шість місяців, а в Єрусалимі царював тридцять і три роки над усім Ізраїлем та Юдою.
2SAM|5|6|І пішов цар та люди його до Єрусалиму на Євусеянина, мешканця того Краю. А той сказав Давидові, говорячи: Ти не ввійдеш сюди, хіба повиганяєш сліпих та кривих! А це значить: Давид ніколи не ввійде сюди!
2SAM|5|7|Та Давид здобув твердиню Сіон, він став Давидовим Містом.
2SAM|5|8|І сказав Давид того дня: Кожен, хто заб'є євусеянина, нехай скине до каналу, а з ним і кривих та сліпих, зненавиджених для Давидової душі. Тому говорять: Сліпий та кривий не ввійде до дому!
2SAM|5|9|І осівся Давид у твердині, і назвав ім'я їй: Давидове Місто. І будував Давид навколо від Мілло й усередині.
2SAM|5|10|І Давид ставав усе більшим, а Господь, Бог Саваот, був із ним.
2SAM|5|11|І послав Хірам, цар тирський, послів до Давида, та кедрового дерева, і теслів, і каменярів для стін, і вони збудували дім для Давида.
2SAM|5|12|І пересвідчився Давид, що Господь поставив його міцно царем над Ізраїлем, і що Він підніс царство його ради народу Свого Ізраїля.
2SAM|5|13|А Давид узяв ще наложниць та жінок з Єрусалиму по виході його з Хеврону, і народилися Давидові ще сини та дочки.
2SAM|5|14|А оце імена народжених йому в Єрусалимі: Шаммуа, і Шовав, і Натан, і Соломон,
2SAM|5|15|і Ївхар, і Елішуа, і Нафеґ, і Яфіа,
2SAM|5|16|і Елішама, і Еліяда, і Еліфалет.
2SAM|5|17|І почули филистимляни, що Давида помазали царем над Ізраїлем, і вийшли всі филистимляни, щоб шукати Давида. І Давид почув про це, і зійшов до твердині.
2SAM|5|18|А филистимляни прийшли та розташувалися в долині Рефаїм.
2SAM|5|19|А Давид запитався Господа, говорячи: Чи виходити мені проти филистимлян? Чи даси їх у мою руку? І Господь відказав до Давида: Виходь, бо справді дам филистимлян у руку твою!
2SAM|5|20|І прийшов Давид до Баал-Пераціму. І побив їх там Давид та й сказав: Господь розірвав ворогів моїх передо мною, як розривають води. Тому він назвав ім'я тому місцю: Баал-Перацім.
2SAM|5|21|І вони полишили там своїх божків, а їх забрав Давид та люди його.
2SAM|5|22|А филистимляни знову прийшли та розташувалися в долині Рефаїм.
2SAM|5|23|І запитався Давид Господа, а Він сказав: Не виходь, оточи їх з-позаду, і прийди до них від бальзамового ліска.
2SAM|5|24|І станеться, коли ти почуєш шелест кроку на верховіттях бальзамового ліска, тоді поспішися, бо то тоді вийшов Господь перед тобою, щоб побити филистимський табір.
2SAM|5|25|І Давид зробив так, як наказав йому Господь, і він побив филистимлян від Ґеви аж туди, кудою йти до Ґезера.
2SAM|6|1|А Давид знову зібрав вибране військо в Ізраїлі, тридцять тисяч.
2SAM|6|2|І встав та й пішов Давид та ввесь народ, що був з ним з Юдиного Баалу, щоб винести звідти Божого ковчега, що над ним кличеться Ім'я, Ім'я Господа Саваота, що замешкує на херувимах.
2SAM|6|3|І вони поставили Божого ковчега на нового воза, і винесли його з Авінадавового дому, що в Ґів'ї. А Узза та Ахйо, сини Авінадавові, провадили того нового воза.
2SAM|6|4|І несли його з Авінадавового дому, що в Ґів'ї, і йшли з ковчегом Божим, а Ахйо йшов перед ковчегом.
2SAM|6|5|А Давид та ввесь Ізраїлів дім грали перед Божим лицем усією силою та піснями, і на цитрах, і на арфах, і на бубнах, на гуслах, і на цимбалах.
2SAM|6|6|І прийшли вони аж до Ґорен-Нахону, а Узза простяг руку до Божого ковчегу, і схопив його, бо зноровилась була худоба.
2SAM|6|7|І запалився Господній гнів на Уззу, і Бог уразив його там за цю провину. І він помер там при Божому ковчезі.
2SAM|6|8|І запалився Давидів гнів за те, що Господь покарав Уззу, і він назвав ім'я тому місцю: Перец-Узза, і так воно зветься аж до цього дня.
2SAM|6|9|І Давид злякався Господа того дня та й сказав: Як увійде до мене Господній ковчег?
2SAM|6|10|І не хотів Давид переносити Господнього ковчега до себе, до Давидового Міста, а скерував його Давид до дому ґатянина Овед-Едома.
2SAM|6|11|І пробував Господній ковчег у домі ґатянина Овед-Едома три місяці, і Господь поблагословив Овед-Едома та ввесь його дім.
2SAM|6|12|І донесено цареві Давидові, говорячи: Господь поблагословив дім Овед-Едома та все, що його, ради ковчегу Божого. І пішов Давид, і виніс Божого ковчега з дому Овед-Едома до Давидового Міста з радістю.
2SAM|6|13|І сталося, коли ті, хто ніс Господнього ковчега, ступали шість кроків, то він приносив у жертву вола та відгодовану штуку худоби.
2SAM|6|14|А Давид танцював перед Господнім лицем зо всієї сили. І Давид був оперезаний лляним ефодом.
2SAM|6|15|І Давид та ввесь Ізраїлів дім несли Господнього ковчега з окриком та з сурмленням сурми.
2SAM|6|16|І сталося, коли Господній ковчег увійшов до Давидового Міста, то Мелхола, Саулова дочка, виглядала через вікно, і побачила царя Давида, що танцював та скакав перед Господнім лицем. І вона погордила ним у серці своєму.
2SAM|6|17|І принесли Господнього ковчега, і поставили його на місці його серед намету, що для нього поставив Давид. І приніс Давид цілопалення перед Господнім лицем та жертву мирну.
2SAM|6|18|А коли Давид скінчив приносити цілопалення та мирні жертви, то він поблагословив народ Іменем Господа Саваота.
2SAM|6|19|І він роздав для всього народу, для всього Ізраїлевого натовпу, від чоловіка й аж до жінки, для кожного по одному буханцеві хліба, по одному кавалкові печеного м'яса та по одному виноградному калачеві. І пішов увесь народ кожен до дому свого.
2SAM|6|20|І вернувся Давид, щоб поблагословити свій дім. І вийшла Мелхола, Саулова дочка, навпроти Давида й сказала: Який славний був сьогодні Ізраїлів цар, що обнажався сьогодні на очах невільниць своїх рабів, як обнажується який з пустунів!
2SAM|6|21|І сказав Давид до Мелхоли: Перед лицем Господа, що вибрав мене над твого батька та над увесь дім його, і наказав мені бути володарем над Господнім народом, над Ізраїлем, буду веселитися перед Господнім лицем!
2SAM|6|22|І коли я буду погорджений ще більш від того, і буду низький у своїх очах, то при невільницях, що ти говорила, і при них я буду шанований!
2SAM|6|23|І в Мелхоли, Саулової дочки, по цьому не було їй дитини аж до дня смерти її.
2SAM|7|1|І сталося, коли цар осів у своєму домі, а Господь дав йому відпочинути від усіх ворогів його навколо,
2SAM|7|2|то цар сказав до пророка Натана: Подивися, я сиджу в кедровому домі, а Божий ковчег знаходиться під завісою!
2SAM|7|3|І сказав Натан до царя: Усе, що в серці твоїм, іди й зроби, бо Господь з тобою.
2SAM|7|4|І сталося тієї ночі, і було Господнє слово до Натана, кажучи:
2SAM|7|5|Іди й скажеш до раба Мого, до Давида: Так сказав Господь: Чи ти збудуєш Мені дім на Моє пробування?
2SAM|7|6|Бо Я не пробував у домі від дня виведення Мого Ізраїлевих синів з Єгипту й аж до цього дня, але ходив у наметі та в шатрі.
2SAM|7|7|Скрізь, де ходив Я поміж Ізраїлевими синами, чи промовив Я хоч слово з яким із Ізраїлевих племен, якому наказав Я пасти народа Мого, Ізраїля, говорячи: Чому не збудували ви Мені кедрового дому?
2SAM|7|8|А тепер так скажеш Моєму рабові Давидові: Так сказав Господь Саваот: Я взяв тебе з пасовиська, як ходив ти за отарою, щоб ти став володарем над народом Моїм, над Ізраїлем.
2SAM|7|9|І був Я з тобою в усьому, де ти ходив, і вигубив Я всіх ворогів твоїх з-перед тебе, і зробив тобі велике ім'я, як ім'я великих на землі.
2SAM|7|10|І встановив Я місце для народу Мого, для Ізраїля, і він пробуватиме на своєму місці, і не буде вже непокоєний, і кривдники не будуть більше гнобити його, як перед тим.
2SAM|7|11|А від того дня, як Я настановив суддів над народом Моїм, Ізраїлем, то Я дав тобі мир від усіх ворогів твоїх. І Господь об'являє тобі, що Господь побудує тобі дім.
2SAM|7|12|Коли виповняться твої дні, і ти ляжеш із своїми батьками, то Я поставлю по тобі насіння твоє, що вийде з утроби твоєї, і зміцню його царство.
2SAM|7|13|Він збудує дім для Ймення Мого, а Я зміцню престола його царства навіки.
2SAM|7|14|Я буду йому за Батька, а він буде Мені за сина. Коли він скривить дорогу свою, то Я покараю його людською палицею та поразами людських синів.
2SAM|7|15|Та милість Моя не відхилиться від нього, як відхилив Я її від Саула, якого Я відкинув перед Тобою.
2SAM|7|16|І буде певним твій дім та царство твоє аж навіки перед тобою. Престол твій буде міцно стояти аж навіки!
2SAM|7|17|Як усі ці слова, як усе це видіння, так говорив Натан до Давида.
2SAM|7|18|Тоді прийшов цар Давид, і сів перед Господнім лицем та й сказав: Хто я, Господи Боже, і що мій дім, що Ти привів мене аж сюди?
2SAM|7|19|Та й це ще було мале в очах Твоїх, Господи Боже, і Ти говорив також про Свого раба в будуччині. А це за законом людським, Господи Боже!
2SAM|7|20|І що ще більше говоритиме Давид Тобі? Та Ти знаєш Свого раба, Господи Боже!
2SAM|7|21|Ради слова Свого та за серцем Своїм Ти зробив усю цю величність, звіщаючи це Своєму рабові.
2SAM|7|22|Тому Ти великий, Господи Боже, бо немає такого, як Ти, і немає Бога, окрім Тебе, згідно з усім, що ми чули своїми ушима.
2SAM|7|23|А який є ще один люд на землі, як Твій народ, Ізраїль, щоб Бог приходив викупити його Собі за народ, і щоб установити йому Своє Ймення, і щоб учинити вам цю величність, та страшні речі для Свого Краю ради народу Свого, якого викупив Собі з Єгипту, від людей та від богів його?
2SAM|7|24|І Ти зміцнив Собі народ Свій, Ізраїля, Собі за народ аж навіки, і Ти, Господи, став для них за Бога.
2SAM|7|25|А тепер, Господи Боже, затверди аж навіки те слово, що Ти говорив про Свого раба та про дім його, і вчини, як Ти говорив!
2SAM|7|26|Нехай буде великим Ім'я Твоє аж навіки, щоб говорити: Господь Саваот Бог над Ізраїлем! А дім Твого раба Давида буде міцно стояти перед лицем Твоїм!
2SAM|7|27|Бо Ти, Господи Саваоте, Боже Ізраїлів, об'явив Своєму рабові, говорячи: Збудую тобі дім, тому раб Твій здобувся на відвагу помолитися до Тебе цією молитвою!
2SAM|7|28|А тепер, Господи Боже, Ти Той Бог, а слова Твої будуть правдою, і Ти говорив Своєму рабові це добро.
2SAM|7|29|А тепер зволь поблагословити дім Свого раба, щоб був навіки перед лицем Твоїм, бо Ти, Господи Боже, говорив це, і від Твого благословення буде поблагословлений навіки дім раба Твого!
2SAM|8|1|І сталося по тому, і побив Давид филистимлян, і поконав їх. І взяв Давид керму влади з руки филистимлян.
2SAM|8|2|І побив він Моава, і переміряв їх шнуром, поклав їх на землю, і відміряв два шнури на побиття, а повен шнур на позоставлення при житті. І стали моавитяни Давидовими рабами, які приносили йому данину.
2SAM|8|3|І побив Давид Ґадад'езера, сина Рехова, царя Цови, коли той ішов був відновити владу свою при річці Ефраті.
2SAM|8|4|І здобув Давид від нього тисячу й сім сотень їздців та двадцять тисяч чоловіка пішого. А коням усіх тих колесниць Давид попідрізував жили, і позоставив із того сто колесниць.
2SAM|8|5|І прийшов Арам дамаський, щоб допомогти Гадад'езерові, цареві Цови, та Давид побив в Арамі двадцять і дві тисячі чоловіка.
2SAM|8|6|І настановив Давид залоги в дамаському Арамі, і став Арам для Давида за рабів, що приносили данину йому, а Господь допомагав Давидові в усьому, де він ходив.
2SAM|8|7|І забрав Давид золоті щити, що були в рабів Ґадад'езера, і приніс їх до Єрусалиму.
2SAM|8|8|А з Бетаху та з Беротаю, міст Гадад'езерових, цар Давид узяв дуже багато міді.
2SAM|8|9|А коли почув Тоі, цар Хамоту, що Давид побив усе військо Гадад'езера,
2SAM|8|10|то Тоі послав свого сина Йорама до царя Давида, щоб повітати його, та щоб поблагословити його за те, що він завжди воював з Гадад'езером та побив його, бо Тоі воював проти Гадад'езера. А в руці його були речі золоті, і речі срібні, і речі мідяні.
2SAM|8|11|Також їх присвятив цар Давид Господеві разом зо сріблом та золотом, що він присвятив був із забраного в усіх народів, яких він здобув:
2SAM|8|12|з Араму, і з Моаву, і з синів Аммона, і з филистимлян, і з Амалика, і зо здобичі Гадад'езера, сина Рехова, царя Цови.
2SAM|8|13|І здобув Давид собі ім'я, коли він вернувся з побиття вісімнадцяти тисяч Араму в Беґе-Мелах.
2SAM|8|14|І він поставив залоги в Едомі, в усьому Едомі поставив залоги. І став увесь Едом за рабів для Давида. І допомагав Господь Давидові в усьому, де він ходив.
2SAM|8|15|І царював Давид над усім Ізраїлем, і чинив Давид суд та справедливість для всього народу свого.
2SAM|8|16|А Йоав, син Церуї, був над військом, а Йосафат, син Ахілудів, був канцлером.
2SAM|8|17|А Садок, син Ахітува, та Ахімелех, син Евіятара, були священики, Серая був писарем.
2SAM|8|18|А Беная, син Єгояди, був над Керетянином та над Пелетянином. А Давидові сини були начальниками царського двору.
2SAM|9|1|І сказав Давид: Чи є ще хто, хто позостався з Саулового дому? Я зроблю йому ласку ради Йонатана.
2SAM|9|2|А при Сауловім домі був раб, а ім'я йому Ціва. І покликали його до Давида, а цар сказав йому: Чи ти Ціва? А той відказав: Раб твій!
2SAM|9|3|І сказав цар: Чи нема вже кого з Саулового дому, щоб я зробив йому Божу ласку? І сказав Ціва до царя: Є ще син Йонатанів, кривий на ноги.
2SAM|9|4|І сказав йому цар: Де він? А Ціва відказав цареві: Ось він у домі Махіра, Амміїлового сина, в Ло-Деварі.
2SAM|9|5|І цар Давид послав, і взяв його з дому Махіра, Амміїлового сина, із Ло-Девару.
2SAM|9|6|І прийшов Мефівошет, син Йонатана, Саулового сина, до Давида, і впав на обличчя своє й поклонився. І Давид сказав: Мефівошете! А той відказав: Ось твій раб!
2SAM|9|7|І сказав йому Давид: Не бійся, бо справді зроблю тобі ласку ради батька твого Йонатана, і зверну тобі все поле твого батька Саула. А ти будеш завжди їсти хліб при моєму столі.
2SAM|9|8|А той уклонився й сказав: Що твій раб, що ти звернувся до такого мертвого пса, як я?
2SAM|9|9|А цар кликнув до Ціви, Саулового слуги, і до нього сказав: Усе, що було Саулове та всього його дому, я дав синові твого пана.
2SAM|9|10|І будеш працювати йому на землі ти й сини твої та раби твої. І будеш приносити з урожаю, і буде хліб для сина твого пана, і він буде його їсти. А Мефівошет, син пана твого, буде завжди їсти хліб при моєму столі. А Ціва мав п'ятнадцять синів та двадцять рабів.
2SAM|9|11|І сказав Ціва до царя: Усе, як накаже мій пан цар своєму рабові, так зробить твій раб. А Мефівошет сказав цар буде їсти при моєму столі, як один із царських синів.
2SAM|9|12|А Мефівошет мав малого сина, а ім'я йому Міха. І всі, хто мешкав у домі Ціви, були раби для Мефівошета.
2SAM|9|13|А Мефівошет сидів в Єрусалимі, бо він завжди їв при царському столі. І він був кривий на обидві свої ноги.
2SAM|10|1|І сталося по тому, і помер цар аммонітський, а замість нього зацарював син його Ганун.
2SAM|10|2|І сказав Давид: Зроблю я ласку Ганунові, Нахашевому синові, як батько його зробив був ласку мені. І послав Давид, щоб його порадувати, щодо батька його, через своїх рабів. І прибули Давидові раби до аммонітського краю.
2SAM|10|3|А аммонітські князі сказали до пана свого Гануна: Чи Давид шанує батька твого в очах твоїх тим, що послав тобі потішителів? Чи ж Давид послав до тебе своїх слуг не на те, щоб оглянули місто та щоб його вивідати, а потім знищити його?
2SAM|10|4|І взяв Ганун Давидових слуг, та й оголив половину їхньої бороди, та обрізав їхню одежу на половину, аж до сидіння їх, та й відпустив їх.
2SAM|10|5|І донесли про це Давидові, а він послав назустріч їм, бо ті мужі були дуже осоромлені. І цар їм сказав: Сидіть в Єрихоні, аж поки відросте вам борода, потім повернетесь.
2SAM|10|6|І побачили аммонітяни, що вони зненавиджені в Давида. І аммонітяни послали й найняли Арам-Бет-Рехову й Арам-Цови, двадцять тисяч піхотинців, та царя Маахи, тисячу чоловіка, і тов'ян дванадцять тисяч чоловіка.
2SAM|10|7|А коли Давид прочув про це, то послав Йоава та все лицарське військо.
2SAM|10|8|І повиходили аммонітяни, і встановилися до бою при вході до брами. А Арам-Цова, і Рехов, і Тов'янин, і Мааха, вони самі були на полі.
2SAM|10|9|І побачив Йоав, що бойовий фронт звернений на нього спереду та позаду, то вибрав Ізраїлевих вибраних, та й установив їх навпроти Арама.
2SAM|10|10|А решту народу дав під руку свого брата Авшая, і встановив навпроти аммонітян,
2SAM|10|11|і сказав: Якщо Арам буде сильніший від мене, то будеш мені на поміч, а якщо аммонітяни будуть сильніші від тебе, то я піду допомагати тобі.
2SAM|10|12|Будь мужній, і станьмо міцно за народ наш та за міста нашого Бога, а Господь нехай зробить, що добре в очах Його!
2SAM|10|13|А коли Йоав та народ, що був із ним, підійшли на бій з Арамом, то ті повтікали перед ним.
2SAM|10|14|А аммонітяни побачили, що втік Арам, то й вони повтікали перед Авішаєм, і ввійшли до міста. І вернувся Йоав від аммонітян і ввійшов до Єрусалиму.
2SAM|10|15|А коли побачив Арам, що він побитий Ізраїлем, то вони позбиралися разом.
2SAM|10|16|І послав Гадад'езер, і вивів Арама, що з другого боку Річки, і ввійшли вони до Геламу. А Шовах, провідник Гадад'езерового війська, був перед ними.
2SAM|10|17|І було донесено Давидові, і він зібрав усього Ізраїля, і перейшов Йордан, та прийшов до Геламу. А Арам установився навпроти Давида, і воював із ним.
2SAM|10|18|І побіг Арам перед Ізраїлем, а Давид повбивав з Араму сім сотень колесниць та сорок тисяч верхівців. І вбив він Шоваха, зверхника війська його, і той там помер.
2SAM|10|19|А коли всі царі, підлеглі Гадад'езера, побачили, що вони побиті Ізраїлем, то замирилися з Ізраїлем, і служили йому. І Арам уже боявся допомагати аммонітянам.
2SAM|11|1|І сталося по року, у час виходу царів на війну, то послав Давид Йоава й своїх слуг із ним, та всього Ізраїля, і вони вигубили аммонітян й облягли Раббу. А Давид сидів в Єрусалимі.
2SAM|11|2|І сталося надвечір, і встав Давид із ложа свого, і проходжувався на даху царського дому. І побачив він із даху жінку, що купалася. А та жінка була дуже вродлива.
2SAM|11|3|І послав Давид, і запитався про ту жінку. А посланий сказав: Таж то Вірсавія, Еліямова дочка, жінка хіттеянина Урії!
2SAM|11|4|І послав Давид посланців, і взяв її. І вона прийшла до нього, і він поклався з нею. А вона очистилася з нечистости своєї, і вернулася до свого дому.
2SAM|11|5|І завагітніла та жінка. І послала вона, і донесла Давидові й сказала: Я завагітніла!
2SAM|11|6|А Давид послав до Йоава: Пошли мені хіттеянина Урію. І Йоав послав Урію до Давида.
2SAM|11|7|І прийшов Урія до нього, а Давид запитався про стан Йоава, і про стан народу, і про стан війни.
2SAM|11|8|І сказав Давид до Урії: Іди до свого дому та обмий свої ноги. І вийшов Урія з царського дому, а за ним понесли гостинця царського.
2SAM|11|9|Та Урія спав при вході до царського дому з усіма слугами пана свого, а до свого дому не пішов.
2SAM|11|10|І донесли Давидові, говорячи: Урія не пішов до дому свого. І сказав Давид до Урії: Чи ж не з дороги ти приходиш? Чому ти не пішов до свого дому?
2SAM|11|11|І сказав Урія до Давида: Ковчег і Ізраїль та Юда сидять у шатрах, а пан мій Йоав та раби мого пана таборують на голому полі. А я піду до свого дому, щоб їсти й пити та лежати зо своєю жінкою? Клянуся життям твоїм та життям душі твоєї, що не зроблю я такої речі!
2SAM|11|12|І сказав Давид до Урії: Позостанься тут і сьогодні, а взавтра я відпущу тебе. І позоставався Урія в Єрусалимі того дня та дня другого.
2SAM|11|13|І покликав його Давид, і той їв та пив перед ним, а він підпоїв його. І вийшов він увечорі, щоб покластися на ложі своїм разом зо слугами пана свого, а до дому свого не пішов.
2SAM|11|14|І сталося ранком, і написав Давид листа до Йоава, і послав через Урію.
2SAM|11|15|А в листі тому він написав так: Поставте Урію напереді найтяжчого бою, і відступіте від нього, щоб він був ударений, і помер.
2SAM|11|16|І сталося, коли Йоав обложував місто, то поставив Урію на те місце, про яке знав, що там хоробрі мужі.
2SAM|11|17|І вийшли люди того міста, і воювали з Йоавом, і впали дехто з народу, із Давидових слуг, і повмирали, також хіттеянин Урія.
2SAM|11|18|І послав Йоав, і доніс Давидові про всі справи того бою.
2SAM|11|19|І наказав він послові, говорячи: Як покінчиш ти оповідати цареві про всі справи того бою,
2SAM|11|20|і буде, якщо ти розгніваєш царя, і він скаже тобі: Чого ви так близько підійшли до міста воювати? Чи ви не знали, що будуть кидати на вас з-над муру?
2SAM|11|21|Хто забив був Авімелеха, Єруббешетового сина? Чи не жінка кинула на нього горішнього каменя від жорен з муру, і він помер у Тевеці? Чого ви близько підійшли до муру? То ти скажеш: Помер також хіттеянин Урія.
2SAM|11|22|І пішов посол і прийшов, і доніс Давидові все, що послав був Йоав.
2SAM|11|23|І сказав посол Давидові: Вони стали сильніші за нас, і вийшли проти нас на поле, та ми були переможцями над ними аж до входу в браму.
2SAM|11|24|А стрільці стріляли на твоїх рабів з муру, і померли дехто з царевих рабів, а також помер твій раб хіттеянин Урія.
2SAM|11|25|І сказав Давид до посла: Так скажеш до Йоава: Нехай не буде злою в очах твоїх ця річ, бо меч пожирає то цього, то того. Підсиль війну свою проти міста, та й розвали його! І підбадьор його, Йоава!
2SAM|11|26|І прочула Урієва жінка, що помер її чоловік Урія, і голосила за своїм чоловіком.
2SAM|11|27|А як минула жалоба, то Давид послав, і забрав її до свого дому, і вона стала йому за жінку, і породила йому сина. Та в Господніх очах була злою та річ, що оце зробив був Давид.
2SAM|12|1|І послав Господь Натана до Давида, а він прийшов до нього та й сказав йому: Два чоловіки були в одному місті, один заможний, а один убогий.
2SAM|12|2|У заможного було дуже багато худоби дрібної та худоби великої.
2SAM|12|3|А вбогий нічого не мав, окрім однієї малої овечки, яку він набув та утримував при житті. І росла вона з ним та з синами його разом, із кавалка хліба його їла й з Келіха його пила, та на лоні його лежала, і була йому як дочка.
2SAM|12|4|І прийшов до багатого чоловіка подорожній, та той жалував узяти з худоби своєї дрібної чи з худоби своєї великої, щоб спорядити їжу для подорожнього, що до нього прийшов, і він узяв овечку того вбогого чоловіка, і спорядив її для чоловіка, що до нього прийшов...
2SAM|12|5|І сильно запалав Давидів гнів на того чоловіка, і він сказав до Натана: Як живий Господь, вартий смерти той чоловік, що чинить таке.
2SAM|12|6|А овечку він оплатить чотирикротно, за те, що зробив таку річ, і за те, що не змилосердився.
2SAM|12|7|І сказав Натан до Давида: Ти той чоловік! Так сказав Господь, Бог Ізраїлів: Я помазав тебе над Ізраїлем, і Я спас тебе з Саулової руки.
2SAM|12|8|І дав тобі дім твого пана, та жінок пана твого на лоно твоє, і дав тобі дім Ізраїля та Юди, а якщо цього мало, то додам тобі ще цього та того.
2SAM|12|9|І чому ти зневажив Господнє слово, і вчинив це зло в очах Його? Хіттеянина Урію вбив ти мечем, а його дружину взяв собі за жінку. А його вбив мечем Аммонових синів.
2SAM|12|10|А тепер не відступить меч від твого дому аж навіки за те, що зневажив ти Мене, і взяв дружину хіттеяника Урії, щоб була тобі за жінку.
2SAM|12|11|Так сказав Господь: Ось Я наведу на тебе зло з твого дому, і заберу жінок твоїх на очах твоїх, і дам ближньому твоєму, а він покладеться з жінками твоїми при світлі цього сонця.
2SAM|12|12|Хоч ти вчинив потаємно, а Я зроблю цю річ перед усім Ізраїлем та перед сонцем.
2SAM|12|13|І сказав Давид до Натана: Згрішив я перед Господом! А Натан сказав до Давида: І Господь зняв твій гріх, не помреш!
2SAM|12|14|Та що ти спонукав зневаження Господа цією річчю, то син твій, народжений тобі, конче помре.
2SAM|12|15|І пішов Натан до свого дому, а Господь уразив дитя, що Давидові породила Урієва жінка, і воно захворіло.
2SAM|12|16|А Давид молив Бога за дитинку, і постив Давид, і входив до кімнати, і ночував, поклавшись на землю.
2SAM|12|17|І прийшли старші його дому до нього, щоб підняти його з землі, та він не хотів, і не підкріпився з ними хлібом.
2SAM|12|18|І сталося сьомого дня, і померло те дитя, а Давидові слуги боялися донести йому, що померло те дитя, бо казали: Ось як була та дитина живою, говорили ми до нього, та не слухав він нашого голосу; а як ми скажемо до нього: Померло це дитя, то ще вчинить щось лихе.
2SAM|12|19|А Давид побачив, що слуги його шепочуться поміж собою, і зрозумів Давид, що померло те дитя. І сказав Давид до своїх слуг: Чи не померло те дитя? А ті відказали: Померло.
2SAM|12|20|І звівся Давид із землі, і помився, і намастився, і змінив свою одежу, і ввійшов до Господнього дому та й поклонився. Потому ввійшов до свого дому, і захотів їсти, і поклали йому хліба, і він їв.
2SAM|12|21|І сказали йому слуги його: Що це за річ, яку ти вчинив? Коли те дитя жило, ти постив та плакав; а як померло те дитя, ти встав та й їв хліб?
2SAM|12|22|А він відказав: Коли те дитя ще жило, я постив та плакав, бо казав: Хто знає, може Господь учинить мені милість, і буде жити дитя те?
2SAM|12|23|А тепер, померло воно. Нащо то я б постив? Чи зможу ще повернути його? Я піду до нього, а воно не вернеться до мене...
2SAM|12|24|І потішив Давид жінку свою Вірсавію, і прийшов до неї, і ліг із нею. І вона вродила сина, а він назвав ім'я йому: Соломон. І Господь полюбив його,
2SAM|12|25|і послав пророка Натана, і той назвав ім'я йому: Єдід'я, ради Господа.
2SAM|12|26|А Йоав воював з Раббою аммонітян, і здобув царське місто.
2SAM|12|27|І послав Йоав послів до Давида, і сказав: Воював я з Раббою, і здобув я місто води.
2SAM|12|28|А тепер збери решту народу, і таборуй біля міста, та здобудь його, щоб не здобув те місто я, і щоб не було воно назване моїм ім'ям.
2SAM|12|29|І зібрав Давид увесь народ, і пішов до Рабби, і воював із нею, та й здобув її.
2SAM|12|30|І взяв він корону з голови їхнього царя, а вага її талант золота, та дорогий камінь, і Давид поклав її на свою голову. І він виніс дуже багато здобичі з того міста.
2SAM|12|31|А народ, що був у ньому, він повиводив, і поклав їх під пилку, і під залізні долота та під залізні сокири, і позаганяв їх до цегельняної печі. І так робив він усім аммонітським містам. І вернувся Давид та ввесь народ до Єрусалиму.
2SAM|13|1|І сталося по тому, мав Авесалом, син Давидів, уродливу сестру, а ім'я їй Тамара. І покохав її Амнон, син Давидів.
2SAM|13|2|І вболівав Амнон так, що він аж захворів через свою сестру Тамару, бо вона була дівчина, і Амнонові здавалося трудно щось їй зробити.
2SAM|13|3|А Амнон мав товариша, а ім'я йому Йонадав, син Шім'ї, Давидового брата. І Йонадав був чоловік дуже хитрий.
2SAM|13|4|І він сказав йому: Чого ти, царевичу, такий марний щоранку? Чи ж не розповіси мені? І сказав йому Амнон: Я кохаю Тамару, сестру брата свого Авесалома.
2SAM|13|5|І сказав йому Йонадав: Ляж на ложі своєму, і вдавай хворого. А коли прийде твій батько, щоб побачити тебе, то скажи йому: Нехай прийде сестра моя Тамара, і нехай підкріпить мене хлібом, і нехай зробить на моїх очах ту їжу, щоб я бачив та їв із руки її.
2SAM|13|6|І поклався Амнон, і вдавав хворого, а цар прийшов побачити його. І сказав Амнон до царя: Нехай прийде сестра моя Тамара, і нехай спече на моїх очах два млинці, і я попоїм з її руки.
2SAM|13|7|І послав Давид до Тамари, до дому, говорячи: Іди до дому твого брата Амнона, і приготов йому їжу.
2SAM|13|8|І прийшла Тамара до дому свого брата Амнона, а він лежить. І взяла вона тіста, і замісила, і приготовила на очах його, та й спекла млинці.
2SAM|13|9|І взяла вона сковорідку, і виложила перед ним, та він відмовився їсти. І сказав Амнон: Випровадь від мене всіх людей. І повиходили від нього всі люди.
2SAM|13|10|І сказав Амнон: Принеси їжу до кімнати, і я з'їм із твоєї руки. І взяла Тамара млинці, що приготовила, та й принесла своєму братові Амнонові до кімнати.
2SAM|13|11|І вона принесла до нього, щоб їв, а він схопив її, та й сказав до неї: Ходи, ляж зо мною, моя сестро!...
2SAM|13|12|А вона йому відказала: Ні, брате мій, не безчесть мене, бо не робиться так в Ізраїлі! Не роби цієї гидоти.
2SAM|13|13|І куди я понесу свою ганьбу? А ти станеш, як один із мерзотників в Ізраїлі. Ти переговори з царем, і він не відмовить віддати мене тобі...
2SAM|13|14|Та він не хотів слухати її голосу. І був він сильніший від неї, і збезчестив її, і лежав із нею...
2SAM|13|15|І по цьому дуже зненавидів її Амнон великою ненавистю, бо ця ненависть, якою він зненавидів її, була більша від любови, якою любив її. І сказав до неї Амнон: Уставай, іди собі...
2SAM|13|16|А вона відказав йому: Через це велике зло, по тому, що зробив ти зо мною, хочеш ще вигнати мене? Та він не хотів її слухати.
2SAM|13|17|І покликав він юнака свого, слугу свого, та й сказав: Виженіть оцю від мене геть, і замкни за нею двері...
2SAM|13|18|А на ній була квітчаста туніка, бо так завжди вбиралися царські дочки, панни. І його слуга випровадив її назовні, і замкнув за нею двері.
2SAM|13|19|А Тамара посипала попелом свою голову, а квітчасту туніку, що була на ній, роздерла, і поклала руку свою на голову свою, і все ходила та голосила...
2SAM|13|20|І сказав до неї брат її Авесалом: Чи брат твій Амнон був із тобою? А тепер, сестро моя, мовчи, брат же твій він! Не бери цієї речі до серця свого... І осіла Тамара, знівечена, у домі брата свого Авесалома.
2SAM|13|21|А цар Давид почув про це все, і сильно розгнівався!
2SAM|13|22|І не говорив Авесалом з Амноном ні про добре, ні про зле, бо Авесалом зненавидів Амнона за те, що той збезчестив сестру його Тамару.
2SAM|13|23|І сталося по двох роках, і мав Авесалом стриження овець у Баал-Хацорі, що при Єфремі, і Авесалом закликав усіх царських синів.
2SAM|13|24|І прийшов Авесалом до царя та й сказав: Ось у раба твого стриження, нехай піде цар та раби його з твоїм рабом.
2SAM|13|25|І сказав цар до Авесалома: Ні, сину мій, не підемо ж ми всі, щоб не бути тобі на тяготу. І той сильно просив його, та він не хотів піти, але поблагословив його.
2SAM|13|26|І сказав Авесалом: А як ні, нехай піде з нами брат мій Амнон! І сказав йому цар: Чого від піде з тобою?
2SAM|13|27|Та Авесалом сильно просив його, і він послав з ним Амнона та всіх царських синів.
2SAM|13|28|А Авесалом загадав юнакам своїм, говорячи: Дивіться, як Амнон звеселіє на серці від вина, то скажу вам: Ударте Амнона! і ви вб'єте його. Не бійтеся, чи ж не я загадав вам? Будьте міцні та відважні!...
2SAM|13|29|І зробили Авесаломові юнаки Амнонові, як загадав був Авесалом. А царські сини повставали, і сіли верхи кожен на мула свого, та й повтікали.
2SAM|13|30|І сталося, були вони ще в дорозі, а вістка прийшла до Давида така: Авесалом повбивав усіх царських синів, і не позосталося з них ні одного...
2SAM|13|31|І цар устав, і роздер шати свої, та й упав на землю, і всі слуги його стояли при ньому з роздертими шатами.
2SAM|13|32|І відповів Йонадав, син Шім'ї, Давидового брата, та й сказав: Нехай не каже мій пан: Усіх юнаків, царських синів, повбивали, бо помер тільки сам Амнон. Бо на наказ Авесалома це було вирішене від дня, як той збезчестив сестру його Тамару.
2SAM|13|33|А тепер нехай мій пан цар не кладе на своє серце такого, говорячи: Усі царські сини повмирали, бо помер тільки сам Амнон.
2SAM|13|34|І Авесалом утік. А юнак вартівник звів свої очі й побачив, аж ось численний народ іде дорогою, що була за ним, від боку гори.
2SAM|13|35|І сказав Йонадав до царя: Ось прийшли царські сини, як слово раба твого, так сталося.
2SAM|13|36|І сталося, як скінчив він говорити, аж ось поприходили царські сини, і піднесли свій голос та й плакали. А також цар та всі слуги його плакали вельми ревним плачем...
2SAM|13|37|А Авесалом утік, і пішов до Талмая, Амміхурового сина, царя ґешурського. А Давид був у жалобі за сином своїм усі ті дні.
2SAM|13|38|А Авесалом утік, і пішов до Ґешуру, і пробув там три роки.
2SAM|13|39|І перестав цар Давид гніватися на Авесалома, бо він був зчасом потішений за Амнона, що помер.
2SAM|14|1|А Йоав, син Церуї, пізнав, що цареве серце прихилилося до Авесалома.
2SAM|14|2|І послав Йоав до Текої, і взяв звідти мудру жінку, та й сказав до неї: Удавай жалобу, і вберись у жалобні шати, і не намащуйся оливою, і будеш, як та жінка, що багато днів у жалобі за померлим.
2SAM|14|3|І прийдеш ти до царя, та й скажеш до нього таке то слово. І Йоав поклав ці слова в її уста.
2SAM|14|4|І говорила та текоїтянка до царя, і впала на обличчя своє на землю, і вклонилася та й сказала: Поможи, царю!
2SAM|14|5|І сказав до неї цар: Що тобі? А та відказала: Та я жінка вдова, а чоловік мій помер.
2SAM|14|6|А в невільниці твоєї двоє синів. І посварилися вони обидва в полі, а рятівника між ними не було, і вдарив один одного, та й убив його.
2SAM|14|7|А ось увесь рід устав на невільницю твою та й кажуть: Видай убійника свого брата, і ми вб'ємо його за душу його брата, якого він убив, і вигубимо також спадкоємця. І погасять вони останню іскру мою, яка позосталася, щоб не лишити моєму чоловікові ані ймення, ані нащадків на поверхні землі...
2SAM|14|8|І сказав цар до тієї жінки: Іди до свого дому, а я накажу про тебе.
2SAM|14|9|І сказала та текоїтянка до царя: На мене, пане мій царю, той гріх, та на дім мого батька, а цар та трон його невинні.
2SAM|14|10|І сказав цар: Того, хто буде говорити на тебе, приведеш його до мене, і він більш уже не займе тебе.
2SAM|14|11|Та вона відказала: Нехай згадає цар Господа, Бога свого, щоб не помножити на згубу месника за кров та щоб вони не погубили мого сина. А він відказав: Як живий Господь, не впаде на землю й волосина сина твого!
2SAM|14|12|І сказала та жінка: Нехай но невільниця твоя скаже слово до свого пана царя! А він відказав: Говори!
2SAM|14|13|І сказала та жінка: А чому ти так думаєш проти Божого народу? Бо цар, коли сказав таке слово, сам себе обвинуватив, бо цар не вертає свого вигнанця.
2SAM|14|14|Бо ми конче помремо, і ми як та вода, вилита на землю, що її не зібрати. Та Бог не знищить душі, і Він задумав не відвернути від Себе відігнаного.
2SAM|14|15|І оце тепер прийшла я сказати панові моєму цареві оцю справу, бо той народ настрашив мене. І сказала твоя невільниця: Нехай скажу я цареві, може виконає цар слово своєї невільниці.
2SAM|14|16|Бо цар вислухає, щоб урятувати свою невільницю з руки того чоловіка, що хоче вигубити мене та мого сина разом із Божого спадку.
2SAM|14|17|І сказала твоя невільниця: Нехай станеться слово мого пана царя на втіху мені, бо мій пан цар як Ангол Божий, і розуміє добре та зле. А Господь, Бог твій, буде з тобою!
2SAM|14|18|А цар відповів та й сказав до тієї жінки: Не заховай передо мною нічого, про що я спитаю тебе. І сказала та жінка: Нехай же говорить пан мій цар!
2SAM|14|19|І цар сказав: Чи не Йоавова рука з тобою в усьому цьому? І відповіла та жінка та й сказала: Як жива душа моя, пане мій царю, не можна відхилитися ані праворуч, ані ліворуч від усього, що говорив мій пан цар, бо твій раб Йоав він наказав мені це, і він уклав в уста твоєї невільниці всі ці слова.
2SAM|14|20|Щоб змінити вигляд тієї справи, раб твій Йоав зробив оцю річ. А пан мій мудрий, як мудрий Божий Ангол, щоб знати про все, що на землі.
2SAM|14|21|І сказав цар до Йоава: Ось зробив ти цю річ, тож піди, поверни того юнака, Авесалома!
2SAM|14|22|І впав Йоав на обличчя своє на землю, і поклонився, та й поблагословив царя. І сказав Йоав: Сьогодні раб твій пізнав, що знайшов ласку в очах твоїх, пане мій царю, бо цар виконав прохання свого раба.
2SAM|14|23|І встав Йоав і пішов до Ґешуру, і привів Авесалома до Єрусалиму.
2SAM|14|24|А цар сказав: Нехай він вернеться до свого дому, але обличчя мого не побачить. І вернувся Авесалом до дому свого, та царського обличчя не бачив.
2SAM|14|25|А такого вродливого мужа, як Авесалом, не було в усьому Ізраїлі, щоб був так дуже хвалений, від стопи ноги його й аж до верху голови його не було в ньому вади.
2SAM|14|26|А коли він голив свою голову, а голив він щороку, бо тяжке було волосся на ньому, тому голив його то важив волосся голови своєї на двісті шеклів царської ваги.
2SAM|14|27|І народилися Авесаломові троє синів та одна дочка, а ім'я їй Тамара. Вона була жінка вродлива з вигляду.
2SAM|14|28|І сидів Авесалом в Єрусалимі два роки часу, а царського обличчя не бачив.
2SAM|14|29|І послав Авесалом до Йоава, щоб послати його до царя, та він не хотів прийти до нього. І послав він іще другий раз, та той не хотів прийти.
2SAM|14|30|І сказав він до своїх слуг: Погляньте на Йоавову ділянку поля, що поруч мого, а в нього там ячмінь, ідіть і підпаліть його огнем. І Авесаломові слуги підпалили ту ділянку поля огнем.
2SAM|14|31|Тоді Йоав устав і прийшов до Авесалома до дому, та й сказав йому: Нащо слуги твої підпалили огнем ту мою ділянку поля?
2SAM|14|32|І сказав Авесалом до Йоава: Я ж посилав до тебе, говорячи: Прийди сюди, і нехай я пошлю тебе до царя сказати: Чого я прийшов із Ґешуру? Добре було б мені ще лишатися там. А тепер нехай я побачу царське обличчя, а якщо є на мені гріх, то нехай уб'є мене...
2SAM|14|33|І прийшов Йоав до царя, і розповів йому те. І покликав він Авесалома, а той прийшов до царя та й поклонився йому обличчям своїм до землі. А цар поцілував Авесалома...
2SAM|15|1|І сталося по тому, і завів собі Авесалом повоза та коні, та п'ятдесят чоловіка, що бігали перед ним.
2SAM|15|2|І вставав Авесалом рано, та й ставав при дорозі до брами. І, бувало, кожного чоловіка, що мав суперечку та йшов до царя на суд, то Авесалом кликав його та й питав: З якого ти міста? І той говорив: З одного з Ізраїлевих племен твій раб.
2SAM|15|3|І говорив до нього Авесалом: Дивися, слова твої добрі та слушні, та в царя нема кому тебе вислухати.
2SAM|15|4|І говорив Авесалом: Коли б мене настановлено суддею в Краю, то до мене приходив би кожен чоловік, що мав би суперечку чи судову справу, а я виправдував би його.
2SAM|15|5|І, бувало, коли хто підходив поклонитися йому, то він простягав свою руку, і хапав його та цілував його.
2SAM|15|6|І робив Авесалом, як ось це, усьому Ізраїлеві, хто приходив на суд до царя. І крав Авесалом серця Ізраїлевих людей!
2SAM|15|7|І сталося в кінці сорока літ, і сказав Авесалом до царя: Піду я та виповню обітницю мою, що я обіцяв був Господеві в Хевроні.
2SAM|15|8|Бо раб твій, коли осів був у Ґешурі в Арамі, склав обітницю, говорячи: Якщо Господь справді поверне мене до Єрусалиму, то я буду служити Господеві.
2SAM|15|9|І сказав йому цар: Іди з миром! І той устав та й пішов до Хеврону.
2SAM|15|10|І порозсилав Авесалом вивідувачів по всіх Ізраїлевих племенах, говорячи: Коли ви почуєте сурмлення сурми, то скажете: Зацарював Авесалом у Хевроні!
2SAM|15|11|А з Авесаломом пішли двісті чоловіка з Єрусалиму, що були покликані; а йшли вони в простоті своїй, і нічого не знали.
2SAM|15|12|І послав Авесалом покликати ґілонянина Ахітофела, Давидового дорадника, з його міста з Ґіло, як він мав приносити жертви. І був то сильний бунт, і народ все змножувався з Авесаломом.
2SAM|15|13|І прийшов вісник до Давида, говорячи: Серце ізраїльтян стало за Авесаломом.
2SAM|15|14|І сказав Давид до всіх своїх слуг, що були з ним в Єрусалимі: Уставайте і втікаймо, а то не зможемо втекти перед Авесаломом. Поспішіть відійти, щоб він не поспішив і не догнав нас, і щоб не було нам від нього лиха, і не побив цього міста вістрям меча.
2SAM|15|15|І сказали цареві царські раби: Усе, що вибере наш пан цар, то при тому твої раби!
2SAM|15|16|І вийшов цар та ввесь його дім пішки, а цар позоставив десять жінок наложниць, щоб стерегли дім.
2SAM|15|17|І вийшов цар та ввесь народ пішки, і стали вони в Бет-Гамерхаку.
2SAM|15|18|А всі його слуги йшли перед ним, а також усі керетяни й усі пелетяни та всі ґатяни, шість сотень чоловіка, що прийшли були пішки з Ґату, ішли перед царем.
2SAM|15|19|А цар сказав до ґатянина Іттая: Чого підеш і ти з нами? Вернися, і сиди з тим царем, бо ти чужий та й вигнанець зо свого місця.
2SAM|15|20|Учора прийшов ти, а сьогодні я мав би турбувати тебе йти з нами? А я йду, куди піду, куди доведеться. Вернися, і забери братів своїх із собою. А Господь учинить тобі милість та правду!
2SAM|15|21|І відповів Іттай до царя та й сказав: Як живий Господь і живий мій пан цар, тільки в тому місці, в якому буде мій пан цар, чи то на смерть, чи то на життя, то там буде твій раб!
2SAM|15|22|І сказав Давид до Іттая: Іди й перейди! І перейшов ґатянин Іттай та всі його люди, та всі діти, що були з ним.
2SAM|15|23|А ввесь той Край плакав ревним голосом, і ввесь народ переходив. А цар переходив потік Кедрон, і ввесь народ переходив дорогою до пустині.
2SAM|15|24|А ось ішли й Садок та всі Левити з ним, що несли ковчега Божого заповіту. І вони поставили Божого ковчега, а Евіятар приносив цілопалення, аж поки ввесь народ не вийшов із міста.
2SAM|15|25|І сказав цар до Садока: Поверни Божого ковчега до міста. Якщо я знайду милість у Господніх очах, і Він поверне мене, то я побачу Його та мешкання Його.
2SAM|15|26|А якщо Він скаже так: Не бажаю тебе, ось я: нехай зробить мені, як добре в очах Його.
2SAM|15|27|І сказав цар до священика Садока: Чи ти бачиш це все? Вернися з миром до міста, а син твій Ахімаац та син Евіятарів Йонатан, обидва ваші сини будуть із вами.
2SAM|15|28|Глядіть, я буду проволікати в степах цієї пустині, аж поки не прийде від вас слово, щоб повідомити мене.
2SAM|15|29|І повернув Садок та Евіятар Божого ковчега до Єрусалиму, та й осілися там.
2SAM|15|30|А Давид сходив узбіччям на гору Оливну, та все плакав. А голова його була покрита, і він ішов босий. А ввесь народ, що був із ним, усі позакривали голову свою, і все йшли та плакали...
2SAM|15|31|А Давидові донесли, говорячи: Ахітофел серед зрадників з Авесаломом. І Давид сказав: Господи, учини ж нерозумною Ахітофелову раду!
2SAM|15|32|І сталося, коли вийшов Давид на верхів'я, де вклоняються Богові, аж ось навпроти нього аркеянин Хушай у роздертій туніці, а порох на його голові.
2SAM|15|33|І сказав йому Давид: Якщо ти підеш зо мною, то будеш мені тягарем.
2SAM|15|34|А якщо вернешся до міста й скажеш Авесаломові: Я буду раб твій, о царю! Я був віддавна рабом батька твого, а тепер я твій раб, то зламаєш мені Ахітофелеву раду.
2SAM|15|35|І чи ж не будуть там із тобою священики Садок та Евіятар? І станеться, усяку річ, яку ти почуєш із царевого дому, розповіси священикам Садокові та Евіятарові.
2SAM|15|36|Ось там із ними двоє їхніх синів: Ахімаац у Садока та Йонатан у Евіятара і ви пошлете через них до мене кожне слово, яке почуєте.
2SAM|15|37|І ввійшов Хушай, Давидів друг, до міста. А Авесалом також увійшов до Єрусалиму.
2SAM|16|1|А коли Давид пройшов трохи з верхів'я, аж ось Ціва, Мефівошетів слуга назустріч йому, та пара в'ючених ослів, а на них двісті хлібів, і сто в'язок родзинок, і сто літніх плодів, та бурдюк вина.
2SAM|16|2|І сказав цар до Ціви: Що це тобі? А Ціва відказав: Ці осли для царського дому на їзду, а хліб та літні плоди на їду юнакам, а вино на пиття змученому в пустині.
2SAM|16|3|І сказав цар: А де син твого пана? А Ціва відказав цареві: Он він сидить в Єрусалимі, бо сказав: Сьогодні Ізраїлів дім поверне мені царство мого батька.
2SAM|16|4|І сказав цар до Ціви: Ось тобі все, що в Мефівошета. А Ціва відказав, уклонившись: Нехай я знайду ласку в очах твоїх, пане мій царю.
2SAM|16|5|І прийшов цар Давид до Бахуріму, аж ось виходить ізвідти чоловік з роду Саулового дому, а ім'я йому Шім'ї, син Ґерин. Він ішов і все проклинав.
2SAM|16|6|І він кидав камінням на Давида та на всіх рабів царя Давида, хоч увесь народ та всі лицарі були на правиці його та на лівиці його.
2SAM|16|7|І отак говорив Шім'ї в прокльоні своїм: Іди, іди геть, кривавий переступнику та чоловіче негідний!
2SAM|16|8|Господь обернув на тебе всю кров Саулового дому, що зацарював ти замість нього. І віддав Господь царство в руку сина твого Авесалома, а ти ось у своєму злі, бо ти кривавий переступник!...
2SAM|16|9|І сказав до царя Авішай, син Церуї: Нащо проклинає цей мертвий пес мого пана царя? Піду я, і зітну йому голову!
2SAM|16|10|А цар відказав: Що обходить це мене та вас, сини Церуїні? Що він проклинає, то це Господь йому сказав: Прокляни Давида! А хто скаже: Нащо ти так зробив?
2SAM|16|11|І сказав Давид до Авішая та до всіх своїх слуг: Ось син мій, що вийшов з утроби моєї, шукає моєї душі, а що вже говорити про цього веніяминівця! Дайте йому спокій, і нехай проклинає, бо так наказав йому зробити Господь!
2SAM|16|12|Може зглянеться Господь над моєю бідою, і поверне мені цього дня добром замість його прокляття...
2SAM|16|13|І йшов Давид та люди його дорогою, а Шім'ї йшов узбіччям гори навпроти нього. І він ішов та все проклинав, і кидав камінням на нього, та порошив порохом.
2SAM|16|14|І прийшов цар та ввесь народ, що був із ним, змучені, і відідхнули там.
2SAM|16|15|А Авесалом та ввесь ізраїльський народ увійшли до Єрусалиму, а з ними Ахітофел.
2SAM|16|16|І сталося, як прийшов аркеянин Хушай, Давидів товариш, до Авесалома, то сказав Хушай до Авесалома: Нехай живе цар, нехай живе цар!
2SAM|16|17|І сказав Авесалом до Хушая: Це така ласка твоя з приятелем твоїм? Чому не пішов ти з своїм приятелем?
2SAM|16|18|І сказав Хушай до Авесалома: Ні, бо кого вибрав Господь та цей народ, та кожен Ізраїлів муж, то я буду його, і з ним позостануся.
2SAM|16|19|А подруге, кому я буду служити? Чи ж не синові його? Як служив я батькові твоєму, так буду й тобі.
2SAM|16|20|І сказав Авесалом до Ахітофела: Дайте пораду, що маємо робити.
2SAM|16|21|І сказав Ахітофел до Авесалома: Прийди до наложниць свого батька, яких він позоставив стерегти дім. І коли почує ввесь Ізраїль, що став ти зненавиджений у свого батька, то зміцняться руки всім, хто з тобою.
2SAM|16|22|І розтягли Авесаломові намета на даху, і Авесалом прийшов до наложниць батька свого на очах усього Ізраїля.
2SAM|16|23|А Ахітофелова порада, яку він радив тими днями, була така певна, як питати про Боже слово, така була Ахітофелова порада і для Давида, і для Авесалома!
2SAM|17|1|І сказав Ахітофел до Авесалома: Виберу я дванадцять тисяч чоловіка, і встану, і поженуся цієї ночі за Давидом.
2SAM|17|2|І нападу я на нього, а він змучений та слабосилий, і він затремтить, і повтікає ввесь народ, що з ним, а я вб'ю й самого царя.
2SAM|17|3|І наверну я ввесь народ до тебе; як не буде чоловіка, якого душі ти шукаєш, то ввесь народ буде мати мир.
2SAM|17|4|І була люба ця річ в очах Авесалома та в очах усіх Ізраїлевих старших.
2SAM|17|5|І сказав Авесалом: Поклич теж аркеянина Хушая, та нехай послухаємо, що в устах його, нехай скаже також він.
2SAM|17|6|І прийшов Хушай до Авесалома, а Авесалом сказав до нього, говорячи: Отак говорив Ахітофел. Чи виконаємо слова його? Якщо ні, говори ти.
2SAM|17|7|І сказав Хушай до Авесалома: Не добра та рада, яку цього разу радив Ахітофел.
2SAM|17|8|І сказав Хушай: Ти знаєш батька свого та людей його, що вони лицарі, та розлючені вони, як медведиця, позбавлена на полі дітей. А батько твій вояк, і не буде ночувати з народом.
2SAM|17|9|Ось тепер він ховається в одній з ям, або в іншому місці. І коли б сталося, що хтось упаде серед них, нападаючих, напочатку, а хтобудь почує та скаже: Сталася поразка в народі, який за Авесаломом,
2SAM|17|10|а хоча б він і хоробрий, якого серце як серце лев'яче, то справді ослабне, бо ввесь Ізраїль знає, що батько твій лицар і хоробрі ті, що з ним.
2SAM|17|11|Тому раджу я: нехай конче збереться до тебе ввесь Ізраїль від Дана й аж до Беер-Шеви, многотою як пісок, що над морем, і ти сам підеш до бою.
2SAM|17|12|І прийдемо ми проти нього в одне з місць, та й нападемо на нього, як падає роса на землю, і не позоставимо ані при нім, ані між усіма людьми, що з ним, ані одного.
2SAM|17|13|А якщо він збереться до якого міста, то ввесь Ізраїль занесе на те місто шнури, та й потягнемо його аж до потоку, так, що не залишиться там ані камінчика.
2SAM|17|14|І сказав Авесалом та всі Ізраїлеві мужі: Ліпша рада аркеянина Хушая від ради Ахітофелової! Бо це Господь наказав зламати добру Ахітофелову раду, щоб Господь приніс зло на Авесалома.
2SAM|17|15|І сказав Хушай до священиків Садока та Евіятара: Так і так радив Ахітофел Авесаломові та Ізраїлевим старшим, а я радив так і так.
2SAM|17|16|А тепер швидко пошліть і донесіть Давидові, говорячи: Не ночуй цієї ночі в степах пустині, але конче перейди на той бік, щоб не був поглинутий цар та ввесь народ, що з ним.
2SAM|17|17|А Йонатан та Ахімаац стояли в Ен-Роґелі. І пішла невільниця й розповіла їм, а вони пішли й донесли цареві Давидові, бо не могли ані показатися, ані ввійти до міста.
2SAM|17|18|Та їх побачив один юнак та й доніс Авесаломові. І вони обидвоє швидко пішли, та й увійшли до дому чоловіка в Бахурімі, що мав колодязя на своїм подвір'ї, і спустилися туди.
2SAM|17|19|А жінка тая взяла й розтягла заслону на верху колодязя, і розложила на ньому зерна, і нічого не було пізнано.
2SAM|17|20|І прийшли Авесаломові раби до тієї жінки до дому та й сказали: Де Ахімаац та Йонатан? А жінка та їм сказала:
2SAM|17|21|І сталося по їхньому відході, вони вийшли з колодязя, і пішли та донесли Давидові. І сказали вони до Давида: Уставайте, і переходьте швидко воду, бо отак радив на вас Ахітофел.
2SAM|17|22|І повставали Давид та ввесь народ, що з ним, та до ранішнього світла перейшли Йордан, і не позосталося ані одного, що не перейшов би Йордану.
2SAM|17|23|А коли Ахітофел побачив, що порада його не виконана, то осідлав осла, і встав та й пішов до свого дому, до свого міста. І він зарядив про дім свій, та й повісився, і помер, і був похований у гробі свого батька...
2SAM|17|24|А Давид прийшов до Маханаїму, а Авесалом перейшов Йордан, він та всі Ізраїлеві мужі із ним.
2SAM|17|25|І Авесалом настановив над військом Амасу замість Йоава. А Амаса був син чоловіка, що ім'я йому Їтра, їзрееліт, який увійшов був до Авіґаїл, дочки Нахашової, сестри Церуї, Йоавиної матері.
2SAM|17|26|І таборував Ізраїль та Авесалом у ґілеадському краї.
2SAM|17|27|І сталося, коли Давид прийшов до Маханаїму, то Шові, Нахашів син з аммонітської Рабби, і Махір, Амміелів син з Ло-Девару, і ґілеадянин Барзіллай з Роґеліму
2SAM|17|28|поприносили постелі, і чаші, і ганчарський посуд, і пшениці, і ячменю, і муки, і праженого зерна,
2SAM|17|29|і меду, і масла, і худобу дрібну, і товщу з худоби великої, для Давида та для народу, що з ним, щоб їли, бо сказали: Цей народ голодний і змучений та спрагнений у пустині.
2SAM|18|1|А Давид переглянув народ, що з ним, і настановив над ними тисячників та сотників.
2SAM|18|2|І послав Давид народ, третину під рукою Йоава, і третину під рукою Авішая, сина Церуї, Йоавового брата, а третину під рукою ґатянина Іттая. І сказав цар до народу: Конче піду також і я з вами!
2SAM|18|3|Та народ сказав: Ти не підеш! Бо якщо ми справді втечемо, вони не звернуть на нас уваги. І якщо половина нас повмирає, вони не звернуть на нас уваги, бо ти як нас десять тисяч. А тепер буде ліпше, як будеш допомагати нам із міста.
2SAM|18|4|І сказав до них цар: Що буде добре в очах ваших, зроблю. І став цар при брамі, а ввесь народ повиходив за сотнями та за тисячами.
2SAM|18|5|А цар наказав Йоавові й Авішаєві та Іттаєві, говорячи: Обережно будьте мені з моїм юнаком Авесаломом! А ввесь народ чув, як цар наказав усім провідникам про Авесалома.
2SAM|18|6|І вийшов народ на поле навперейми Ізраїля, і був бій в Єфремовому лісі.
2SAM|18|7|І був побитий там Ізраїлів народ Давидовими рабами. І була там того дня велика поразка, полягло двадцять тисяч!
2SAM|18|8|І поширився там бій по всій тій землі, і того дня більш народу пожер ліс, ніж поїв меч.
2SAM|18|9|І спіткався Авесалом із Давидовими рабами, а Авесалом їхав на мулі. І підбіг мул під гущавину великого дуба, а його волосся заплуталося в дубі, і він опинився між небом та між землею, а мул, що під ним, перебіг...
2SAM|18|10|І побачив це один чоловік, і доніс Йоаву та й сказав: Ось я бачив Авесалома, що висить на дубі.
2SAM|18|11|І сказав Йоав до чоловіка, що доносив йому: Ось ти бачив, а чому ти не вразив його там на землі, а я дав би був тобі десять шеклів срібла та одного пояса.
2SAM|18|12|І сказав той чоловік до Йоава: А коли б я важив на руці своїй навіть тисячу шеклів срібла, не простягну своєї руки на царського сина, бо ми чули на власні вуха, що цар наказав тобі й Авішаєві та Іттаєві, говорячи: Збережіть мені мого юнака Авесалома!
2SAM|18|13|Або коли б я допустився в душі своїй неправди, а всяка річ не затаїться перед царем! то й ти став би проти мене.
2SAM|18|14|І сказав Йоав: Не буду отак зволікати з тобою! І він узяв три стрілі в руку свою, і вбив їх у серце Авесалома, що ще живий висів на середині дуба...
2SAM|18|15|І оточили його десять юнаків, Йоавові зброєноші, і вдарили Авесалома, та й убили його...
2SAM|18|16|І засурмив Йоав у сурму, а народ повернувся з погоні за Ізраїлем, бо Йоав стримав народ.
2SAM|18|17|І взяли вони Авесалома, та й кинули його в лісі до великої ями, і накидали над ним дуже велику могилу з каміння, а ввесь Ізраїль повтікав кожен до намету свого.
2SAM|18|18|А Авесалом узяв був і поставив собі ще за життя свого пам'ятника, що в царській долині, бо він казав: Нема в мене сина, щоб згадувати про ймення моє. І він назвав пам'ятникові ім'я на своє ім'я. І звалось його: Яд-Авесалом, і так зветься він аж до цього дня.
2SAM|18|19|А Ахімаац, Садоків син, сказав: Побіжу я й сповіщу цареві, що Господь визволив його від руки його ворогів.
2SAM|18|20|І сказав йому Йоав: Не ти вісник цього дня, а сповістиш іншого дня. А цього дня не сповістиш тому, що це ж царський син помер.
2SAM|18|21|І сказав Йоав до кушита: Іди, донеси цареві, що ти бачив. А кушит уклонився Йоавові, та й побіг.
2SAM|18|22|А Ахімаац, син Садока, знову сказав до Йоава: А нехай буде, що буде! Побіжу й я за кушитом! Йоав же відказав: Пощо ти побіжиш, мій сину, коли нема доброї вістки?
2SAM|18|23|А нехай буде, що буде, побіжу! І той сказав йому: Біжи! І побіг Ахімаац дорогою рівнини, і випередив кушита.
2SAM|18|24|А Давид сидів між двома брамами. А вартівник пішов на дах брами на мур, і звів свої очі та й побачив, аж ось біжить самітний чоловік.
2SAM|18|25|І кликнув вартівник, і доніс цареві. А цар сказав: Якщо він сам, вістка в устах його! А чоловік усе йшов та зближався.
2SAM|18|26|І побачив вартівник іншого чоловіка, що біг. І кликнув вартівник до сторожа брами й сказав: Ось біжить самітний чоловік. А цар сказав: І цей зо звісткою!
2SAM|18|27|І сказав вартівник: Я бачу біг першого, як біг Ахімааца, Садокового сина. А цар сказав: То чоловік добрий, і приходить з доброю звісткою.
2SAM|18|28|І кликнув Ахімаац, і сказав до царя: Мир! І вклонився він цареві своїм обличчям до землі та й сказав: Благословенний Господь, Бог твій, що видав людей, які піднесли були руку свою проти мого пана царя!
2SAM|18|29|А цар сказав: Чи гаразд із моїм юнаком Авесаломом? І сказав Ахімаац: Я бачив велике замішання, коли Йоав посилав царського раба та мене, твойого раба, та я не знаю, що то...
2SAM|18|30|І сказав цар: Відійди набік, стань отут. І той відійшов набік та й став.
2SAM|18|31|Аж ось приходить кушит. І сказав кушит: Нехай прийме звістку мій пан цар, бо сьогодні визволив тебе Господь від руки всіх повстаючих на тебе.
2SAM|18|32|І сказав цар до кушита: Чи гаразд із моїм юнаком Авесаломом? І сказав кушит: Нехай станетья, як тому юнакові, ворогам мого пана царя та всім, що повстали на тебе на зло!...
2SAM|18|33|(19-1) І затремтів цар, і вийшов на горішній поверх брами, та й заплакав. А коли йшов, то так говорив: Сину мій, Авесаломе, сину мій! Сину мій, Авесаломе! О, якби я був помер замість тебе, Авесаломе! Сину мій, сину мій!...
2SAM|19|1|(19-2) А Йоаву донесено: Ось цар плаче, і зачав жалобу по Авесаломові.
2SAM|19|2|(19-3) І того дня ця перемога обернулася на жалобу для всього народу, бо того дня народ почув, що казали: Засмутився цар за своїм сином!
2SAM|19|3|(19-4) І прокрадався народ того дня, щоб увійти до міста, як прокрадається народ, засоромлений своєю втечею з бою...
2SAM|19|4|(19-5) А цар закрив своє обличчя. І голосив цар сильним голосом: Сину мій, Авесаломе! Авесаломе, сину мій! Сину мій!...
2SAM|19|5|(19-6) І прийшов Йоав до дому царя, та й сказав: Сьогодні ти засоромив обличчя всіх своїх рабів, які сьогодні врятували життя твоє, і життя синів твоїх та дочок твоїх, і життя жінок твоїх, і життя наложниць твоїх,
2SAM|19|6|(19-7) через те, що ти любиш тих, хто тебе ненавидить, і ненавидиш тих, хто тебе любить, бож сьогодні ти виявив, що нема в тебе вождів ані слуг. Бо сьогодні я знаю, що коли б Авесалом був живий, а ми всі сьогодні були мертві, то тоді це було б любе в очах твоїх...
2SAM|19|7|(19-8) А тепер устань, і говори до серця своїх рабів. Бо присягаю Господом, якщо ти не вийдеш, то цієї ночі ніхто не буде ночувати з тобою, і це буде тобі гірше за всяке зло, що приходило на тебе від молодости твоєї аж дотепер!
2SAM|19|8|(19-9) І цар устав та й засів у брамі, а всьому народові донесли, говорячи: Ось цар сидить у брамі! І посходився ввесь народ перед царське обличчя, а Ізраїль повтікав кожен до своїх наметів.
2SAM|19|9|(19-10) І сперечався ввесь народ по всіх Ізраїлевих племенах, говорячи: Цар урятував нас від руки всіх наших ворогів, він же врятував нас із руки филистимлян, а тепер утік із краю перед Авесаломом.
2SAM|19|10|(19-11) А Авесалом, якого ми помазали були над собою, помер на війні. А тепер чого ви зволікаєте щоб вернути царя?
2SAM|19|11|(19-12) І цар Давид послав до священиків, до Садока та до Евіятара, говорячи: Говоріть так до Юдиних старших: Чого ви будете останніми, щоб вернути царя до його дому? А слово всього Ізраїля прийшло вже до царя, до його дому.
2SAM|19|12|(19-13) Ви браття мої, ви кість моя та тіло моє! І чого ви будете останніми, щоб вернути царя?
2SAM|19|13|(19-14) А Амасі скажете: Чи ж ти не кість моя та не тіло моє? Нехай так зробить мені Бог, і нехай ще додасть, якщо ти не будеш у мене вождем війська по всі дні замість Йоава.
2SAM|19|14|(19-15) І прихилив він серце всіх Юдиних мужів, як одного чоловіка. І послали вони до царя: Вернися ти та всі твої слуги!
2SAM|19|15|(19-16) І вернувся цар, і прийшов аж до Йордану, а Юда прийшов до Ґілґалу назустріч цареві, щоб перепровадити царя через Йордан.
2SAM|19|16|(19-17) А Шім'ї, Ґерин син, Веніяминівець, що з Бахуріму, поспішив і зійшов з Юдиними мужами на зустріч царя Давида.
2SAM|19|17|(19-18) І з ним було тисяча чоловіка з Веніямина, та Ціва, слуга Саулового дому, і п'ятнадцятеро синів його та двадцятеро його рабів із ним. І вони перейшли Йордан перед царем.
2SAM|19|18|(19-19) І перейшов порон, щоб перепровадити царський дім та зробити, що було добре в очах його. А Шім'ї, Ґерин син, упав перед царем, як той переходив Йордан,
2SAM|19|19|(19-20) та й цареві сказав: Нехай пан не порахує мені переступу, і не пам'ятай, що раб твій провинився був того дня, коли мій пан цар вийшов був з Єрусалиму, щоб цар не поклав це до серця свого!
2SAM|19|20|(19-21) Бо раб твій знає, що згрішив він, і ось я прийшов сьогодні з усього Йосипового дому перший, щоб вийти зустріти мого пана царя.
2SAM|19|21|(19-22) А Авішай, син Церуїн, відповів та й сказав: Чи ж не буде забитий Шім'ї за те, що проклинав Господнього помазанця?
2SAM|19|22|(19-23) А Давид відказав: Що вам до мене, сини Церуїні, що ви сьогодні стаєте мені за сатану? Чи сьогодні буде забитий хто в Ізраїлі? Хіба ж я не знаю, що сьогодні я цар над Ізраїлем?
2SAM|19|23|(19-24) А до Шім'ї цар сказав: Не помреш! І заприсягнув йому цар.
2SAM|19|24|(19-25) І зійшов спіткати царя й Мефівошет, онук Саулів. А він не оправляв ніг своїх і не оправляв вуса свого, і не оправляв своєї одежі від дня, як цар вийшов, аж до дня, коли він вернувся з миром.
2SAM|19|25|(19-26) І сталося, коли прийшов він до Єрусалиму зустріти царя, то сказав йому цар: Чому ти не пішов зо мною, Мефівошете?
2SAM|19|26|(19-27) А той відказав: Пане мій царю, раб мій обманив мене! Бо я, раб твій, сказав: осідлаю собі осла, і сяду на нього, та й поїду з царем, бо раб твій кульгавий.
2SAM|19|27|(19-28) Та він очернив раба твого перед паном моїм царем. А мій пан цар, немов Божий Ангол, тому зроби, що добре в очах твоїх!
2SAM|19|28|(19-29) Бож хіба ввесь дім батька мого не був вартий смерти перед моїм паном царем? Та ти вмістив раба свого серед їдців свого столу. І яке ж я маю право скаржитися перед царем?
2SAM|19|29|(19-30) І сказав йому цар: Пощо ти говориш іще оці свої слова? Я сказав: ти та Ціва поділите поле.
2SAM|19|30|(19-31) І сказав Мефівошет до царя: Нехай він візьме навіть усе по тому, коли мій пан, цар прийшов із миром до дому свого!.
2SAM|19|31|(19-32) А ґілеадянин Барзіллай зійшов з Роґеліму, і перейшов з царем Йордан, щоб провести його за Йордан.
2SAM|19|32|(19-33) А Барзіллай був дуже старий, віку восьмидесяти літ. І він годував царя, як той сидів був у Маханаїмі, бо він був дуже заможна людина.
2SAM|19|33|(19-34) І сказав цар до Барзіллая: Перейди зо мною, і я буду годувати тебе при собі в Єрусалимі.
2SAM|19|34|(19-35) І сказав Барзіллай до царя: Скільки ще часу життя мого, що я піду з царем до Єрусалиму?
2SAM|19|35|(19-36) Я сьогодні віку восьмидесяти літ. Чи можу я розпізнавати між добрим та злим? Чи розкуштує твій раб, що буду їсти та що буду пити? Чи послухаю я ще голосу співаків та співачок? І пощо буде ще раб твій тягарем для свого пана царя?
2SAM|19|36|(19-37) Трохи перейде твій раб із царем за Йордан. І чого цар висвідчує мені оце?
2SAM|19|37|(19-38) Нехай раб твій вернеться, і нехай помре у своєму місті при гробі батька свого та своєї матері. А ось раб твій, син мій Кімган перейде з паном моїм, із царем, а ти зроби йому, що добре в очах твоїх.
2SAM|19|38|(19-39) І сказав цар: Кімган перейде зо мною, а я зроблю йому, що миле в очах твоїх. І все, що вибереш у мене, я зроблю тобі!
2SAM|19|39|(19-40) І ввесь народ перейшов Йордан, перейшов і цар. І цар поцілував Барзіллая, та й поблагословив його, і той вернувся на своє місце.
2SAM|19|40|(19-41) І перейшов цар до Ґілґалу, а з ним перейшов Кімган та ввесь Юдин народ, і вони перепровадили царя, а також перейшла половина Ізраїлевого народу.
2SAM|19|41|(19-42) Аж ось усі ізраїльтяни прийшли до царя. І сказали вони цареві: Чому вкрали тебе наші браття, люди Юдині, і перепровадили царя та його дім через Йордан, та всіх Давидових людей з ним?
2SAM|19|42|(19-43) І відповіли всі Юдині люди Ізраїлеві: Бо близький цар до нас! І чого то запалився тобі гнів на цю річ? Чи справді з'їли ми що в царя? Чи теж справді він роздав нам які дарунки?
2SAM|19|43|(19-44) І відповіли ізраїльтяни юдеям та й сказали: Нас десять частин у царя, а також і в Давида ми ліпші від вас. Чому ж ви злегковажили нас? Хіба ж не нам було перше слово, щоб вернути царя? Але слово юдеїв було гостріше від слова ізраїльтян.
2SAM|20|1|І трапився там негідний чоловік, а ім'я йому Шева, син Біхрі, веніяминівець. І засурмив він у сурму та й сказав: Немає нам частки в Давиді, і нема нам спадщини у сина Єссеєвого! Ізраїлю, усі до наметів своїх!
2SAM|20|2|І пішов кожен ізраїльтянин від Давида за Шевою, сином Біхрі, а юдеянин позостався при своєму цареві від Йордану й аж до Єрусалиму.
2SAM|20|3|І прийшов Давид до свого дому в Єрусалим. І взяв цар десять жінок наложниць, яких настановив був пильнувати дім, та й віддав їх до дому сторожі; і він їх годував, але до них не приходив. І були вони ув'язнені аж до дня своєї смерти, удівство за життя чоловіка.
2SAM|20|4|І сказав цар до Амаси: Склич мені юдеян у три дні, а ти стань отут!
2SAM|20|5|І пішов Амаса, щоб скликати Юду, та спізнився від означеного часу, про який він умовився.
2SAM|20|6|І сказав Давид до Авішая: Тепер Шева, син Біхрі, зробить нам зло більше від Авесалома. Візьми ти слуг свого пана, та й поженися за ним, щоб він не знайшов собі твердинних міст, і не щез із наших очей.
2SAM|20|7|І вийшли за ним Йоавові люди, і керетянин, і пелетянин та всі лицарі, і повиходили вони з Єрусалиму, щоб гнатися за Шевою, сином Біхрі.
2SAM|20|8|Вони були при великому камені, що в Ґів'оні, а Амаса вийшов проти них. А Йоав був зодягнений в шату свою, а ній пояс із мечем, прип'ятим на стегні його в піхві, з якої легко виходив і входив.
2SAM|20|9|І сказав Йоав до Амаси: Чи гаразд тобі, брате мій? І Йоав узяв правою рукою Амасу за бороду, щоб поцілувати його.
2SAM|20|10|А Амаса не остерігся меча, що був у Йоавовій руці. І той ударив його ним у живіт, і вилив нутро його на землю, і не повторив йому, а той помер... І Йоав та брат його Авішай гналися за Шевою, сином Біхрі.
2SAM|20|11|А один з Йоавових слуг став над ним та й говорив: Хто жадає Йоава, і хто за Давида, за Йоавом!
2SAM|20|12|А Амасу валявся в крові на середині битої дороги. І побачив той чоловік, що ввесь народ став, то стягнув Амасу з битої дороги на поле, і накинув на нього одежину, бо бачив, що кожен приходив до нього та ставав.
2SAM|20|13|Як був він стягнений з битої дороги, пішов кожен чоловік за Йоавом, щоб гнатися за Шевою, сином Біхрі.
2SAM|20|14|А той перейшов серед усіх Ізраїлевих племен до Авелу та до Бет-Маахи, і серед усіх береян, і були вони зібрані, і теж пішли за ним.
2SAM|20|15|А Йоавові люди прийшли й облягли його в Авелі Бет-Маахи, і насипали при місті вала, що стояв на передмур'ї. А ввесь народ, що був з Йоавом, заходився завалити мура.
2SAM|20|16|І покликала мудра жінка з міста: Слухайте, слухайте, скажіть но Йоавові: Підійди сюди, й я буду говорити до тебе!
2SAM|20|17|І він підійшов до неї, а та жінка сказала: Чи ти Йоав? А він відказав: Я. І вона сказала йому: Послухай слів своєї невільниці!. А він відказав: Я слухаю.
2SAM|20|18|І сказала вона, говорячи: Колись треба було переговорювати, а саме, конче запитатися в Авелі, і так закінчили б справу.
2SAM|20|19|Я із спокійних та вірних міст Ізраїля, ти ж шукаєш погубити місто та матерів серед Ізраїля. Пощо ти нищиш спадщину Господню?
2SAM|20|20|А Йоав відповів та й сказав: Борони Боже, борони мене, Боже! Присягаю, що не знищу й не вигублю!
2SAM|20|21|Це не так, бо чоловік з Єфремових гір, Шева, син Біхрі, ім'я йому, підніс свою руку на царя на Давида. Дайте його самого, й я піду від міста. І сказала та жінка до Йоава: Ось голову його кинуть тобі через мур!
2SAM|20|22|І пішла та жінка до всього народу в своїй мудрості, і відрубали голову Шеви, сина Біхрі, та й кинули до Йоава. А той засурмив у сурму, і розійшлися від міста кожен до наметів своїх. А Йоав вернувся в Єрусалим до царя.
2SAM|20|23|І став Йоав над усім Ізраїлевим військом, а Беная, син Єгоядин, над керітянином та над пелетянином;
2SAM|20|24|а Адорам над даниною, а Йосафат, син Ахілудів, був канцлером;
2SAM|20|25|а Сева писарем, а Садок та Евіятар священиками.
2SAM|20|26|А також яірянин Іра був священиком у Давида.
2SAM|21|1|І був голод за днів Давида три роки, рік за роком. І шукав Давид Господнього лиця, а Господь сказав: Кров на Саула та на його дім за те, що повбивав він ґів'онітян.
2SAM|21|2|І покликав цар ґів'онітян та й сказав їм про це. А ґів'онітяни, вони не з Ізраїлевих синів, а з останку амореянина, а Ізраїлеві сини були присягнули їм. Та Саул шукав, щоб повбивати їх через свою горливість для синів Ізраїля та Юди.
2SAM|21|3|І сказав Давид до ґів'онітян: Що я зроблю вам і чим надолужу, щоб ви поблагословили Господню спадщину?
2SAM|21|4|І сказали йому ґів'онітяни: Не треба нам ані срібла, ані золота від Саула та від дому його, і не треба нам забивати чоловіка в Ізраїлі. А він сказав: Що ви скажете, зроблю вам.
2SAM|21|5|І сказали вони до царя: Чоловік той, що вигубив нас, і що замишляв на нас, щоб нас винищити, щоб ми не стали в усій Ізраїлевій границі,
2SAM|21|6|нехай буде нам дано семеро мужа з синів його, і ми повішаємо їх для Господа в Ґів'аті Саула, Господнього вибранця. А цар сказав: Я дам.
2SAM|21|7|Та змилосердився цар над Мефівошетом, сином Йонатана, Саулового сина, через Господню присягу, що була поміж ними, між Давидом та між Йонатаном, Сауловим сином.
2SAM|21|8|І взяв цар двох синів Ріцпи, дочки Айї, яких вона породила Саулові, Армонія та Мефівошета, і п'ятьох синів Мелхоли, Саулової дочки, що вона породила Адріїлові, синові мехолатянина Барзіллая,
2SAM|21|9|та й дав їх у руку ґів'онітян, і вони повішали їх на горі перед Господнім лицем. І впали семеро разом, а були вони побиті в перших днях жнив, коли початок жнив ячменю.
2SAM|21|10|А Ріцпа, дочка Айїна, взяла веретище, і простягла його собі на скелі, і була там від початку жнив аж поки не зійшли на них води з неба, і не дала вона спочити на них птаству небесному вдень, а польовій звірині вночі...
2SAM|21|11|І було донесено Давидові, що зробила Ріцпа, Айїна дочка, Саулова наложниця.
2SAM|21|12|А Давид пішов, і взяв кості Саула та кості сина його Йонатана від господарів ґілеадського Явешу, що викрали були їх із майдану Бет-Шану що їх повісили там филистимляни того дня, коли филистимляни побили Саула в Ґілбоа.
2SAM|21|13|І виніс він звідти кості Саула та кості сина його Йонатана, і зібрали кості повішаних.
2SAM|21|14|І поховали кості Саула та сина його Йонатана в Веніяминовому краї, в Целі, в гробі батька його Кіша. І зробили все, що наказав був цар, і потому Бог був ублаганий Краєм.
2SAM|21|15|І була ще війна филистимлян з Ізраїлем. І зійшов Давид та з ним слуги його, і воювали з филистимлянами. І змучився Давид.
2SAM|21|16|І був Ішбі в Нові, що з нащадків Рафи, а вага його списа три сотні шеклів міді, і оперезаний він був новою зброєю. І він сказав, щоб забити Давида.
2SAM|21|17|Та поміг йому Авішай, син Церуїн, і він ударив филистимлянина, та й забив його. Тоді Давидові люди присягли йому, говорячи: Ти не вийдеш уже з нами на війну, і не погасиш Ізраїлевого світильника!
2SAM|21|18|І сталося потім, і була ще війна в Нові з филистимлянами. Тоді хушанин Сіббехай побив Сафа, що з нащадків Рафи.
2SAM|21|19|І була ще війна в Нові з филистимлянами, і віфлеємець Елханан, син Яаре, і побив ґатянина Ґоліята, а держак списа його був, як ткацький вал.
2SAM|21|20|І була ще війна в Ґаті. А там чоловік великого зросту, що мав на руках та на ногах по шість пальців, числом двадцять і чотири. Також і він був народжений тому Рафі.
2SAM|21|21|І зневажав він Ізраїля, та вбив його Йонатан, син Шім'ї, Давидового брата!
2SAM|21|22|Четверо тих були народжені тому Рафі в Ґаті, і попадали вони від руки Давида та від руки його слуг.
2SAM|22|1|І промовив Давид до Господа слова оцієї пісні того дня, як Господь урятував був його з руки всіх його ворогів та з долоні Саулової,
2SAM|22|2|та й сказав: Господь моя скеля й твердиня моя, і для мене Спаситель Він мій!
2SAM|22|3|Мій Бог моя скеля, сховаюсь я в ній, Він щит мій і ріг, Він спасіння мого, Він башта моя та моє пристановище! Спасителю мій, Ти врятуєш мене від насилля!
2SAM|22|4|Я кличу: Преславний Господь, і я визволений від своїх ворогів!
2SAM|22|5|Бо хвилі смертельні мене оточили, потоки велійяала лякають мене.
2SAM|22|6|Тенета шеолу мене оточили, а пастки смертельні мене попередили!
2SAM|22|7|В тісноті своїй кличу до Господа, і до Бога свого я волаю, І Він почує мій голос із храму Свого, і в ушах Його зойк мій.
2SAM|22|8|Захиталась земля й затремтіла, затряслися й хитались небесні підвалини, бо Він запалився від гніву!
2SAM|22|9|з ніздер Його бухнув дим, з Його ж уст пожирущий огонь, запаливсь жар від Нього!
2SAM|22|10|Він небо простяг і спустився, а хмара густа під ногами Його.
2SAM|22|11|Усівся Він на херувима й летів, і явився на вітряних крилах.
2SAM|22|12|А навколо Себе поклав темряву, мов куріні, збір води, густі хмари високі.
2SAM|22|13|Від блиску, що був перед Ним, запалилось вугілля горюче.
2SAM|22|14|Господь загримів у небесах, і Свій голос Всевишній подав.
2SAM|22|15|Він послав Свої стріли та їх розпорошив, послав блискавку й їх побентежив.
2SAM|22|16|І показалися річища водні, і відкрились основи вселенної, від свару Твойого, о Господи, від подиху вітру із ніздер Його.
2SAM|22|17|Він послав із високости, узяв Він мене, витяг мене з вод великих.
2SAM|22|18|Він мене врятував від мойого потужного ворога, від моїх ненависників, бо сильніші від мене вони.
2SAM|22|19|Напали на мене вони в день нещастя мого, та Господь був моїм опертям.
2SAM|22|20|І на місце широке Він вивів мене, Він мене врятував, бо вподобав мене!
2SAM|22|21|Нехай Господь зробить мені по моїй справедливості, хай заплатить мені згідно з чистістю рук моїх!
2SAM|22|22|Бо беріг я дороги Господні, і від Бога свойого я не відступив,
2SAM|22|23|бо всі Його присуди передо мною, постанови ж Його, не вступлюся від них!
2SAM|22|24|І був я Йому непорочним, і стерігся своєї провини.
2SAM|22|25|Господь заплатив був мені по моїй справедливості, за чистотою моєю перед очима Його.
2SAM|22|26|З справедливим Ти справедливо поводишся, із чесним по-чесному,
2SAM|22|27|із чистим поводишся чисто, а з лукавим за лукавством його!
2SAM|22|28|І народ із біди Ти спасаєш, а очі Твої на зухвалих, яких Ти принижуєш.
2SAM|22|29|Бо світильник Ти, Господи, мій, і освітить Господь мою темряву!
2SAM|22|30|Бо з Тобою поб'ю я ворожого відділа, із Богом своїм проберусь через мур!
2SAM|22|31|Бог непорочна дорога Його, слово Господнє очищене, щит Він для всіх, хто вдається до Нього!
2SAM|22|32|Бо хто Бог, окрім Господа? І хто скеля, крім нашого Бога?
2SAM|22|33|Бог сильне моє пристановище, і дорогу мою Непорочний вивідував.
2SAM|22|34|Він чинить ноги мої, як оленячі, і ставить мене на висотах моїх,
2SAM|22|35|Мої руки навчає до бою, і на рамена мої лука мідяного напинає.
2SAM|22|36|І дав Ти мені щит спасіння Свого, і чинить великим мене Твоя поміч!
2SAM|22|37|Ти чиниш широким мій крок підо мною, і стопи мої не спіткнуться.
2SAM|22|38|Жену я своїх ворогів, і повигублюю їх, і не вернуся, аж поки не винищу їх!
2SAM|22|39|Я їх повигублюю й їх потрощу, і не встануть вони, і повпадають під ноги мої.
2SAM|22|40|Ти ж для бою мене підперізуєш силою, валиш під мене моїх ворохобників.
2SAM|22|41|Повернув Ти плечима до мене моїх ворогів, моїх ненависників, й я їх понищу!
2SAM|22|42|Озирались вони та немає спасителя, кликали до Господа і не відповів їм!
2SAM|22|43|І я їх зітру, як той порох землі, як болото на вулицях їх розітру й розтопчу їх!
2SAM|22|44|Ти ж від бунту народу мойого мене бережеш, на голову люду мене стережеш, мені будуть служити народи, яких я й не знав!
2SAM|22|45|Передо мною чужинці підлещуються, на вістку про мене слухняні мені.
2SAM|22|46|В'януть чужинці, і тремтять у твердинях своїх.
2SAM|22|47|Живий Господь, і благословенна будь, Скеле моя, і нехай піднесеться Бог скелі спасіння мого!
2SAM|22|48|Бог, що помсти за мене дає, і що народи під мене познижував,
2SAM|22|49|що рятує мене від моїх ворогів, Ти звеличив мене над повстанців на мене, спасаєш мене від насильника!
2SAM|22|50|Тому то хвалю Тебе, Господи, серед народів, Іменню Твоєму співаю!
2SAM|22|51|Ти башта спасіння Свойого царя, і милість вчиняєш Своєму помазанцеві, Давиду й насінню його аж навіки!
2SAM|23|1|А оце останні Давидові слова: Слово Давида, сина Єссеєвого, і слово мужа високопоставленого, помазаного Богом Якововим, і солодкого піснотворця Ізраїлевого.
2SAM|23|2|Дух Господній говорить в мені, а слово Його на моїм язику!
2SAM|23|3|Сказав Бог Ізраїлів, Скеля Ізраїлева говорила мені: пануючий серед людей, справедливий панує у Божім страху!
2SAM|23|4|І він буде, як світло поранку безхмарного, коли сонце виходить уранці, як з блиску трава виростає з землі по дощі!
2SAM|23|5|Чи мій дім не такий перед Богом? Вічного бо заповіта в усьому мені там укладено і він стережеться, бо він усе спасіння моє й усе жадання! Хіба Він не дасть, щоб він виріс?
2SAM|23|6|А нечестивий, як терен, відкинений, і вони всі, бо рукою його не беруть.
2SAM|23|7|А хто хоче до них доторкнутись, нехай запасеться залізом чи держаком списа, і на місці своїм огнем будуть попалені!
2SAM|23|8|А оце імена Давидових лицарів: Йошев-Башшевет, тахкемонець, голова ґвардії, він вимахував своїм держаком одним разом на вісім сотень побитих.
2SAM|23|9|По ньому Елеазар, син Додо, сина Ахохі, був серед трьох лицарів з Давидом. Коли филистимляни зневажали ізраїльтян, що зібралися там на війну, і повтікали всі ізраїльтяни,
2SAM|23|10|він устав, та й ударив на филистимлян, аж змучилася рука його, і приліпилася рука його до меча. І зробив Господь велике спасіння того дня, а народ вертався за ним тільки на грабування.
2SAM|23|11|А по ньому Шамма, син Аґе, гарарянин. І зібралися филистимляни до Лехи, а там була ділянка поля, повна сочевиці, а народ повтікав перед филистимлянами.
2SAM|23|12|І став він посередині тієї ділянки та й врятував її, а филистимлян побив. І зробив Господь велике спасіння.
2SAM|23|13|І зійшли троє з тридцяти напочатку, і прийшли в жнива до Давида, до твердині Адуллам. А громада филистимлян таборувала в долині Рефаїм.
2SAM|23|14|Давид же тоді був у твердині, а залога филистимська була тоді в Віфлеємі.
2SAM|23|15|І спрагнув Давид та й сказав: Хто напоїть мене водою з криниці, що в брамі?
2SAM|23|16|І продерлися ці три лицарі до филистимського табору, і зачерпнули води з віфлеємської криниці, що в брамі. І вони винесли, і принесли до Давида, та він не схотів її пити, і вилив її для Господа,
2SAM|23|17|та й сказав: Борони мене, Господи, чинити таке! Чи я буду пити кров тих мужів, що ходили, наражаючи життям своїм? І не хотів він пити її... Оце зробили три ці лицарі.
2SAM|23|18|А Авішай, брат Йоава, Церуїного сина, він голова цих тридцяти. І він вимахував своїм списом над трьома сотнями, що побив. І він мав славу серед тих трьох.
2SAM|23|19|Із тих тридцятьох він був найбільше поважаний, і став він їм за провідника. А до тих трьох не належав.
2SAM|23|20|А Беная, син Єгоядин, син хороброго мужа, багаточинний, з Кавцеїлу, побив двох синів Аріїла моавського. І він зійшов, і забив лева в середині ями сніжного дня.
2SAM|23|21|Також побив він одного єгиптянина, мужа поставного, а в руці цього єгиптянина був спис. І зійшов він до нього з києм, і видер списа з руки того єгиптянина, та й убив його списом його.
2SAM|23|22|Оце зробив Беная, син Єгоядин, і його слава була серед тих трьох лицарів.
2SAM|23|23|З тих тридцяти він був поважніший, а до тих трьох не належав. І Давид призначив його до своєї таємної ради.
2SAM|23|24|Асаїл, Йоавів брат, серед тих тридцяти; Елханан, син Додів, із Віфлеєму;
2SAM|23|25|Шамма хародянин, Еліка хародянин,
2SAM|23|26|Хелец цалтянин; Іра, син Іквешів, текоїтянин;
2SAM|23|27|Авіезер аннетотянин, Мевуннай хушатянин,
2SAM|23|28|Цалмон ахохянин, Магарай нетофатянин,
2SAM|23|29|Хелев, син Баанин, нетофатянин; Іттай, син Ріваїв, міґґів'атянин, сини Веніяминові;
2SAM|23|30|Беная пір'ятонянин, Гіддай з Нахале-Ґаашу,
2SAM|23|31|Аві-Алвон арватянин, Азмавет бархум'янин,
2SAM|23|32|Ел'яхба шаалвонянин, сини Яшемові, Йонатан,
2SAM|23|33|Шамма гарарянин; Ахіам, син Шарарів, арарянин;
2SAM|23|34|Еліфелет, син Ахасбаїв, сина маахатянина; Еліям, син Ахітофелів, ґіллонянин;
2SAM|23|35|Хецрав кармелянин, Паарай арб'янин,
2SAM|23|36|Їґ'ал, син Натанів, з Цови; Бані ґадянин,
2SAM|23|37|Целек аммонеянин; Нахарай бееротянин, зброєноша Йоава, сина Церуїного;
2SAM|23|38|Іра їтрянин, Ґарев їтрянин,
2SAM|23|39|Урія хіттянин, усіх тридцять і сім.
2SAM|24|1|І знову запалився Господній гнів на Ізраїля, і намовив сатана Давида проти них, говорячи: Іди, перелічи Ізраїля та Юду!
2SAM|24|2|І сказав цар до Йоава, вождя війська, що з ним: Перемандруй серед усіх Ізраїлевих племен від Дану аж до Беер-Шеви, і перелічіть народ, і я пізнаю число цього народу.
2SAM|24|3|І сказав Йоав до царя: Нехай же Господь, Бог твій, додасть до народу в сто раз стільки, скільки є, а очі мого пана, царя, бачать. Та нащо пан мій, цар, уподобав собі таку річ?
2SAM|24|4|Та цареве слово до Йоава та на військових провідників перемогло. І вийшов Йоав та військові провідники від царя, щоб перелічити Ізраїлів народ.
2SAM|24|5|І перейшли вони Йордан, і таборували в Ароері, з правого боку міста, що лежить в середині долини Ґаду та при Язері.
2SAM|24|6|І прийшли вони до Ґілеаду та до краю Тахтім-Ходші. І прийшли до Дан-Яану, і навколо до Сидону.
2SAM|24|7|І прийшли вони до твердині Цор й до всіх міст хіввеянина та ханаанеянина, і вийшли до Юдиного Неґеву, до Беер-Шеви.
2SAM|24|8|І мандрували вони по цілому краю, і прийшли в кінці дев'яти місяців та двадцяти днів до Єрусалиму.
2SAM|24|9|І дав Йоав цареві число переліку народу. І було Ізраїля вісімсот тисяч сильних мужів, що витягають меча, а Юдиного мужа п'ятьсот тисяч чоловіка.
2SAM|24|10|І збентежилося Давидове серце, як перелічив він народ. І сказав Давид до Господа: Я дуже згрішив, що зробив це! А тепер, Господи, відсунь же провину Свого раба, бо я дуже немудро вчинив!...
2SAM|24|11|І встав Давид рано вранці, а Господнє слово було до пророка Ґада, Давидового прозорливця, говорячи:
2SAM|24|12|Іди, та й скажеш Давидові: Так сказав Господь: Три карі кладу Я на тебе, вибери собі одну з них, і Я зроблю її тобі.
2SAM|24|13|І прийшов Ґад до Давида, і розповів йому та й до нього сказав: Чи прийдуть тобі сім літ голоду в твоїм краї, чи теж три місяці твого втікання перед ворогами твоїми, а вони тебе гнатимуть, чи теж буде три дні моровиця в твоїм Краї? Подумай тепер та й ріши, яке слово верну я Тому, Хто послав мене.
2SAM|24|14|І сказав Давид до Ґада: Сильно скорблю я! Нехай же впадемо ми до Господньої руки, бо велике Його милосердя, а в руку людську нехай я не впаду!...
2SAM|24|15|І дав Господь моровицю в Ізраїлі від ранку й аж до часу умовлення, і померло з народу від Дану й аж до Беер-Шеви сімдесят тисяч чоловіка...
2SAM|24|16|І простяг той Ангол свою руку на Єрусалима, щоб вигубити його, та Господь пожалував щодо того зла. І сказав Він до Ангола, що вигубляв серед народу: Забагато тепер, попусти свою руку! А Ангол Господній був при тоці євусеянина Аравни.
2SAM|24|17|І сказав Давид до Господа, коли побачив того Ангола, що побивав серед народу, і проказав: Я ось згрішив, і пішов проти Закону. А ці вівці, що зробили вони? Нехай же рука Твоя буде на мені та на домі батька мого!...
2SAM|24|18|І прийшов того дня Ґад до Давида, та й сказав йому: Устань, постав Господеві жертівника на току євусеянина Аравни.
2SAM|24|19|І пішов Давид за словами Ґадовими, як наказав був Господь.
2SAM|24|20|І виглянув Аравна, і побачив царя та його слуг, що йдуть до нього. І вийшов Аравна, і вклонився цареві обличчям своїм до землі.
2SAM|24|21|І сказав Аравна: Чого прийшов пан мій, цар, до свого раба? А Давид відказав: Купити від тебе цього тока, щоб збудувати жертівника для Господа, і буде стримана зараза від народу.
2SAM|24|22|І сказав Аравна до Давида: Нехай пан мій, цар, візьме, і нехай принесе жертву, що добре в очах його. Дивися, ось худоба на цілопалення, а молотілки та ярма на дрова.
2SAM|24|23|Усе віддає Аравна, о царю, цареві. І сказав Аравна до царя: Господь, Бог твій, нехай уподобає Собі тебе!
2SAM|24|24|І сказав цар до Аравни: Ні, бо тільки куплю від тебе за ціну, і не принесу дармо цілопалень Господеві, Богові моєму. І купив Давид тока й худобу за срібло п'ятидесяти шеклів.
2SAM|24|25|І Давид збудував там жертівника для Господа, і приніс цілопалення та мирні жертви. І Господь був ублаганий для Краю, і була стримана зараза від Ізраїля.
