1THESS|1|1|Paul, Silvanus, and Timothy, To the church of the Thessalonians in God the Father and the Lord Jesus Christ: Grace to you and peace.
1THESS|1|2|We give thanks to God always for all of you, constantly mentioning you in our prayers,
1THESS|1|3|remembering before our God and Father your work of faith and labor of love and steadfastness of hope in our Lord Jesus Christ.
1THESS|1|4|For we know, brothers loved by God, that he has chosen you,
1THESS|1|5|because our gospel came to you not only in word, but also in power and in the Holy Spirit and with full conviction. You know what kind of men we proved to be among you for your sake.
1THESS|1|6|And you became imitators of us and of the Lord, for you received the word in much affliction, with the joy of the Holy Spirit,
1THESS|1|7|so that you became an example to all the believers in Macedonia and in Achaia.
1THESS|1|8|For not only has the word of the Lord sounded forth from you in Macedonia and Achaia, but your faith in God has gone forth everywhere, so that we need not say anything.
1THESS|1|9|For they themselves report concerning us the kind of reception we had among you, and how you turned to God from idols to serve the living and true God,
1THESS|1|10|and to wait for his Son from heaven, whom he raised from the dead, Jesus who delivers us from the wrath to come.
1THESS|2|1|For you yourselves know, brothers, that our coming to you was not in vain.
1THESS|2|2|But though we had already suffered and been shamefully treated at Philippi, as you know, we had boldness in our God to declare to you the gospel of God in the midst of much conflict.
1THESS|2|3|For our appeal does not spring from error or impurity or any attempt to deceive,
1THESS|2|4|but just as we have been approved by God to be entrusted with the gospel, so we speak, not to please man, but to please God who tests our hearts.
1THESS|2|5|For we never came with words of flattery, as you know, nor with a pretext for greed- God is witness.
1THESS|2|6|Nor did we seek glory from people, whether from you or from others, though we could have made demands as apostles of Christ.
1THESS|2|7|But we were gentle among you, like a nursing mother taking care of her own children.
1THESS|2|8|So, being affectionately desirous of you, we were ready to share with you not only the gospel of God but also our own selves, because you had become very dear to us.
1THESS|2|9|For you remember, brothers, our labor and toil: we worked night and day, that we might not be a burden to any of you, while we proclaimed to you the gospel of God.
1THESS|2|10|You are witnesses, and God also, how holy and righteous and blameless was our conduct toward you believers.
1THESS|2|11|For you know how, like a father with his children,
1THESS|2|12|we exhorted each one of you and encouraged you and charged you to walk in a manner worthy of God, who calls you into his own kingdom and glory.
1THESS|2|13|And we also thank God constantly for this, that when you received the word of God, which you heard from us, you accepted it not as the word of men but as what it really is, the word of God, which is at work in you believers.
1THESS|2|14|For you, brothers, became imitators of the churches of God in Christ Jesus that are in Judea. For you suffered the same things from your own countrymen as they did from the Jews,
1THESS|2|15|who killed both the Lord Jesus and the prophets, and drove us out, and displease God and oppose all mankind
1THESS|2|16|by hindering us from speaking to the Gentiles that they might be saved- so as always to fill up the measure of their sins. But God's wrath has come upon them at last!
1THESS|2|17|But since we were torn away from you, brothers, for a short time, in person not in heart, we endeavored the more eagerly and with great desire to see you face to face,
1THESS|2|18|because we wanted to come to you- I, Paul, again and again- but Satan hindered us.
1THESS|2|19|For what is our hope or joy or crown of boasting before our Lord Jesus at his coming? Is it not you?
1THESS|2|20|For you are our glory and joy.
1THESS|3|1|Therefore when we could bear it no longer, we were willing to be left behind at Athens alone,
1THESS|3|2|and we sent Timothy, our brother and God's coworker in the gospel of Christ, to establish and exhort you in your faith,
1THESS|3|3|that no one be moved by these afflictions. For you yourselves know that we are destined for this.
1THESS|3|4|For when we were with you, we kept telling you beforehand that we were to suffer affliction, just as it has come to pass, and just as you know.
1THESS|3|5|For this reason, when I could bear it no longer, I sent to learn about your faith, for fear that somehow the tempter had tempted you and our labor would be in vain.
1THESS|3|6|But now that Timothy has come to us from you, and has brought us the good news of your faith and love and reported that you always remember us kindly and long to see us, as we long to see you-
1THESS|3|7|for this reason, brothers, in all our distress and affliction we have been comforted about you through your faith.
1THESS|3|8|For now we live, if you are standing fast in the Lord.
1THESS|3|9|For what thanksgiving can we return to God for you, for all the joy that we feel for your sake before our God,
1THESS|3|10|as we pray most earnestly night and day that we may see you face to face and supply what is lacking in your faith?
1THESS|3|11|Now may our God and Father himself, and our Lord Jesus, direct our way to you,
1THESS|3|12|and may the Lord make you increase and abound in love for one another and for all, as we do for you,
1THESS|3|13|so that he may establish your hearts blameless in holiness before our God and Father, at the coming of our Lord Jesus with all his saints.
1THESS|4|1|Finally, then, brothers, we ask and urge you in the Lord Jesus, that as you received from us how you ought to live and to please God, just as you are doing, that you do so more and more.
1THESS|4|2|For you know what instructions we gave you through the Lord Jesus.
1THESS|4|3|For this is the will of God, your sanctification: that you abstain from sexual immorality;
1THESS|4|4|that each one of you know how to control his own body in holiness and honor,
1THESS|4|5|not in the passion of lust like the Gentiles who do not know God;
1THESS|4|6|that no one transgress and wrong his brother in this matter, because the Lord is an avenger in all these things, as we told you beforehand and solemnly warned you.
1THESS|4|7|For God has not called us for impurity, but in holiness.
1THESS|4|8|Therefore whoever disregards this, disregards not man but God, who gives his Holy Spirit to you.
1THESS|4|9|Now concerning brotherly love you have no need for anyone to write to you, for you yourselves have been taught by God to love one another,
1THESS|4|10|for that indeed is what you are doing to all the brothers throughout Macedonia. But we urge you, brothers, to do this more and more,
1THESS|4|11|and to aspire to live quietly, and to mind your own affairs, and to work with your hands, as we instructed you,
1THESS|4|12|so that you may live properly before outsiders and be dependent on no one.
1THESS|4|13|But we do not want you to be uninformed, brothers, about those who are asleep, that you may not grieve as others do who have no hope.
1THESS|4|14|For since we believe that Jesus died and rose again, even so, through Jesus, God will bring with him those who have fallen asleep.
1THESS|4|15|For this we declare to you by a word from the Lord, that we who are alive, who are left until the coming of the Lord, will not precede those who have fallen asleep.
1THESS|4|16|For the Lord himself will descend from heaven with a cry of command, with the voice of an archangel, and with the sound of the trumpet of God. And the dead in Christ will rise first.
1THESS|4|17|Then we who are alive, who are left, will be caught up together with them in the clouds to meet the Lord in the air, and so we will always be with the Lord.
1THESS|4|18|Therefore encourage one another with these words.
1THESS|5|1|Now concerning the times and the seasons, brothers, you have no need to have anything written to you.
1THESS|5|2|For you yourselves are fully aware that the day of the Lord will come like a thief in the night.
1THESS|5|3|While people are saying, "There is peace and security," then sudden destruction will come upon them as labor pains come upon a pregnant woman, and they will not escape.
1THESS|5|4|But you are not in darkness, brothers, for that day to surprise you like a thief.
1THESS|5|5|For you are all children of light, children of the day. We are not of the night or of the darkness.
1THESS|5|6|So then let us not sleep, as others do, but let us keep awake and be sober.
1THESS|5|7|For those who sleep, sleep at night, and those who get drunk, are drunk at night.
1THESS|5|8|But since we belong to the day, let us be sober, having put on the breastplate of faith and love, and for a helmet the hope of salvation.
1THESS|5|9|For God has not destined us for wrath, but to obtain salvation through our Lord Jesus Christ,
1THESS|5|10|who died for us so that whether we are awake or asleep we might live with him.
1THESS|5|11|Therefore encourage one another and build one another up, just as you are doing.
1THESS|5|12|We ask you, brothers, to respect those who labor among you and are over you in the Lord and admonish you,
1THESS|5|13|and to esteem them very highly in love because of their work. Be at peace among yourselves.
1THESS|5|14|And we urge you, brothers, admonish the idle, encourage the fainthearted, help the weak, be patient with them all.
1THESS|5|15|See that no one repays anyone evil for evil, but always seek to do good to one another and to everyone.
1THESS|5|16|Rejoice always,
1THESS|5|17|pray without ceasing,
1THESS|5|18|give thanks in all circumstances; for this is the will of God in Christ Jesus for you.
1THESS|5|19|Do not quench the Spirit.
1THESS|5|20|Do not despise prophecies,
1THESS|5|21|but test everything; hold fast what is good.
1THESS|5|22|Abstain from every form of evil.
1THESS|5|23|Now may the God of peace himself sanctify you completely, and may your whole spirit and soul and body be kept blameless at the coming of our Lord Jesus Christ.
1THESS|5|24|He who calls you is faithful; he will surely do it.
1THESS|5|25|Brothers, pray for us.
1THESS|5|26|Greet all the brothers with a holy kiss.
1THESS|5|27|I put you under oath before the Lord to have this letter read to all the brothers.
1THESS|5|28|The grace of our Lord Jesus Christ be with you.
