OBAD|1|1|The vision of Obadiah. Thus saith the Lord GOD concerning Edom; We have heard a rumour from the LORD, and an ambassador is sent among the heathen, Arise ye, and let us rise up against her in battle.
OBAD|1|2|Behold, I have made thee small among the heathen: thou art greatly despised.
OBAD|1|3|The pride of thine heart hath deceived thee, thou that dwellest in the clefts of the rock, whose habitation is high; that saith in his heart, Who shall bring me down to the ground?
OBAD|1|4|Though thou exalt thyself as the eagle, and though thou set thy nest among the stars, thence will I bring thee down, saith the LORD.
OBAD|1|5|If thieves came to thee, if robbers by night, (how art thou cut off!) would they not have stolen till they had enough? if the grapegatherers came to thee, would they not leave some grapes?
OBAD|1|6|How are the things of Esau searched out! how are his hidden things sought up!
OBAD|1|7|All the men of thy confederacy have brought thee even to the border: the men that were at peace with thee have deceived thee, and prevailed against thee; that they eat thy bread have laid a wound under thee: there is none understanding in him.
OBAD|1|8|Shall I not in that day, saith the LORD, even destroy the wise men out of Edom, and understanding out of the mount of Esau?
OBAD|1|9|And thy mighty men, O Teman, shall be dismayed, to the end that every one of the mount of Esau may be cut off by slaughter.
OBAD|1|10|For thy violence against thy brother Jacob shame shall cover thee, and thou shalt be cut off for ever.
OBAD|1|11|In the day that thou stoodest on the other side, in the day that the strangers carried away captive his forces, and foreigners entered into his gates, and cast lots upon Jerusalem, even thou wast as one of them.
OBAD|1|12|But thou shouldest not have looked on the day of thy brother in the day that he became a stranger; neither shouldest thou have rejoiced over the children of Judah in the day of their destruction; neither shouldest thou have spoken proudly in the day of distress.
OBAD|1|13|Thou shouldest not have entered into the gate of my people in the day of their calamity; yea, thou shouldest not have looked on their affliction in the day of their calamity, nor have laid hands on their substance in the day of their calamity;
OBAD|1|14|Neither shouldest thou have stood in the crossway, to cut off those of his that did escape; neither shouldest thou have delivered up those of his that did remain in the day of distress.
OBAD|1|15|For the day of the LORD is near upon all the heathen: as thou hast done, it shall be done unto thee: thy reward shall return upon thine own head.
OBAD|1|16|For as ye have drunk upon my holy mountain, so shall all the heathen drink continually, yea, they shall drink, and they shall swallow down, and they shall be as though they had not been.
OBAD|1|17|But upon mount Zion shall be deliverance, and there shall be holiness; and the house of Jacob shall possess their possessions.
OBAD|1|18|And the house of Jacob shall be a fire, and the house of Joseph a flame, and the house of Esau for stubble, and they shall kindle in them, and devour them; and there shall not be any remaining of the house of Esau; for the LORD hath spoken it.
OBAD|1|19|And they of the south shall possess the mount of Esau; and they of the plain the Philistines: and they shall possess the fields of Ephraim, and the fields of Samaria: and Benjamin shall possess Gilead.
OBAD|1|20|And the captivity of this host of the children of Israel shall possess that of the Canaanites, even unto Zarephath; and the captivity of Jerusalem, which is in Sepharad, shall possess the cities of the south.
OBAD|1|21|And saviours shall come up on mount Zion to judge the mount of Esau; and the kingdom shall be the LORD's.
