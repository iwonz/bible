DAN|1|1|In the third year of the reign of Jehoiakim king of Judah, Nebuchadnezzar king of Babylon came to Jerusalem and besieged it.
DAN|1|2|And the Lord delivered Jehoiakim king of Judah into his hand, along with some of the articles from the temple of God. These he carried off to the temple of his god in Babylonia and put in the treasure house of his god.
DAN|1|3|Then the king ordered Ashpenaz, chief of his court officials, to bring in some of the Israelites from the royal family and the nobility-
DAN|1|4|young men without any physical defect, handsome, showing aptitude for every kind of learning, well informed, quick to understand, and qualified to serve in the king's palace. He was to teach them the language and literature of the Babylonians.
DAN|1|5|The king assigned them a daily amount of food and wine from the king's table. They were to be trained for three years, and after that they were to enter the king's service.
DAN|1|6|Among these were some from Judah: Daniel, Hananiah, Mishael and Azariah.
DAN|1|7|The chief official gave them new names: to Daniel, the name Belteshazzar; to Hananiah, Shadrach; to Mishael, Meshach; and to Azariah, Abednego.
DAN|1|8|But Daniel resolved not to defile himself with the royal food and wine, and he asked the chief official for permission not to defile himself this way.
DAN|1|9|Now God had caused the official to show favor and sympathy to Daniel,
DAN|1|10|but the official told Daniel, "I am afraid of my lord the king, who has assigned your food and drink. Why should he see you looking worse than the other young men your age? The king would then have my head because of you."
DAN|1|11|Daniel then said to the guard whom the chief official had appointed over Daniel, Hananiah, Mishael and Azariah,
DAN|1|12|"Please test your servants for ten days: Give us nothing but vegetables to eat and water to drink.
DAN|1|13|Then compare our appearance with that of the young men who eat the royal food, and treat your servants in accordance with what you see."
DAN|1|14|So he agreed to this and tested them for ten days.
DAN|1|15|At the end of the ten days they looked healthier and better nourished than any of the young men who ate the royal food.
DAN|1|16|So the guard took away their choice food and the wine they were to drink and gave them vegetables instead.
DAN|1|17|To these four young men God gave knowledge and understanding of all kinds of literature and learning. And Daniel could understand visions and dreams of all kinds.
DAN|1|18|At the end of the time set by the king to bring them in, the chief official presented them to Nebuchadnezzar.
DAN|1|19|The king talked with them, and he found none equal to Daniel, Hananiah, Mishael and Azariah; so they entered the king's service.
DAN|1|20|In every matter of wisdom and understanding about which the king questioned them, he found them ten times better than all the magicians and enchanters in his whole kingdom.
DAN|1|21|And Daniel remained there until the first year of King Cyrus.
DAN|2|1|In the second year of his reign, Nebuchadnezzar had dreams; his mind was troubled and he could not sleep.
DAN|2|2|So the king summoned the magicians, enchanters, sorcerers and astrologers to tell him what he had dreamed. When they came in and stood before the king,
DAN|2|3|he said to them, "I have had a dream that troubles me and I want to know what it means. "
DAN|2|4|Then the astrologers answered the king in Aramaic, "O king, live forever! Tell your servants the dream, and we will interpret it."
DAN|2|5|The king replied to the astrologers, "This is what I have firmly decided: If you do not tell me what my dream was and interpret it, I will have you cut into pieces and your houses turned into piles of rubble.
DAN|2|6|But if you tell me the dream and explain it, you will receive from me gifts and rewards and great honor. So tell me the dream and interpret it for me."
DAN|2|7|Once more they replied, "Let the king tell his servants the dream, and we will interpret it."
DAN|2|8|Then the king answered, "I am certain that you are trying to gain time, because you realize that this is what I have firmly decided:
DAN|2|9|If you do not tell me the dream, there is just one penalty for you. You have conspired to tell me misleading and wicked things, hoping the situation will change. So then, tell me the dream, and I will know that you can interpret it for me."
DAN|2|10|The astrologers answered the king, "There is not a man on earth who can do what the king asks! No king, however great and mighty, has ever asked such a thing of any magician or enchanter or astrologer.
DAN|2|11|What the king asks is too difficult. No one can reveal it to the king except the gods, and they do not live among men."
DAN|2|12|This made the king so angry and furious that he ordered the execution of all the wise men of Babylon.
DAN|2|13|So the decree was issued to put the wise men to death, and men were sent to look for Daniel and his friends to put them to death.
DAN|2|14|When Arioch, the commander of the king's guard, had gone out to put to death the wise men of Babylon, Daniel spoke to him with wisdom and tact.
DAN|2|15|He asked the king's officer, "Why did the king issue such a harsh decree?" Arioch then explained the matter to Daniel.
DAN|2|16|At this, Daniel went in to the king and asked for time, so that he might interpret the dream for him.
DAN|2|17|Then Daniel returned to his house and explained the matter to his friends Hananiah, Mishael and Azariah.
DAN|2|18|He urged them to plead for mercy from the God of heaven concerning this mystery, so that he and his friends might not be executed with the rest of the wise men of Babylon.
DAN|2|19|During the night the mystery was revealed to Daniel in a vision. Then Daniel praised the God of heaven
DAN|2|20|and said: "Praise be to the name of God for ever and ever; wisdom and power are his.
DAN|2|21|He changes times and seasons; he sets up kings and deposes them. He gives wisdom to the wise and knowledge to the discerning.
DAN|2|22|He reveals deep and hidden things; he knows what lies in darkness, and light dwells with him.
DAN|2|23|I thank and praise you, O God of my fathers: You have given me wisdom and power, you have made known to me what we asked of you, you have made known to us the dream of the king."
DAN|2|24|Then Daniel went to Arioch, whom the king had appointed to execute the wise men of Babylon, and said to him, "Do not execute the wise men of Babylon. Take me to the king, and I will interpret his dream for him."
DAN|2|25|Arioch took Daniel to the king at once and said, "I have found a man among the exiles from Judah who can tell the king what his dream means."
DAN|2|26|The king asked Daniel (also called Belteshazzar), "Are you able to tell me what I saw in my dream and interpret it?"
DAN|2|27|Daniel replied, "No wise man, enchanter, magician or diviner can explain to the king the mystery he has asked about,
DAN|2|28|but there is a God in heaven who reveals mysteries. He has shown King Nebuchadnezzar what will happen in days to come. Your dream and the visions that passed through your mind as you lay on your bed are these:
DAN|2|29|"As you were lying there, O king, your mind turned to things to come, and the revealer of mysteries showed you what is going to happen.
DAN|2|30|As for me, this mystery has been revealed to me, not because I have greater wisdom than other living men, but so that you, O king, may know the interpretation and that you may understand what went through your mind.
DAN|2|31|"You looked, O king, and there before you stood a large statue-an enormous, dazzling statue, awesome in appearance.
DAN|2|32|The head of the statue was made of pure gold, its chest and arms of silver, its belly and thighs of bronze,
DAN|2|33|its legs of iron, its feet partly of iron and partly of baked clay.
DAN|2|34|While you were watching, a rock was cut out, but not by human hands. It struck the statue on its feet of iron and clay and smashed them.
DAN|2|35|Then the iron, the clay, the bronze, the silver and the gold were broken to pieces at the same time and became like chaff on a threshing floor in the summer. The wind swept them away without leaving a trace. But the rock that struck the statue became a huge mountain and filled the whole earth.
DAN|2|36|"This was the dream, and now we will interpret it to the king.
DAN|2|37|You, O king, are the king of kings. The God of heaven has given you dominion and power and might and glory;
DAN|2|38|in your hands he has placed mankind and the beasts of the field and the birds of the air. Wherever they live, he has made you ruler over them all. You are that head of gold.
DAN|2|39|"After you, another kingdom will rise, inferior to yours. Next, a third kingdom, one of bronze, will rule over the whole earth.
DAN|2|40|Finally, there will be a fourth kingdom, strong as iron-for iron breaks and smashes everything-and as iron breaks things to pieces, so it will crush and break all the others.
DAN|2|41|Just as you saw that the feet and toes were partly of baked clay and partly of iron, so this will be a divided kingdom; yet it will have some of the strength of iron in it, even as you saw iron mixed with clay.
DAN|2|42|As the toes were partly iron and partly clay, so this kingdom will be partly strong and partly brittle.
DAN|2|43|And just as you saw the iron mixed with baked clay, so the people will be a mixture and will not remain united, any more than iron mixes with clay.
DAN|2|44|"In the time of those kings, the God of heaven will set up a kingdom that will never be destroyed, nor will it be left to another people. It will crush all those kingdoms and bring them to an end, but it will itself endure forever.
DAN|2|45|This is the meaning of the vision of the rock cut out of a mountain, but not by human hands-a rock that broke the iron, the bronze, the clay, the silver and the gold to pieces. "The great God has shown the king what will take place in the future. The dream is true and the interpretation is trustworthy."
DAN|2|46|Then King Nebuchadnezzar fell prostrate before Daniel and paid him honor and ordered that an offering and incense be presented to him.
DAN|2|47|The king said to Daniel, "Surely your God is the God of gods and the Lord of kings and a revealer of mysteries, for you were able to reveal this mystery."
DAN|2|48|Then the king placed Daniel in a high position and lavished many gifts on him. He made him ruler over the entire province of Babylon and placed him in charge of all its wise men.
DAN|2|49|Moreover, at Daniel's request the king appointed Shadrach, Meshach and Abednego administrators over the province of Babylon, while Daniel himself remained at the royal court.
DAN|3|1|King Nebuchadnezzar made an image of gold, ninety feet high and nine feet wide, and set it up on the plain of Dura in the province of Babylon.
DAN|3|2|He then summoned the satraps, prefects, governors, advisers, treasurers, judges, magistrates and all the other provincial officials to come to the dedication of the image he had set up.
DAN|3|3|So the satraps, prefects, governors, advisers, treasurers, judges, magistrates and all the other provincial officials assembled for the dedication of the image that King Nebuchadnezzar had set up, and they stood before it.
DAN|3|4|Then the herald loudly proclaimed, "This is what you are commanded to do, O peoples, nations and men of every language:
DAN|3|5|As soon as you hear the sound of the horn, flute, zither, lyre, harp, pipes and all kinds of music, you must fall down and worship the image of gold that King Nebuchadnezzar has set up.
DAN|3|6|Whoever does not fall down and worship will immediately be thrown into a blazing furnace."
DAN|3|7|Therefore, as soon as they heard the sound of the horn, flute, zither, lyre, harp and all kinds of music, all the peoples, nations and men of every language fell down and worshiped the image of gold that King Nebuchadnezzar had set up.
DAN|3|8|At this time some astrologers came forward and denounced the Jews.
DAN|3|9|They said to King Nebuchadnezzar, "O king, live forever!
DAN|3|10|You have issued a decree, O king, that everyone who hears the sound of the horn, flute, zither, lyre, harp, pipes and all kinds of music must fall down and worship the image of gold,
DAN|3|11|and that whoever does not fall down and worship will be thrown into a blazing furnace.
DAN|3|12|But there are some Jews whom you have set over the affairs of the province of Babylon-Shadrach, Meshach and Abednego-who pay no attention to you, O king. They neither serve your gods nor worship the image of gold you have set up."
DAN|3|13|Furious with rage, Nebuchadnezzar summoned Shadrach, Meshach and Abednego. So these men were brought before the king,
DAN|3|14|and Nebuchadnezzar said to them, "Is it true, Shadrach, Meshach and Abednego, that you do not serve my gods or worship the image of gold I have set up?
DAN|3|15|Now when you hear the sound of the horn, flute, zither, lyre, harp, pipes and all kinds of music, if you are ready to fall down and worship the image I made, very good. But if you do not worship it, you will be thrown immediately into a blazing furnace. Then what god will be able to rescue you from my hand?"
DAN|3|16|Shadrach, Meshach and Abednego replied to the king, "O Nebuchadnezzar, we do not need to defend ourselves before you in this matter.
DAN|3|17|If we are thrown into the blazing furnace, the God we serve is able to save us from it, and he will rescue us from your hand, O king.
DAN|3|18|But even if he does not, we want you to know, O king, that we will not serve your gods or worship the image of gold you have set up."
DAN|3|19|Then Nebuchadnezzar was furious with Shadrach, Meshach and Abednego, and his attitude toward them changed. He ordered the furnace heated seven times hotter than usual
DAN|3|20|and commanded some of the strongest soldiers in his army to tie up Shadrach, Meshach and Abednego and throw them into the blazing furnace.
DAN|3|21|So these men, wearing their robes, trousers, turbans and other clothes, were bound and thrown into the blazing furnace.
DAN|3|22|The king's command was so urgent and the furnace so hot that the flames of the fire killed the soldiers who took up Shadrach, Meshach and Abednego,
DAN|3|23|and these three men, firmly tied, fell into the blazing furnace.
DAN|3|24|Then King Nebuchadnezzar leaped to his feet in amazement and asked his advisers, "Weren't there three men that we tied up and threw into the fire?" They replied, "Certainly, O king."
DAN|3|25|He said, "Look! I see four men walking around in the fire, unbound and unharmed, and the fourth looks like a son of the gods."
DAN|3|26|Nebuchadnezzar then approached the opening of the blazing furnace and shouted, "Shadrach, Meshach and Abednego, servants of the Most High God, come out! Come here!" So Shadrach, Meshach and Abednego came out of the fire,
DAN|3|27|and the satraps, prefects, governors and royal advisers crowded around them. They saw that the fire had not harmed their bodies, nor was a hair of their heads singed; their robes were not scorched, and there was no smell of fire on them.
DAN|3|28|Then Nebuchadnezzar said, "Praise be to the God of Shadrach, Meshach and Abednego, who has sent his angel and rescued his servants! They trusted in him and defied the king's command and were willing to give up their lives rather than serve or worship any god except their own God.
DAN|3|29|Therefore I decree that the people of any nation or language who say anything against the God of Shadrach, Meshach and Abednego be cut into pieces and their houses be turned into piles of rubble, for no other god can save in this way."
DAN|3|30|Then the king promoted Shadrach, Meshach and Abednego in the province of Babylon.
DAN|4|1|King Nebuchadnezzar, To the peoples, nations and men of every language, who live in all the world: May you prosper greatly!
DAN|4|2|It is my pleasure to tell you about the miraculous signs and wonders that the Most High God has performed for me.
DAN|4|3|How great are his signs, how mighty his wonders! His kingdom is an eternal kingdom; his dominion endures from generation to generation.
DAN|4|4|I, Nebuchadnezzar, was at home in my palace, contented and prosperous.
DAN|4|5|I had a dream that made me afraid. As I was lying in my bed, the images and visions that passed through my mind terrified me.
DAN|4|6|So I commanded that all the wise men of Babylon be brought before me to interpret the dream for me.
DAN|4|7|When the magicians, enchanters, astrologers and diviners came, I told them the dream, but they could not interpret it for me.
DAN|4|8|Finally, Daniel came into my presence and I told him the dream. (He is called Belteshazzar, after the name of my god, and the spirit of the holy gods is in him.)
DAN|4|9|I said, "Belteshazzar, chief of the magicians, I know that the spirit of the holy gods is in you, and no mystery is too difficult for you. Here is my dream; interpret it for me.
DAN|4|10|These are the visions I saw while lying in my bed: I looked, and there before me stood a tree in the middle of the land. Its height was enormous.
DAN|4|11|The tree grew large and strong and its top touched the sky; it was visible to the ends of the earth.
DAN|4|12|Its leaves were beautiful, its fruit abundant, and on it was food for all. Under it the beasts of the field found shelter, and the birds of the air lived in its branches; from it every creature was fed.
DAN|4|13|"In the visions I saw while lying in my bed, I looked, and there before me was a messenger, a holy one, coming down from heaven.
DAN|4|14|He called in a loud voice: 'Cut down the tree and trim off its branches; strip off its leaves and scatter its fruit. Let the animals flee from under it and the birds from its branches.
DAN|4|15|But let the stump and its roots, bound with iron and bronze, remain in the ground, in the grass of the field. "'Let him be drenched with the dew of heaven, and let him live with the animals among the plants of the earth.
DAN|4|16|Let his mind be changed from that of a man and let him be given the mind of an animal, till seven times pass by for him.
DAN|4|17|"'The decision is announced by messengers, the holy ones declare the verdict, so that the living may know that the Most High is sovereign over the kingdoms of men and gives them to anyone he wishes and sets over them the lowliest of men.'
DAN|4|18|"This is the dream that I, King Nebuchadnezzar, had. Now, Belteshazzar, tell me what it means, for none of the wise men in my kingdom can interpret it for me. But you can, because the spirit of the holy gods is in you."
DAN|4|19|Then Daniel (also called Belteshazzar) was greatly perplexed for a time, and his thoughts terrified him. So the king said, "Belteshazzar, do not let the dream or its meaning alarm you." Belteshazzar answered, "My lord, if only the dream applied to your enemies and its meaning to your adversaries!
DAN|4|20|The tree you saw, which grew large and strong, with its top touching the sky, visible to the whole earth,
DAN|4|21|with beautiful leaves and abundant fruit, providing food for all, giving shelter to the beasts of the field, and having nesting places in its branches for the birds of the air-
DAN|4|22|you, O king, are that tree! You have become great and strong; your greatness has grown until it reaches the sky, and your dominion extends to distant parts of the earth.
DAN|4|23|"You, O king, saw a messenger, a holy one, coming down from heaven and saying, 'Cut down the tree and destroy it, but leave the stump, bound with iron and bronze, in the grass of the field, while its roots remain in the ground. Let him be drenched with the dew of heaven; let him live like the wild animals, until seven times pass by for him.'
DAN|4|24|"This is the interpretation, O king, and this is the decree the Most High has issued against my lord the king:
DAN|4|25|You will be driven away from people and will live with the wild animals; you will eat grass like cattle and be drenched with the dew of heaven. Seven times will pass by for you until you acknowledge that the Most High is sovereign over the kingdoms of men and gives them to anyone he wishes.
DAN|4|26|The command to leave the stump of the tree with its roots means that your kingdom will be restored to you when you acknowledge that Heaven rules.
DAN|4|27|Therefore, O king, be pleased to accept my advice: Renounce your sins by doing what is right, and your wickedness by being kind to the oppressed. It may be that then your prosperity will continue."
DAN|4|28|All this happened to King Nebuchadnezzar.
DAN|4|29|Twelve months later, as the king was walking on the roof of the royal palace of Babylon,
DAN|4|30|he said, "Is not this the great Babylon I have built as the royal residence, by my mighty power and for the glory of my majesty?"
DAN|4|31|The words were still on his lips when a voice came from heaven, "This is what is decreed for you, King Nebuchadnezzar: Your royal authority has been taken from you.
DAN|4|32|You will be driven away from people and will live with the wild animals; you will eat grass like cattle. Seven times will pass by for you until you acknowledge that the Most High is sovereign over the kingdoms of men and gives them to anyone he wishes."
DAN|4|33|Immediately what had been said about Nebuchadnezzar was fulfilled. He was driven away from people and ate grass like cattle. His body was drenched with the dew of heaven until his hair grew like the feathers of an eagle and his nails like the claws of a bird.
DAN|4|34|At the end of that time, I, Nebuchadnezzar, raised my eyes toward heaven, and my sanity was restored. Then I praised the Most High; I honored and glorified him who lives forever. His dominion is an eternal dominion; his kingdom endures from generation to generation.
DAN|4|35|All the peoples of the earth are regarded as nothing. He does as he pleases with the powers of heaven and the peoples of the earth. No one can hold back his hand or say to him: "What have you done?"
DAN|4|36|At the same time that my sanity was restored, my honor and splendor were returned to me for the glory of my kingdom. My advisers and nobles sought me out, and I was restored to my throne and became even greater than before.
DAN|4|37|Now I, Nebuchadnezzar, praise and exalt and glorify the King of heaven, because everything he does is right and all his ways are just. And those who walk in pride he is able to humble.
DAN|5|1|King Belshazzar gave a great banquet for a thousand of his nobles and drank wine with them.
DAN|5|2|While Belshazzar was drinking his wine, he gave orders to bring in the gold and silver goblets that Nebuchadnezzar his father had taken from the temple in Jerusalem, so that the king and his nobles, his wives and his concubines might drink from them.
DAN|5|3|So they brought in the gold goblets that had been taken from the temple of God in Jerusalem, and the king and his nobles, his wives and his concubines drank from them.
DAN|5|4|As they drank the wine, they praised the gods of gold and silver, of bronze, iron, wood and stone.
DAN|5|5|Suddenly the fingers of a human hand appeared and wrote on the plaster of the wall, near the lampstand in the royal palace. The king watched the hand as it wrote.
DAN|5|6|His face turned pale and he was so frightened that his knees knocked together and his legs gave way.
DAN|5|7|The king called out for the enchanters, astrologers and diviners to be brought and said to these wise men of Babylon, "Whoever reads this writing and tells me what it means will be clothed in purple and have a gold chain placed around his neck, and he will be made the third highest ruler in the kingdom."
DAN|5|8|Then all the king's wise men came in, but they could not read the writing or tell the king what it meant.
DAN|5|9|So King Belshazzar became even more terrified and his face grew more pale. His nobles were baffled.
DAN|5|10|The queen, hearing the voices of the king and his nobles, came into the banquet hall. "O king, live forever!" she said. "Don't be alarmed! Don't look so pale!
DAN|5|11|There is a man in your kingdom who has the spirit of the holy gods in him. In the time of your father he was found to have insight and intelligence and wisdom like that of the gods. King Nebuchadnezzar your father-your father the king, I say-appointed him chief of the magicians, enchanters, astrologers and diviners.
DAN|5|12|This man Daniel, whom the king called Belteshazzar, was found to have a keen mind and knowledge and understanding, and also the ability to interpret dreams, explain riddles and solve difficult problems. Call for Daniel, and he will tell you what the writing means."
DAN|5|13|So Daniel was brought before the king, and the king said to him, "Are you Daniel, one of the exiles my father the king brought from Judah?
DAN|5|14|I have heard that the spirit of the gods is in you and that you have insight, intelligence and outstanding wisdom.
DAN|5|15|The wise men and enchanters were brought before me to read this writing and tell me what it means, but they could not explain it.
DAN|5|16|Now I have heard that you are able to give interpretations and to solve difficult problems. If you can read this writing and tell me what it means, you will be clothed in purple and have a gold chain placed around your neck, and you will be made the third highest ruler in the kingdom."
DAN|5|17|Then Daniel answered the king, "You may keep your gifts for yourself and give your rewards to someone else. Nevertheless, I will read the writing for the king and tell him what it means.
DAN|5|18|"O king, the Most High God gave your father Nebuchadnezzar sovereignty and greatness and glory and splendor.
DAN|5|19|Because of the high position he gave him, all the peoples and nations and men of every language dreaded and feared him. Those the king wanted to put to death, he put to death; those he wanted to spare, he spared; those he wanted to promote, he promoted; and those he wanted to humble, he humbled.
DAN|5|20|But when his heart became arrogant and hardened with pride, he was deposed from his royal throne and stripped of his glory.
DAN|5|21|He was driven away from people and given the mind of an animal; he lived with the wild donkeys and ate grass like cattle; and his body was drenched with the dew of heaven, until he acknowledged that the Most High God is sovereign over the kingdoms of men and sets over them anyone he wishes.
DAN|5|22|"But you his son, O Belshazzar, have not humbled yourself, though you knew all this.
DAN|5|23|Instead, you have set yourself up against the Lord of heaven. You had the goblets from his temple brought to you, and you and your nobles, your wives and your concubines drank wine from them. You praised the gods of silver and gold, of bronze, iron, wood and stone, which cannot see or hear or understand. But you did not honor the God who holds in his hand your life and all your ways.
DAN|5|24|Therefore he sent the hand that wrote the inscription.
DAN|5|25|"This is the inscription that was written: Mene, Mene, Tekel, Parsin
DAN|5|26|"This is what these words mean: Mene: God has numbered the days of your reign and brought it to an end.
DAN|5|27|Tekel: You have been weighed on the scales and found wanting.
DAN|5|28|Peres: Your kingdom is divided and given to the Medes and Persians."
DAN|5|29|Then at Belshazzar's command, Daniel was clothed in purple, a gold chain was placed around his neck, and he was proclaimed the third highest ruler in the kingdom.
DAN|5|30|That very night Belshazzar, king of the Babylonians, was slain,
DAN|5|31|and Darius the Mede took over the kingdom, at the age of sixty-two.
DAN|6|1|It pleased Darius to appoint 120 satraps to rule throughout the kingdom,
DAN|6|2|with three administrators over them, one of whom was Daniel. The satraps were made accountable to them so that the king might not suffer loss.
DAN|6|3|Now Daniel so distinguished himself among the administrators and the satraps by his exceptional qualities that the king planned to set him over the whole kingdom.
DAN|6|4|At this, the administrators and the satraps tried to find grounds for charges against Daniel in his conduct of government affairs, but they were unable to do so. They could find no corruption in him, because he was trustworthy and neither corrupt nor negligent.
DAN|6|5|Finally these men said, "We will never find any basis for charges against this man Daniel unless it has something to do with the law of his God."
DAN|6|6|So the administrators and the satraps went as a group to the king and said: "O King Darius, live forever!
DAN|6|7|The royal administrators, prefects, satraps, advisers and governors have all agreed that the king should issue an edict and enforce the decree that anyone who prays to any god or man during the next thirty days, except to you, O king, shall be thrown into the lions' den.
DAN|6|8|Now, O king, issue the decree and put it in writing so that it cannot be altered-in accordance with the laws of the Medes and Persians, which cannot be repealed."
DAN|6|9|So King Darius put the decree in writing.
DAN|6|10|Now when Daniel learned that the decree had been published, he went home to his upstairs room where the windows opened toward Jerusalem. Three times a day he got down on his knees and prayed, giving thanks to his God, just as he had done before.
DAN|6|11|Then these men went as a group and found Daniel praying and asking God for help.
DAN|6|12|So they went to the king and spoke to him about his royal decree: "Did you not publish a decree that during the next thirty days anyone who prays to any god or man except to you, O king, would be thrown into the lions' den?" The king answered, "The decree stands-in accordance with the laws of the Medes and Persians, which cannot be repealed."
DAN|6|13|Then they said to the king, "Daniel, who is one of the exiles from Judah, pays no attention to you, O king, or to the decree you put in writing. He still prays three times a day."
DAN|6|14|When the king heard this, he was greatly distressed; he was determined to rescue Daniel and made every effort until sundown to save him.
DAN|6|15|Then the men went as a group to the king and said to him, "Remember, O king, that according to the law of the Medes and Persians no decree or edict that the king issues can be changed."
DAN|6|16|So the king gave the order, and they brought Daniel and threw him into the lions' den. The king said to Daniel, "May your God, whom you serve continually, rescue you!"
DAN|6|17|A stone was brought and placed over the mouth of the den, and the king sealed it with his own signet ring and with the rings of his nobles, so that Daniel's situation might not be changed.
DAN|6|18|Then the king returned to his palace and spent the night without eating and without any entertainment being brought to him. And he could not sleep.
DAN|6|19|At the first light of dawn, the king got up and hurried to the lions' den.
DAN|6|20|When he came near the den, he called to Daniel in an anguished voice, "Daniel, servant of the living God, has your God, whom you serve continually, been able to rescue you from the lions?"
DAN|6|21|Daniel answered, "O king, live forever!
DAN|6|22|My God sent his angel, and he shut the mouths of the lions. They have not hurt me, because I was found innocent in his sight. Nor have I ever done any wrong before you, O king."
DAN|6|23|The king was overjoyed and gave orders to lift Daniel out of the den. And when Daniel was lifted from the den, no wound was found on him, because he had trusted in his God.
DAN|6|24|At the king's command, the men who had falsely accused Daniel were brought in and thrown into the lions' den, along with their wives and children. And before they reached the floor of the den, the lions overpowered them and crushed all their bones.
DAN|6|25|Then King Darius wrote to all the peoples, nations and men of every language throughout the land: "May you prosper greatly!
DAN|6|26|"I issue a decree that in every part of my kingdom people must fear and reverence the God of Daniel. "For he is the living God and he endures forever; his kingdom will not be destroyed, his dominion will never end.
DAN|6|27|He rescues and he saves; he performs signs and wonders in the heavens and on the earth. He has rescued Daniel from the power of the lions."
DAN|6|28|So Daniel prospered during the reign of Darius and the reign of Cyrus the Persian.
DAN|7|1|In the first year of Belshazzar king of Babylon, Daniel had a dream, and visions passed through his mind as he was lying on his bed. He wrote down the substance of his dream.
DAN|7|2|Daniel said: "In my vision at night I looked, and there before me were the four winds of heaven churning up the great sea.
DAN|7|3|Four great beasts, each different from the others, came up out of the sea.
DAN|7|4|"The first was like a lion, and it had the wings of an eagle. I watched until its wings were torn off and it was lifted from the ground so that it stood on two feet like a man, and the heart of a man was given to it.
DAN|7|5|"And there before me was a second beast, which looked like a bear. It was raised up on one of its sides, and it had three ribs in its mouth between its teeth. It was told, 'Get up and eat your fill of flesh!'
DAN|7|6|"After that, I looked, and there before me was another beast, one that looked like a leopard. And on its back it had four wings like those of a bird. This beast had four heads, and it was given authority to rule.
DAN|7|7|"After that, in my vision at night I looked, and there before me was a fourth beast-terrifying and frightening and very powerful. It had large iron teeth; it crushed and devoured its victims and trampled underfoot whatever was left. It was different from all the former beasts, and it had ten horns.
DAN|7|8|"While I was thinking about the horns, there before me was another horn, a little one, which came up among them; and three of the first horns were uprooted before it. This horn had eyes like the eyes of a man and a mouth that spoke boastfully.
DAN|7|9|"As I looked, "thrones were set in place, and the Ancient of Days took his seat. His clothing was as white as snow; the hair of his head was white like wool. His throne was flaming with fire, and its wheels were all ablaze.
DAN|7|10|A river of fire was flowing, coming out from before him. Thousands upon thousands attended him; ten thousand times ten thousand stood before him. The court was seated, and the books were opened.
DAN|7|11|"Then I continued to watch because of the boastful words the horn was speaking. I kept looking until the beast was slain and its body destroyed and thrown into the blazing fire.
DAN|7|12|(The other beasts had been stripped of their authority, but were allowed to live for a period of time.)
DAN|7|13|"In my vision at night I looked, and there before me was one like a son of man, coming with the clouds of heaven. He approached the Ancient of Days and was led into his presence.
DAN|7|14|He was given authority, glory and sovereign power; all peoples, nations and men of every language worshiped him. His dominion is an everlasting dominion that will not pass away, and his kingdom is one that will never be destroyed.
DAN|7|15|"I, Daniel, was troubled in spirit, and the visions that passed through my mind disturbed me.
DAN|7|16|I approached one of those standing there and asked him the true meaning of all this. "So he told me and gave me the interpretation of these things:
DAN|7|17|'The four great beasts are four kingdoms that will rise from the earth.
DAN|7|18|But the saints of the Most High will receive the kingdom and will possess it forever-yes, for ever and ever.'
DAN|7|19|"Then I wanted to know the true meaning of the fourth beast, which was different from all the others and most terrifying, with its iron teeth and bronze claws-the beast that crushed and devoured its victims and trampled underfoot whatever was left.
DAN|7|20|I also wanted to know about the ten horns on its head and about the other horn that came up, before which three of them fell-the horn that looked more imposing than the others and that had eyes and a mouth that spoke boastfully.
DAN|7|21|As I watched, this horn was waging war against the saints and defeating them,
DAN|7|22|until the Ancient of Days came and pronounced judgment in favor of the saints of the Most High, and the time came when they possessed the kingdom.
DAN|7|23|"He gave me this explanation: 'The fourth beast is a fourth kingdom that will appear on earth. It will be different from all the other kingdoms and will devour the whole earth, trampling it down and crushing it.
DAN|7|24|The ten horns are ten kings who will come from this kingdom. After them another king will arise, different from the earlier ones; he will subdue three kings.
DAN|7|25|He will speak against the Most High and oppress his saints and try to change the set times and the laws. The saints will be handed over to him for a time, times and half a time.
DAN|7|26|"'But the court will sit, and his power will be taken away and completely destroyed forever.
DAN|7|27|Then the sovereignty, power and greatness of the kingdoms under the whole heaven will be handed over to the saints, the people of the Most High. His kingdom will be an everlasting kingdom, and all rulers will worship and obey him.'
DAN|7|28|"This is the end of the matter. I, Daniel, was deeply troubled by my thoughts, and my face turned pale, but I kept the matter to myself."
DAN|8|1|In the third year of King Belshazzar's reign, I, Daniel, had a vision, after the one that had already appeared to me.
DAN|8|2|In my vision I saw myself in the citadel of Susa in the province of Elam; in the vision I was beside the Ulai Canal.
DAN|8|3|I looked up, and there before me was a ram with two horns, standing beside the canal, and the horns were long. One of the horns was longer than the other but grew up later.
DAN|8|4|I watched the ram as he charged toward the west and the north and the south. No animal could stand against him, and none could rescue from his power. He did as he pleased and became great.
DAN|8|5|As I was thinking about this, suddenly a goat with a prominent horn between his eyes came from the west, crossing the whole earth without touching the ground.
DAN|8|6|He came toward the two-horned ram I had seen standing beside the canal and charged at him in great rage.
DAN|8|7|I saw him attack the ram furiously, striking the ram and shattering his two horns. The ram was powerless to stand against him; the goat knocked him to the ground and trampled on him, and none could rescue the ram from his power.
DAN|8|8|The goat became very great, but at the height of his power his large horn was broken off, and in its place four prominent horns grew up toward the four winds of heaven.
DAN|8|9|Out of one of them came another horn, which started small but grew in power to the south and to the east and toward the Beautiful Land.
DAN|8|10|It grew until it reached the host of the heavens, and it threw some of the starry host down to the earth and trampled on them.
DAN|8|11|It set itself up to be as great as the Prince of the host; it took away the daily sacrifice from him, and the place of his sanctuary was brought low.
DAN|8|12|Because of rebellion, the host of the saints and the daily sacrifice were given over to it. It prospered in everything it did, and truth was thrown to the ground.
DAN|8|13|Then I heard a holy one speaking, and another holy one said to him, "How long will it take for the vision to be fulfilled-the vision concerning the daily sacrifice, the rebellion that causes desolation, and the surrender of the sanctuary and of the host that will be trampled underfoot?"
DAN|8|14|He said to me, "It will take 2,300 evenings and mornings; then the sanctuary will be reconsecrated."
DAN|8|15|While I, Daniel, was watching the vision and trying to understand it, there before me stood one who looked like a man.
DAN|8|16|And I heard a man's voice from the Ulai calling, "Gabriel, tell this man the meaning of the vision."
DAN|8|17|As he came near the place where I was standing, I was terrified and fell prostrate. "Son of man," he said to me, "understand that the vision concerns the time of the end."
DAN|8|18|While he was speaking to me, I was in a deep sleep, with my face to the ground. Then he touched me and raised me to my feet.
DAN|8|19|He said: "I am going to tell you what will happen later in the time of wrath, because the vision concerns the appointed time of the end.
DAN|8|20|The two-horned ram that you saw represents the kings of Media and Persia.
DAN|8|21|The shaggy goat is the king of Greece, and the large horn between his eyes is the first king.
DAN|8|22|The four horns that replaced the one that was broken off represent four kingdoms that will emerge from his nation but will not have the same power.
DAN|8|23|"In the latter part of their reign, when rebels have become completely wicked, a stern-faced king, a master of intrigue, will arise.
DAN|8|24|He will become very strong, but not by his own power. He will cause astounding devastation and will succeed in whatever he does. He will destroy the mighty men and the holy people.
DAN|8|25|He will cause deceit to prosper, and he will consider himself superior. When they feel secure, he will destroy many and take his stand against the Prince of princes. Yet he will be destroyed, but not by human power.
DAN|8|26|"The vision of the evenings and mornings that has been given you is true, but seal up the vision, for it concerns the distant future."
DAN|8|27|I, Daniel, was exhausted and lay ill for several days. Then I got up and went about the king's business. I was appalled by the vision; it was beyond understanding.
DAN|9|1|In the first year of Darius son of Ahasuerus (a Mede by descent), who was made ruler over the Babylonian kingdom-
DAN|9|2|in the first year of his reign, I, Daniel, understood from the Scriptures, according to the word of the LORD given to Jeremiah the prophet, that the desolation of Jerusalem would last seventy years.
DAN|9|3|So I turned to the Lord God and pleaded with him in prayer and petition, in fasting, and in sackcloth and ashes.
DAN|9|4|I prayed to the LORD my God and confessed: "O Lord, the great and awesome God, who keeps his covenant of love with all who love him and obey his commands,
DAN|9|5|we have sinned and done wrong. We have been wicked and have rebelled; we have turned away from your commands and laws.
DAN|9|6|We have not listened to your servants the prophets, who spoke in your name to our kings, our princes and our fathers, and to all the people of the land.
DAN|9|7|"Lord, you are righteous, but this day we are covered with shame-the men of Judah and people of Jerusalem and all Israel, both near and far, in all the countries where you have scattered us because of our unfaithfulness to you.
DAN|9|8|O LORD, we and our kings, our princes and our fathers are covered with shame because we have sinned against you.
DAN|9|9|The Lord our God is merciful and forgiving, even though we have rebelled against him;
DAN|9|10|we have not obeyed the LORD our God or kept the laws he gave us through his servants the prophets.
DAN|9|11|All Israel has transgressed your law and turned away, refusing to obey you. "Therefore the curses and sworn judgments written in the Law of Moses, the servant of God, have been poured out on us, because we have sinned against you.
DAN|9|12|You have fulfilled the words spoken against us and against our rulers by bringing upon us great disaster. Under the whole heaven nothing has ever been done like what has been done to Jerusalem.
DAN|9|13|Just as it is written in the Law of Moses, all this disaster has come upon us, yet we have not sought the favor of the LORD our God by turning from our sins and giving attention to your truth.
DAN|9|14|The LORD did not hesitate to bring the disaster upon us, for the LORD our God is righteous in everything he does; yet we have not obeyed him.
DAN|9|15|"Now, O Lord our God, who brought your people out of Egypt with a mighty hand and who made for yourself a name that endures to this day, we have sinned, we have done wrong.
DAN|9|16|O Lord, in keeping with all your righteous acts, turn away your anger and your wrath from Jerusalem, your city, your holy hill. Our sins and the iniquities of our fathers have made Jerusalem and your people an object of scorn to all those around us.
DAN|9|17|"Now, our God, hear the prayers and petitions of your servant. For your sake, O Lord, look with favor on your desolate sanctuary.
DAN|9|18|Give ear, O God, and hear; open your eyes and see the desolation of the city that bears your Name. We do not make requests of you because we are righteous, but because of your great mercy.
DAN|9|19|O Lord, listen! O Lord, forgive! O Lord, hear and act! For your sake, O my God, do not delay, because your city and your people bear your Name."
DAN|9|20|While I was speaking and praying, confessing my sin and the sin of my people Israel and making my request to the LORD my God for his holy hill-
DAN|9|21|while I was still in prayer, Gabriel, the man I had seen in the earlier vision, came to me in swift flight about the time of the evening sacrifice.
DAN|9|22|He instructed me and said to me, "Daniel, I have now come to give you insight and understanding.
DAN|9|23|As soon as you began to pray, an answer was given, which I have come to tell you, for you are highly esteemed. Therefore, consider the message and understand the vision:
DAN|9|24|"Seventy 'sevens' are decreed for your people and your holy city to finish transgression, to put an end to sin, to atone for wickedness, to bring in everlasting righteousness, to seal up vision and prophecy and to anoint the most holy.
DAN|9|25|"Know and understand this: From the issuing of the decree to restore and rebuild Jerusalem until the Anointed One, the ruler, comes, there will be seven 'sevens,' and sixty-two 'sevens.' It will be rebuilt with streets and a trench, but in times of trouble.
DAN|9|26|After the sixty-two 'sevens,' the Anointed One will be cut off and will have nothing. The people of the ruler who will come will destroy the city and the sanctuary. The end will come like a flood: War will continue until the end, and desolations have been decreed.
DAN|9|27|He will confirm a covenant with many for one 'seven.' In the middle of the 'seven' he will put an end to sacrifice and offering. And on a wing of the temple he will set up an abomination that causes desolation, until the end that is decreed is poured out on him. "
DAN|10|1|In the third year of Cyrus king of Persia, a revelation was given to Daniel (who was called Belteshazzar). Its message was true and it concerned a great war. The understanding of the message came to him in a vision.
DAN|10|2|At that time I, Daniel, mourned for three weeks.
DAN|10|3|I ate no choice food; no meat or wine touched my lips; and I used no lotions at all until the three weeks were over.
DAN|10|4|On the twenty-fourth day of the first month, as I was standing on the bank of the great river, the Tigris,
DAN|10|5|I looked up and there before me was a man dressed in linen, with a belt of the finest gold around his waist.
DAN|10|6|His body was like chrysolite, his face like lightning, his eyes like flaming torches, his arms and legs like the gleam of burnished bronze, and his voice like the sound of a multitude.
DAN|10|7|I, Daniel, was the only one who saw the vision; the men with me did not see it, but such terror overwhelmed them that they fled and hid themselves.
DAN|10|8|So I was left alone, gazing at this great vision; I had no strength left, my face turned deathly pale and I was helpless.
DAN|10|9|Then I heard him speaking, and as I listened to him, I fell into a deep sleep, my face to the ground.
DAN|10|10|A hand touched me and set me trembling on my hands and knees.
DAN|10|11|He said, "Daniel, you who are highly esteemed, consider carefully the words I am about to speak to you, and stand up, for I have now been sent to you." And when he said this to me, I stood up trembling.
DAN|10|12|Then he continued, "Do not be afraid, Daniel. Since the first day that you set your mind to gain understanding and to humble yourself before your God, your words were heard, and I have come in response to them.
DAN|10|13|But the prince of the Persian kingdom resisted me twenty-one days. Then Michael, one of the chief princes, came to help me, because I was detained there with the king of Persia.
DAN|10|14|Now I have come to explain to you what will happen to your people in the future, for the vision concerns a time yet to come."
DAN|10|15|While he was saying this to me, I bowed with my face toward the ground and was speechless.
DAN|10|16|Then one who looked like a man touched my lips, and I opened my mouth and began to speak. I said to the one standing before me, "I am overcome with anguish because of the vision, my lord, and I am helpless.
DAN|10|17|How can I, your servant, talk with you, my lord? My strength is gone and I can hardly breathe."
DAN|10|18|Again the one who looked like a man touched me and gave me strength.
DAN|10|19|"Do not be afraid, O man highly esteemed," he said. "Peace! Be strong now; be strong." When he spoke to me, I was strengthened and said, "Speak, my lord, since you have given me strength."
DAN|10|20|So he said, "Do you know why I have come to you? Soon I will return to fight against the prince of Persia, and when I go, the prince of Greece will come;
DAN|10|21|but first I will tell you what is written in the Book of Truth. (No one supports me against them except Michael, your prince.
DAN|11|1|And in the first year of Darius the Mede, I took my stand to support and protect him.)
DAN|11|2|"Now then, I tell you the truth: Three more kings will appear in Persia, and then a fourth, who will be far richer than all the others. When he has gained power by his wealth, he will stir up everyone against the kingdom of Greece.
DAN|11|3|Then a mighty king will appear, who will rule with great power and do as he pleases.
DAN|11|4|After he has appeared, his empire will be broken up and parceled out toward the four winds of heaven. It will not go to his descendants, nor will it have the power he exercised, because his empire will be uprooted and given to others.
DAN|11|5|"The king of the South will become strong, but one of his commanders will become even stronger than he and will rule his own kingdom with great power.
DAN|11|6|After some years, they will become allies. The daughter of the king of the South will go to the king of the North to make an alliance, but she will not retain her power, and he and his power will not last. In those days she will be handed over, together with her royal escort and her father and the one who supported her.
DAN|11|7|"One from her family line will arise to take her place. He will attack the forces of the king of the North and enter his fortress; he will fight against them and be victorious.
DAN|11|8|He will also seize their gods, their metal images and their valuable articles of silver and gold and carry them off to Egypt. For some years he will leave the king of the North alone.
DAN|11|9|Then the king of the North will invade the realm of the king of the South but will retreat to his own country.
DAN|11|10|His sons will prepare for war and assemble a great army, which will sweep on like an irresistible flood and carry the battle as far as his fortress.
DAN|11|11|"Then the king of the South will march out in a rage and fight against the king of the North, who will raise a large army, but it will be defeated.
DAN|11|12|When the army is carried off, the king of the South will be filled with pride and will slaughter many thousands, yet he will not remain triumphant.
DAN|11|13|For the king of the North will muster another army, larger than the first; and after several years, he will advance with a huge army fully equipped.
DAN|11|14|"In those times many will rise against the king of the South. The violent men among your own people will rebel in fulfillment of the vision, but without success.
DAN|11|15|Then the king of the North will come and build up siege ramps and will capture a fortified city. The forces of the South will be powerless to resist; even their best troops will not have the strength to stand.
DAN|11|16|The invader will do as he pleases; no one will be able to stand against him. He will establish himself in the Beautiful Land and will have the power to destroy it.
DAN|11|17|He will determine to come with the might of his entire kingdom and will make an alliance with the king of the South. And he will give him a daughter in marriage in order to overthrow the kingdom, but his plans will not succeed or help him.
DAN|11|18|Then he will turn his attention to the coastlands and will take many of them, but a commander will put an end to his insolence and will turn his insolence back upon him.
DAN|11|19|After this, he will turn back toward the fortresses of his own country but will stumble and fall, to be seen no more.
DAN|11|20|"His successor will send out a tax collector to maintain the royal splendor. In a few years, however, he will be destroyed, yet not in anger or in battle.
DAN|11|21|"He will be succeeded by a contemptible person who has not been given the honor of royalty. He will invade the kingdom when its people feel secure, and he will seize it through intrigue.
DAN|11|22|Then an overwhelming army will be swept away before him; both it and a prince of the covenant will be destroyed.
DAN|11|23|After coming to an agreement with him, he will act deceitfully, and with only a few people he will rise to power.
DAN|11|24|When the richest provinces feel secure, he will invade them and will achieve what neither his fathers nor his forefathers did. He will distribute plunder, loot and wealth among his followers. He will plot the overthrow of fortresses-but only for a time.
DAN|11|25|"With a large army he will stir up his strength and courage against the king of the South. The king of the South will wage war with a large and very powerful army, but he will not be able to stand because of the plots devised against him.
DAN|11|26|Those who eat from the king's provisions will try to destroy him; his army will be swept away, and many will fall in battle.
DAN|11|27|The two kings, with their hearts bent on evil, will sit at the same table and lie to each other, but to no avail, because an end will still come at the appointed time.
DAN|11|28|The king of the North will return to his own country with great wealth, but his heart will be set against the holy covenant. He will take action against it and then return to his own country.
DAN|11|29|"At the appointed time he will invade the South again, but this time the outcome will be different from what it was before.
DAN|11|30|Ships of the western coastlands will oppose him, and he will lose heart. Then he will turn back and vent his fury against the holy covenant. He will return and show favor to those who forsake the holy covenant.
DAN|11|31|"His armed forces will rise up to desecrate the temple fortress and will abolish the daily sacrifice. Then they will set up the abomination that causes desolation.
DAN|11|32|With flattery he will corrupt those who have violated the covenant, but the people who know their God will firmly resist him.
DAN|11|33|"Those who are wise will instruct many, though for a time they will fall by the sword or be burned or captured or plundered.
DAN|11|34|When they fall, they will receive a little help, and many who are not sincere will join them.
DAN|11|35|Some of the wise will stumble, so that they may be refined, purified and made spotless until the time of the end, for it will still come at the appointed time.
DAN|11|36|"The king will do as he pleases. He will exalt and magnify himself above every god and will say unheard-of things against the God of gods. He will be successful until the time of wrath is completed, for what has been determined must take place.
DAN|11|37|He will show no regard for the gods of his fathers or for the one desired by women, nor will he regard any god, but will exalt himself above them all.
DAN|11|38|Instead of them, he will honor a god of fortresses; a god unknown to his fathers he will honor with gold and silver, with precious stones and costly gifts.
DAN|11|39|He will attack the mightiest fortresses with the help of a foreign god and will greatly honor those who acknowledge him. He will make them rulers over many people and will distribute the land at a price.
DAN|11|40|"At the time of the end the king of the South will engage him in battle, and the king of the North will storm out against him with chariots and cavalry and a great fleet of ships. He will invade many countries and sweep through them like a flood.
DAN|11|41|He will also invade the Beautiful Land. Many countries will fall, but Edom, Moab and the leaders of Ammon will be delivered from his hand.
DAN|11|42|He will extend his power over many countries; Egypt will not escape.
DAN|11|43|He will gain control of the treasures of gold and silver and all the riches of Egypt, with the Libyans and Nubians in submission.
DAN|11|44|But reports from the east and the north will alarm him, and he will set out in a great rage to destroy and annihilate many.
DAN|11|45|He will pitch his royal tents between the seas at the beautiful holy mountain. Yet he will come to his end, and no one will help him.
DAN|12|1|"At that time Michael, the great prince who protects your people, will arise. There will be a time of distress such as has not happened from the beginning of nations until then. But at that time your people-everyone whose name is found written in the book-will be delivered.
DAN|12|2|Multitudes who sleep in the dust of the earth will awake: some to everlasting life, others to shame and everlasting contempt.
DAN|12|3|Those who are wise will shine like the brightness of the heavens, and those who lead many to righteousness, like the stars for ever and ever.
DAN|12|4|But you, Daniel, close up and seal the words of the scroll until the time of the end. Many will go here and there to increase knowledge."
DAN|12|5|Then I, Daniel, looked, and there before me stood two others, one on this bank of the river and one on the opposite bank.
DAN|12|6|One of them said to the man clothed in linen, who was above the waters of the river, "How long will it be before these astonishing things are fulfilled?"
DAN|12|7|The man clothed in linen, who was above the waters of the river, lifted his right hand and his left hand toward heaven, and I heard him swear by him who lives forever, saying, "It will be for a time, times and half a time. When the power of the holy people has been finally broken, all these things will be completed."
DAN|12|8|I heard, but I did not understand. So I asked, "My lord, what will the outcome of all this be?"
DAN|12|9|He replied, "Go your way, Daniel, because the words are closed up and sealed until the time of the end.
DAN|12|10|Many will be purified, made spotless and refined, but the wicked will continue to be wicked. None of the wicked will understand, but those who are wise will understand.
DAN|12|11|"From the time that the daily sacrifice is abolished and the abomination that causes desolation is set up, there will be 1,290 days.
DAN|12|12|Blessed is the one who waits for and reaches the end of the 1,335 days.
DAN|12|13|"As for you, go your way till the end. You will rest, and then at the end of the days you will rise to receive your allotted inheritance."
