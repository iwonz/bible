HEB|1|1|Long ago, at many times and in many ways, God spoke to our fathers by the prophets,
HEB|1|2|but in these last days he has spoken to us by his Son, whom he appointed the heir of all things, through whom also he created the world.
HEB|1|3|He is the radiance of the glory of God and the exact imprint of his nature, and he upholds the universe by the word of his power. After making purification for sins, he sat down at the right hand of the Majesty on high,
HEB|1|4|having become as much superior to angels as the name he has inherited is more excellent than theirs.
HEB|1|5|For to which of the angels did God ever say, "You are my Son, today I have begotten you"? Or again, "I will be to him a father, and he shall be to me a son"?
HEB|1|6|And again, when he brings the firstborn into the world, he says, "Let all God's angels worship him."
HEB|1|7|Of the angels he says, "He makes his angels winds, and his ministers a flame of fire."
HEB|1|8|But of the Son he says, "Your throne, O God, is forever and ever, the scepter of uprightness is the scepter of your kingdom.
HEB|1|9|You have loved righteousness and hated wickedness; therefore God, your God, has anointed you with the oil of gladness beyond your companions."
HEB|1|10|And, "You, Lord, laid the foundation of the earth in the beginning, and the heavens are the work of your hands;
HEB|1|11|they will perish, but you remain; they will all wear out like a garment,
HEB|1|12|like a robe you will roll them up, like a garment they will be changed. But you are the same, and your years will have no end."
HEB|1|13|And to which of the angels has he ever said, "Sit at my right hand until I make your enemies a footstool for your feet"?
HEB|1|14|Are they not all ministering spirits sent out to serve for the sake of those who are to inherit salvation?
HEB|2|1|Therefore we must pay much closer attention to what we have heard, lest we drift away from it.
HEB|2|2|For since the message declared by angels proved to be reliable and every transgression or disobedience received a just retribution,
HEB|2|3|how shall we escape if we neglect such a great salvation? It was declared at first by the Lord, and it was attested to us by those who heard,
HEB|2|4|while God also bore witness by signs and wonders and various miracles and by gifts of the Holy Spirit distributed according to his will.
HEB|2|5|Now it was not to angels that God subjected the world to come, of which we are speaking.
HEB|2|6|It has been testified somewhere, "What is man, that you are mindful of him, or the son of man, that you care for him?
HEB|2|7|You made him for a little while lower than the angels; you have crowned him with glory and honor,
HEB|2|8|putting everything in subjection under his feet." Now in putting everything in subjection to him, he left nothing outside his control. At present, we do not yet see everything in subjection to him.
HEB|2|9|But we see him who for a little while was made lower than the angels, namely Jesus, crowned with glory and honor because of the suffering of death, so that by the grace of God he might taste death for everyone.
HEB|2|10|For it was fitting that he, for whom and by whom all things exist, in bringing many sons to glory, should make the founder of their salvation perfect through suffering.
HEB|2|11|For he who sanctifies and those who are sanctified all have one origin. That is why he is not ashamed to call them brothers,
HEB|2|12|saying, "I will tell of your name to my brothers; in the midst of the congregation I will sing your praise."
HEB|2|13|And again, "I will put my trust in him." And again, "Behold, I and the children God has given me."
HEB|2|14|Since therefore the children share in flesh and blood, he himself likewise partook of the same things, that through death he might destroy the one who has the power of death, that is, the devil,
HEB|2|15|and deliver all those who through fear of death were subject to lifelong slavery.
HEB|2|16|For surely it is not angels that he helps, but he helps the offspring of Abraham.
HEB|2|17|Therefore he had to be made like his brothers in every respect, so that he might become a merciful and faithful high priest in the service of God, to make propitiation for the sins of the people.
HEB|2|18|For because he himself has suffered when tempted, he is able to help those who are being tempted.
HEB|3|1|Therefore, holy brothers, you who share in a heavenly calling, consider Jesus, the apostle and high priest of our confession,
HEB|3|2|who was faithful to him who appointed him, just as Moses also was faithful in all God's house.
HEB|3|3|For Jesus has been counted worthy of more glory than Moses- as much more glory as the builder of a house has more honor than the house itself.
HEB|3|4|(For every house is built by someone, but the builder of all things is God.)
HEB|3|5|Now Moses was faithful in all God's house as a servant, to testify to the things that were to be spoken later,
HEB|3|6|but Christ is faithful over God's house as a son. And we are his house if indeed we hold fast our confidence and our boasting in our hope.
HEB|3|7|Therefore, as the Holy Spirit says, "Today, if you hear his voice,
HEB|3|8|do not harden your hearts as in the rebellion, on the day of testing in the wilderness,
HEB|3|9|where your fathers put me to the test and saw my works
HEB|3|10|for forty years. Therefore I was provoked with that generation, and said, 'They always go astray in their heart; they have not known my ways.'
HEB|3|11|As I swore in my wrath, 'They shall not enter my rest.'"
HEB|3|12|Take care, brothers, lest there be in any of you an evil, unbelieving heart, leading you to fall away from the living God.
HEB|3|13|But exhort one another every day, as long as it is called "today," that none of you may be hardened by the deceitfulness of sin.
HEB|3|14|For we share in Christ, if indeed we hold our original confidence firm to the end.
HEB|3|15|As it is said, "Today, if you hear his voice, do not harden your hearts as in the rebellion."
HEB|3|16|For who were those who heard and yet rebelled? Was it not all those who left Egypt led by Moses?
HEB|3|17|And with whom was he provoked for forty years? Was it not with those who sinned, whose bodies fell in the wilderness?
HEB|3|18|And to whom did he swear that they would not enter his rest, but to those who were disobedient?
HEB|3|19|So we see that they were unable to enter because of unbelief.
HEB|4|1|Therefore, while the promise of entering his rest still stands, let us fear lest any of you should seem to have failed to reach it.
HEB|4|2|For good news came to us just as to them, but the message they heard did not benefit them, because they were not united by faith with those who listened.
HEB|4|3|For we who have believed enter that rest, as he has said, "As I swore in my wrath, 'They shall not enter my rest,'" although his works were finished from the foundation of the world.
HEB|4|4|For he has somewhere spoken of the seventh day in this way: "And God rested on the seventh day from all his works."
HEB|4|5|And again in this passage he said, "They shall not enter my rest."
HEB|4|6|Since therefore it remains for some to enter it, and those who formerly received the good news failed to enter because of disobedience,
HEB|4|7|again he appoints a certain day, "Today," saying through David so long afterward, in the words already quoted, "Today, if you hear his voice, do not harden your hearts."
HEB|4|8|For if Joshua had given them rest, God would not have spoken of another day later on.
HEB|4|9|So then, there remains a Sabbath rest for the people of God,
HEB|4|10|for whoever has entered God's rest has also rested from his works as God did from his.
HEB|4|11|Let us therefore strive to enter that rest, so that no one may fall by the same sort of disobedience.
HEB|4|12|For the word of God is living and active, sharper than any two-edged sword, piercing to the division of soul and of spirit, of joints and of marrow, and discerning the thoughts and intentions of the heart.
HEB|4|13|And no creature is hidden from his sight, but all are naked and exposed to the eyes of him to whom we must give account.
HEB|4|14|Since then we have a great high priest who has passed through the heavens, Jesus, the Son of God, let us hold fast our confession.
HEB|4|15|For we do not have a high priest who is unable to sympathize with our weaknesses, but one who in every respect has been tempted as we are, yet without sin.
HEB|4|16|Let us then with confidence draw near to the throne of grace, that we may receive mercy and find grace to help in time of need.
HEB|5|1|For every high priest chosen from among men is appointed to act on behalf of men in relation to God, to offer gifts and sacrifices for sins.
HEB|5|2|He can deal gently with the ignorant and wayward, since he himself is beset with weakness.
HEB|5|3|Because of this he is obligated to offer sacrifice for his own sins just as he does for those of the people.
HEB|5|4|And no one takes this honor for himself, but only when called by God, just as Aaron was.
HEB|5|5|So also Christ did not exalt himself to be made a high priest, but was appointed by him who said to him, "You are my Son, today I have begotten you";
HEB|5|6|as he says also in another place, "You are a priest forever, after the order of Melchizedek."
HEB|5|7|In the days of his flesh, Jesus offered up prayers and supplications, with loud cries and tears, to him who was able to save him from death, and he was heard because of his reverence.
HEB|5|8|Although he was a son, he learned obedience through what he suffered.
HEB|5|9|And being made perfect, he became the source of eternal salvation to all who obey him,
HEB|5|10|being designated by God a high priest after the order of Melchizedek.
HEB|5|11|About this we have much to say, and it is hard to explain, since you have become dull of hearing.
HEB|5|12|For though by this time you ought to be teachers, you need someone to teach you again the basic principles of the oracles of God. You need milk, not solid food,
HEB|5|13|for everyone who lives on milk is unskilled in the word of righteousness, since he is a child.
HEB|5|14|But solid food is for the mature, for those who have their powers of discernment trained by constant practice to distinguish good from evil.
HEB|6|1|Therefore let us leave the elementary doctrine of Christ and go on to maturity, not laying again a foundation of repentance from dead works and of faith toward God,
HEB|6|2|and of instruction about washings, the laying on of hands, the resurrection of the dead, and eternal judgment.
HEB|6|3|And this we will do if God permits.
HEB|6|4|For it is impossible to restore again to repentance those who have once been enlightened, who have tasted the heavenly gift, and have shared in the Holy Spirit,
HEB|6|5|and have tasted the goodness of the word of God and the powers of the age to come,
HEB|6|6|if they then fall away, since they are crucifying once again the Son of God to their own harm and holding him up to contempt.
HEB|6|7|For land that has drunk the rain that often falls on it, and produces a crop useful to those for whose sake it is cultivated, receives a blessing from God.
HEB|6|8|But if it bears thorns and thistles, it is worthless and near to being cursed, and its end is to be burned.
HEB|6|9|Though we speak in this way, yet in your case, beloved, we feel sure of better things- things that belong to salvation.
HEB|6|10|For God is not so unjust as to overlook your work and the love that you showed for his sake in serving the saints, as you still do.
HEB|6|11|And we desire each one of you to show the same earnestness to have the full assurance of hope until the end,
HEB|6|12|so that you may not be sluggish, but imitators of those who through faith and patience inherit the promises.
HEB|6|13|For when God made a promise to Abraham, since he had no one greater by whom to swear, he swore by himself,
HEB|6|14|saying, "Surely I will bless you and multiply you."
HEB|6|15|And thus Abraham, having patiently waited, obtained the promise.
HEB|6|16|For people swear by something greater than themselves, and in all their disputes an oath is final for confirmation.
HEB|6|17|So when God desired to show more convincingly to the heirs of the promise the unchangeable character of his purpose, he guaranteed it with an oath,
HEB|6|18|so that by two unchangeable things, in which it is impossible for God to lie, we who have fled for refuge might have strong encouragement to hold fast to the hope set before us.
HEB|6|19|We have this as a sure and steadfast anchor of the soul, a hope that enters into the inner place behind the curtain,
HEB|6|20|where Jesus has gone as a forerunner on our behalf, having become a high priest forever after the order of Melchizedek.
HEB|7|1|For this Melchizedek, king of Salem, priest of the Most High God, met Abraham returning from the slaughter of the kings and blessed him,
HEB|7|2|and to him Abraham apportioned a tenth part of everything. He is first, by translation of his name, king of righteousness, and then he is also king of Salem, that is, king of peace.
HEB|7|3|He is without father or mother or genealogy, having neither beginning of days nor end of life, but resembling the Son of God he continues a priest forever.
HEB|7|4|See how great this man was to whom Abraham the patriarch gave a tenth of the spoils!
HEB|7|5|And those descendants of Levi who receive the priestly office have a commandment in the law to take tithes from the people, that is, from their brothers, though these also are descended from Abraham.
HEB|7|6|But this man who does not have his descent from them received tithes from Abraham and blessed him who had the promises.
HEB|7|7|It is beyond dispute that the inferior is blessed by the superior.
HEB|7|8|In the one case tithes are received by mortal men, but in the other case, by one of whom it is testified that he lives.
HEB|7|9|One might even say that Levi himself, who receives tithes, paid tithes through Abraham,
HEB|7|10|for he was still in the loins of his ancestor when Melchizedek met him.
HEB|7|11|Now if perfection had been attainable through the Levitical priesthood (for under it the people received the law), what further need would there have been for another priest to arise after the order of Melchizedek, rather than one named after the order of Aaron?
HEB|7|12|For when there is a change in the priesthood, there is necessarily a change in the law as well.
HEB|7|13|For the one of whom these things are spoken belonged to another tribe, from which no one has ever served at the altar.
HEB|7|14|For it is evident that our Lord was descended from Judah, and in connection with that tribe Moses said nothing about priests.
HEB|7|15|This becomes even more evident when another priest arises in the likeness of Melchizedek,
HEB|7|16|who has become a priest, not on the basis of a legal requirement concerning bodily descent, but by the power of an indestructible life.
HEB|7|17|For it is witnessed of him, "You are a priest forever, after the order of Melchizedek."
HEB|7|18|On the one hand, a former commandment is set aside because of its weakness and uselessness
HEB|7|19|(for the law made nothing perfect); but on the other hand, a better hope is introduced, through which we draw near to God.
HEB|7|20|And it was not without an oath. For those who formerly became priests were made such without an oath,
HEB|7|21|but this one was made a priest with an oath by the one who said to him: "The Lord has sworn and will not change his mind, 'You are a priest forever.'"
HEB|7|22|This makes Jesus the guarantor of a better covenant.
HEB|7|23|The former priests were many in number, because they were prevented by death from continuing in office,
HEB|7|24|but he holds his priesthood permanently, because he continues forever.
HEB|7|25|Consequently, he is able to save to the uttermost those who draw near to God through him, since he always lives to make intercession for them.
HEB|7|26|For it was indeed fitting that we should have such a high priest, holy, innocent, unstained, separated from sinners, and exalted above the heavens.
HEB|7|27|He has no need, like those high priests, to offer sacrifices daily, first for his own sins and then for those of the people, since he did this once for all when he offered up himself.
HEB|7|28|For the law appoints men in their weakness as high priests, but the word of the oath, which came later than the law, appoints a Son who has been made perfect forever.
HEB|8|1|Now the point in what we are saying is this: we have such a high priest, one who is seated at the right hand of the throne of the Majesty in heaven,
HEB|8|2|a minister in the holy places, in the true tent that the Lord set up, not man.
HEB|8|3|For every high priest is appointed to offer gifts and sacrifices; thus it is necessary for this priest also to have something to offer.
HEB|8|4|Now if he were on earth, he would not be a priest at all, since there are priests who offer gifts according to the law.
HEB|8|5|They serve a copy and shadow of the heavenly things. For when Moses was about to erect the tent, he was instructed by God, saying, "See that you make everything according to the pattern that was shown you on the mountain."
HEB|8|6|But as it is, Christ has obtained a ministry that is as much more excellent than the old as the covenant he mediates is better, since it is enacted on better promises.
HEB|8|7|For if that first covenant had been faultless, there would have been no occasion to look for a second.
HEB|8|8|For he finds fault with them when he says: "Behold, the days are coming, declares the Lord, when I will establish a new covenant with the house of Israel and with the house of Judah,
HEB|8|9|not like the covenant that I made with their fathers on the day when I took them by the hand to bring them out of the land of Egypt. For they did not continue in my covenant, and so I showed no concern for them, declares the Lord.
HEB|8|10|For this is the covenant that I will make with the house of Israel after those days, declares the Lord: I will put my laws into their minds, and write them on their hearts, and I will be their God, and they shall be my people.
HEB|8|11|And they shall not teach, each one his neighbor and each one his brother, saying, 'Know the Lord,' for they shall all know me, from the least of them to the greatest.
HEB|8|12|For I will be merciful toward their iniquities, and I will remember their sins no more."
HEB|8|13|In speaking of a new covenant, he makes the first one obsolete. And what is becoming obsolete and growing old is ready to vanish away.
HEB|9|1|Now even the first covenant had regulations for worship and an earthly place of holiness.
HEB|9|2|For a tent was prepared, the first section, in which were the lampstand and the table and the bread of the Presence. It is called the Holy Place.
HEB|9|3|Behind the second curtain was a second section called the Most Holy Place,
HEB|9|4|having the golden altar of incense and the ark of the covenant covered on all sides with gold, in which was a golden urn holding the manna, and Aaron's staff that budded, and the tablets of the covenant.
HEB|9|5|Above it were the cherubim of glory overshadowing the mercy seat. Of these things we cannot now speak in detail.
HEB|9|6|These preparations having thus been made, the priests go regularly into the first section, performing their ritual duties,
HEB|9|7|but into the second only the high priest goes, and he but once a year, and not without taking blood, which he offers for himself and for the unintentional sins of the people.
HEB|9|8|By this the Holy Spirit indicates that the way into the holy places is not yet opened as long as the first section is still standing
HEB|9|9|(which is symbolic for the present age). According to this arrangement, gifts and sacrifices are offered that cannot perfect the conscience of the worshiper,
HEB|9|10|but deal only with food and drink and various washings, regulations for the body imposed until the time of reformation.
HEB|9|11|But when Christ appeared as a high priest of the good things that have come, then through the greater and more perfect tent (not made with hands, that is, not of this creation)
HEB|9|12|he entered once for all into the holy places, not by means of the blood of goats and calves but by means of his own blood, thus securing an eternal redemption.
HEB|9|13|For if the sprinkling of defiled persons with the blood of goats and bulls and with the ashes of a heifer sanctifies for the purification of the flesh,
HEB|9|14|how much more will the blood of Christ, who through the eternal Spirit offered himself without blemish to God, purify our conscience from dead works to serve the living God.
HEB|9|15|Therefore he is the mediator of a new covenant, so that those who are called may receive the promised eternal inheritance, since a death has occurred that redeems them from the transgressions committed under the first covenant.
HEB|9|16|For where a will is involved, the death of the one who made it must be established.
HEB|9|17|For a will takes effect only at death, since it is not in force as long as the one who made it is alive.
HEB|9|18|Therefore not even the first covenant was inaugurated without blood.
HEB|9|19|For when every commandment of the law had been declared by Moses to all the people, he took the blood of calves and goats, with water and scarlet wool and hyssop, and sprinkled both the book itself and all the people,
HEB|9|20|saying, "This is the blood of the covenant that God commanded for you."
HEB|9|21|And in the same way he sprinkled with the blood both the tent and all the vessels used in worship.
HEB|9|22|Indeed, under the law almost everything is purified with blood, and without the shedding of blood there is no forgiveness of sins.
HEB|9|23|Thus it was necessary for the copies of the heavenly things to be purified with these rites, but the heavenly things themselves with better sacrifices than these.
HEB|9|24|For Christ has entered, not into holy places made with hands, which are copies of the true things, but into heaven itself, now to appear in the presence of God on our behalf.
HEB|9|25|Nor was it to offer himself repeatedly, as the high priest enters the holy places every year with blood not his own,
HEB|9|26|for then he would have had to suffer repeatedly since the foundation of the world. But as it is, he has appeared once for all at the end of the ages to put away sin by the sacrifice of himself.
HEB|9|27|And just as it is appointed for man to die once, and after that comes judgment,
HEB|9|28|so Christ, having been offered once to bear the sins of many, will appear a second time, not to deal with sin but to save those who are eagerly waiting for him.
HEB|10|1|For since the law has but a shadow of the good things to come instead of the true form of these realities, it can never, by the same sacrifices that are continually offered every year, make perfect those who draw near.
HEB|10|2|Otherwise, would they not have ceased to be offered, since the worshipers, having once been cleansed, would no longer have any consciousness of sin?
HEB|10|3|But in these sacrifices there is a reminder of sin every year.
HEB|10|4|For it is impossible for the blood of bulls and goats to take away sins.
HEB|10|5|Consequently, when Christ came into the world, he said, "Sacrifices and offerings you have not desired, but a body have you prepared for me;
HEB|10|6|in burnt offerings and sin offerings you have taken no pleasure.
HEB|10|7|Then I said, 'Behold, I have come to do your will, O God, as it is written of me in the scroll of the book.'"
HEB|10|8|When he said above, "You have neither desired nor taken pleasure in sacrifices and offerings and burnt offerings and sin offerings" (these are offered according to the law),
HEB|10|9|then he added, "Behold, I have come to do your will." He abolishes the first in order to establish the second.
HEB|10|10|And by that will we have been sanctified through the offering of the body of Jesus Christ once for all.
HEB|10|11|And every priest stands daily at his service, offering repeatedly the same sacrifices, which can never take away sins.
HEB|10|12|But when Christ had offered for all time a single sacrifice for sins, he sat down at the right hand of God,
HEB|10|13|waiting from that time until his enemies should be made a footstool for his feet.
HEB|10|14|For by a single offering he has perfected for all time those who are being sanctified.
HEB|10|15|And the Holy Spirit also bears witness to us; for after saying,
HEB|10|16|"This is the covenant that I will make with them after those days, declares the Lord: I will put my laws on their hearts, and write them on their minds,"
HEB|10|17|then he adds, "I will remember their sins and their lawless deeds no more."
HEB|10|18|Where there is forgiveness of these, there is no longer any offering for sin.
HEB|10|19|Therefore, brothers, since we have confidence to enter the holy places by the blood of Jesus,
HEB|10|20|by the new and living way that he opened for us through the curtain, that is, through his flesh,
HEB|10|21|and since we have a great priest over the house of God,
HEB|10|22|let us draw near with a true heart in full assurance of faith, with our hearts sprinkled clean from an evil conscience and our bodies washed with pure water.
HEB|10|23|Let us hold fast the confession of our hope without wavering, for he who promised is faithful.
HEB|10|24|And let us consider how to stir up one another to love and good works,
HEB|10|25|not neglecting to meet together, as is the habit of some, but encouraging one another, and all the more as you see the Day drawing near.
HEB|10|26|For if we go on sinning deliberately after receiving the knowledge of the truth, there no longer remains a sacrifice for sins,
HEB|10|27|but a fearful expectation of judgment, and a fury of fire that will consume the adversaries.
HEB|10|28|Anyone who has set aside the law of Moses dies without mercy on the evidence of two or three witnesses.
HEB|10|29|How much worse punishment, do you think, will be deserved by the one who has spurned the Son of God, and has profaned the blood of the covenant by which he was sanctified, and has outraged the Spirit of grace?
HEB|10|30|For we know him who said, "Vengeance is mine; I will repay." And again, "The Lord will judge his people."
HEB|10|31|It is a fearful thing to fall into the hands of the living God.
HEB|10|32|But recall the former days when, after you were enlightened, you endured a hard struggle with sufferings,
HEB|10|33|sometimes being publicly exposed to reproach and affliction, and sometimes being partners with those so treated.
HEB|10|34|For you had compassion on those in prison, and you joyfully accepted the plundering of your property, since you knew that you yourselves had a better possession and an abiding one.
HEB|10|35|Therefore do not throw away your confidence, which has a great reward.
HEB|10|36|For you have need of endurance, so that when you have done the will of God you may receive what is promised.
HEB|10|37|For, "Yet a little while, and the coming one will come and will not delay;
HEB|10|38|but my righteous one shall live by faith, and if he shrinks back, my soul has no pleasure in him."
HEB|10|39|But we are not of those who shrink back and are destroyed, but of those who have faith and preserve their souls.
HEB|11|1|Now faith is the assurance of things hoped for, the conviction of things not seen.
HEB|11|2|For by it the people of old received their commendation.
HEB|11|3|By faith we understand that the universe was created by the word of God, so that what is seen was not made out of things that are visible.
HEB|11|4|By faith Abel offered to God a more acceptable sacrifice than Cain, through which he was commended as righteous, God commending him by accepting his gifts. And through his faith, though he died, he still speaks.
HEB|11|5|By faith Enoch was taken up so that he should not see death, and he was not found, because God had taken him. Now before he was taken he was commended as having pleased God.
HEB|11|6|And without faith it is impossible to please him, for whoever would draw near to God must believe that he exists and that he rewards those who seek him.
HEB|11|7|By faith Noah, being warned by God concerning events as yet unseen, in reverent fear constructed an ark for the saving of his household. By this he condemned the world and became an heir of the righteousness that comes by faith.
HEB|11|8|By faith Abraham obeyed when he was called to go out to a place that he was to receive as an inheritance. And he went out, not knowing where he was going.
HEB|11|9|By faith he went to live in the land of promise, as in a foreign land, living in tents with Isaac and Jacob, heirs with him of the same promise.
HEB|11|10|For he was looking forward to the city that has foundations, whose designer and builder is God.
HEB|11|11|By faith Sarah herself received power to conceive, even when she was past the age, since she considered him faithful who had promised.
HEB|11|12|Therefore from one man, and him as good as dead, were born descendants as many as the stars of heaven and as many as the innumerable grains of sand by the seashore.
HEB|11|13|These all died in faith, not having received the things promised, but having seen them and greeted them from afar, and having acknowledged that they were strangers and exiles on the earth.
HEB|11|14|For people who speak thus make it clear that they are seeking a homeland.
HEB|11|15|If they had been thinking of that land from which they had gone out, they would have had opportunity to return.
HEB|11|16|But as it is, they desire a better country, that is, a heavenly one. Therefore God is not ashamed to be called their God, for he has prepared for them a city.
HEB|11|17|By faith Abraham, when he was tested, offered up Isaac, and he who had received the promises was in the act of offering up his only son,
HEB|11|18|of whom it was said, "Through Isaac shall your offspring be named."
HEB|11|19|He considered that God was able even to raise him from the dead, from which, figuratively speaking, he did receive him back.
HEB|11|20|By faith Isaac invoked future blessings on Jacob and Esau.
HEB|11|21|By faith Jacob, when dying, blessed each of the sons of Joseph, bowing in worship over the head of his staff.
HEB|11|22|By faith Joseph, at the end of his life, made mention of the exodus of the Israelites and gave directions concerning his bones.
HEB|11|23|By faith Moses, when he was born, was hidden for three months by his parents, because they saw that the child was beautiful, and they were not afraid of the king's edict.
HEB|11|24|By faith Moses, when he was grown up, refused to be called the son of Pharaoh's daughter,
HEB|11|25|choosing rather to be mistreated with the people of God than to enjoy the fleeting pleasures of sin.
HEB|11|26|He considered the reproach of Christ greater wealth than the treasures of Egypt, for he was looking to the reward.
HEB|11|27|By faith he left Egypt, not being afraid of the anger of the king, for he endured as seeing him who is invisible.
HEB|11|28|By faith he kept the Passover and sprinkled the blood, so that the Destroyer of the firstborn might not touch them.
HEB|11|29|By faith the people crossed the Red Sea as if on dry land, but the Egyptians, when they attempted to do the same, were drowned.
HEB|11|30|By faith the walls of Jericho fell down after they had been encircled for seven days.
HEB|11|31|By faith Rahab the prostitute did not perish with those who were disobedient, because she had given a friendly welcome to the spies.
HEB|11|32|And what more shall I say? For time would fail me to tell of Gideon, Barak, Samson, Jephthah, of David and Samuel and the prophets-
HEB|11|33|who through faith conquered kingdoms, enforced justice, obtained promises, stopped the mouths of lions,
HEB|11|34|quenched the power of fire, escaped the edge of the sword, were made strong out of weakness, became mighty in war, put foreign armies to flight.
HEB|11|35|Women received back their dead by resurrection. Some were tortured, refusing to accept release, so that they might rise again to a better life.
HEB|11|36|Others suffered mocking and flogging, and even chains and imprisonment.
HEB|11|37|They were stoned, they were sawn in two, they were killed with the sword. They went about in skins of sheep and goats, destitute, afflicted, mistreated-
HEB|11|38|of whom the world was not worthy- wandering about in deserts and mountains, and in dens and caves of the earth.
HEB|11|39|And all these, though commended through their faith, did not receive what was promised,
HEB|11|40|since God had provided something better for us, that apart from us they should not be made perfect.
HEB|12|1|Therefore, since we are surrounded by so great a cloud of witnesses, let us also lay aside every weight, and sin which clings so closely, and let us run with endurance the race that is set before us,
HEB|12|2|looking to Jesus, the founder and perfecter of our faith, who for the joy that was set before him endured the cross, despising the shame, and is seated at the right hand of the throne of God.
HEB|12|3|Consider him who endured from sinners such hostility against himself, so that you may not grow weary or fainthearted.
HEB|12|4|In your struggle against sin you have not yet resisted to the point of shedding your blood.
HEB|12|5|And have you forgotten the exhortation that addresses you as sons? "My son, do not regard lightly the discipline of the Lord, nor be weary when reproved by him.
HEB|12|6|For the Lord disciplines the one he loves, and chastises every son whom he receives."
HEB|12|7|It is for discipline that you have to endure. God is treating you as sons. For what son is there whom his father does not discipline?
HEB|12|8|If you are left without discipline, in which all have participated, then you are illegitimate children and not sons.
HEB|12|9|Besides this, we have had earthly fathers who disciplined us and we respected them. Shall we not much more be subject to the Father of spirits and live?
HEB|12|10|For they disciplined us for a short time as it seemed best to them, but he disciplines us for our good, that we may share his holiness.
HEB|12|11|For the moment all discipline seems painful rather than pleasant, but later it yields the peaceful fruit of righteousness to those who have been trained by it.
HEB|12|12|Therefore lift your drooping hands and strengthen your weak knees,
HEB|12|13|and make straight paths for your feet, so that what is lame may not be put out of joint but rather be healed.
HEB|12|14|Strive for peace with everyone, and for the holiness without which no one will see the Lord.
HEB|12|15|See to it that no one fails to obtain the grace of God; that no "root of bitterness" springs up and causes trouble, and by it many become defiled;
HEB|12|16|that no one is sexually immoral or unholy like Esau, who sold his birthright for a single meal.
HEB|12|17|For you know that afterward, when he desired to inherit the blessing, he was rejected, for he found no chance to repent, though he sought it with tears.
HEB|12|18|For you have not come to what may be touched, a blazing fire and darkness and gloom and a tempest
HEB|12|19|and the sound of a trumpet and a voice whose words made the hearers beg that no further messages be spoken to them.
HEB|12|20|For they could not endure the order that was given, "If even a beast touches the mountain, it shall be stoned."
HEB|12|21|Indeed, so terrifying was the sight that Moses said, "I tremble with fear."
HEB|12|22|But you have come to Mount Zion and to the city of the living God, the heavenly Jerusalem, and to innumerable angels in festal gathering,
HEB|12|23|and to the assembly of the firstborn who are enrolled in heaven, and to God, the judge of all, and to the spirits of the righteous made perfect,
HEB|12|24|and to Jesus, the mediator of a new covenant, and to the sprinkled blood that speaks a better word than the blood of Abel.
HEB|12|25|See that you do not refuse him who is speaking. For if they did not escape when they refused him who warned them on earth, much less will we escape if we reject him who warns from heaven.
HEB|12|26|At that time his voice shook the earth, but now he has promised, "Yet once more I will shake not only the earth but also the heavens."
HEB|12|27|This phrase, "Yet once more," indicates the removal of things that are shaken- that is, things that have been made- in order that the things that cannot be shaken may remain.
HEB|12|28|Therefore let us be grateful for receiving a kingdom that cannot be shaken, and thus let us offer to God acceptable worship, with reverence and awe,
HEB|12|29|for our God is a consuming fire.
HEB|13|1|Let brotherly love continue.
HEB|13|2|Do not neglect to show hospitality to strangers, for thereby some have entertained angels unawares.
HEB|13|3|Remember those who are in prison, as though in prison with them, and those who are mistreated, since you also are in the body.
HEB|13|4|Let marriage be held in honor among all, and let the marriage bed be undefiled, for God will judge the sexually immoral and adulterous.
HEB|13|5|Keep your life free from love of money, and be content with what you have, for he has said, "I will never leave you nor forsake you."
HEB|13|6|So we can confidently say, "The Lord is my helper; I will not fear; what can man do to me?"
HEB|13|7|Remember your leaders, those who spoke to you the word of God. Consider the outcome of their way of life, and imitate their faith.
HEB|13|8|Jesus Christ is the same yesterday and today and forever.
HEB|13|9|Do not be led away by diverse and strange teachings, for it is good for the heart to be strengthened by grace, not by foods, which have not benefited those devoted to them.
HEB|13|10|We have an altar from which those who serve the tent have no right to eat.
HEB|13|11|For the bodies of those animals whose blood is brought into the holy places by the high priest as a sacrifice for sin are burned outside the camp.
HEB|13|12|So Jesus also suffered outside the gate in order to sanctify the people through his own blood.
HEB|13|13|Therefore let us go to him outside the camp and bear the reproach he endured.
HEB|13|14|For here we have no lasting city, but we seek the city that is to come.
HEB|13|15|Through him then let us continually offer up a sacrifice of praise to God, that is, the fruit of lips that acknowledge his name.
HEB|13|16|Do not neglect to do good and to share what you have, for such sacrifices are pleasing to God.
HEB|13|17|Obey your leaders and submit to them, for they are keeping watch over your souls, as those who will have to give an account. Let them do this with joy and not with groaning, for that would be of no advantage to you.
HEB|13|18|Pray for us, for we are sure that we have a clear conscience, desiring to act honorably in all things.
HEB|13|19|I urge you the more earnestly to do this in order that I may be restored to you the sooner.
HEB|13|20|Now may the God of peace who brought again from the dead our Lord Jesus, the great shepherd of the sheep, by the blood of the eternal covenant,
HEB|13|21|equip you with everything good that you may do his will, working in us that which is pleasing in his sight, through Jesus Christ, to whom be glory forever and ever. Amen.
HEB|13|22|I appeal to you, brothers, bear with my word of exhortation, for I have written to you briefly.
HEB|13|23|You should know that our brother Timothy has been released, with whom I shall see you if he comes soon.
HEB|13|24|Greet all your leaders and all the saints. Those who come from Italy send you greetings.
HEB|13|25|Grace be with all of you.
