NAH|1|1|An oracle concerning Nineveh. The book of the vision of Nahum the Elkoshite.
NAH|1|2|The LORD is a jealous and avenging God; the LORD takes vengeance and is filled with wrath. The LORD takes vengeance on his foes and maintains his wrath against his enemies.
NAH|1|3|The LORD is slow to anger and great in power; the LORD will not leave the guilty unpunished. His way is in the whirlwind and the storm, and clouds are the dust of his feet.
NAH|1|4|He rebukes the sea and dries it up; he makes all the rivers run dry. Bashan and Carmel wither and the blossoms of Lebanon fade.
NAH|1|5|The mountains quake before him and the hills melt away. The earth trembles at his presence, the world and all who live in it.
NAH|1|6|Who can withstand his indignation? Who can endure his fierce anger? His wrath is poured out like fire; the rocks are shattered before him.
NAH|1|7|The LORD is good, a refuge in times of trouble. He cares for those who trust in him,
NAH|1|8|but with an overwhelming flood he will make an end of Nineveh; he will pursue his foes into darkness.
NAH|1|9|Whatever they plot against the LORD he will bring to an end; trouble will not come a second time.
NAH|1|10|They will be entangled among thorns and drunk from their wine; they will be consumed like dry stubble.
NAH|1|11|From you, O Nineveh, has one come forth who plots evil against the LORD and counsels wickedness.
NAH|1|12|This is what the LORD says: "Although they have allies and are numerous, they will be cut off and pass away. Although I have afflicted you, O Judah, I will afflict you no more.
NAH|1|13|Now I will break their yoke from your neck and tear your shackles away."
NAH|1|14|The LORD has given a command concerning you, Nineveh: "You will have no descendants to bear your name. I will destroy the carved images and cast idols that are in the temple of your gods. I will prepare your grave, for you are vile."
NAH|1|15|Look, there on the mountains, the feet of one who brings good news, who proclaims peace! Celebrate your festivals, O Judah, and fulfill your vows. No more will the wicked invade you; they will be completely destroyed.
NAH|2|1|An attacker advances against you, Nineveh. Guard the fortress, watch the road, brace yourselves, marshal all your strength!
NAH|2|2|The LORD will restore the splendor of Jacob like the splendor of Israel, though destroyers have laid them waste and have ruined their vines.
NAH|2|3|The shields of his soldiers are red; the warriors are clad in scarlet. The metal on the chariots flashes on the day they are made ready; the spears of pine are brandished.
NAH|2|4|The chariots storm through the streets, rushing back and forth through the squares. They look like flaming torches; they dart about like lightning.
NAH|2|5|He summons his picked troops, yet they stumble on their way. They dash to the city wall; the protective shield is put in place.
NAH|2|6|The river gates are thrown open and the palace collapses.
NAH|2|7|It is decreed that the city be exiled and carried away. Its slave girls moan like doves and beat upon their breasts.
NAH|2|8|Nineveh is like a pool, and its water is draining away. "Stop! Stop!" they cry, but no one turns back.
NAH|2|9|Plunder the silver! Plunder the gold! The supply is endless, the wealth from all its treasures!
NAH|2|10|She is pillaged, plundered, stripped! Hearts melt, knees give way, bodies tremble, every face grows pale.
NAH|2|11|Where now is the lions' den, the place where they fed their young, where the lion and lioness went, and the cubs, with nothing to fear?
NAH|2|12|The lion killed enough for his cubs and strangled the prey for his mate, filling his lairs with the kill and his dens with the prey.
NAH|2|13|"I am against you," declares the LORD Almighty. "I will burn up your chariots in smoke, and the sword will devour your young lions. I will leave you no prey on the earth. The voices of your messengers will no longer be heard."
NAH|3|1|Woe to the city of blood, full of lies, full of plunder, never without victims!
NAH|3|2|The crack of whips, the clatter of wheels, galloping horses and jolting chariots!
NAH|3|3|Charging cavalry, flashing swords and glittering spears! Many casualties, piles of dead, bodies without number, people stumbling over the corpses-
NAH|3|4|all because of the wanton lust of a harlot, alluring, the mistress of sorceries, who enslaved nations by her prostitution and peoples by her witchcraft.
NAH|3|5|"I am against you," declares the LORD Almighty. "I will lift your skirts over your face. I will show the nations your nakedness and the kingdoms your shame.
NAH|3|6|I will pelt you with filth, I will treat you with contempt and make you a spectacle.
NAH|3|7|All who see you will flee from you and say, 'Nineveh is in ruins-who will mourn for her?' Where can I find anyone to comfort you?"
NAH|3|8|Are you better than Thebes, situated on the Nile, with water around her? The river was her defense, the waters her wall.
NAH|3|9|Cush and Egypt were her boundless strength; Put and Libya were among her allies.
NAH|3|10|Yet she was taken captive and went into exile. Her infants were dashed to pieces at the head of every street. Lots were cast for her nobles, and all her great men were put in chains.
NAH|3|11|You too will become drunk; you will go into hiding and seek refuge from the enemy.
NAH|3|12|All your fortresses are like fig trees with their first ripe fruit; when they are shaken, the figs fall into the mouth of the eater.
NAH|3|13|Look at your troops- they are all women! The gates of your land are wide open to your enemies; fire has consumed their bars.
NAH|3|14|Draw water for the siege, strengthen your defenses! Work the clay, tread the mortar, repair the brickwork!
NAH|3|15|There the fire will devour you; the sword will cut you down and, like grasshoppers, consume you. Multiply like grasshoppers, multiply like locusts!
NAH|3|16|You have increased the number of your merchants till they are more than the stars of the sky, but like locusts they strip the land and then fly away.
NAH|3|17|Your guards are like locusts, your officials like swarms of locusts that settle in the walls on a cold day- but when the sun appears they fly away, and no one knows where.
NAH|3|18|O king of Assyria, your shepherds slumber; your nobles lie down to rest. Your people are scattered on the mountains with no one to gather them.
NAH|3|19|Nothing can heal your wound; your injury is fatal. Everyone who hears the news about you claps his hands at your fall, for who has not felt your endless cruelty?
