MAL|1|1|Oraculum. Verbum Domini ad Israel in manu Malachiae.
MAL|1|2|" Dilexi vos, dicit Dominus, et dixistis: "In quo dilexisti nos?". Nonne frater erat Esau Iacob?, dicit Dominus; et dilexi Iacob,
MAL|1|3|Esau autem odio habui et posui montes eius in solitudinem et hereditatem eius thoibus deserti.
MAL|1|4|Quod si dixerit Edom: "Destructi sumus, sed revertentes aedificabimus, quae destructa sunt", haec dicit Dominus exercituum: Isti aedificabunt, et ego destruam; et vocabuntur 'Termini impietatis' et 'Populus, cui iratus est Dominus usque in aeternum'.
MAL|1|5|Et oculi vestri videbunt, et vos dicetis: "Magnificatus est Dominus ultra terminos Israel".
MAL|1|6|Filius honorat patrem, et servus dominum suum. Si ergo pater ego sum, ubi est honor meus? Et si Dominus ego sum, ubi est timor meus?, dicit Dominus exercituum ad vos, o sacerdotes, qui despicitis nomen meum et dicitis: "In quo despeximus nomen tuum?".
MAL|1|7|Offertis super altare meum panem pollutum et dicitis: "In quo polluimus te?". In eo quod dicitis: "Mensa Domini contemptibilis est".
MAL|1|8|Si offeratis caecum ad immolandum, nonne malum est? Et si offeratis claudum et languidum, nonne malum est? Offer illud duci tuo, si placuerit ei, aut si susceperit faciem tuam!, dicit Dominus exercituum.
MAL|1|9|Sed nunc deprecamini vultum Dei, ut misereatur vestri! De manu enim vestra factum est hoc. Num suscipiet facies vestras?, dicit Dominus exercituum.
MAL|1|10|Quis est in vobis, qui claudat ostia, ne incendatis altare meum gratuito? Non est mihi voluntas in vobis, dicit Dominus exercituum; et munus non suscipiam de manu vestra.
MAL|1|11|Ab ortu enim solis usque ad occasum magnum est nomen meum in gentibus, et in omni loco sacrificatur et offertur nomini meo oblatio munda, quia magnum nomen meum in gentibus, dicit Dominus exercituum.
MAL|1|12|Vos autem polluistis illud in eo quod dicitis: "Mensa Domini contaminata est, et contemptibilis esca eius".
MAL|1|13|Et dicitis: "Quantus labor!", et despicitis illam, dicit Dominus exercituum. Et infertis de rapinis claudum et languidum et infertis sicut munus. Numquid suscipiam illud de manu vestra?, dicit Dominus.
MAL|1|14|Maledictus dolosus, qui habet in grege suo masculum et votum faciens immolat debile Domino. Quia Rex magnus ego, dicit Dominus exercituum, et nomen meum horribile in gentibus.
MAL|2|1|Et nunc ad vos mandatum hoc, o sacerdotes.
MAL|2|2|Si nolueritis audi re et si nolueritis ponere super cor, ut detis gloriam nomini meo, ait Dominus exercituum, mittam in vos maledictionem et maledicam benedictionibus vestris; et maledicam illis, quoniam non posuistis super cor.
MAL|2|3|Ecce ego abscindam vobis brachiumet dispergam stercus super vultum vestrum,stercus sollemnitatum vestrarum,et assumet vos secum;
MAL|2|4|et scietis quia misi ad vos mandatum istud,ut esset pactum meum cum Levi,dicit Dominus exercituum.
MAL|2|5|Pactum meum fuit cum eo vitae et pacis,et dedi haec ei simul cum timore, et timuit meet a facie nominis mei pavebat.
MAL|2|6|Lex veritatis fuit in ore eius,et iniquitas non est inventa in labiis eius;in pace et in aequitate ambulavit mecumet multos avertit ab iniquitate.
MAL|2|7|Labia enim sacerdotis custodiunt scientiam,et legem requirunt ex ore eius,quia angelus Domini exercituum est.
MAL|2|8|Vos autem recessistis de viaet scandalizastis plurimos in lege;irritum fecistis pactum Levi,dicit Dominus exercituum;
MAL|2|9|propter quod et ego dedi voscontemptibiles et humiles omnibus populis,sicut non servastis vias measet accepistis personam in lege.
MAL|2|10|Numquid non pater unus omnium nostrum? Numquid non Deus unus creavit nos? Quare ergo dolum facit unusquisque nostrum cum fratre suo, violans pactum patrum nostrorum?
MAL|2|11|Dolum fecit Iuda, et abominatio facta est in Israel et in Ierusalem, quia contaminavit Iuda sanctuarium Domini, quod diligit, et accepit uxorem filiam dei alieni.
MAL|2|12|Disperdet Dominus virum, qui fecerit hoc, filium et nepotem, de tabernaculis Iacob et de offerentibus munus Domino exercituum.
MAL|2|13|Et hoc rursum facitis: operitis lacrimis altare Domini, fletu et mugitu, ita ut non respiciam ultra ad sacrificium nec accipiam placabile quid de manu vestra;
MAL|2|14|et dicitis: "Quam ob causam?". Quia Dominus testificatus est inter te et uxorem adulescentiae tuae, cui tu factus es infidelis; et haec particeps tua et uxor foederis tui.
MAL|2|15|Nonne unitatem fecit carnis et spiritus? Et quid unitas quaerit nisi semen a Deo? Custodite ergo spiritum vestrum; et uxori adulescentiae tuae noli esse infidelis.
MAL|2|16|Si quis odio dimittit, dicit Dominus, Deus Israel, operit iniquitas vestimentum eius, dicit Dominus exercituum. Custodite spiritum vestrum et nolite esse infideles.
MAL|2|17|Laborare facitis Dominum in sermonibus vestris et dicitis: "In quo eum facimus laborare?". In eo quod dicitis: "Omnis, qui facit malum, bonus est in conspectu Domini, et tales ei placent" aut: "Ubi est Deus iudicii?".
MAL|3|1|Ecce ego mittam angelum meum, et praeparabit viam an te faciem meam; et statim veniet ad templum suum Dominator, quem vos quaeritis, et angelus testamenti, quem vos vultis. Ecce venit, dicit Dominus exercituum;
MAL|3|2|et quis poterit sustinere diem adventus eius, et quis stabit, cum apparebit? Ipse enim quasi ignis conflans et quasi herba fullonum;
MAL|3|3|et sedebit conflans et emundans argentum et purgabit filios Levi et colabit eos quasi aurum et quasi argentum, et erunt Domino offerentes sacrificia in iustitia.
MAL|3|4|Et placebit Domino sacrificium Iudae et Ierusalem sicut diebus pristinis et sicut annis antiquis.
MAL|3|5|Et accedam ad vos in iudicio; et ero testis velox maleficis et adulteris et periuris et, qui opprimunt mercennarios, viduas et pupillos et flectunt ius peregrinorum nec timuerunt me, dicit Dominus exercituum.
MAL|3|6|Ego enim Dominus et non mutatus sum;sed vos, filii lacob, nondum ad finem pervenistis.
MAL|3|7|A diebus enim patrum vestrorumrecessistis a praeceptis legitimis meis et non custodistis ea.Revertimini ad me,et revertar ad vos,dicit Dominus exercituum.Et dicitis: "In quo revertemur?".
MAL|3|8|Numquid homo potest defraudare Deum?Sed vos defraudatis me.Et dicitis: "In quo defraudavimus te?".In decimis et in primitiis.
MAL|3|9|Maledictione vos maledicti estis,quia me vos defraudatis, gens tota.
MAL|3|10|Inferte omnem decimam in horreum,et sit cibus in domo mea;et probate me super hoc,dicit Dominus exercituum:si non aperuero vobis cataractas caeliet effudero vobis benedictionem usque ad abundantiam
MAL|3|11|et increpabo pro vobis devorantem,et non corrumpet fructum terrae,nec erit sterilis vobis vinea in agro,dicit Dominus exercituum.
MAL|3|12|Et beatos vos dicent omnes gentes;eritis enim vos terra desiderabilis,dicit Dominus exercituum.
MAL|3|13|Invaluerunt super me verba vestra, dicit Dominus;
MAL|3|14|et dicitis: "Quid locuti sumus contra te?". Dicitis: "Vanum est servire Deo; et, quod emolumentum, quia custodivimus praecepta eius et quia ambulavimus tristes coram Domino exercituum?
MAL|3|15|Ergo nunc beatos dicimus arrogantes; siquidem aedificati sunt facientes impietatem et tentaverunt Deum et salvi facti sunt".
MAL|3|16|Tunc locuti sunt timentes Dominum, unusquisque cum proximo suo. Et attendit Dominus et audivit; et scriptus est liber memorabilium coram eo timentibus Dominum et cogitantibus nomen eius.
MAL|3|17|Erunt mihi, ait Dominus exercituum, in die, qua ego facio in peculium; et parcam eis, sicut parcit vir filio suo servienti sibi.
MAL|4|1|Rursum videbitis quid sit inter iustum et impium, inter servientem Deo et non servientem ei.
MAL|4|2|Ecce enim dies veniet succensa quasi caminus; et erunt omnes superbi et omnes facientes impietatem stipula; et inflammabit eos dies veniens, dicit Dominus exercituum, quae non derelinquet eis radicem et ramum.
MAL|4|3|Et orietur vobis timentibus nomen meum sol iustitiae et sanitas in pennis eius; et egrediemini et salietis sicut vituli saginati
MAL|4|4|et calcabitis impios, cum fuerint cinis sub planta pedum vestrorum in die, quam ego facio, dicit Dominus exercituum.
MAL|4|5|Mementote legis Moysi servi mei,cui mandaviin Horeb ad omnem Israelpraecepta et iudicia.
MAL|4|6|Ecce ego mittam vobisEliam prophetam,antequam veniat dies Dominimagnus et horribilis;
MAL|4|7|et convertet cor patrum ad filioset cor filiorum ad patres eorum,ne veniam et percutiamterram anathemate "
