LUKE|1|1|Через те, що багато-хто брались складати оповість про справи, які стались між нами,
LUKE|1|2|як нам ті розповіли, хто спочатку були самовидцями й слугами Слова,
LUKE|1|3|тому й я, все від першої хвилі докладно розвідавши, забажав описати за порядком для тебе, високодостойний Теофіле,
LUKE|1|4|щоб пізнав ти істоту науки, якої навчився.
LUKE|1|5|За днів царя юдейського Ірода був один священик, на ім'я Захарій, з денної черги Авія, та дружина його із дочок Ааронових, а ім'я їй Єлисавета.
LUKE|1|6|І обоє вони були праведні перед Богом, бездоганно сповняючи заповіді й постанови Господні.
LUKE|1|7|А дитини не мали вони, бо Єлисавета неплідна була, та й віку старого обоє були.
LUKE|1|8|І ось раз, як у порядку своєї черги він служив перед Богом,
LUKE|1|9|за звичаєм священства, жеребком йому випало до Господнього храму ввійти й покадити.
LUKE|1|10|Під час же кадіння вся безліч народу молилась знадвору.
LUKE|1|11|І з'явивсь йому Ангол Господній, ставши праворуч кадильного жертівника.
LUKE|1|12|І стривоживсь Захарій, побачивши, і острах на нього напав.
LUKE|1|13|А Ангол до нього промовив: Не бійся, Захаріє, бо почута молитва твоя, і дружина твоя Єлисавета сина породить тобі, ти ж даси йому ймення Іван.
LUKE|1|14|І він буде на радість та втіху тобі, і з його народження багато-хто втішаться.
LUKE|1|15|Бо він буде великий у Господа, ні вина, ні п'янкого напою не питиме, і наповниться Духом Святим ще з утроби своєї матері.
LUKE|1|16|І багато синів із Ізраїля він наверне до їхнього Господа Бога.
LUKE|1|17|І він сам перед Ним буде йти в духу й силі Іллі, щоб серця батьків привернути до дітей, і неслухняних до мудрости праведних, щоб готових людей спорядити для Господа.
LUKE|1|18|І промовив Захарій до Ангола: Із чого пізнаю я це? Я ж старий, та й дружина моя вже похилого віку...
LUKE|1|19|А Ангол прорік йому в відповідь: Я Гавриїл, що стою перед Богом; мене послано, щоб говорити з тобою, і звістити тобі про цю Добру Новину.
LUKE|1|20|І замовкнеш ось ти, і говорити не зможеш аж до дня, коли станеться це, за те, що ти віри не йняв був словам моїм, які збудуться часу свого!
LUKE|1|21|А люди чекали Захарія, та й дивувались, чого забаривсь він у храмі.
LUKE|1|22|Коли ж вийшов, не міг говорити до них, і вони зрозуміли, що видіння він бачив у храмі. А він тільки знаки їм давав, і залишився німий...
LUKE|1|23|І як дні його служби скінчились, він вернувся до дому свого.
LUKE|1|24|А після тих днів зачала його дружина Єлисавета, і таїлась п'ять місяців, кажучи:
LUKE|1|25|Так для мене Господь учинив за тих днів, коли зглянувся Він, щоб зняти наругу мою між людьми!
LUKE|1|26|А шостого місяця від Бога був посланий Ангол Гавриїл у галілейське місто, що йому на ім'я Назарет,
LUKE|1|27|до діви, що заручена з мужем була, на ім'я йому Йосип, із дому Давидового, а ім'я діві Марія.
LUKE|1|28|І, ввійшовши до неї, промовив: Радій, благодатная, Господь із тобою! Ти благословенна між жонами!
LUKE|1|29|Вона ж затривожилась словом, та й стала роздумувати, що б то значило це привітання.
LUKE|1|30|А Ангол промовив до неї: Не бійся, Маріє, бо в Бога благодать ти знайшла!
LUKE|1|31|І ось ти в утробі зачнеш, і Сина породиш, і даси Йому ймення Ісус.
LUKE|1|32|Він же буде Великий, і Сином Всевишнього званий, і Господь Бог дасть Йому престола Його батька Давида.
LUKE|1|33|І повік царюватиме Він у домі Якова, і царюванню Його не буде кінця.
LUKE|1|34|А Марія озвалась до Ангола: Як же станеться це, коли мужа не знаю?...
LUKE|1|35|І Ангол промовив у відповідь їй: Дух Святий злине на тебе, і Всевишнього сила обгорне тебе, через те то й Святе, що народиться, буде Син Божий!
LUKE|1|36|А ото твоя родичка Єлисавета і вона зачала в своїй старості сина, і оце шостий місяць для неї, яку звуть неплідною.
LUKE|1|37|Бо для Бога нема неможливої жадної речі!
LUKE|1|38|А Марія промовила: Я ж Господня раба: нехай буде мені згідно з словом твоїм! І відійшов Ангол від неї.
LUKE|1|39|Тими днями зібралась Марія й пішла, поспішаючи, у гірську околицю, у місто Юдине.
LUKE|1|40|І ввійшла вона в дім Захарія, та й поздоровила Єлисавету.
LUKE|1|41|Коли ж Єлисавета зачула Маріїн привіт, затріпотала дитина в утробі її. І Єлисавета наповнилась Духом Святим,
LUKE|1|42|і скрикнула голосом гучним, та й прорекла: Благословенна Ти між жонами, і благословенний Плід утроби твоєї!
LUKE|1|43|І звідкіля мені це, що до мене прийшла мати мого Господа?
LUKE|1|44|Бо як тільки в вухах моїх голос привіту твого забринів, від радощів затріпотала дитина в утробі моїй!
LUKE|1|45|Блаженна ж та, що повірила, бо сповниться проречене їй від Господа!
LUKE|1|46|А Марія промовила: Величає душа моя Господа,
LUKE|1|47|і радіє мій дух у Бозі, Спасі моїм,
LUKE|1|48|що зглянувся Він на покору Своєї раби, бо ось від часу цього всі роди мене за блаженну вважатимуть,
LUKE|1|49|бо велике вчинив мені Потужний! Його ж Імення святе,
LUKE|1|50|і милість Його з роду в рід на тих, хто боїться Його!
LUKE|1|51|Він показує міць Свого рамена, розпорошує тих, хто пишається думкою серця свого!
LUKE|1|52|Він могутніх скидає з престолів, підіймає покірливих,
LUKE|1|53|удовольняє голодних добром, а багатих пускає ні з чим!
LUKE|1|54|Пригорнув Він Ізраїля, Свого слугу, щоб милість згадати,
LUKE|1|55|як прорік був Він нашим отцям, Аврааму й насінню його аж повіки!
LUKE|1|56|І залишалась у неї Марія щось місяців зо три, та й вернулась до дому свого.
LUKE|1|57|А Єлисаветі настав час родити, і сина вона породила.
LUKE|1|58|І почули сусіди й родина її, що Господь Свою милість велику на неї послав, та й утішалися разом із нею.
LUKE|1|59|І сталося восьмого дня, прийшли, щоб обрізати дитя, і хотіли назвати його йменням батька його Захарій.
LUKE|1|60|І озвалася мати його та й сказала: Ні, нехай названий буде Іван!
LUKE|1|61|А до неї сказали: Таж у родині твоїй нема жадного, який названий був тим ім'ям!
LUKE|1|62|І кивали до батька його, як хотів би назвати його?
LUKE|1|63|Попросивши ж табличку, написав він слова: Іван імення йому. І всі дивувались.
LUKE|1|64|І в тій хвилі уста та язик розв'язались йому, і він став говорити, благословляючи Бога!
LUKE|1|65|І страх обгорнув усіх їхніх сусідів, і по всіх верховинах юдейських пронеслася чутка про це все...
LUKE|1|66|А всі, що почули, розважали у серці своїм та казали: Чим то буде дитина оця?... І Господня рука була з нею.
LUKE|1|67|Його ж батько Захарій наповнився Духом Святим, та й став пророкувати й казати:
LUKE|1|68|Благословенний Господь, Бог Ізраїлів, що зглянувся й визволив люд Свій!
LUKE|1|69|Він ріг спасіння підніс нам у домі Давида, Свого слуги,
LUKE|1|70|як був заповів відвіку устами святих пророків Своїх,
LUKE|1|71|що від ворогів наших визволить нас, та з руки всіх наших ненависників,
LUKE|1|72|що вчинить Він милість нашим отцям, і буде пригадувати Свій святий заповіт,
LUKE|1|73|що дотримає й нам ту присягу, якою Він присягавсь Авраамові, отцю нашому,
LUKE|1|74|щоб ми, визволившись із руки ворогів, служили безстрашно Йому
LUKE|1|75|у святості й праведності перед Ним по всі дні життя нашого.
LUKE|1|76|Ти ж, дитино, станеш пророком Всевишнього, бо будеш ходити перед Господом, щоб дорогу Йому приготувати,
LUKE|1|77|щоб народу Його дати пізнати спасіння у відпущенні їхніх гріхів,
LUKE|1|78|через велике милосердя нашого Бога, що ним Схід із висоти нас відвідав,
LUKE|1|79|щоб світити всім тим, хто перебуває в темряві й тіні смертельній, щоб спрямувати наші ноги на дорогу миру!
LUKE|1|80|А дитина росла, і скріплялась на дусі, і перебувала в пустинях до дня свого з'явлення перед Ізраїлем.
LUKE|2|1|І трапилося тими днями, вийшов наказ царя Августа переписати всю землю.
LUKE|2|2|Цей перепис перший відбувся тоді, коли владу над Сирією мав Квіріній.
LUKE|2|3|І всі йшли записатися, кожен у місто своє.
LUKE|2|4|Пішов теж і Йосип із Галілеї, із міста Назарету, до Юдеї, до міста Давидового, що зветься Віфлеєм, бо походив із дому та з роду Давидового,
LUKE|2|5|щоб йому записатись із Марією, із ним зарученою, що була вагітна.
LUKE|2|6|І сталось, як були вони там, то настав їй день породити.
LUKE|2|7|І породила вона свого Первенця Сина, і Його сповила, і до ясел поклала Його, бо в заїзді місця не стало для них...
LUKE|2|8|А в тій стороні були пастухи, які пильнували на полі, і нічної пори вартували отару свою.
LUKE|2|9|Аж ось Ангол Господній з'явивсь коло них, і слава Господня осяяла їх. І вони перестрашились страхом великим...
LUKE|2|10|Та Ангол промовив до них: Не лякайтесь, бо я ось благовіщу вам радість велику, що станеться людям усім.
LUKE|2|11|Бо сьогодні в Давидовім місті народився для вас Спаситель, Який є Христос Господь.
LUKE|2|12|А ось вам ознака: Дитину сповиту ви знайдете, що в яслах лежатиме.
LUKE|2|13|І ось раптом з'явилася з Анголом сила велика небесного війська, що Бога хвалили й казали:
LUKE|2|14|Слава Богу на висоті, і на землі мир, у людях добра воля!
LUKE|2|15|І сталось, коли Анголи відійшли від них в небо, пастухи зачали говорити один одному: Ходім до Віфлеєму й побачмо, що сталося там, про що сповістив нас Господь.
LUKE|2|16|І прийшли, поспішаючи, і знайшли там Марію та Йосипа, та Дитинку, що в яслах лежала.
LUKE|2|17|А побачивши, розповіли про все те, що про Цю Дитину було їм звіщено.
LUKE|2|18|І всі, хто почув, дивувались тому, що їм пастухи говорили...
LUKE|2|19|А Марія оці всі слова зберігала, розважаючи, у серці своїм.
LUKE|2|20|Пастухи ж повернулись, прославляючи й хвалячи Бога за все, що почули й побачили, так як їм було сказано.
LUKE|2|21|Коли ж виповнились вісім день, щоб обрізати Його, то Ісусом назвали Його, як був Ангол назвав, перше ніж Він в утробі зачався.
LUKE|2|22|А коли за Законом Мойсея минулися дні їхнього очищення, то до Єрусалиму принесли Його, щоб поставити Його перед Господом,
LUKE|2|23|як у Законі Господнім написано: Кожне дитя чоловічої статі, що розкриває утробу, має бути посвячене Господу,
LUKE|2|24|і щоб жертву скласти, як у Законі Господньому сказано, пару горличат або двоє голубенят.
LUKE|2|25|І ото був в Єрусалимі один чоловік, йому ймення Семен, людина праведна та благочестива, що потіхи чекав для Ізраїля. І Святий Дух був на ньому.
LUKE|2|26|І від Духа Святого йому було звіщено смерти не бачити, перше ніж побачить Христа Господнього.
LUKE|2|27|І Дух у храм припровадив його. І як внесли Дитину Ісуса батьки, щоб за Нього вчинити звичаєм законним,
LUKE|2|28|тоді взяв він на руки Його, хвалу Богу віддав та й промовив:
LUKE|2|29|Нині відпускаєш раба Свого, Владико, за словом Твоїм із миром,
LUKE|2|30|бо побачили очі мої Спасіння Твоє,
LUKE|2|31|яке Ти приготував перед всіма народами,
LUKE|2|32|Світло на просвіту поганам і на славу народу Твого Ізраїля!
LUKE|2|33|І дивувалися батько Його й мати тим, що про Нього було розповіджене.
LUKE|2|34|А Семен їх поблагословив та й прорік до Марії, Його матері: Ось призначений Цей багатьом на падіння й уставання в Ізраїлі, і на знак сперечання,
LUKE|2|35|і меч душу прошиє самій же тобі, щоб відкрились думки сердець багатьох!
LUKE|2|36|Була й Анна пророчиця, дочка Фануїлова з племени Асирового, вона дожила до глибокої старости, живши з мужем сім років від свого дівування,
LUKE|2|37|удова років вісімдесяти й чотирьох, що не відлучалась від храму, служачи Богові вдень і вночі постами й молитвами.
LUKE|2|38|І години тієї вона надійшла, Бога славила та говорила про Нього всім, хто визволення Єрусалиму чекав.
LUKE|2|39|А як виконали за Законом Господнім усе, то вернулись вони в Галілею, до міста свого Назарету.
LUKE|2|40|А Дитина росла та зміцнялася духом, набираючись мудрости. І благодать Божа на Ній пробувала.
LUKE|2|41|А батьки Його щорічно ходили до Єрусалиму на свято Пасхи.
LUKE|2|42|І коли мав Він дванадцять років, вони за звичаєм на свято пішли.
LUKE|2|43|Як дні ж свята скінчились були, і вертались вони, молодий Ісус в Єрусалимі лишився, а Йосип та мати Його не знали того.
LUKE|2|44|Вони думали, що Він із подорожніми йде; пройшли день дороги, та й стали шукати Його поміж родичами та знайомими.
LUKE|2|45|Але, не знайшовши, вернулися в Єрусалим, та й шукали Його.
LUKE|2|46|І сталось, що третього дня відшукали у храмі Його, як сидів серед учителів, і вислухував їх, і запитував їх.
LUKE|2|47|Усі ж, хто слухав Його, дивувалися розумові та Його відповідям.
LUKE|2|48|І як вони Його вгледіли, то здивувались, а мати сказала до Нього: Дитино, чому так Ти зробив нам? Ось Твій батько та я із журбою шукали Тебе...
LUKE|2|49|А Він їм відказав: Чого ж ви шукали Мене? Хіба ви не знали, що повинно Мені бути в тому, що належить Моєму Отцеві?
LUKE|2|50|Та не зрозуміли вони того слова, що Він їм говорив.
LUKE|2|51|І пішов Він із ними, і прибув у Назарет, і був їм слухняний. А мати Його зберігала оці всі слова в своїм серці.
LUKE|2|52|А Ісус зростав мудрістю, і віком та благодаттю, у Бога й людей.
LUKE|3|1|У п'ятнадцятий рік панування Тиверія кесаря, коли Понтій Пилат панував над Юдеєю, коли в Галілеї тетрархом був Ірод, а Пилип, його брат, був тетрархом Ітуреї й землі Трахонітської, за тетрарха Лісанія в Авіліні,
LUKE|3|2|за первосвящеників Анни й Кайяфи було Боже слово в пустині Іванові, сину Захарія.
LUKE|3|3|І він перейшов усю землю Йорданську, проповідуючи хрищення покаяння для прощення гріхів,
LUKE|3|4|як написано в книзі пророцтва пророка Ісаї: Голос того, хто кличе: У пустині готуйте дорогу для Господа, рівняйте стежки Йому!
LUKE|3|5|Нехай кожна долина наповниться, гора ж кожна та пригорок знизиться, що нерівне, нехай випростовується, а дороги вибоїсті стануть гладенькі,
LUKE|3|6|і кожна людина побачить Боже спасіння!
LUKE|3|7|А Іван говорив до людей, хто приходив, христитися в нього: Роде зміїний, хто навчив вас тікати від гніву майбутнього?
LUKE|3|8|Отож, учиніть гідний плід покаяння. І не починайте казати в собі: Маємо батька Авраама. Бо кажу вам, що Бог може піднести дітей Авраамові з цього каміння.
LUKE|3|9|Бо вже он до коріння дерев і сокира прикладена: кожне ж дерево, що доброго плоду не родить, буде зрубане та до огню буде вкинене.
LUKE|3|10|А люди питали його й говорили: Що ж нам робити?
LUKE|3|11|І сказав він у відповідь їм: У кого дві сорочці, нехай дасть немаючому; а хто має поживу, нехай робить так само.
LUKE|3|12|І приходили й митники, щоб христитись від нього, і питали його: Учителю, що ми маємо робити?
LUKE|3|13|А він їм казав: Не стягайте нічого над те, що вам звелено.
LUKE|3|14|Питали ж його й вояки й говорили: А нам що робити? І він їм відповів: Нікого не кривдьте, ані не оскаржайте фальшиво, удовольняйтесь платнею своєю.
LUKE|3|15|Коли ж усі люди чекали, і в серцях своїх думали всі про Івана, чи то він не Христос,
LUKE|3|16|Іван відповідав усім, кажучи: Я хрищу вас водою, але йде ось Потужніший за мене, що Йому розв'язати ремінця від Його взуття я негідний, Він христитиме вас Святим Духом й огнем!
LUKE|3|17|У руці Своїй має Він віячку, і перечистить Свій тік: пшеницю збере до засіків Своїх, а полову попалить ув огні невгасимім.
LUKE|3|18|Тож багато навчав він і іншого, звіщаючи Добру Новину народові.
LUKE|3|19|А Ірод тетрарх, що Іван докоряв йому за Іродіяду, дружину брата свого, і за все зло, яке заподіяв був Ірод,
LUKE|3|20|до всього додав іще й те, що Івана замкнув до в'язниці.
LUKE|3|21|І сталося, як христились усі люди, і як Ісус, охристившись, молився, розкрилося небо,
LUKE|3|22|і Дух Святий злинув на Нього в тілесному вигляді, як голуб, і голос із неба почувся, що мовив: Ти Син Мій Улюблений, що Я вподобав Тебе!
LUKE|3|23|А Сам Ісус, розпочинаючи, мав років із тридцять, бувши, як думано, сином Йосипа, Ілія,
LUKE|3|24|сина Маттатового, сина Левіїного, сина Мелхіїного, сина Яннаєвого, сина Йосипового,
LUKE|3|25|сина Маттатієвого, сина Амосова, сина Наумового, сина Еслієвого, сина Наггеєвого,
LUKE|3|26|сина Маатового, сина Маттатієвого, сина Семенієвого, сина Йосихового, сина Йодаєвого,
LUKE|3|27|сина Йоананового, сина Рисаєвого, сина Зоровавелевого, сина Салатіїлового, сина Нирієвого,
LUKE|3|28|сина Мелхієвого, сина Аддієвого, сина Косамового, сина Елмадамового, сина Ірового,
LUKE|3|29|сина Ісуєвого, сина Еліезерового, сина Йоримового, сина Маттатієвого, сина Левієвого,
LUKE|3|30|сина Семенового, сина Юдиного, сина Йосипового, сина Йонамового, сина Еліякимового,
LUKE|3|31|сина Мелеаєвого, сина Меннаєвого, сина Маттатаєвого, сина Натамового, сина Давидового,
LUKE|3|32|сина Єссеєвого, сина Йовидового, сина Воозового, сина Салаєвого, сина Наассонового,
LUKE|3|33|сина Амінадавого, сина Адмінієвого, сина Арнієвого, сина Есромового, сина Фаресового, сина Юдиного,
LUKE|3|34|сина Яковлевого, сина Ісакового, сина Авраамового, сина Тариного, сина Нахорового,
LUKE|3|35|сина Серухового, сина Рагавового, сина Фалекового, сина Еверового, сина Салиного,
LUKE|3|36|сина Каїнамового, сина Арфаксадового, сина Симового, сина Ноєвого, сина Ламехового,
LUKE|3|37|сина Матусалового, сина Енохового, сина Яретового, сина Малелеїлового, сина Каїнамового,
LUKE|3|38|сина Еносового, сина Ситового, сина Адамового, Сином Божим.
LUKE|4|1|А Ісус, повний Духа Святого, вернувсь з-над Йордану, і Дух на пустиню Його попровадив.
LUKE|4|2|Сорок день там диявол Його спокушав, і за тих днів Він нічого не їв, а коли закінчились вони, то вкінці зголоднів.
LUKE|4|3|І диявол до Нього сказав: Якщо Ти Син Божий, скажи цьому каменеві, щоб хлібом він став!
LUKE|4|4|А Ісус відповів йому: Написано: Не хлібом самим буде жити людина, але кожним Словом Божим!
LUKE|4|5|І він вивів Його на гору високу, і за хвилину часу показав Йому всі царства на світі.
LUKE|4|6|І диявол сказав Йому: Я дам Тобі всю оцю владу та їхню славу, бо мені це передане, і я даю, кому хочу, її.
LUKE|4|7|Тож коли Ти поклонишся передо мною, то все буде Твоє!
LUKE|4|8|І промовив Ісус йому в відповідь: Написано: Господеві Богові своєму вклоняйся, і служи Одному Йому!
LUKE|4|9|І повів Його в Єрусалим, і на наріжнику храму поставив, та й каже Йому: Як Ти Син Божий, кинься звідси додолу!
LUKE|4|10|Бо написано: Він накаже про Тебе Своїм Анголам, щоб Тебе берегли!
LUKE|4|11|і: Вони на руках понесуть Тебе, щоб коли не спіткнув Ти об камінь Своєї ноги!
LUKE|4|12|А Ісус відказав йому в відповідь: Сказано: Не спокушай Господа Бога свого!
LUKE|4|13|І диявол, скінчивши все цеє спокушування, відійшов від Нього до часу.
LUKE|4|14|А Ісус у силі Духа вернувся до Галілеї, і чутка про Нього рознеслась по всій тій країні.
LUKE|4|15|І Він їх навчав по їхніх синагогах, і всі Його славили.
LUKE|4|16|І прибув Він до Назарету, де був вихований. І звичаєм Своїм Він прийшов дня суботнього до синагоги, і встав, щоб читати.
LUKE|4|17|І подали Йому книгу пророка Ісаї. Розгорнувши ж Він книгу, знайшов місце, де було так написано:
LUKE|4|18|На Мені Дух Господній, бо Мене Він помазав, щоб Добру Новину звіщати вбогим. Послав Він Мене проповідувати полоненим визволення, а незрячим прозріння, відпустити на волю помучених,
LUKE|4|19|щоб проповідувати рік Господнього змилування.
LUKE|4|20|І, книгу згорнувши, віддав службі й сів. А очі всіх у синагозі звернулись на Нього.
LUKE|4|21|І почав Він до них говорити: Сьогодні збулося Писання, яке ви почули!
LUKE|4|22|І всі Йому стверджували й дивувались словам благодаті, що линули з уст Його. І казали вони: Чи ж то Він не син Йосипів?
LUKE|4|23|Він же промовив до них: Ви Мені конче скажете приказку: Лікарю, уздоров самого себе! Учини те й тут, у вітчизні Своїй, що сталося чули ми у Капернаумі.
LUKE|4|24|І сказав Він: Поправді кажу вам: Жаден пророк не буває приємний у вітчизні своїй.
LUKE|4|25|Та правдиво кажу вам: Багато вдовиць перебувало за днів Іллі серед Ізраїля, коли на три роки й шість місяців небо було зачинилося, так що голод великий настав був по всій тій землі,
LUKE|4|26|а Ілля не до жадної з них не був посланий, тільки в Сарепту Сидонську до овдовілої жінки.
LUKE|4|27|І багато було прокажених за Єлисея пророка в Ізраїлі, але жаден із них не очистився, крім Неємана сиріянина.
LUKE|4|28|І всі в синагозі, почувши оце, переповнились гнівом.
LUKE|4|29|І, вставши, вони Його вигнали за місто, і повели аж до краю гори, на якій їхнє місто було побудоване, щоб скинути додолу Його...
LUKE|4|30|Але Він перейшов серед них, і віддалився.
LUKE|4|31|І прийшов Він у Капернаум, галілейське місто, і там їх навчав по суботах.
LUKE|4|32|І дивувались науці Його, бо слово Його було владне.
LUKE|4|33|І був чоловік у синагозі, що мав духа нечистого демона, і він закричав гучним голосом:
LUKE|4|34|Ах, що нам до Тебе, Ісусе Назарянине? Ти прийшов погубити нас. Я знаю Тебе, хто Ти, Божий Святий...
LUKE|4|35|А Ісус заборонив йому, кажучи: Замовчи, і вийди з нього! І, кинувши демон того насередину, вийшов із нього, нічого йому не пошкодивши.
LUKE|4|36|І всіх жах обгорнув, і питали вони один одного, кажучи: Що то за наука, що духам нечистим наказує з владою й силою, і виходять вони?...
LUKE|4|37|І неслася чутка про Нього по всіх місцях краю.
LUKE|4|38|А як вийшов Він із синагоги, увійшов у дім Симона. Теща ж Симонова в великій гарячці лежала. І просили за неї Його.
LUKE|4|39|І, ставши над нею, Він заборонив тій гарячці, і вона полишила її. І, зараз уставши, теща їм прислуговувала.
LUKE|4|40|Коли ж сонце заходило, то всі, хто мав яких хворих на різні недуги, до Нього приводили їх. Він же клав Свої руки на кожного з них, та їх уздоровляв.
LUKE|4|41|Із багатьох же виходили й демони, кричачи та говорячи: Ти Син Божий! Та Він їм забороняв, і не давав говорити, що знали вони, що Христос Він.
LUKE|4|42|Коли ж настав день, Він вийшов, і подавсь до самотнього місця. А люди шукали Його. І прийшовши до Нього, Його затримували, щоб від них не відходив.
LUKE|4|43|Він же промовив до них: І іншим містам Я повинен звіщати Добру Новину про Боже Царство, бо на те Мене послано.
LUKE|4|44|І Він проповідував по синагогах Галілеї.
LUKE|5|1|І сталось, як тиснувся натовп до Нього, щоб почути Слово Боже, Він стояв біля озера Генісаретського.
LUKE|5|2|І Він побачив два човни, що стояли край озера. А рибалки, відійшовши від них, полоскали невода.
LUKE|5|3|І Він увійшов до одного з човнів, що був Симонів, і просив, щоб він трохи відплив від землі. І Він сів, та й навчав народ із човна.
LUKE|5|4|А коли перестав Він навчати, промовив до Симона: Попливи на глибінь, і закиньте на полов свій невід.
LUKE|5|5|А Симон сказав Йому в відповідь: Наставнику, цілу ніч ми працювали, і не вловили нічого, та за словом Твоїм укину невода.
LUKE|5|6|А зробивши оце, вони безліч риби набрали і їхній невід почав прориватись...
LUKE|5|7|І кивали вони до товаришів, що були в другім човні, щоб прийшли помогти їм. Ті прийшли, та й наповнили обидва човни, аж стали вони потопати.
LUKE|5|8|А як Симон Петро це побачив, то припав до колін Ісусових, кажучи: Господи, вийди від мене, бо я грішна людина!
LUKE|5|9|Бо від полову риби, що зловили вони, обгорнув жах його та й усіх, хто з ним був,
LUKE|5|10|також Якова й Івана, синів Зеведеєвих, що були спільниками Симона. І сказав Ісус Симонові: Не лякайсь, від цього часу ти будеш ловити людей!
LUKE|5|11|І вони повитягали на землю човни, покинули все, та й пішли вслід за Ним.
LUKE|5|12|А як Він перебував в одному з міст, ось один чоловік, увесь укритий проказою, Ісуса побачивши, упав ницьма, та й благав Його, кажучи: Господи, коли хочеш, Ти можеш очистити мене!
LUKE|5|13|А Він руку простяг, доторкнувся до нього й сказав: Хочу, будь чистий! І зараз із нього проказа зійшла...
LUKE|5|14|І звелів Він йому не казати нікому про це. Але йди, покажися священикові, і принеси за своє очищення, як Мойсей наказав, на свідчення їм.
LUKE|5|15|А чутка про Нього ще більше пішла, і багато народу приходило слухати та вздоровлятись від Нього з недугів своїх.
LUKE|5|16|Він же відходив на місце самотнє й молився.
LUKE|5|17|І сталось одного із днів, коли Він навчав, і сиділи фарисеї й законовчителі, що посходилися зо всіх сіл Галілеї й Юдеї та з Єрусалиму, а сила Господня готова була вздоровляти їх,
LUKE|5|18|і ось люди на ложі принесли чоловіка, що розслаблений був, і намагалися внести його, і перед Ним покласти.
LUKE|5|19|Не знайшовши ж кудою пронести його з-за народу, злізли на дім, і крізь стелю спустили із ложем його на середину перед Ісуса.
LUKE|5|20|І, побачивши їхню віру, сказав Він йому: Чоловіче, прощаються тобі гріхи твої!
LUKE|5|21|А книжники та фарисеї почали міркувати й казати: Хто ж Оцей, що богозневагу говорить? Хто може прощати гріхи, окрім Бога Самого?...
LUKE|5|22|Відчувши ж Ісус думки їхні, промовив у відповідь їм: Що міркуєте ви в серцях ваших?
LUKE|5|23|Що легше: сказати: Прощаються тобі гріхи твої, чи сказати: Уставай та й ходи?
LUKE|5|24|Але щоб ви знали, що Син Людський має владу на землі прощати гріхи, тож каже Він розслабленому: Кажу Я тобі: Уставай, візьми ложе своє, та й іди у свій дім!
LUKE|5|25|І той зараз устав перед ними, узявши те, на чому лежав, і пішов у свій дім, прославляючи Бога.
LUKE|5|26|І всіх жах обгорнув, і славили Бога вони. І переповнились страхом, говорячи: Дивні речі сьогодні ми бачили!...
LUKE|5|27|Після цього ж Він вийшов, і побачив митника, на ймення Левія, що сидів на митниці, та й промовив йому: Іди за Мною!
LUKE|5|28|І, покинувши все, той устав, і пішов услід за Ним.
LUKE|5|29|І справив Левій у своїм домі велику гостину для Нього. І був натовп великий митників й інших, що сиділи з Ним при столі.
LUKE|5|30|Фарисеї ж та книжники їхні нарікали на Нього, та учням Його говорили: Чому з митниками та із грішниками ви їсте та п'єте?
LUKE|5|31|А Ісус відповів і промовив до них: Лікаря не потребують здорові, а слабі.
LUKE|5|32|Не прийшов Я, щоб праведних кликати до покаяння, а грішних.
LUKE|5|33|Вони ж відказали до Нього: Чому учні Іванові часто постять та моляться, також і фарисейські, а Твої споживають та п'ють?
LUKE|5|34|Ісус же промовив до них: Чи ж ви можете змусити, щоб постили гості весільні, поки з ними ще є молодий?
LUKE|5|35|Але прийдуть ті дні, коли заберуть молодого від них, тоді й постити будуть тих днів...
LUKE|5|36|Розповів же і приказку їм: Ніхто латки з одежі нової в одежу стару не вставляє, а то подере й нову, а латка з нової старій не надасться.
LUKE|5|37|І ніхто не вливає вина молодого в старі бурдюки, а то попрориває вино молоде бурдюки, і вино розіллється, і бурдюки пропадуть.
LUKE|5|38|Але треба вливати вино молоде до нових бурдюків.
LUKE|5|39|І ніхто, старе пивши, молодого не схоче, бо каже: Старе ліпше!
LUKE|6|1|І сталось, як Він переходив ланами, у суботу, Його учні зривали колосся та їли, розтерши руками.
LUKE|6|2|А деякі з фарисеїв сказали: Нащо робите те, чого не годиться робити в суботу?
LUKE|6|3|І промовив Ісус їм у відповідь: Хіба ви не читали того, що зробив був Давид, коли сам зголоднів, також ті, хто був із ним?
LUKE|6|4|Як він увійшов був до Божого дому, і, взявши хліби показні, яких їсти не можна було, тільки самим священикам, споживав, і дав тим, хто був із ним?
LUKE|6|5|І сказав Він до них: Син Людський Господь і суботі!
LUKE|6|6|І сталось, як в іншу суботу зайшов Він до синагоги й навчав, знаходився там чоловік, що правиця йому була всохла.
LUKE|6|7|А книжники та фарисеї вважали, чи в суботу того не вздоровить, щоб знайти проти Нього оскарження.
LUKE|6|8|А Він знав думки їхні, і сказав чоловікові, що мав суху руку: Підведися, і стань посередині! Той підвівся і став.
LUKE|6|9|Ісус же промовив до них: Запитаю Я вас: Що годиться в суботу робити добре, чи робити лихе, душу спасти, чи згубити?
LUKE|6|10|І, позирнувши на всіх них, сказав чоловікові: Простягни свою руку! Той зробив, і рука його стала здорова!
LUKE|6|11|А вони переповнились лютістю, і один з одним змовлялись, що робити з Ісусом?...
LUKE|6|12|І сталось, що часу того Він вийшов на гору молитися, і перебув цілу ніч на молитві до Бога.
LUKE|6|13|А коли настав день, покликав Він учнів Своїх, і обрав із них Дванадцятьох, яких і апостолами Він назвав:
LUKE|6|14|Симона, якого й Петром Він назвав, і Андрія, брата його, Якова й Івана, Пилипа й Варфоломія,
LUKE|6|15|Матвія й Хому, Якова Алфієвого й Симона, званого Зилотом,
LUKE|6|16|Юду Якового, й Юду Іскаріотського, що й зрадником став.
LUKE|6|17|Як зійшов Він із ними, то спинився на рівному місці, також натовп густий Його учнів, і безліч людей з усієї Юдеї та з Єрусалиму, і з приморського Тиру й Сидону,
LUKE|6|18|що посходилися, щоб послухати Його та вздоровитися із недугів своїх, також ті, хто від духів нечистих страждав, і вони вздоровлялися.
LUKE|6|19|Увесь же народ намагався бодай доторкнутись до Нього, бо від Нього виходила сила, і всіх вздоровляла.
LUKE|6|20|А Він, звівши очі на учнів Своїх, говорив: Блаженні убогі, Царство Боже бо ваше.
LUKE|6|21|Блаженні голодні тепер, бо ви нагодовані будете. Блаженні засмучені зараз, бо втішитесь ви.
LUKE|6|22|Блаженні ви будете, коли люди зненавидять вас, і коли проженуть вас, і ганьбитимуть, і знеславлять, як зле, ім'я ваше за Людського Сина.
LUKE|6|23|Радійте того дня й веселіться, нагорода бо ваша велика на небесах. Бо так само чинили пророкам батьки їхні.
LUKE|6|24|Горе ж вам, багатіям, бо втіху свою ви вже маєте.
LUKE|6|25|Горе вам, тепер ситим, бо зазнаєте голоду ви. Горе вам, що тепер потішаєтеся, бо будете ви сумувати та плакати.
LUKE|6|26|Горе вам, як усі люди про вас говоритимуть добре, бо так само чинили фальшивим пророкам батьки їхні!
LUKE|6|27|А вам, хто слухає, Я кажу: Любіть своїх ворогів, добро робіть тим, хто ненавидить вас.
LUKE|6|28|Благословляйте тих, хто вас проклинає, і моліться за тих, хто кривду вам чинить.
LUKE|6|29|Хто вдарить тебе по щоці, підстав йому й другу, а хто хоче плаща твого взяти, не забороняй і сорочки.
LUKE|6|30|І кожному, хто в тебе просить подай, а від того, хто твоє забирає, назад не жадай.
LUKE|6|31|І як бажаєте, щоб вам люди чинили, так само чиніть їм і ви.
LUKE|6|32|А коли любите тих, хто любить вас, яка вам за те ласка? Люблять бо й грішники тих, хто їх любить.
LUKE|6|33|І коли добре чините тим, хто добро чинить вам, яка вам за те ласка? Бо те саме і грішники роблять.
LUKE|6|34|А коли позичаєте тим, що й від них сподіваєтесь взяти, яка вам за те ласка? Позичають бо й грішники грішникам, щоб одержати стільки ж.
LUKE|6|35|Тож любіть своїх ворогів, робіть добро, позичайте, не ждучи нічого назад, і ваша за це нагорода великою буде, і синами Всевишнього станете ви, добрий бо Він до невдячних і злих!
LUKE|6|36|Будьте ж милосердні, як і Отець ваш милосердний!
LUKE|6|37|Також не судіть, щоб не суджено й вас; і не осуджуйте, щоб і вас не осуджено; прощайте, то простять і вам.
LUKE|6|38|Давайте і дадуть вам; мірою доброю, натоптаною, струснутою й переповненою вам у подолок дадуть. Бо якою ви мірою міряєте, такою відміряють вам.
LUKE|6|39|Розповів також приказку їм: Чи ж може водити сліпого сліпий? Хіба не обидва в яму впадуть?
LUKE|6|40|Учень не більший за вчителя; але, удосконалившись, кожен буде, як учитель його.
LUKE|6|41|Чого ж в оці брата свого ти заскалку бачиш, колоди ж у власному оці не чуєш?
LUKE|6|42|Як ти можеш сказати до брата свого: Давай, брате, я заскалку вийму із ока твого, сам колоди, що в оці твоїм, не вбачаючи? Лицеміре, вийми перше колоду із власного ока, а потім побачиш, як вийняти заскалку з ока брата твого!
LUKE|6|43|Нема доброго дерева, що родило б злий плід, ані дерева злого, що родило б плід добрий.
LUKE|6|44|Кожне ж дерево з плоду свого пізнається. Не збирають бо фіґ із тернини, винограду ж на глоду не рвуть.
LUKE|6|45|Добра людина із доброї скарбниці серця добре виносить, а лиха із лихої виносить лихе. Бо чим серце наповнене, те говорять уста його!
LUKE|6|46|Що звете ви Мене: Господи, Господи, та не робите того, що Я говорю?
LUKE|6|47|Скажу вам, до кого подібний усякий, хто до Мене приходить та слів Моїх слухає, і виконує їх:
LUKE|6|48|Той подібний тому чоловікові, що, будуючи дім, він глибоко викопав, і основу на камінь поклав. Коли ж злива настала, вода кинулася на той дім, та однак не змогла захитати його, бо збудований добре він був!
LUKE|6|49|А хто слухає та не виконує, той подібний тому чоловікові, що свій дім збудував на землі без основи. І наперла на нього ріка, і зараз упав він, і велика була того дому руїна!
LUKE|7|1|А коли Він скінчив усі слова Свої до народу, що слухав Його, то ввійшов у Капернаум.
LUKE|7|2|У одного ж сотника тяжко раб занедужав, що був дорогий йому, і вмирати вже мав.
LUKE|7|3|А коли про Ісуса почув, то послав він до Нього юдейських старших, і благав Його, щоб прийшов, і вздоровив раба його.
LUKE|7|4|Вони ж прибули до Ісуса, та й ревно благали Його й говорили: Він достойний, щоб Ти це зробив йому.
LUKE|7|5|Бо він любить народ наш, та й для нас синагогу поставив.
LUKE|7|6|І пішов Ісус із ними. І коли недалеко від дому вже був, сотник друзів послав, щоб сказати Йому: Не турбуйся, о Господи, бо я недостойний, щоб зайшов Ти під стріху мою.
LUKE|7|7|Тому то й себе не вважав я за гідного, щоб до Тебе прийти. Та промов тільки слово, і раб мій одужає.
LUKE|7|8|Бо й я людина підвладна, і вояків під собою я маю; і одному кажу: піди, то йде він, а тому: прийди, і приходить, а своєму рабові: зроби теє і зробить.
LUKE|7|9|Почувши ж таке, Ісус здивувався йому, і, звернувшись до натовпу, що йшов слідком за Ним, промовив: Кажу вам: навіть серед Ізраїля Я не знайшов був такої великої віри!
LUKE|7|10|А коли посланці повернулись додому, то знайшли, що одужав той раб!
LUKE|7|11|І сталось, наступного дня Він відправивсь у місто, що зветься Наїн, а з Ним ішли учні Його та багато народу.
LUKE|7|12|І ось, як до брами міської наблизився Він, виносили вмерлого, одинака в своєї матері, що вдовою була. І з нею був натовп великий із міста.
LUKE|7|13|Як Господь же побачив її, то змилосердивсь над нею, і до неї промовив: Не плач!
LUKE|7|14|І Він підійшов, і доторкнувся до мар, носії ж зупинились. Тоді Він сказав: Юначе, кажу тобі: встань!
LUKE|7|15|І мертвий устав, і почав говорити. І його Він віддав його матері.
LUKE|7|16|А всіх острах пройняв, і Бога хвалили вони й говорили: Великий Пророк з'явився між нами, і зглянувся Бог над народом Своїм!
LUKE|7|17|І розійшлася ця чутка про Нього по цілій Юдеї, і по всій тій країні.
LUKE|7|18|Про все ж те сповістили Івана учні його. І покликав Іван двох із учнів своїх,
LUKE|7|19|і послав їх до Господа з запитом: Чи Ти Той, Хто має прийти, чи чекати нам Іншого?
LUKE|7|20|А мужі, прийшовши до Нього, сказали: Іван Христитель послав нас до Тебе, питаючи: Чи Ти Той, Хто має прийти, чи чекати нам Іншого?
LUKE|7|21|А саме тоді багатьох уздоровив був Він від недугів і мук, і від духів злих, і сліпим багатьом вернув зір.
LUKE|7|22|І промовив Ісус їм у відповідь: Ідіть, і перекажіть Іванові, що ви бачили й чули: Сліпі прозрівають, криві ходять, очищуються слабі на проказу, і чують глухі, воскресають померлі, убогим звіщається Добра Новина.
LUKE|7|23|І блаженний, хто через Мене спокуси не матиме!
LUKE|7|24|А коли відійшли посланці Іванові, Він почав говорити про Івана народові: На що ви дивитись ходили в пустиню? Чи на очерет, що вітер гойдає його?
LUKE|7|25|Та на що ви дивитись ходили? Може на чоловіка, у м'які шати одягненого? Аджеж ті, хто одягається славно, і розкішно живе, по палатах царських.
LUKE|7|26|На що ж ви ходили дивитись? На пророка? Так, кажу вам, навіть більше, аніж на пророка.
LUKE|7|27|Це той, що про нього написано: Ось перед обличчя Твоє посилаю Свого посланця, який перед Тобою дорогу Твою приготує!
LUKE|7|28|Кажу вам: Між народженими від жінок нема більшого понад Івана. Та найменший у Божому Царстві той більший за нього.
LUKE|7|29|І всі люди, що слухали, і митники визнали Божу волю за слушну, і охристились Івановим хрищенням.
LUKE|7|30|А фарисеї й законники відкинули Божу волю про себе, і не христились від нього.
LUKE|7|31|І промовив Господь: До кого ж уподоблю людей цього роду? І до кого подібні вони?
LUKE|7|32|Подібні вони до дітей, що на ринку сидять й один одного кличуть та кажуть: Ми вам грали були, а ви не танцювали, ми співали вам жалібно, та не плакали ви...
LUKE|7|33|Бо прийшов Іван Христитель, що хліба не їсть і вина не п'є, а ви кажете: Має він демона.
LUKE|7|34|Прийшов же Син Людський, що їсть і п'є, а ви кажете: Чоловік Цей ласун і п'яниця, Він приятель митників і грішників.
LUKE|7|35|І виправдалася мудрість усіма своїми ділами.
LUKE|7|36|А один із фарисеїв просив Його, щоб спожив Він із ним. І, прийшовши до дому того фарисея, Він сів при столі.
LUKE|7|37|І ось жінка одна, що була в місті, грішниця, як дізналась, що, Він у фарисеєвім домі засів при столі, алябастрову пляшечку мира принесла,
LUKE|7|38|і, припавши до ніг Його ззаду, плачучи, почала обливати слізьми Йому ноги, і волоссям своїм витирала, ноги Йому цілувала та миром мастила...
LUKE|7|39|Побачивши це, фарисей, що покликав Його, міркував собі, кажучи: Коли б був Він пророк, Він би знав, хто ото й яка жінка до Нього торкається, бож то грішниця!
LUKE|7|40|І озвався Ісус та й говорить до нього: Маю, Симоне, дещо сказати тобі. А той відказав: Кажи, Учителю.
LUKE|7|41|І промовив Ісус: Були два боржники в одного вірителя; один був винен п'ятсот динаріїв, а другий п'ятдесят.
LUKE|7|42|Як вони ж не могли заплатити, простив він обом. Скажи ж, котрий із них більше полюбить його?
LUKE|7|43|Відповів Симон, говорячи: Думаю, той, кому більше простив. І сказав Він йому: Розсудив ти правдиво.
LUKE|7|44|І, обернувшись до жінки, Він промовив до Симона: Чи ти бачиш цю жінку? Я прибув у твій дім, ти на ноги Мої не подав і води, а вона окропила слізьми Мої ноги й обтерла волоссям своїм.
LUKE|7|45|Поцілунку не дав ти Мені, а вона, відколи ввійшов Я, Мої ноги цілує невпинно.
LUKE|7|46|Голови ти Моєї оливою не намастив, а вона миром ноги мої намастила...
LUKE|7|47|Ось тому говорю Я тобі: Численні гріхи її прощені, бо багато вона полюбила. Кому ж мало прощається, такий мало любить.
LUKE|7|48|А до неї промовив: Прощаються тобі гріхи!
LUKE|7|49|А ті, що сиділи з Ним при столі, почали гомоніти про себе: Хто ж це Такий, що прощає й гріхи?
LUKE|7|50|А до жінки сказав Він: Твоя віра спасла тебе, іди з миром собі!
LUKE|8|1|І сталось, що Він після того проходив містами та селами, проповідуючи та звіщаючи Добру Новину про Боже Царство. Із ним Дванадцять були,
LUKE|8|2|та дехто з жінок, що були вздоровлені від злих духів і хвороб: Марія, Магдалиною звана, що з неї сім демонів вийшло,
LUKE|8|3|і Іванна, дружина Худзи, урядника Іродового, і Сусанна, і інших багато, що маєтком своїм їм служили.
LUKE|8|4|І, як зібралось багато народу, і з міста до Нього поприходили, то Він промовляти став притчею.
LUKE|8|5|Ось вийшов сіяч, щоб посіяти зерно своє. І, як сіяв, упало одне край дороги, і було повитоптуване, а птахи небесні його повидзьобували.
LUKE|8|6|Друге ж упало на ґрунт кам'янистий, і, зійшовши, усохло, не мало бо вогкости.
LUKE|8|7|А інше упало між терен, і вигнався терен, і його поглушив.
LUKE|8|8|Інше ж упало на добрую землю, і, зійшовши, уродило стокротно. Це сказавши, закликав: Хто має вуха, щоб слухати, нехай слухає!
LUKE|8|9|Запитали ж Його Його учні, говорячи: Що визначає ця притча?
LUKE|8|10|А Він відказав: Вам дано пізнати таємниці Божого Царства, а іншим у притчах, щоб дивились вони і не бачили, слухали і не розуміли.
LUKE|8|11|Ось що означає ця притча: Зерно це Боже Слово.
LUKE|8|12|А котрі край дороги, це ті, хто слухає, але потім приходить диявол, і забирає слово з їхнього серця, щоб не ввірували й не спаслися вони.
LUKE|8|13|А що на кам'янистому ґрунті, це ті, хто тільки почує, то слово приймає з радістю; та кореня не мають вони, вірують дочасно, і за час випробовування відпадають.
LUKE|8|14|А що впало між терен, це ті, хто слухає слово, але, ходячи, бувають придушені клопотами, та багатством, та життьовими розкошами, і плоду вони не дають.
LUKE|8|15|А те, що на добрій землі, це оті, хто як слово почує, береже його в щирому й доброму серці, і плід приносять вони в терпеливості.
LUKE|8|16|А світла засвіченого ніхто не покриває посудиною, і не ставить під ліжко, але ставить його на свічник, щоб бачили світло, хто входить.
LUKE|8|17|Немає нічого захованого, що не виявиться, ні таємного, що воно не пізнається, і не вийде наяв.
LUKE|8|18|Тож пильнуйте, як слухаєте! Бо хто має, то дасться йому, хто ж не має, забереться від нього і те, що, здається йому, ніби має.
LUKE|8|19|До Нього ж прийшли були мати й брати Його, та через народ не могли доступитись до Нього.
LUKE|8|20|І сповістили Йому: Твоя мати й брати Твої он стоять осторонь, і бажають побачити Тебе.
LUKE|8|21|А Він відповів і промовив до них: Моя мати й брати Мої це ті, хто слухає Боже Слово, і виконує!
LUKE|8|22|І сталось, одного з тих днів увійшов Він до човна, а з Ним Його учні. І сказав Він до них: Переплиньмо на другий бік озера. І відчалили.
LUKE|8|23|А коли вони плинули, Він заснув. І знялася на озері буря велика, аж вода заливати їх стала, і були в небезпеці вони.
LUKE|8|24|І вони підійшли, і розбудили Його та й сказали: Учителю, Учителю, гинемо! Він же встав, наказав бурі й хвилям, і вони вщухнули, і тиша настала!
LUKE|8|25|А до них Він сказав: Де ж ваша віра? І дивувались вони, перестрашені, і говорили один до одного: Хто ж це такий, що вітрам і воді Він наказує, а вони Його слухають?
LUKE|8|26|І вони припливли до землі Гадаринської, що навпроти Галілеї.
LUKE|8|27|І, як на землю Він вийшов, перестрів Його один чоловік із міста, що довгі роки мав він демонів, не вдягався в одежу, і мешкав не в домі, а в гробах.
LUKE|8|28|А коли він Ісуса побачив, то закричав, поваливсь перед Ним, і голосом гучним закликав: Що до мене Тобі, Ісусе, Сину Бога Всевишнього? Благаю Тебе, не муч мене!
LUKE|8|29|Бо звелів Він нечистому духові вийти з людини. Довгий час він хапав був його, і в'язали його ланцюгами й кайданами, і стерегли його, але він розривав ланцюги, і демон гнав по пустині його.
LUKE|8|30|А Ісус запитався його: Як тобі на ім'я? І той відказав: Леґіон, бо багато ввійшло в нього демонів.
LUKE|8|31|І благали Його, щоб Він їм не звелів іти в безодню.
LUKE|8|32|Пасся ж там на горі гурт великий свиней. І просилися демони ті, щоб дозволив піти їм у них. І дозволив Він їм.
LUKE|8|33|А як демони вийшли з того чоловіка, то в свиней увійшли. І череда кинулась із кручі до озера, і потопилась.
LUKE|8|34|Пастухи ж, як побачили теє, що сталось, повтікали, та в місті й по селах звістили.
LUKE|8|35|І вийшли побачити, що сталось. І прийшли до Ісуса й знайшли, що той чоловік, що демони вийшли із нього, сидів при ногах Ісусових вдягнений та при умі, і полякались...
LUKE|8|36|Самовидці ж їм розповіли, як видужав той біснуватий.
LUKE|8|37|І ввесь народ Гадаринського краю став благати Його, щоб пішов Він від них, великий бо страх обгорнув їх. Він же до човна ввійшов і вернувся.
LUKE|8|38|А той чоловік, що демони вийшли із нього, став благати Його, щоб бути при Ньому. Та Він відпустив його, кажучи:
LUKE|8|39|Вернися до дому свого, і розповіж, які речі великі вчинив тобі Бог! І той пішов, і по цілому місту звістив, які речі великі для нього Ісус учинив!
LUKE|8|40|А коли повернувся Ісус, то люди Його прийняли, бо всі чекали Його.
LUKE|8|41|Аж ось прийшов муж, Яір на ім'я, що був старшим синагоги. Він припав до Ісусових ніг, та й став благати Його завітати до дому його.
LUKE|8|42|Бо він мав одиначку дочку, років десь із дванадцять, і вмирала вона. А коли Він ішов, народ тиснув Його.
LUKE|8|43|А жінка одна, що дванадцять років хворою на кровотечу була, що ніхто вздоровити не міг її,
LUKE|8|44|підійшовши ззаду, доторкнулась до краю одежі Його, і хвилі тієї спинилася їй кровотеча!
LUKE|8|45|А Ісус запитав: Хто доторкнувся до Мене? Коли ж відмовлялися всі, то Петро відказав: Учителю, народ коло Тебе он товпиться й тисне.
LUKE|8|46|Ісус же промовив: Доторкнувсь хтось до Мене, бо Я відчув силу, що вийшла з Мене...
LUKE|8|47|А жінка, побачивши, що вона не втаїлась, трясучись, підійшла та й упала перед Ним, і призналася перед усіма людьми, чому доторкнулась до Нього, і як хвилі тієї одужала.
LUKE|8|48|Він же промовив до неї: Дочко, твоя віра спасла тебе; іди з миром собі!
LUKE|8|49|Як Він ще промовляв, приходить ось від старшини синагоги один та й говорить: Дочка твоя вмерла, не турбуй же Вчителя!
LUKE|8|50|Ісус же, почувши, йому відповів: Не лякайсь, тільки віруй, і буде спасена вона.
LUKE|8|51|Прийшовши ж до дому, не пустив Він нікого з Собою ввійти, крім Петра, та Івана, та Якова, та батька дівчати, та матері.
LUKE|8|52|А всі плакали та голосили за нею... Він же промовив: Не плачте, не вмерла вона, але спить!
LUKE|8|53|І насміхалися з Нього, бо знали, що вмерла вона.
LUKE|8|54|А Він узяв за руку її та й скрикнув, говорячи: Дівчатко, вставай!
LUKE|8|55|І вернувся їй дух, і хвилі тієї вона ожила... І звелів дать їй їсти.
LUKE|8|56|І здивувались батьки її. А Він наказав їм нікому не розповідати, що сталось.
LUKE|9|1|І скликав Він Дванадцятьох, і дав їм силу та владу над усіма демонами, і вздоровляти недуги.
LUKE|9|2|І послав їх проповідувати Царство Боже та вздоровляти недужих.
LUKE|9|3|І промовив до них: Не беріть нічого в дорогу: ані палиці, ані торби, ні хліба, ні срібла, ані майте по двоє убрань.
LUKE|9|4|І в який дім увійдете, зоставайтеся там, і звідти відходьте.
LUKE|9|5|А як хто вас не прийме, то, виходячи з міста того, обтрусіть від ніг ваших порох на свідчення супроти них.
LUKE|9|6|І вийшли вони, та й ходили по селах, звіщаючи Добру Новину та всюди вздоровляючи.
LUKE|9|7|А Ірод тетрарх прочув усе, що сталось було, і вагався, бо дехто казали, що Іван це із мертвих устав,
LUKE|9|8|а інші, що Ілля то з'явився, а знов інші, що ожив це один із стародавніх пророків.
LUKE|9|9|Тоді Ірод сказав: Іванові стяв я голову; хто ж Оцей, що я чую про Нього речі такі? І він намагався побачити Його.
LUKE|9|10|А коли повернулись апостоли, вони розповіли Йому, що зробили. І Він їх узяв, та й пішов самотою на місце безлюдне, біля міста, що зветься Віфсаіда.
LUKE|9|11|А як люди довідалися, то пішли вслід за Ним. І Він їх прийняв, і розповідав їм про Боже Царство, та тих уздоровляв, хто потребував уздоровлення.
LUKE|9|12|А день став схилятися. І Дванадцятеро підійшли та й сказали Йому: Відпусти вже людей, нехай вони йдуть у довколишні села й оселі спочити й здобути поживи, бо ми тут у місці безлюдному!
LUKE|9|13|А Він їм сказав: Дайте їсти їм ви. Вони ж відказали: Немає в нас більше, як п'ятеро хліба й дві рибі. Хіба підемо та купимо поживи для всього народу цього.
LUKE|9|14|Бо було чоловіків десь тисяч із п'ять. І сказав Він до учнів Своїх: Розсадіть їх рядами по п'ятидесяти.
LUKE|9|15|І зробили отак, і всіх їх розсадили.
LUKE|9|16|І Він узяв п'ять хлібів та дві рибі, споглянув на небо, поблагословив їх, і поламав, і дав учням, щоб клали народові.
LUKE|9|17|І всі їли й наситились! А з кусків позосталих зібрали дванадцять кошів...
LUKE|9|18|І сталось, як насамоті Він молився, з Ним учні були. І спитав Він їх, кажучи: За кого Мене люди вважають?
LUKE|9|19|Вони ж відповіли та сказали: За Івана Христителя, а ті за Іллю, а інші, що воскрес один із давніх пророків.
LUKE|9|20|А Він запитав їх: А ви за кого Мене маєте? Петро ж відповів та сказав: За Христа Божого!
LUKE|9|21|Він же їм заказав, і звелів не казати нікому про це.
LUKE|9|22|І сказав Він: Синові Людському треба багато страждати, і Його відцураються старші, і первосвященики, і книжники, і буде Він убитий, але третього дня Він воскресне!
LUKE|9|23|А до всіх Він промовив: Коли хоче хто йти вслід за Мною, хай зречеться самого себе, і хай візьме щоденно свого хреста, та й за Мною йде.
LUKE|9|24|Бо хто хоче душу свою зберегти, той погубить її, а хто ради Мене згубить душу свою, той її збереже.
LUKE|9|25|Яка ж користь людині, що здобуде ввесь світ, але занапастить чи згубить себе?
LUKE|9|26|Бо хто буде Мене та Моєї науки соромитися, того посоромиться також Син Людський, як прийде у славі Своїй, і Отчій, і святих Анголів.
LUKE|9|27|Правдиво ж кажу вам, що деякі з тут-о приявних не скуштують смерти, аж поки не побачать Царства Божого.
LUKE|9|28|І сталось після оцих слів днів за вісім, узяв Він Петра, і Івана, і Якова, та й пішов помолитись на гору.
LUKE|9|29|І коли Він молився, то вигляд лиця Його переобразився, а одежа Його стала біла й блискуча.
LUKE|9|30|І ось два мужі з Ним розмовляли, були то Мойсей та Ілля,
LUKE|9|31|що з'явилися в славі, і говорили про кінець Його, який в Єрусалимі Він мав докінчити.
LUKE|9|32|А Петро та приявні з ним були зморені сном, але, пробудившись, бачили славу Його й обох мужів, що стояли при Ньому.
LUKE|9|33|І сталось, як із Ним розлучались вони, то промовив Петро до Ісуса: Учителю, добре нам бути отут! Поставмо ж отут три шатрі: задля Тебе одне, і Мойсею одне, і одне для Іллі! Він не знав, що говорить...
LUKE|9|34|А як він говорив це, насунула хмара та їх заслонила. І вони полякались, як стали ті входити в хмару.
LUKE|9|35|І почувся ось голос із хмари, який промовляв: Це Син Мій Улюблений, Його слухайтеся!
LUKE|9|36|А коли оцей голос лунав, Ісус Сам позостався. А вони промовчали, і нікому нічого тих днів не казали, що бачили.
LUKE|9|37|А наступного дня, як спустились з гори, перестрів Його натовп великий.
LUKE|9|38|І закричав ось один чоловік із народу й сказав: Учителю, благаю Тебе, зглянься над сином моїм, бо одинак він у мене!
LUKE|9|39|А ото дух хапає його, і він нагло кричить, і трясе ним, аж той піну пускає. І, вимучивши він його, насилу відходить.
LUKE|9|40|І учнів Твоїх я благав його вигнати, та вони не змогли.
LUKE|9|41|А Ісус відповів і промовив: О, роде невірний й розбещений, доки буду Я з вами, і терпітиму вас? Приведи свого сина сюди!
LUKE|9|42|А як той іще йшов, демон кинув його та затряс. Та Ісус заказав тому духу нечистому, і вздоровив дитину, і віддав її батькові її.
LUKE|9|43|І всі дивувалися величі Божій! А як усі дивувались усьому, що чинив був Ісус, Він промовив до учнів Своїх:
LUKE|9|44|Вкладіть до вух своїх ці ось слова: Людський Син буде виданий людям до рук...
LUKE|9|45|Проте не зрозуміли вони цього слова, було бо закрите від них, щоб його не збагнули, та боялись Його запитати про це слово.
LUKE|9|46|І прийшло їм на думку: хто б найбільший з них був?
LUKE|9|47|А Ісус, думку серця їх знавши, узяв дитину, і поставив її біля Себе.
LUKE|9|48|І промовив до них: Як хто прийме дитину оцю в Ім'я Моє, Мене він приймає, а як хто Мене прийме, приймає Того, Хто послав Мене. Хто бо найменший між вами всіма, той великий!
LUKE|9|49|А Іван відповів і сказав: Учителю, ми бачили одного чоловіка, що Ім'ям Твоїм демонів виганяв, і ми заборонили йому, бо він з нами не ходить.
LUKE|9|50|Ісус же йому відказав: Не забороняйте, бо хто не проти вас, той за вас!
LUKE|9|51|І сталось, коли дні вознесення Його наближались, Він постановив піти в Єрусалим.
LUKE|9|52|І Він посланців вислав перед Собою. І пішли вони, та й прибули до села самарянського, щоб ночівлю Йому приготовити.
LUKE|9|53|А ті не прийняли Його, бо йшов Він у напрямі Єрусалиму.
LUKE|9|54|Як побачили ж те учні Яків й Іван, то сказали: Господи, хочеш, то ми скажемо, щоб огонь зійшов з неба та винищив їх, як і Ілля був зробив.
LUKE|9|55|А Він обернувся до них, їм докорив та й сказав: Ви не знаєте, якого ви духа.
LUKE|9|56|Бо Син Людський прийшов не губить душі людські, а спасати! І пішли вони в інше село.
LUKE|9|57|І сталось, як дорогою йшли, сказав був до Нього один: Я піду за Тобою, хоч би куди Ти пішов.
LUKE|9|58|Ісус же йому відказав: Мають нори лисиці, а гнізда небесні пташки, Син же Людський не має ніде й голови прихилити!
LUKE|9|59|І промовив до другого Він: Іди за Мною. А той відказав: Дозволь мені перше піти, і батька свого поховати.
LUKE|9|60|Він же йому відказав: Зостав мертвим ховати мерців своїх. А ти йди та звіщай Царство Боже.
LUKE|9|61|А інший сказав був: Господи, я піду за Тобою, та дозволь мені перш попрощатись із своїми домашніми.
LUKE|9|62|Ісус же промовив до нього: Ніхто з тих, хто кладе свою руку на плуга та назад озирається, не надається до Божого Царства!
LUKE|10|1|Після того призначив Господь і інших Сімдесят, і послав їх по двох перед Себе до кожного міста та місця, куди Сам мав іти.
LUKE|10|2|І промовив до них: Хоч жниво велике, та робітників мало; тож благайте Господаря жнива, щоб робітників вислав на жниво Своє.
LUKE|10|3|Ідіть! Оце посилаю Я вас, як ягнят між вовки.
LUKE|10|4|Не носіть ні калитки, ні торби, ні сандаль, і не вітайте в дорозі нікого.
LUKE|10|5|Як до дому ж якого ви ввійдете, то найперше кажіть: Мир дому цьому!
LUKE|10|6|І коли син миру там буде, то спочине на ньому ваш мир, коли ж ні до вас вернеться.
LUKE|10|7|Зоставайтеся ж у домі тім самім, споживайте та пийте, що є в них, бо вартий робітник своєї заплати. Не ходіть з дому в дім.
LUKE|10|8|А як прийдете в місто яке, і вас приймуть, споживайте, що вам подадуть.
LUKE|10|9|Уздоровлюйте хворих, що в нім, промовляйте до них: Наблизилося Царство Боже до вас!
LUKE|10|10|А як прийдете в місто яке, і вас не приймуть, то вийдіть на вулиці його та й кажіть:
LUKE|10|11|Ми обтрушуємо вам навіть порох, що прилип до нас із вашого міста. Та знайте оце, що наблизилося Царство Боже!
LUKE|10|12|Кажу вам: того дня легше буде содомлянам, аніж місту тому!
LUKE|10|13|Горе тобі, Хоразіне, горе тобі, Віфсаїдо! Бо коли б то у Тирі й Сидоні були відбулися ті чуда, що сталися в вас, то давно б вони покаялися в волосяниці та в попелі!
LUKE|10|14|Але на суді відрадніш буде Тиру й Сидону, як вам...
LUKE|10|15|А ти, Капернауме, що до неба піднісся, аж до аду ти зійдеш!
LUKE|10|16|Хто слухає вас Мене слухає, хто ж погорджує вами погорджує Мною, хто ж погорджує Мною погорджує Тим, Хто послав Мене.
LUKE|10|17|А ті Сімдесят повернулися з радістю, кажучи: Господи, навіть демони коряться нам у Ім'я Твоє!
LUKE|10|18|Він же промовив до них: Я бачив того сатану, що з неба спадав, немов блискавка.
LUKE|10|19|Ось Я владу вам дав наступати на змій та скорпіонів, і на всю силу ворожу, і ніщо вам не зашкодить.
LUKE|10|20|Та не тіштеся тим, що вам коряться духи, але тіштесь, що ваші ймення записані в небі!
LUKE|10|21|Того часу Ісус звеселився був Духом Святим і промовив: Прославляю Тебе, Отче, Господи неба й землі, що втаїв Ти оце від премудрих і розумних, та його немовлятам відкрив. Так, Отче, бо Тобі так було до вподоби!
LUKE|10|22|Передав Мені все Мій Отець. І не знає ніхто, хто є Син, тільки Отець, і хто Отець тільки Син, та кому Син захоче відкрити.
LUKE|10|23|І, звернувшись до учнів, наодинці їм сказав: Блаженні ті очі, що бачать, що бачите ви!
LUKE|10|24|Кажу ж вам, що багато пророків і царів бажали побачити, що бачите ви та й не бачили, і почути, що чуєте ви і не чули!
LUKE|10|25|І підвівсь ось законник один, і сказав, Його випробовуючи: Учителю, що робити мені, щоб вічне життя осягнути?
LUKE|10|26|Він же йому відказав: Що в Законі написано, як ти читаєш?
LUKE|10|27|А той відповів і сказав: Люби Господа Бога свого всім серцем своїм, і всією душею своєю, і всією силою своєю, і всім своїм розумом, і свого ближнього, як самого себе.
LUKE|10|28|Він же йому відказав: Правильно ти відповів. Роби це, і будеш жити.
LUKE|10|29|А той бажав сам себе виправдати, та й сказав до Ісуса: А хто то мій ближній?
LUKE|10|30|А Ісус відповів і промовив: Один чоловік ішов з Єрусалиму до Єрихону, і попався розбійникам, що обдерли його, і завдали йому рани, та й утекли, покинувши ледве живого його.
LUKE|10|31|Проходив випадком тією дорогою священик один, побачив його, і проминув.
LUKE|10|32|Так само й Левит надійшов на те місце, поглянув, і теж проминув.
LUKE|10|33|Проходив же там якийсь самарянин, та й натрапив на нього, і, побачивши, змилосердився.
LUKE|10|34|І він підійшов, і обв'язав йому рани, наливши оливи й вина. Потому його посадив на худобину власну, і приставив його до гостиниці, та й клопотався про нього.
LUKE|10|35|А другого дня, від'їжджавши, вийняв він два динарії, та й дав їх господареві й проказав: Заопікуйся ним, а як більше що витратиш, заплачу тобі, як вернуся.
LUKE|10|36|Котрий же з цих трьох на думку твою був ближній тому, хто попався розбійникам?
LUKE|10|37|А він відказав: Той, хто вчинив йому милість. Ісус же сказав йому: Іди, і роби так і ти!
LUKE|10|38|І сталось, коли вони йшли, Він прийшов до одного села. Одна ж жінка, Марта їй на ім'я, прийняла Його в дім свій.
LUKE|10|39|Була ж в неї сестра, що звалась Марія; вона сіла в ногах у Ісуса, та й слухала слова Його.
LUKE|10|40|А Марта великою послугою клопоталась, а спинившись, сказала: Господи, чи байдуже Тобі, що на мене саму полишила служити сестра моя? Скажи ж їй, щоб мені помогла.
LUKE|10|41|Господь же промовив у відповідь їй: Марто, Марто, турбуєшся й журишся ти про багато чого,
LUKE|10|42|а потрібне одне. Марія ж обрала найкращу частку, яка не відбереться від неї...
LUKE|11|1|І сталось, як молився Він у місці одному, і коли перестав, озвався до Нього один із Його учнів: Господи, навчи нас молитися, як і Іван навчив своїх учнів.
LUKE|11|2|Він же промовив до них: Коли молитеся, говоріть: Отче наш, що єси на небесах! Нехай святиться Ім'я Твоє, нехай прийде Царство Твоє, нехай буде воля Твоя, як на небі, так і на землі.
LUKE|11|3|Хліба нашого насущного дай нам на кожний день.
LUKE|11|4|І прости нам наші гріхи, бо й самі ми прощаємо кожному боржникові нашому. І не введи нас у випробовування, але визволи нас від лукавого!
LUKE|11|5|І сказав Він до них: Хто з вас матиме приятеля, і піде до нього опівночі, і скаже йому: Позич мені, друже, три хліби,
LUKE|11|6|бо прийшов із дороги до мене мій приятель, я ж не маю, що дати йому.
LUKE|11|7|А той із середини в відповідь скаже: Не роби мені клопоту, уже замкнені двері, і мої діти зо мною на ліжкові. Не можу я встати та дати тобі.
LUKE|11|8|Кажу вам: коли він не встане, і не дасть ради дружби йому, то за докучання його він устане та й дасть йому, скільки той потребує.
LUKE|11|9|І Я вам кажу: просіть, і буде вам дано, шукайте і знайдете, стукайте і відчинять вам!
LUKE|11|10|Бо кожен, хто просить одержує, хто шукає знаходить, а тому, хто стукає відчинять.
LUKE|11|11|І котрий з вас, батьків, як син хліба проситиме, подасть йому каменя? Або, як проситиме риби, замість риби подасть йому гадину?
LUKE|11|12|Або, як яйця він проситиме, дасть йому скорпіона?
LUKE|11|13|Отож, коли ви, бувши злі, потрапите добрі дари своїм дітям давати, скільки ж більше Небесний Отець подасть Духа Святого всім тим, хто проситиме в Нього?
LUKE|11|14|Раз вигонив Він демона, який був німий. І коли демон вийшов, німий заговорив. А народ дивувався.
LUKE|11|15|А деякі з них гомоніли: Виганяє Він демонів силою Вельзевула, князя демонів...
LUKE|11|16|А інші, випробовуючи, хотіли від Нього ознаки із неба.
LUKE|11|17|Він же знав думки їхні, і промовив до них: Кожне царство, само проти себе поділене, запустіє, і дім на дім упаде.
LUKE|11|18|А коли й сатана поділився сам супроти себе, як стоятиме царство його? А ви кажете, що Вельзевулом вигоню Я демонів.
LUKE|11|19|Коли ж Вельзевулом вигоню Я демонів, то чим виганяють їх ваші сини? Тому вони стануть вам суддями.
LUKE|11|20|А коли перстом Божим вигоню Я демонів, то справді прийшло до вас Боже Царство.
LUKE|11|21|Коли сильний збройно свій двір стереже, то в безпеці маєток його.
LUKE|11|22|Коли ж дужчий від нього його нападе й переможе, то всю зброю йому забере, на яку покладався був той, і роздасть свою здобич.
LUKE|11|23|Хто не зо Мною, той проти Мене; і хто не збирає зо Мною, той розкидає!
LUKE|11|24|Коли дух нечистий виходить з людини, то блукає місцями безвідними, відпочинку шукаючи, але, не знаходячи, каже: Вернуся до хати своєї, звідки я вийшов.
LUKE|11|25|А як вернеться він, то хату знаходить заметену й прибрану.
LUKE|11|26|Тоді він іде та й приводить сімох інших духів, лютіших за себе, і входять вони та й живуть там. І буде останнє людині тій гірше за перше!
LUKE|11|27|І сталось, як Він це говорив, одна жінка з народу свій голос піднесла й сказала до Нього: Блаженна утроба, що носила Тебе, і груди, що Ти ссав їх!
LUKE|11|28|А Він відказав: Так. Блаженні ж і ті, хто слухає Божого Слова і його береже!
LUKE|11|29|А як люди збиралися, Він почав промовляти: Рід цей рід лукавий: він ознаки шукає, та ознаки йому не дадуть, крім ознаки пророка Йони.
LUKE|11|30|Бо як Йона ознакою був для ніневітян, так буде й Син Людський для роду цього.
LUKE|11|31|Цариця південна на суд стане з мужами роду цього, і їх засудить, бо вона з кінця світу прийшла Соломонову мудрість послухати. А тут ось Хтось більший, аніж Соломон!
LUKE|11|32|Ніневітяни стануть на суд із цим родом, і засудять його, вони бо покаялися через Йонину проповідь. А тут ось Хтось більший, ніж Йона!
LUKE|11|33|Засвіченого світильника ніхто в сховок не ставить, ані під посудину, але на свічник, щоб бачили світло, хто входить.
LUKE|11|34|Око твоє то світильник для тіла; тому, як око твоє буде дуже, то й усе тіло твоє буде світле. А коли б твоє око нездатне було, то й усе тіло твоє буде темне.
LUKE|11|35|Отож, уважай, щоб те світло, що в тобі, не сталося темрявою!
LUKE|11|36|Бо коли твоє тіло все світле, і не має жадної темної частини, то все буде світле, неначе б світильник осяяв блиском тебе.
LUKE|11|37|Коли Він говорив, то один фарисей став благати Його пообідати в нього. Він же прийшов та й сів при столі.
LUKE|11|38|Фарисей же, побачивши це, здивувався, що перед обідом Він перш не обмився.
LUKE|11|39|Господь же промовив до нього: Тепер ви, фарисеї, он чистите зовнішність кухля та миски, а ваше нутро повне здирства та кривди!
LUKE|11|40|Нерозумні, чи ж Той, Хто створив оте зовнішнє, не створив Він і внутрішнє?
LUKE|11|41|Тож милостиню подавайте з унутрішнього, і ось все буде вам чисте.
LUKE|11|42|Горе вам, фарисеям, бо ви десятину даєте з м'яти та рути й усякого зілля, але обминаєте суд та Божу любов; це треба робити, і того не лишати!
LUKE|11|43|Горе вам, фарисеям, що любите перші лавки в синагогах та привіти на ринках!
LUKE|11|44|Горе вам, бо ви як гроби непомітні, люди ж ходять по них і не знають того...
LUKE|11|45|Озвався ж один із законників, і каже Йому: Учителю, кажучи це, Ти і нас ображаєш!
LUKE|11|46|А Він відказав: Горе й вам, законникам, бо ви на людей тягарі накладаєте, які важко носити, а самі й одним пальцем своїм не доторкуєтесь тягарів!
LUKE|11|47|Горе вам, бо надгробки пророкам ви ставите, ваші ж батьки були їх повбивали...
LUKE|11|48|Так, визнаєте ви й хвалите вчинки батьків своїх: бо вони їх повбивали, а ви їм надгробки будуєте!
LUKE|11|49|Через те й мудрість Божа сказала: Я пошлю їм пророків й апостолів, вони ж декого з них повбивають, а декого виженуть,
LUKE|11|50|щоб на роді оцім відомстилася кров усіх пророків, що пролита від створення світу,
LUKE|11|51|від крови Авеля аж до крови Захарія, що загинув між жертівником і храмом! Так, кажу вам, відомститься це все на цім роді!
LUKE|11|52|Горе вам, законникам, бо взяли ви ключа розуміння: самі не ввійшли, і тим, хто хотів увійти, боронили!
LUKE|11|53|А коли Він виходив ізвідти, стали книжники та фарисеї сильно тиснути та від Нього допитуватись про багато речей,
LUKE|11|54|вони чатували на Нього, щоб зловити що з уст Його (і щоб оскаржити Його).
LUKE|12|1|Того часу, як зібралися десятитисячні натовпи народу, аж топтали вони один одного, Він почав промовляти перш до учнів Своїх: Стережіться розчини фарисейської, що є лицемірство!
LUKE|12|2|Бо немає нічого захованого, що не відкриється, ні таємного, що не виявиться.
LUKE|12|3|Тому все, що казали ви потемки, при світлі почується, що ж шептали на вухо в коморах, на дахах проповідане буде.
LUKE|12|4|Кажу ж вам, Своїм друзям: Не бійтеся тих, хто тіло вбиває, а потім більш нічого не може вчинити!
LUKE|12|5|Але вкажу вам, кого треба боятися: Бійтесь того, хто має владу, убивши, укинути в геєнну. Так, кажу вам: Того бійтеся!
LUKE|12|6|Чи ж не п'ять горобців продають за два гроші? Та проте перед Богом із них ні один не забутий.
LUKE|12|7|Але навіть волосся вам на голові пораховане все. Не бійтесь: вартніші ви за багатьох горобців!
LUKE|12|8|Кажу ж вам: Кожного, хто перед людьми Мене визнає, того визнає й Син Людський перед Анголами Божими.
LUKE|12|9|Хто ж Мене відцурається перед людьми, того відцураються перед Анголами Божими.
LUKE|12|10|І кожному, хто скаже слово на Людського Сина, йому проститься; а хто зневажатиме Духа Святого, не проститься.
LUKE|12|11|А коли вас водитимуть до синагог, і до урядів, і до влад, не турбуйтеся, як або що відповідати чи що говорити,
LUKE|12|12|Дух бо Святий вас навчить тієї години, що потрібно казати!
LUKE|12|13|І озвався до Нього один із народу: Учителю, скажи братові моєму, щоб він спадщиною поділився зо мною.
LUKE|12|14|А Він відказав йому: Чоловіче, хто поставив над вами Мене за суддю або за подільника?
LUKE|12|15|І промовив до них: Глядіть, остерігайтеся всякої зажерливости, бо життя чоловіка не залежить від достатку маєтку його.
LUKE|12|16|І Він розповів їм притчу, говорячи: В одного багача гойно нива вродила була.
LUKE|12|17|І міркував він про себе й казав: Що робити, що не маю куди зібрати плодів своїх?
LUKE|12|18|І сказав: Оце я зроблю, порозвалюю клуні свої, і просторніші поставлю, і позбираю туди пашню свою всю та свій достаток.
LUKE|12|19|І скажу я душі своїй: Душе, маєш багато добра, на багато років складеного. Спочивай, їж та пий, і веселися!
LUKE|12|20|Бог же до нього прорік: Нерозумний, ночі цієї ось душу твою зажадають від тебе, і кому позостанеться те, що ти був наготовив?...
LUKE|12|21|Так буває і з тим, хто збирає для себе, та не багатіє в Бога.
LUKE|12|22|І промовив Він учням Своїм: Через це кажу вам: Не журіться про життя, що ви будете їсти, і ні про тіло, у що ви зодягнетеся.
LUKE|12|23|Бо більше від їжі життя, а тіло від одягу.
LUKE|12|24|Погляньте на гайвороння, що не сіють, не жнуть, нема в них комори, ні клуні, проте Бог їх годує. Скільки ж більше за птахів ви варті!
LUKE|12|25|Хто ж із вас, коли журиться, добавити зможе до зросту свого бодай ліктя одного?
LUKE|12|26|Тож коли ви й найменшого не подолаєте, то чого ж ви про інше клопочетеся?
LUKE|12|27|Погляньте на ті он лілеї, як вони не прядуть, ані тчуть. Але говорю вам, що й сам Соломон у всій славі своїй не вдягався отак, як одна з них!
LUKE|12|28|І коли он траву, що сьогодні на полі, а взавтра до печі вкидається, Бог так зодягає, скільки ж краще зодягне Він вас, маловірні!
LUKE|12|29|І не шукайте, що будете їсти, чи що будете пити, і не клопочіться.
LUKE|12|30|Бо всього цього й люди світу оцього шукають, Отець же ваш знає, що того вам потрібно.
LUKE|12|31|Шукайте отож Його Царства, а це вам додасться!
LUKE|12|32|Не лякайся, черідко мала, бо сподобалося Отцю вашому дати вам Царство.
LUKE|12|33|Продавайте достатки свої та милостиню подавайте. Робіть калитки собі не старіючі, невичерпний скарб той у небі, куди не закрадається злодій, і міль де не точить.
LUKE|12|34|Бо де скарб ваш, там буде й серце ваше!
LUKE|12|35|Нехай підперезані будуть вам стегна, а світла ручні позасвічувані!
LUKE|12|36|І будьте подібними до людей, що очікують пана свого, коли вернеться він із весілля, щоб, як прийде й застукає, відчинити негайно йому.
LUKE|12|37|Блаженні раби ті, що пан, коли прийде, то знайде, що пильнують вони! Поправді кажу вам: підпережеться він і їх посадовить, і, підійшовши, буде їм послуговувати.
LUKE|12|38|І коли прийде о другій чи прийде о третій сторожі, та знайде так само, блаженні вони!
LUKE|12|39|Знайте ж це, що коли б знав господар, о котрій то годині підкрадеться злодій, то він пильнував би, і свого б дому не дав підкопати.
LUKE|12|40|Тому будьте готові і ви, бо прийде Син Людський тієї години, коли ви не думаєте!
LUKE|12|41|Озвався ж Петро: Господи, чи до нас кажеш притчу оцю, чи до всіх?
LUKE|12|42|А Господь відказав: Хто ж тоді вірний і мудрий домоправитель, що пан настановить його над своїми челядниками, щоб давати харч визначену своєчасно?
LUKE|12|43|Блаженний той раб, що пан його прийде та знайде, що робить він так!
LUKE|12|44|Поправді кажу вам, що над всім маєтком своїм він поставить його.
LUKE|12|45|А коли раб той скаже у серці своїм: Забариться пан мій прийти, і зачне бити слуг та служниць, їсти та пити та напиватися,
LUKE|12|46|то прийде раба того пан за дня, якого він не сподівається, і о годині, якої не знає, і розітне його пополовині, і визначить долю йому з невірними!
LUKE|12|47|А раб той, що знав волю свого господаря, але не приготував, ані не вчинив згідно волі його, буде тяжко побитий.
LUKE|12|48|Хто ж не знав, а вчинив каригідне, буде мало він битий. Тож від кожного, кому дано багато, багато від нього й жадатимуть. А кому багато повірено, від того ще більше жадатимуть.
LUKE|12|49|Я прийшов огонь кинути на землю, і як Я прагну, щоб він уже запалав!
LUKE|12|50|Я ж маю христитися хрищенням, і як Я мучуся, поки те сповниться!
LUKE|12|51|Чи ви думаєте, що прийшов Я мир дати на землю? Ні, кажу вам, але поділ!
LUKE|12|52|Віднині бо п'ятеро в домі одному поділені будуть: троє супроти двох, і двоє супроти трьох.
LUKE|12|53|Стане батько на сина, а син проти батька, мати проти дочки, а дочка проти матері, свекруха навпроти невістки своєї, а невістка навпроти свекрухи!...
LUKE|12|54|Промовив же Він і до народу: Як побачите хмару, що з заходу суне, то кажете зараз: Зближається дощ, і так і буває.
LUKE|12|55|А коли віє вітер південний, то кажете: Буде спекота, і буває.
LUKE|12|56|Лицеміри, лице неба й землі розпізнати ви вмієте, чому ж не розпізнаєте часу цього?
LUKE|12|57|Чого ж і самі по собі ви не судите, що справедливе?
LUKE|12|58|Бо коли до уряду ти йдеш зо своїм супротивником, попильнуй з ним залагодити по дорозі, щоб тебе до судді не потяг він, а суддя щоб прислужникові не віддав тебе, а прислужник щоб не посадив до в'язниці тебе.
LUKE|12|59|Поправді кажу тобі: Не вийдеш ізвідти, поки не віддаси й останнього шеляга!
LUKE|13|1|Того часу прийшли були дехто, та й розповіли Йому про галілеян, що їхню кров Пилат змішав був із їхніми жертвами.
LUKE|13|2|Ісус же сказав їм у відповідь: Чи ви думаєте, що оці галілеяни, що так постраждали, грішніші були від усіх галілеян?
LUKE|13|3|Ні, кажу вам; та коли не покаєтеся, то загинете всі так!
LUKE|13|4|Або ті вісімнадцять, що башта на них завалилась була в Сілоамі й побила їх, чи думаєте, що ті винні були більш за всіх, що в Єрусалимі живуть?
LUKE|13|5|Ні, кажу вам; та коли не покаєтеся, то загинете всі так!
LUKE|13|6|І Він розповів оцю притчу: Один чоловік у своїм винограднику мав посаджене фіґове дерево. І прийшов він шукати на ньому плоду, але не знайшов.
LUKE|13|7|І сказав винареві: Оце третій рік, відколи приходжу шукати плоду на цім фіґовім дереві, але не знаходжу; зрубай його, нащо й землю марнує воно?
LUKE|13|8|А той йому в відповідь каже: Позостав його, пане, і на цей рік, аж поки його обкопаю довкола, і обкладу його гноєм,
LUKE|13|9|чи року наступного плоду не вродить воно. Коли ж ні, то зрубаєш його.
LUKE|13|10|І навчав Він в одній з синагог у суботу.
LUKE|13|11|І ось там була одна жінка, що вісімнадцять років мала духа немочі, і була скорчена, і не могла ніяк випростатись.
LUKE|13|12|А Ісус, як побачив її, то покликав до Себе. І сказав їй: Жінко, звільнена ти від недуги своєї.
LUKE|13|13|І Він руки на неї поклав, і вона зараз випросталась, і стала славити Бога!
LUKE|13|14|Озвався ж старший синагоги, обурений, що Ісус уздоровив у суботу, і сказав до народу: Є шість день, коли працювати належить, приходьте тоді та вздоровлюйтеся, а не дня суботнього.
LUKE|13|15|А Господь відповів і промовив до нього: Лицеміре, хіба ж не відв'язує кожен із вас у суботу свого вола чи осла від ясел, і не веде напоїти?
LUKE|13|16|Чи ж цю дочку Авраамову, яку сатана був зв'язав вісімнадцять ось років, не належить звільнити її суботнього дня від цих пут?
LUKE|13|17|А як Він говорив це, засоромилися всі Його супротивники. І тішився ввесь народ всіма славними вчинками, які Він чинив!
LUKE|13|18|Він же промовив: До чого подібне Царство Боже, і до чого його прирівняю?
LUKE|13|19|Подібне воно до гірчичного зерна, що взяв чоловік і посіяв його в своїм саді. І воно виросло, і деревом стало, і кублилось птаство небесне на віттях його.
LUKE|13|20|І знову сказав Він: Із чим порівняю Я Божеє Царство?
LUKE|13|21|Подібне до розчини, що її бере жінка, і кладе на три мірки муки, аж поки все вкисне.
LUKE|13|22|І проходив містами та селами Він і навчав, до Єрусалиму простуючи.
LUKE|13|23|І озвався до Нього один: Господи, хіба буде мало спасених? А Він відказав їм:
LUKE|13|24|Силкуйтеся ввійти тісними ворітьми, бо кажу вам, багато-хто будуть намагатися ввійти, та не зможуть!
LUKE|13|25|Як устане Господар та двері замкне, ви зачнете вистоювати ізнадвору, та стукати в двері й казати: Господи, відчини нам! А Він вам у відповідь скаже: Не знаю Я вас, звідки ви!
LUKE|13|26|Тоді станете ви говорити: Ми їли й пили перед Тобою і на вулицях наших навчав Ти...
LUKE|13|27|А Він вам відкаже: Говорю вам, не знаю Я, звідки ви. Відійдіть від Мене всі, хто чинить неправду!
LUKE|13|28|Буде плач там і скрегіт зубів, як побачите ви Авраама, та Ісака та Якова, та пророків усіх в Царстві Божім, себе ж вигнаних геть...
LUKE|13|29|І прийдуть інші від сходу й заходу, і півночі й півдня, і при столі в Царстві Божім засядуть!
LUKE|13|30|І ось, є останні, що стануть за перших, і є перші, що стануть останніми!
LUKE|13|31|Тієї години підійшли дехто з фарисеїв, і сказали Йому: Вийди собі, і піди звідси, хоче бо Ірод убити Тебе...
LUKE|13|32|А Він відказав їм: Ідіть і скажіть тому лисові: Ось демонів Я виганяю, і чиню вздоровлення, сьогодні та взавтра, а третього дня закінчу.
LUKE|13|33|Однак, Мені треба ходити сьогодні та взавтра, і часу найближчого, бо згинути не може пророк поза Єрусалимом.
LUKE|13|34|Єрусалиме, Єрусалиме, що вбиваєш пророків та каменуєш посланих до тебе! Скільки раз Я хотів позбирати дітей твоїх, як та квочка збирає під крила курчаток своїх, та ви не захотіли!
LUKE|13|35|Ось ваш дім зостається порожній для вас! Говорю бо Я вам: Ви мене не побачите, аж поки не настане, що скажете: Благословенний, Хто йде в Господнє Ім'я!
LUKE|14|1|І сталось, що Він у суботу ввійшов був до дому одного з фарисейських старшин, щоб хліба спожити, а вони назирали за Ним.
LUKE|14|2|І ото перед Ним був один чоловік, слабий на водянку.
LUKE|14|3|Ісус же озвався й сказав до законників та фарисеїв: Чи вздоровляти в суботу годиться чи ні?
LUKE|14|4|Вони ж мовчали. А Він, доторкнувшись, уздоровив його та відпустив...
LUKE|14|5|І сказав Він до них: Коли осел або віл котрогось із вас упаде до криниці, то хіба він не витягне зараз його дня суботнього?
LUKE|14|6|І вони не могли відповісти на це.
LUKE|14|7|А як Він спостеріг, як вони собі перші місця вибирали, то сказав до запрошених притчу:
LUKE|14|8|Коли хто покличе тебе на весілля, не сідай на першому місці, щоб не трапився хто поважніший за тебе з покликаних,
LUKE|14|9|і щоб той, хто покликав тебе та його, не прийшов і тобі не сказав: Поступися цьому місцем! І тоді ти із соромом станеш займати місце останнє...
LUKE|14|10|Але як ти будеш запрошений, то приходь, і сідай на останньому місці, щоб той, хто покликав тебе, підійшов і сказав тобі: Приятелю, сідай вище! Тоді буде честь тобі перед покликаними з тобою.
LUKE|14|11|Хто бо підноситься буде впокорений, а хто впокоряється той піднесеться.
LUKE|14|12|А тому, хто Його був покликав, сказав Він: Коли ти справляєш обід чи вечерю, не клич друзів своїх, ні братів своїх, ані своїх родичів, ні сусідів багатих, щоб так само й вони коли не запросили тебе, і буде взаємна відплата тобі.
LUKE|14|13|Але, як справляєш гостину, клич убогих, калік, кривих та сліпих,
LUKE|14|14|і будеш блаженний, бо не мають вони чим віддати тобі, віддасться ж тобі за воскресіння праведних!
LUKE|14|15|Як почув це один із отих, що сиділи з Ним при столі, то до Нього сказав: Блаженний, хто хліб споживатиме в Божому Царстві!
LUKE|14|16|Він же промовив до нього: Один чоловік спорядив був велику вечерю, і запросив багатьох.
LUKE|14|17|І послав він свого раба часу вечері сказати запрошеним: Ідіть, бо вже все наготовано.
LUKE|14|18|І зараз усі почали відмовлятися. Перший сказав йому: Поле купив я, і маю потребу піти та оглянути його. Прошу тебе, вибач мені!
LUKE|14|19|А другий сказав: Я купив собі п'ять пар волів, і йду спробувати їх. Прошу тебе, вибач мені!
LUKE|14|20|І знов інший сказав: Одружився ось я, і через те я не можу прибути.
LUKE|14|21|І вернувся той раб і панові своєму про все розповів. Розгнівавсь господар тоді, та й сказав до свого раба: Піди швидко на вулиці та на завулки міські, і приведи сюди вбогих, і калік, і сліпих, і кривих.
LUKE|14|22|І згодом раб повідомив: Пане, сталося так, як звелів ти, та місця є ще.
LUKE|14|23|І сказав пан рабові: Піди на дороги й на загороди, та й силуй прийти, щоб наповнився дім мій.
LUKE|14|24|Кажу бо я вам, що жаден із запрошених мужів тих не покуштує моєї вечері... Бо багато покликаних, та вибраних мало!
LUKE|14|25|Ішло ж з Ним багато людей. І, звернувшись, сказав Він до них:
LUKE|14|26|Коли хто приходить до Мене, і не зненавидить свого батька та матері, і дружини й дітей, і братів і сестер, а до того й своєї душі, той не може буть учнем Моїм!
LUKE|14|27|І хто свого хреста не несе, і не йде вслід за Мною, той не може бути учнем Моїм!
LUKE|14|28|Хто бо з вас, коли башту поставити хоче, перше не сяде й видатків не вирахує, чи має потрібне на виконання,
LUKE|14|29|щоб, коли покладе він основу, але докінчити не зможе, усі, хто побачить, не стали б сміятися з нього,
LUKE|14|30|говорячи: Чоловік цей почав будувати, але докінчити не міг...
LUKE|14|31|Або який цар, ідучи на війну супроти царя іншого, перше не сяде порадитися, чи спроможен він із десятьма тисячами стріти того, хто йде з двадцятьма тисячами проти нього?
LUKE|14|32|Коли ж ні, то, як той ще далеко, шле посольство до нього та й просить про мир.
LUKE|14|33|Так ото й кожен із вас, який не зречеться усього, що має, не може бути учнем Моїм.
LUKE|14|34|Сіль добра річ. Коли ж сіль несолоною стане, чим приправити її?
LUKE|14|35|Ні на землю, ні на гній не потрібна вона, її геть викидають. Хто має вуха, щоб слухати, нехай слухає!
LUKE|15|1|Наближались до Нього всі митники й грішники, щоб послухати Його.
LUKE|15|2|Фарисеї ж та книжники нарікали й казали: Приймає Він грішників та з ними їсть.
LUKE|15|3|А Він їм розповів оцю притчу, говорячи:
LUKE|15|4|Котрий з вас чоловік, мавши сотню овець і загубивши одну з них, не покине в пустині тих дев'ятидесяти й дев'яти, та й не піде шукати загинулої, аж поки не знайде її?
LUKE|15|5|А знайшовши, кладе на рамена свої та радіє.
LUKE|15|6|І, прийшовши додому, скликає він друзів і сусідів, та й каже до них: Радійте зо мною, бо знайшов я вівцю свою тую загублену.
LUKE|15|7|Говорю вам, що так само на небі радітимуть більш за одного грішника, що кається, аніж за дев'ятдесятьох і дев'ятьох праведників, що не потребують покаяння!...
LUKE|15|8|Або яка жінка, що має десять драхм, коли згубить драхму одну, не засвічує світла, і не мете хати, і не шукає уважно, аж поки не знайде?
LUKE|15|9|А знайшовши, кличе приятельок та сусідок та каже: Радійте зо мною, бо знайшла я загублену драхму!
LUKE|15|10|Так само, кажу вам, радість буває в Божих Анголів за одного грішника, який кається.
LUKE|15|11|І Він оповів: У чоловіка одного було два сини.
LUKE|15|12|І молодший із них сказав батькові: Дай мені, батьку, належну частину маєтку! І той поділив поміж ними маєток.
LUKE|15|13|А по небагатьох днях зібрав син молодший усе, та й подавсь до далекого краю, і розтратив маєток свій там, живучи марнотратно.
LUKE|15|14|А як він усе прожив, настав голод великий у тім краї, і він став бідувати.
LUKE|15|15|І пішов він тоді і пристав до одного з мешканців тієї землі, а той вислав його на поля свої пасти свиней.
LUKE|15|16|І бажав він наповнити шлунка свого хоч стручками, що їли їх свині, та ніхто не давав їх йому.
LUKE|15|17|Тоді він спам'ятався й сказав: Скільки в батька мого наймитів мають хліба аж надмір, а я отут з голоду гину!
LUKE|15|18|Устану, і піду я до батька свого, та й скажу йому: Прогрішився я, отче, против неба та супроти тебе...
LUKE|15|19|Недостойний я вже зватись сином твоїм; прийми ж мене, як одного з своїх наймитів...
LUKE|15|20|І, вставши, пішов він до батька свого. А коли він далеко ще був, його батько вгледів його, і переповнився жалем: і побіг він, і кинувсь на шию йому, і зачав цілувати його!
LUKE|15|21|І озвався до нього той син: Прогрішився я, отче, против неба та супроти тебе, і недостойний вже зватися сином твоїм...
LUKE|15|22|А батько рабам своїм каже: Принесіть негайно одежу найкращу, і його зодягніть, і персня подайте на руку йому, а сандалі на ноги.
LUKE|15|23|Приведіть теля відгодоване та заколіть, будемо їсти й радіти,
LUKE|15|24|бо цей син мій був мертвий і ожив, був пропав і знайшовся! І почали веселитись вони.
LUKE|15|25|А син старший його був на полі. І коли він ішов й наближався до дому, почув музики та танці.
LUKE|15|26|І покликав одного зо слуг, та й спитав: Що це таке?
LUKE|15|27|А той каже йому: То вернувся твій брат, і твій батько звелів заколоти теля відгодоване, бож здоровим його він прийняв.
LUKE|15|28|І розгнівався той, і ввійти не хотів. Тоді вийшов батько його й став просити його.
LUKE|15|29|А той відповів і до батька сказав: Ото, стільки років служу я тобі, і ніколи наказу твого не порушив, ти ж ніколи мені й козеняти не дав, щоб із приятелями своїми потішився я...
LUKE|15|30|Коли ж син твій вернувся оцей, що проїв твій маєток із блудницями, ти для нього звелів заколоти теля відгодоване...
LUKE|15|31|І сказав він йому: Ти завжди зо мною, дитино, і все моє то твоє!
LUKE|15|32|Веселитись та тішитись треба було, бо цей брат твій був мертвий і ожив, був пропав і знайшовся!
LUKE|16|1|Оповів же Він й учням Своїм: Один чоловік був багатий, і мав управителя, що оскаржений був перед ним, ніби він переводить маєток його.
LUKE|16|2|І він покликав його, і до нього сказав: Що це чую про тебе? Дай звіт про своє управительство, бо більше не зможеш рядити.
LUKE|16|3|І управитель почав міркувати собі: Що я маю робити, коли пан управительство відійме від мене? Копати не можу, просити соромлюсь.
LUKE|16|4|Знаю, що я зроблю, щоб мене прийняли до домів своїх, коли буду я скинений із управительства.
LUKE|16|5|І закликав він нарізно кожного з боржників свого пана, та й питається першого: Скільки винен ти панові моєму?
LUKE|16|6|А той відказав: Сто кадок оливи. І сказав він йому: Візьми ось розписку свою, швидко сідай та й пиши: п'ятдесят.
LUKE|16|7|А потім питається другого: А ти скільки винен? І той відказав: Сто кірців пшениці. І сказав він йому: Візьми ось розписку свою й напиши: вісімдесят.
LUKE|16|8|І пан похвалив управителя цього невірного, що він мудро вчинив. Бо сини цього світу в своїм поколінні мудріші, аніж сини світла.
LUKE|16|9|І Я вам кажу: Набувайте друзів собі від багатства неправедного, щоб, коли проминеться воно, прийняли вас до вічних осель.
LUKE|16|10|Хто вірний в найменшому, і в великому вірний; і хто несправедливий в найменшому, і в великому несправедливий.
LUKE|16|11|Отож, коли в несправедливім багатстві ви не були вірні, хто вам правдиве довірить?
LUKE|16|12|І коли ви в чужому не були вірні, хто ваше вам дасть?
LUKE|16|13|Жаден раб не може служить двом панам, бо або одного зненавидить, а другого буде любити, або буде триматись одного, а другого знехтує. Не можете Богові й мамоні служити!
LUKE|16|14|Чули все це й фарисеї, що були сріблолюбці, та й стали сміятися з Нього.
LUKE|16|15|Він же промовив до них: Ви себе видаєте за праведних перед людьми, але ваші серця знає Бог. Що бо високе в людей, те перед Богом гидота.
LUKE|16|16|Закон і Пророки були до Івана; відтоді Царство Боже благовіститься, і кожен силкується втиснутись в нього.
LUKE|16|17|Легше небо й земля проминеться, аніж одна риса з Закону загине.
LUKE|16|18|Кожен, хто дружину свою відпускає, і бере собі іншу, той чинить перелюб. І хто побереться з тією, яку хто відпустив, той чинить перелюб.
LUKE|16|19|Один чоловік був багатий, і зодягався в порфіру й віссон, і щоденно розкішно бенкетував.
LUKE|16|20|Був і вбогий один, на ім'я йому Лазар, що лежав у воріт його, струпами вкритий,
LUKE|16|21|і бажав годуватися кришками, що зо столу багатого падали; пси ж приходили й рани лизали йому...
LUKE|16|22|Та ось сталось, що вбогий умер, і на Авраамове лоно віднесли його Анголи. Умер же й багатий, і його поховали.
LUKE|16|23|І, терплячи муки в аду, звів він очі свої, та й побачив здаля Авраама та Лазаря на лоні його.
LUKE|16|24|І він закричав та сказав: Змилуйся, отче Аврааме, надо мною, і пошли мені Лазаря, нехай умочить у воду кінця свого пальця, і мого язика прохолодить, бо я мучуся в полум'ї цім!...
LUKE|16|25|Авраам же промовив: Згадай, сину, що ти вже прийняв за життя свого добре своє, а Лазар так само лихе; тепер він тут тішиться, а ти мучишся.
LUKE|16|26|А крім того всього, поміж нами та вами велика безодня поставлена, так що ті, що хочуть, переходити не можуть ізвідси до вас, ані не переходять ізвідти до нас.
LUKE|16|27|А він відказав: Отож, отче, благаю тебе, щоб його ти послав у дім батька мого,
LUKE|16|28|бо п'ятьох братів маю, хай він їм засвідчить, щоб і вони не прийшли на це місце страждання!
LUKE|16|29|Авраам же сказав: Вони мають Мойсея й Пророків, нехай слухають їх!
LUKE|16|30|А він відказав: Ні ж бо, отче Аврааме, але коли прийде хто з мертвих до них, то покаються.
LUKE|16|31|Йому ж він відказав: Як Мойсея й Пророків не слухають, то коли хто й із мертвих воскресне, не йнятимуть віри!
LUKE|17|1|І сказав Він до учнів Своїх: Неможливо, щоб спокуси не мали прийти; але горе тому, через кого приходять вони!
LUKE|17|2|Краще б такому було, коли б жорно млинове на шию йому почепити та й кинути в море, аніж щоб спокусив він одного з малих цих!
LUKE|17|3|Уважайте на себе! Коли провиниться твій брат, докори йому, а коли він покається, то вибач йому.
LUKE|17|4|І хоча б сім раз денно він провинивсь проти тебе, і сім раз звернувся до тебе, говорячи: Каюся, вибач йому!
LUKE|17|5|І сказали апостоли Господу: Додай Ти нам віри!
LUKE|17|6|А Господь відказав: Коли б мали ви віру, хоч як зерно гірчичне, і сказали шовковиці цій: Вирвися з коренем і посадися до моря, то й послухала б вас!
LUKE|17|7|Хто ж із вас, мавши раба, що оре чи пасе, скаже йому, як він вернеться з поля: Негайно йди та сідай до столу?
LUKE|17|8|Але чи ж не скаже йому: Приготуй що вечеряти, і підпережись, і мені прислуговуй, аж поки я їстиму й питиму, а потому ти сам будеш їсти та пити?
LUKE|17|9|Чи ж він дякує тому рабові, що наказане виконав?
LUKE|17|10|Так і ви, коли зробите все вам наказане, то кажіть: Ми нікчемні раби, бо зробили лиш те, що повинні зробити були!
LUKE|17|11|І сталось, коли Він ішов до Єрусалиму, то проходив поміж Самарією та Галілеєю.
LUKE|17|12|І, коли входив до одного села, перестріли Його десять мужів, слабих на проказу, що стали здалека.
LUKE|17|13|І голос піднесли вони та й казали: Ісусе, Наставнику, змилуйсь над нами!
LUKE|17|14|І, побачивши їх, Він промовив до них: Підіть і покажіться священикам! І сталось, коли вони йшли, то очистились...
LUKE|17|15|Один же з них, як побачив, що видужав, то вернувся, і почав гучним голосом славити Бога.
LUKE|17|16|І припав він обличчям до ніг Його, складаючи дяку Йому. А то самарянин був...
LUKE|17|17|Ісус же промовив у відповідь: Чи не десять очистилось, а дев'ять же де?
LUKE|17|18|Чому не вернулись вони хвалу Богові віддати, крім цього чужинця?
LUKE|17|19|І сказав Він йому: Підведися й іди: твоя віра спасла тебе!
LUKE|17|20|А як фарисеї спитали Його, коли Царство Божеє прийде, то Він їм відповів і сказав: Царство Боже не прийде помітно,
LUKE|17|21|і не скажуть: Ось тут, або: Там. Бо Божеє Царство всередині вас!
LUKE|17|22|І сказав Він до учнів: Прийдуть дні, коли побажаєте бачити один з днів Сина Людського, та не побачите...
LUKE|17|23|І скажуть до вас: Ось тут, чи: Ось там, не йдіть, і за ним не біжіть!
LUKE|17|24|Бо як блискавка, блиснувши, світить із одного краю під небом до другого краю під небом, так буде Свого дня й Син Людський.
LUKE|17|25|А перше належить багато страждати Йому, і відцурається рід цей від Нього...
LUKE|17|26|І, як було за днів Ноєвих, то буде так само й за днів Сина Людського:
LUKE|17|27|їли, пили, женилися, заміж виходили, аж до того дня, коли Ной увійшов до ковчегу; прийшов же потоп, і всіх вигубив.
LUKE|17|28|Так само, як було за днів Лотових: їли, пили, купували, продавали, садили, будували;
LUKE|17|29|того ж дня, як Лот вийшов із Содому, огонь із сіркою з неба линув, і всіх погубив.
LUKE|17|30|Так буде й того дня, як Син Людський з'явиться!
LUKE|17|31|Хто буде того дня на домі, а речі його будуть у домі, нехай їх забрати не злазить. Хто ж на полі, так само нехай назад не вертається,
LUKE|17|32|пам'ятайте про Лотову дружину!
LUKE|17|33|Хто дбатиме зберегти свою душу, той погубить її, а коли хто погубить, той оживить її.
LUKE|17|34|Кажу вам: удвох будуть ночі тієї на одному ліжкові: один візьметься, а другий полишиться.
LUKE|17|35|Дві молотимуть разом, одна візьметься, а друга полишиться.
LUKE|17|36|Двоє будуть на полі, один візьметься, а другий полишиться!
LUKE|17|37|І казали вони Йому в відповідь: Де, Господи? А Він відказав їм: Де труп, там зберуться й орли...
LUKE|18|1|І Він розповів їм і притчу про те, що треба молитися завжди, і не занепадати духом,
LUKE|18|2|говорячи: У місті якомусь суддя був один, що Бога не боявся, і людей не соромився.
LUKE|18|3|У тому ж місті вдова перебувала, що до нього ходила й казала: Оборони мене від мого супротивника!
LUKE|18|4|Але він довгий час не хотів. А згодом сказав сам до себе: Хоч і Бога я не боюся, і людей не соромлюся,
LUKE|18|5|але через те, що вдовиця оця докучає мені, то візьму в оборону її, щоб вона без кінця не ходила, і не докучала мені.
LUKE|18|6|І промовив Господь: Чи чуєте, що говорить суддя цей неправедний?
LUKE|18|7|А чи ж Бог в оборону не візьме обраних Своїх, що голосять до Нього день і ніч, хоч і бариться Він щодо них?
LUKE|18|8|Кажу вам, що Він їм незабаром подасть оборону! Та Син Людський, як прийде, чи Він на землі знайде віру?...
LUKE|18|9|А для деяких, що були себе певні, що вони ніби праведні, і за ніщо мали інших, Він притчу оцю розповів.
LUKE|18|10|Два чоловіки до храму ввійшли помолитись, один фарисей, а другий був митник.
LUKE|18|11|Фарисей, ставши, так молився про себе: Дякую, Боже, Тобі, що я не такий, як інші люди: здирщики, неправедні, перелюбні, або як цей митник.
LUKE|18|12|Я пощу два рази на тиждень, даю десятину з усього, що тільки надбаю!
LUKE|18|13|А митник здалека стояв, та й очей навіть звести до неба не смів, але бив себе в груди й казав: Боже, будь милостивий до мене грішного!...
LUKE|18|14|Говорю вам, що цей повернувся до дому свого більш виправданий, аніж той. Бо кожен, хто підноситься, буде понижений, хто ж понижається, той піднесеться.
LUKE|18|15|До Нього ж приносили й немовлят, щоб до них доторкнувся, а учні, побачивши, їм докоряли.
LUKE|18|16|А Ісус їх покликав та й каже: Пустіте дітей, щоб до Мене приходили, і не забороняйте їм, бо таких Царство Боже.
LUKE|18|17|Поправді кажу вам: Хто Божого Царства не прийме, як дитя, той у нього не ввійде!
LUKE|18|18|І запитався Його один із начальників, говорячи: Учителю Добрий, що робити мені, щоб вспадкувати вічне життя?
LUKE|18|19|Ісус же йому відказав: Чого звеш Мене Добрим? Ніхто не є Добрий, тільки Сам Бог!
LUKE|18|20|Знаєш заповіді: Не чини перелюбу, не вбивай, не кради, не свідкуй неправдиво, шануй свого батька та матір.
LUKE|18|21|А він відказав: Усе це я виконав від юнацтва свого!
LUKE|18|22|Як почув це Ісус, то промовив до нього: Одного тобі ще бракує: Розпродай усе, що ти маєш, і вбогим роздай, і матимеш скарб свій на небі. Вертайся тоді, та й іди вслід за Мною!
LUKE|18|23|А він, коли почув це, то засумував, бо був вельми багатий.
LUKE|18|24|Як побачив Ісус, що той засумував, то промовив: Як тяжко багатим увійти в Царство Боже!
LUKE|18|25|Бо верблюдові легше пройти через голчине вушко, ніж багатому в Божеє Царство ввійти...
LUKE|18|26|Ті ж, що чули, спитали: Хто ж тоді може спастися?
LUKE|18|27|А Він відповів: Неможливеє людям можливе для Бога!
LUKE|18|28|І промовив Петро: От усе ми покинули, та й пішли за Тобою слідом.
LUKE|18|29|А Ісус відказав їм: Поправді кажу вам: Немає такого, щоб покинув свій дім, або дружину, чи братів, чи батьків, чи дітей ради Божого Царства,
LUKE|18|30|і не одержав би значно більш цього часу, а в віці наступнім життя вічне.
LUKE|18|31|І, взявши Дванадцятьох, промовив до них: Оце в Єрусалим ми йдемо, і все здійсниться, що писали Пророки про Людського Сина.
LUKE|18|32|Бо Він виданий буде поганам, і буде осміяний, і покривджений, і опльований,
LUKE|18|33|і, збичувавши, уб'ють Його, але третього дня Він воскресне!
LUKE|18|34|Та з цього нічого вони не збагнули, і ця річ перед ними закрита була, і сказаного вони не розуміли.
LUKE|18|35|І сталось, як Він наближався був до Єрихону, один невидющий сидів при дорозі й просив.
LUKE|18|36|А коли він прочув, що проходить народ, то спитався: Що це таке?
LUKE|18|37|А йому відказали, що проходить Ісус Назарянин.
LUKE|18|38|І став він кричати й казати: Ісусе, Сину Давидів, змилуйся надо мною!
LUKE|18|39|А ті, що попереду йшли, сварились на нього, щоб він замовк, а він іще більше кричав: Сину Давидів, змилуйся надо мною!
LUKE|18|40|І спинився Ісус, і привести його до Себе звелів. А коли той наблизивсь до Нього, то Він запитався його:
LUKE|18|41|Що ти хочеш, щоб зробив Я тобі? А той відповів: Господи, нехай стану видющим!
LUKE|18|42|Ісус же до нього сказав. Стань видющий! Твоя віра спасла тебе!
LUKE|18|43|І зараз видющим той став, і пішов вслід за Ним, прославляючи Бога. А всі люди, бачивши це, віддали хвалу Богові.
LUKE|19|1|І, ввійшовши Ісус, переходив через Єрихон.
LUKE|19|2|І ось чоловік, що звався Закхей, він був старший над митниками, і був багатий,
LUKE|19|3|бажав бачити Ісуса, хто Він, але з-за народу не міг, бо малий був на зріст.
LUKE|19|4|І, забігши вперед, він виліз на фіґове дерево, щоб бачити Його, бо Він мав побіч нього проходити.
LUKE|19|5|А коли на це місце Ісус підійшов, то поглянув угору до нього й промовив: Закхею, зійди зараз додолу, бо сьогодні потрібно Мені бути в домі твоїм!
LUKE|19|6|І той зараз додолу ізліз, і прийняв Його з радістю.
LUKE|19|7|А всі, як побачили це, почали нарікати, і казали: Він до грішного мужа в гостину зайшов!
LUKE|19|8|Став же Закхей та й промовив до Господа: Господи, половину маєтку свого я віддам ось убогим, а коли кого скривдив був чим, верну вчетверо.
LUKE|19|9|Ісус же промовив до нього: Сьогодні на дім цей спасіння прийшло, бо й він син Авраамів.
LUKE|19|10|Син бо Людський прийшов, щоб знайти та спасти, що загинуло!
LUKE|19|11|Коли ж вони слухали це, розповів Він іще одну притчу, бо Він був недалеко від Єрусалиму, вони ж думали, що об'явиться Боже Царство тепер.
LUKE|19|12|Отож Він сказав: Один чоловік, роду славного, відправлявся в далеку країну, щоб царство прийняти й вернутись.
LUKE|19|13|І покликав він десятьох своїх рабів, дав їм десять мін, і сказав їм: Торгуйте, аж поки вернуся.
LUKE|19|14|Та його громадяни його ненавиділи, і послали посланців услід за ним, кажучи: Не хочемо, щоб він був над нами царем.
LUKE|19|15|І сталось, коли він вернувся, як царство прийняв, то звелів поскликати рабів, яким срібло роздав, щоб довідатися, хто що набув.
LUKE|19|16|І перший прийшов і сказав: Пане, міна твоя принесла десять мін.
LUKE|19|17|І відказав він йому: Гаразд, рабе добрий! Ти в малому був вірний, володій десятьма містами.
LUKE|19|18|І другий прийшов і сказав: Пане, твоя міна п'ять мін принесла.
LUKE|19|19|Він же сказав і тому: Будь і ти над п'ятьма містами.
LUKE|19|20|І ще інший прийшов і сказав: Пане, ось міна твоя, що я мав її сховану в хустці.
LUKE|19|21|Я бо боявся тебе, ти ж бо людина жорстока: береш, чого не поклав, і жнеш, чого не посіяв.
LUKE|19|22|І відказав той йому: Устами твоїми, злий рабе, суджу я тебе! Ти знав, що я жорстока людина, беру, чого не поклав, і жну, чого не посіяв.
LUKE|19|23|Чому ж не віддав ти міняльникам срібла мого, і я, повернувшись, узяв би своє із прибутком?
LUKE|19|24|І сказав він присутнім: Візьміть міну від нього, та дайте тому, хто десять мін має.
LUKE|19|25|І відказали йому: Пане, він десять мін має.
LUKE|19|26|Говорю бо я вам: Кожному, хто має, то дасться йому, хто ж не має, забереться від нього і те, що він має.
LUKE|19|27|А тих ворогів моїх, які не хотіли, щоб царював я над ними, приведіте сюди, і на очах моїх їх повбивайте.
LUKE|19|28|А як це оповів, Він далі пішов, простуючи в Єрусалим.
LUKE|19|29|І ото, як наблизився до Вітфагії й Віфанії, на горі, що Оливною зветься, Він двох учнів послав,
LUKE|19|30|наказуючи: Ідіть у село, яке перед вами; увійшовши до нього, знайдете прив'язане осля, що на нього ніколи ніхто із людей не сідав. Відв'яжіть його, і приведіть.
LUKE|19|31|Коли ж вас хто спитає: Нащо відв'язуєте?, відкажіть тому так: Господь потребує його.
LUKE|19|32|Посланці ж відійшли, і знайшли, як Він їм був сказав.
LUKE|19|33|А коли осля стали відв'язувати, хазяї його їх запитали: Нащо осля ви відв'язуєте?
LUKE|19|34|Вони ж відказали: Господь потребує його.
LUKE|19|35|І вони привели до Ісуса його, і, поклавши одежу свою на осля, посадили Ісуса.
LUKE|19|36|Коли ж Він їхав, вони простилали одежу свою по дорозі.
LUKE|19|37|А як Він наближався вже до сходу з гори Оливної, то ввесь натовп учнів, радіючи, почав гучним голосом Бога хвалити за всі чуда, що бачили,
LUKE|19|38|кажучи: Благословенний Цар, що йде у Господнє Ім'я! Мир на небесах, і слава на висоті!
LUKE|19|39|А деякі фарисеї з народу сказали до Нього: Учителю, заборони Своїм учням!
LUKE|19|40|А Він їм промовив у відповідь: Кажу вам, що коли ці замовкнуть, то каміння кричатиме!
LUKE|19|41|І коли Він наблизився, і місто побачив, то заплакав за ним,
LUKE|19|42|і сказав: О, якби й ти хоч цього дня пізнало, що потрібне для миру тобі! Та тепер від очей твоїх сховане це.
LUKE|19|43|Бо прийдуть на тебе ті дні, і твої вороги тебе валом оточать, і обляжуть тебе, і стиснуть тебе звідусюди.
LUKE|19|44|І зрівняють з землею тебе, і поб'ють твої діти в тобі, і не позоставлять у тобі каменя на камені, бо не зрозуміло ти часу відвідин твоїх...
LUKE|19|45|А коли Він у храм увійшов, то почав виганяти продавців,
LUKE|19|46|до них кажучи: Написано: Дім Мій дім молитви, а ви з нього зробили печеру розбійників.
LUKE|19|47|І Він кожного дня у храмі навчав. А первосвященики й книжники й найважніші з народу шукали, щоб Його погубити,
LUKE|19|48|але не знаходили, що вчинити Йому, бо ввесь народ горнувся до Нього та слухав Його.
LUKE|20|1|І сталось одного з тих днів, як навчав Він у храмі людей, та Добру Новину звіщав, прийшли первосвященики й книжники з старшими,
LUKE|20|2|та й до Нього промовили, кажучи: Скажи нам, якою владою Ти чиниш оце? Або хто Тобі владу цю дав?
LUKE|20|3|І промовив до них Він у відповідь: Запитаю й Я вас одну річ, і відповідайте Мені:
LUKE|20|4|Іванове хрищення з неба було, чи від людей?
LUKE|20|5|Вони ж міркували собі й говорили: Коли скажемо: З неба, відкаже: Чого ж ви йому не повірили?
LUKE|20|6|А як скажемо: Від людей, то всі люди камінням поб'ють нас, бо були переконані, що Іван то пророк.
LUKE|20|7|І вони відповіли, що не знають, ізвідки...
LUKE|20|8|А Ісус відказав їм: То й Я не скажу вам, якою владою Я це чиню.
LUKE|20|9|І Він розповідати почав людям притчу оцю. Один чоловік насадив виноградника, і віддав його винарям, та й відбув на час довший.
LUKE|20|10|А певного часу послав він раба до своїх винарів, щоб дали йому частку з плодів виноградника. Та побили його винарі, і відіслали ні з чим.
LUKE|20|11|І знову послав він до них раба іншого, а вони й того збили й зневажили, та й відіслали ні з чим.
LUKE|20|12|І послав він ще третього, а вони й того зранили й вигнали.
LUKE|20|13|Сказав тоді пан виноградника: Що маю робити? Пошлю свого сина улюбленого, може його посоромляться...
LUKE|20|14|Винарі ж, як його вгледіли, міркували собі та казали: Це спадкоємець; ходім, замордуймо його, щоб спадщина наша була.
LUKE|20|15|І вони його вивели за виноградника, та й убили... Що ж зробить їм пан виноградника?
LUKE|20|16|Він прийде та й вигубить цих винарів, виноградника ж іншим віддасть. Слухачі ж повіли: Нехай цього не станеться!
LUKE|20|17|А Він глянув на них та й сказав: Що ж оце, що написане: Камінь, що його будівничі відкинули, той наріжним став каменем!
LUKE|20|18|Кожен, хто впаде на цей камінь розіб'ється, а на кого він сам упаде, то розчавить його.
LUKE|20|19|А книжники й первосвященики руки на Нього хотіли накласти тієї години, але побоялись народу. Бо вони розуміли, що про них Він цю притчу сказав.
LUKE|20|20|І вони слідкували за Ним, і підіслали підглядачів, які праведних із себе вдавали, щоб зловити на слові Його, і Його видати урядові й владі намісника.
LUKE|20|21|І вони запитали Його та сказали: Учителю, знаємо ми, що Ти добре говориш і навчаєш, і не дивишся на обличчя, але наставляєш на Божу дорогу правдиво.
LUKE|20|22|Чи годиться давати податок для кесаря, чи ні?
LUKE|20|23|Знаючи ж їхню хитрість, сказав Він до них: Чого ви Мене випробовуєте?
LUKE|20|24|Покажіте динарія Мені. Чий образ і напис він має? Вони відказали: Кесарів.
LUKE|20|25|А Він їм відказав: Тож віддайте кесареве кесареві, а Богові Боже!
LUKE|20|26|І не могли вони перед людьми зловити на слові Його. І дивувались вони з Його відповіді, та й замовкли.
LUKE|20|27|І підійшли дехто із саддукеїв, що твердять, ніби немає воскресіння, і запитали Його,
LUKE|20|28|та сказали: Учителю, Мойсей написав нам: Як умре кому брат, який має дружину, а помре бездітний, то нехай його брат візьме дружину, і відновить насіння для брата свого.
LUKE|20|29|Було ж сім братів. І перший, узявши дружину, бездітний умер.
LUKE|20|30|І другий узяв був ту дружину, та й той вмер бездітний.
LUKE|20|31|І третій узяв був її, так само й усі семеро, і вони дітей не позоставили, та й повмирали.
LUKE|20|32|А по всіх умерла й жінка.
LUKE|20|33|А в воскресінні котрому із них вона дружиною буде? Бо семеро мали за дружину її.
LUKE|20|34|Ісус же промовив у відповідь їм: Женяться й заміж виходять сини цього віку.
LUKE|20|35|А ті, що будуть достойні того віку й воскресіння з мертвих, не будуть ні женитись, ні заміж виходити,
LUKE|20|36|ні вмерти вже не можуть, бо рівні вони Анголам, і вони сини Божі, синами воскресіння бувши.
LUKE|20|37|А що мертві встають, то й Мойсей показав при кущі, коли він назвав Господа Богом Авраамовим, і Богом Ісаковим, і Богом Якововим.
LUKE|20|38|Бог же не є Богом мертвих, а живих, бо всі в Нього живуть.
LUKE|20|39|Дехто ж із книжників відповіли та сказали: Учителю, Ти добре сказав!
LUKE|20|40|І вже не насмілювалися питати Його ні про що.
LUKE|20|41|І сказав Він до них: Як то кажуть, що Христос син Давидів?
LUKE|20|42|Таж Давид сам говорить у книзі Псалмів: Промовив Господь Господеві моєму: сядь праворуч Мене,
LUKE|20|43|поки не покладу Я Твоїх ворогів підніжком ногам Твоїм!
LUKE|20|44|Отже, Давид Його Господом зве, як же Він йому син?
LUKE|20|45|І, як увесь народ слухав, Він промовив до учнів Своїх:
LUKE|20|46|Стережіться книжників, що хочуть у довгих одежах ходити, і люблять привіти на ринках, і перші лавки в синагогах, і перші місця на бенкетах,
LUKE|20|47|що вдовині хати поїдають, і моляться довго напоказ, вони тяжче осудження приймуть!
LUKE|21|1|І поглянув Він угору, і побачив заможних, що кидали дари свої до скарбниці.
LUKE|21|2|Побачив і вбогу вдовицю одну, що дві лепті туди вона вкинула.
LUKE|21|3|І сказав Він: Поправді кажу вам, що ця вбога вдовиця вкинула більше за всіх!
LUKE|21|4|Бо всі клали від лишка свого в дар Богові, а вона поклала з убозтва свого ввесь прожиток, що мала...
LUKE|21|5|Коли ж дехто казав про храм, що прикрашений дорогоцінним камінням та дарами, тоді Він прорік:
LUKE|21|6|Надійдуть ті дні, коли з того, що бачите, не зостанеться й каменя на камені, який не зруйнується...
LUKE|21|7|І запитали Його та сказали: Учителю, коли ж оце станеться? І, яка буде ознака, коли має початися це?
LUKE|21|8|Він же промовив: Стережіться, щоб вас хто не звів. Бо багато-хто прийдуть в Ім'я Моє, кажучи: Це Я, і Час наблизився. Та за ними не йдіть!
LUKE|21|9|І, як про війни та розрухи почуєте ви, не лякайтесь, бо перш статись належить тому. Але це не кінець ще.
LUKE|21|10|Тоді промовляв Він до них: Повстане народ на народ, і царство на царство.
LUKE|21|11|І будуть землетруси великі та голод, та помір місцями, і страшні та великі ознаки на небі.
LUKE|21|12|Але перед усім тим накладуть на вас руки свої, і переслідувати будуть, і видаватимуть вас у синагоги й в'язниці, і поведуть вас до царів та правителів через Ім'я Моє.
LUKE|21|13|Але це стане вам на свідоцтво.
LUKE|21|14|Отож, покладіть у серця свої наперед не гадати, що будете відповідати,
LUKE|21|15|бо дам Я вам мову та мудрість, що не зможуть противитись чи суперечити їй всі противники ваші.
LUKE|21|16|І будуть вас видавати і батьки, і брати, і рідня, і друзі, а декому з вас заподіють і смерть.
LUKE|21|17|І за Ім'я Моє будуть усі вас ненавидіти.
LUKE|21|18|Але й волосина вам із голови не загине!
LUKE|21|19|Терпеливістю вашою душі свої ви здобудете.
LUKE|21|20|А коли ви побачите Єрусалим, військом оточений, тоді знайте, що до нього наблизилося спустошення.
LUKE|21|21|Тоді ті, хто в Юдеї, нехай у гори втікають; хто ж у середині міста, нехай вийдуть; хто ж в околицях, хай не вертаються в нього!
LUKE|21|22|Бо то будуть дні помсти, щоб виконалося все написане.
LUKE|21|23|Горе ж вагітним та тим, хто годує грудьми, у ті дні, бо буде велика нужда на землі та гнів над цим людом!
LUKE|21|24|І поляжуть під гострим мечем, і заберуть до неволі поміж усі народи, і погани топтатимуть Єрусалим, аж поки не скінчиться час тих поган...
LUKE|21|25|І будуть ознаки на сонці, і місяці, і зорях, і тривога людей на землі, і збентеження від шуму моря та хвиль,
LUKE|21|26|коли люди будуть мертвіти від страху й чекання того, що йде на ввесь світ, бо сили небесні порушаться.
LUKE|21|27|І побачать тоді Сина Людського, що йтиме на хмарах із силою й великою славою!
LUKE|21|28|Коли ж стане збуватися це, то випростуйтесь, і підійміть свої голови, бо зближається ваше визволення!
LUKE|21|29|І розповів Він їм притчу: Погляньте на фіґове дерево, і на всілякі дерева:
LUKE|21|30|як вони вже розпукуються, то, бачивши це, самі знаєте, що близько вже літо.
LUKE|21|31|Так і ви, як побачите, що діється це, то знайте, що Боже Царство вже близько!
LUKE|21|32|Поправді кажу вам: Не перейде цей рід, аж усе оце станеться.
LUKE|21|33|Небо й земля проминуться, але не минуться слова Мої!
LUKE|21|34|Уважайте ж на себе, щоб ваші серця не обтяжувалися ненажерством та п'янством, і життєвими клопотами, і щоб день той на вас не прийшов несподівано,
LUKE|21|35|немов сітка; бо він прийде на всіх, що живуть на поверхні всієї землі.
LUKE|21|36|Тож пильнуйте, і кожного часу моліться, щоб змогли ви уникнути всього того, що має відбутись, та стати перед Сином Людським!
LUKE|21|37|За дня ж Він у храмі навчав, а на ніч виходив та перебував на горі, що зветься Оливна.
LUKE|21|38|А зранку всі люди до Нього приходили в храм, щоб послухати Його.
LUKE|22|1|Наближалося ж свято Опрісноків, що Пасхою зветься.
LUKE|22|2|А первосвященики й книжники стали шукати, як би вбити Його, та боялись народу...
LUKE|22|3|Сатана ж увійшов у Юду, званого Іскаріот, одного з Дванадцятьох.
LUKE|22|4|І він пішов, і почав умовлятися з первосвящениками та начальниками, як він видасть Його.
LUKE|22|5|Ті ж зраділи, і погодилися дати йому срібняків.
LUKE|22|6|І він обіцяв, і шукав відповідного часу, щоб їм видати Його без народу...
LUKE|22|7|І настав день Опрісноків, коли пасху приносити в жертву належало.
LUKE|22|8|І послав Він Петра та Івана, говорячи: Підіть, і приготуйте нам пасху, щоб її спожили ми.
LUKE|22|9|А вони запитали Його: Де Ти хочеш, щоб ми приготували?
LUKE|22|10|А Він їм відказав: Ось, як будете входити в місто, стріне вас чоловік, воду несучи у глекові, ідіть за ним аж до дому, куди він увійде.
LUKE|22|11|І скажіть до господаря дому: Учитель питає тебе: Де кімната, в якій споживу зо Своїми учнями пасху?
LUKE|22|12|І він вам покаже велику горницю вистелену: там приготуйте.
LUKE|22|13|І вони відійшли, і знайшли, як Він їм говорив, і зачали там готувати пасху.
LUKE|22|14|А коли настав час, сів до столу, і апостоли з Ним.
LUKE|22|15|І промовив до них: Я дуже бажав спожити цю пасху із вами, перш ніж муки прийму.
LUKE|22|16|Бо кажу вам, що вже споживати не буду її, поки сповниться в Божому Царстві вона.
LUKE|22|17|Узявши ж чашу, і вчинивши подяку, Він промовив: Візьміть її, і поділіть між собою.
LUKE|22|18|Кажу ж вам, що віднині не питиму Я від оцього плоду виноградного, доки Божеє Царство не прийде.
LUKE|22|19|Узявши ж хліб і вчинивши подяку, поламав і дав їм, проказуючи: Це тіло Моє, що за вас віддається. Це чиніть на спомин про Мене!
LUKE|22|20|По вечері так само ж і чашу, говорячи: Оця чаша Новий Заповіт у Моїй крові, що за вас проливається.
LUKE|22|21|Та однак, за столом ось зо Мною рука Мого зрадника.
LUKE|22|22|Бо Син Людський іде, як призначено; але горе тому чоловікові, хто Його видає!
LUKE|22|23|А вони почали між собою питати, котрий з них мав би це вчинити?
LUKE|22|24|І сталось між ними й змагання, котрий з них уважатися має за більшого.
LUKE|22|25|Він же промовив до них: Царі народів панують над ними, а ті, що ними володіють, доброчинцями звуться.
LUKE|22|26|Але не так ви: хто найбільший між вами, нехай буде, як менший, а начальник як службовець.
LUKE|22|27|Бо хто більший: чи той, хто сидить при столі, чи хто прислуговує? Чи не той, хто сидить при столі? А Я серед вас, як службовець.
LUKE|22|28|Ви ж оті, що перетривали зо Мною в спокусах Моїх,
LUKE|22|29|і Я вам заповітую Царство, як Отець Мій Мені заповів,
LUKE|22|30|щоб ви в Царстві Моїм споживали й пили за столом Моїм, і щоб ви на престолах засіли судити дванадцять племен Ізраїлевих.
LUKE|22|31|І промовив Господь: Симоне, Симоне, ось сатана жадав вас, щоб вас пересіяти, мов ту пшеницю.
LUKE|22|32|Я ж молився за тебе, щоб не зменшилась віра твоя; ти ж колись, як навернешся, зміцни браттю свою!
LUKE|22|33|А той відказав Йому: Господи, я з Тобою готовий іти до в'язниці й на смерть!
LUKE|22|34|Він же прорік: Говорю тобі, Петре, півень не заспіває сьогодні, як ти тричі зречешся, що не знаєш Мене...
LUKE|22|35|І Він їм сказав: Як Я вас посилав без калитки, і без торби, і без сандаль, чи вам бракувало чого? Вони ж відказали: Нічого.
LUKE|22|36|А тепер каже їм хто має калитку, нехай візьме, теж і торбу; хто ж не має, нехай продасть одіж свою та й купить меча.
LUKE|22|37|Говорю бо Я вам, що виконатися на Мені має й це ось написане: До злочинців Його зараховано. Бо те, що про Мене, виконується.
LUKE|22|38|І сказали вони: Господи, ось тут два мечі. А Він їм відказав: Досить!
LUKE|22|39|І Він вийшов, і пішов за звичаєм на гору Оливну. А за Ним пішли учні Його.
LUKE|22|40|А прийшовши на місце, сказав їм: Моліться, щоб не впасти в спокусу.
LUKE|22|41|А Він Сам, відійшовши від них, як докинути каменем, на коліна припав та й молився,
LUKE|22|42|благаючи: Отче, як волієш, пронеси мимо Мене цю чашу! Та проте не Моя, а Твоя нехай станеться воля!...
LUKE|22|43|І Ангол із неба з'явився до Нього, і додавав Йому сили.
LUKE|22|44|А як був у смертельній тривозі, ще пильніш Він молився. І піт Його став, немов каплі крови, що спливали на землю...
LUKE|22|45|І, підвівшись з молитви, Він до учнів прийшов, і знайшов їх, що спали з журби...
LUKE|22|46|І промовив до них: Чого ви спите? Уставайте й моліться, щоб не впасти в спокусу!
LUKE|22|47|І, коли Він іще говорив, ось народ з'явився, і один із Дванадцятьох, що Юдою зветься, ішов перед ними. І він підійшов до Ісуса, щоб поцілувати Його. Бо він знака їм дав був: кого я поцілую, то Він!
LUKE|22|48|Ісус же промовив до нього: Чи оце поцілунком ти, Юдо, видаєш Сина Людського?
LUKE|22|49|А ті, що були з Ним, як побачили, що має статись, сказали Йому: Господи, чи мечем нам не вдарити?
LUKE|22|50|І, один із них рубонув раба первосвященикового, та й відтяв праве вухо йому.
LUKE|22|51|Та Ісус відізвався й сказав: Лишіть, уже досить! І, доторкнувшись до вуха його, уздоровив його.
LUKE|22|52|А до первосвящеників і влади сторожі храму та старших, що прийшли проти Нього, промовив Ісус: Немов на розбійника вийшли з мечами та киями...
LUKE|22|53|Як щоденно Я з вами у храмі бував, не піднесли на Мене ви рук. Та це ваша година тепер, і влада темряви...
LUKE|22|54|А схопивши Його, повели й привели у дім первосвященика. Петро ж здалека йшов слідкома.
LUKE|22|55|Як розклали ж огонь серед двору, і вкупі сиділи, сидів і Петро поміж ними.
LUKE|22|56|А служниця одна його вгледіла, як сидів коло світла, і, придивившись до нього, сказала: І цей був із Ним!
LUKE|22|57|І відрікся від Нього він, твердячи: Не знаю я, жінко, Його!
LUKE|22|58|Незабаром же другий побачив його та й сказав: І ти від отих. А Петро відказав: Ні, чоловіче!...
LUKE|22|59|І як часу минуло з годину, хтось інший твердив і казав: Поправді, і цей був із Ним, бо він галілеянин.
LUKE|22|60|А Петро відказав: Чоловіче, не відаю, про що ти говориш... І зараз, як іще говорив він, півень заспівав.
LUKE|22|61|І Господь обернувся й подививсь на Петра. А Петро згадав слово Господнє, як сказав Він йому: Перше, ніж заспіває півень, відречешся ти тричі від Мене.
LUKE|22|62|І, вийшовши звідти, він гірко заплакав!
LUKE|22|63|А люди, які ув'язнили Ісуса, знущалися з Нього та били.
LUKE|22|64|І, закривши Його, вони били Його по обличчі, і питали Його, приговорюючи: Пророкуй, хто то вдарив Тебе?
LUKE|22|65|І багато інших богозневаг говорили на Нього вони...
LUKE|22|66|А коли настав день, то зібралися старші народу, первосвященики й книжники, і повели Його в синедріон свій,
LUKE|22|67|і казали: Коли Ти Христос, скажи нам. А Він їм відповів: Коли Я вам скажу, не повірите ви.
LUKE|22|68|А коли й поспитаю вас Я, не дасте Мені відповіді.
LUKE|22|69|Незабаром Син Людський сидітиме по правиці сили Божої!
LUKE|22|70|Тоді всі запитали: То Ти Божий Син? А Він їм відповів: Самі кажете ви, що то Я...
LUKE|22|71|А вони відказали: Нащо потрібні ще свідки для нас? Бо ми чули самі з Його уст!
LUKE|23|1|І знялися всі їхні збори, і повели до Пилата Його.
LUKE|23|2|І зачали оскаржати Його й говорити: Ми ствердили, що Цей ворохобить народ наш, і забороняє податок давати кесареві, та й говорить, що Він, Христос Цар.
LUKE|23|3|І Пилат запитав Його, кажучи: Чи Ти Цар Юдейський? А Він відказав йому в відповідь: Сам ти кажеш...
LUKE|23|4|І Пилат сказав первосвященикам та до народу: Я не знаходжу жадної провини в Цій Людині.
LUKE|23|5|А вони намагались, говорячи: Він бунтує народ, навчаючи в усій Юдеї, від Галілеї почавши аж посі.
LUKE|23|6|А Пилат, вчувши про Галілею, спитав: Хіба Він галілеянин?
LUKE|23|7|І, дізнавшись, що Він із влади Ірода, відіслав Його Іродові, бо той в Єрусалимі також перебував тими днями.
LUKE|23|8|Коли ж Ірод побачив Ісуса, то дуже зрадів, бо він від давнього часу бажав Його бачити, багато за Нього чував, і сподівався побачити чудо яке, що буває від Нього.
LUKE|23|9|І багато питався Його, та нічого не відповідав Він йому.
LUKE|23|10|І стояли тут первосвященики й книжники, та завзято Його оскаржали.
LUKE|23|11|Тоді Ірод із військом своїм ізневажив Його й насміявся, зодягнувши Його в яснобілу одіж, і відіслав до Пилата Його.
LUKE|23|12|І того дня стали Ірод із Пилатом за приятелів між собою, бо давніш ворожнеча між ними була.
LUKE|23|13|А Пилат скликав первосвящеників, і старшин, і народ,
LUKE|23|14|і промовив до них: Привели ви мені Чоловіка Цього, як того, що бунтує народ. А ось я перед вами розвідав, і не знаходжу в Людині Оцій ані однієї провини такої, про що ви оскаржаєте.
LUKE|23|15|Також Ірод, бо він відіслав Його нам. І ось нічого, що на смерть заслуговувало б, Він не вчинив.
LUKE|23|16|Отже я покараю Його й відпущу.
LUKE|23|17|Бо повинен був їм відпустити одного на свято.
LUKE|23|18|А народ став кричати й казати: Візьми Цього, відпусти ж нам Варавву!
LUKE|23|19|А той за повстання одне, яке сталося в місті, і за вбивство посаджений був до в'язниці.
LUKE|23|20|І знову сказав їм Пилат, хотячи відпустити Ісуса.
LUKE|23|21|Та кричали вони й говорили: Розіпни, розіпни Його!
LUKE|23|22|Він же втретє промовив до них: Яке ж зло вчинив Він? Я нічого, що на смерть заслуговувало б, на Нім не знайшов. Отже я покараю Його й відпущу.
LUKE|23|23|А вони сильним криком свого домагалися, та вимагали розп'ясти Його. І взяв гору крик їхній та первосвящеників.
LUKE|23|24|І Пилат присудив, щоб було, як просили вони:
LUKE|23|25|відпустив їм Варавву, посадженого за повстання та вбивство в в'язницю, за якого просили вони, а Ісуса віддав їхній волі...
LUKE|23|26|І як Його повели, то схопили якогось Симона із Кірінеї, що з поля вертався, і поклали на нього хреста, щоб він ніс за Ісусом!
LUKE|23|27|А за Ним ішов натовп великий людей і жінок, які плакали та голосили за Ним.
LUKE|23|28|А Ісус обернувся до них та й промовив: Дочки єрусалимські, не ридайте за Мною, за собою ридайте й за дітьми своїми!
LUKE|23|29|Бо ось дні настають, коли скажуть: Блаженні неплідні, та утроби, які не родили, і груди, що не годували...
LUKE|23|30|Тоді стануть казати горам: Поспадайте на нас, а узгір'ям: Покрийте нас!
LUKE|23|31|Бо коли таке роблять зеленому дереву, то що буде сухому?
LUKE|23|32|І вели з Ним також двох злочинників інших, щоб убити.
LUKE|23|33|А коли прибули на те місце, що звуть Череповище, розп'яли тут Його та злочинників, одного праворуч, а одного ліворуч.
LUKE|23|34|Ісус же промовив: Отче, відпусти їм, бо не знають, що чинять вони!... А як Його одіж ділили, то кидали жереба.
LUKE|23|35|А люди стояли й дивились... Насміхалися з ними й старшини, говорячи: Він інших спасав, нехай Сам Себе визволить, коли Він Христос, Божий Обранець!
LUKE|23|36|І вояки глузували з Нього: приступаючи, оцет Йому подавали,
LUKE|23|37|і казали: Коли Цар Ти Юдейський, спаси Себе Сам!
LUKE|23|38|Був же й напис над Ним письмом грецьким, латинським і гебрейським написаний: Це Цар Юдейський.
LUKE|23|39|А один із розп'ятих злочинників став зневажати Його й говорити: Чи Ти не Христос? То спаси Себе й нас!
LUKE|23|40|Обізвався ж той другий, і докоряв йому, кажучи: Чи не боїшся ти Бога, коли й сам на те саме засуджений?
LUKE|23|41|Але ми справедливо засуджені, і належну заплату за вчинки свої беремо, Цей же жадного зла не вчинив.
LUKE|23|42|І сказав до Ісуса: Спогадай мене, Господи, коли прийдеш у Царство Своє!
LUKE|23|43|І промовив до нього Ісус: Поправді кажу тобі: ти будеш зо Мною сьогодні в раю!
LUKE|23|44|Наближалася шоста година, і темрява стала по цілій землі аж до години дев'ятої...
LUKE|23|45|І сонце затьмилось, і в храмі завіса роздерлась надвоє...
LUKE|23|46|І, скрикнувши голосом гучним, промовив Ісус: Отче, у руки Твої віддаю Свого духа! І це прорікши, Він духа віддав...
LUKE|23|47|Коли ж сотник побачив, що сталось, він Бога прославив, говорячи: Дійсно праведний був Чоловік Цей!
LUKE|23|48|І ввесь натовп, який зійшовсь на видовище це, як побачив, що сталось, бив у груди себе та вертався...
LUKE|23|49|Усі ж знайомі Його й ті жінки, що прийшли були з Ним із Галілеї, здалека стояли й дивились на це...
LUKE|23|50|І ось муж, на ім'я йому Йосип, що був радником синедріону, людина шановна і праведна,
LUKE|23|51|не пристав він до ради та чину їх, із Ариматеї, юдейського міста, що й сам сподівався Божого Царства,
LUKE|23|52|цей прийшов до Пилата, і тіла Ісусового став просити.
LUKE|23|53|І Йосип, знявши Його, обгорнув плащаницею, і поклав Його в гробі, що в скелі був висічений, і що в ньому ніколи ніхто не лежав.
LUKE|23|54|День той був Приготування, і наставала субота.
LUKE|23|55|А жінки, що прийшли були з Ним із Галілеї, ішли слідом, і вони бачили гроба, і як покладене тіло Його.
LUKE|23|56|Повернувшись, вони наготували пахощів і мира, а в суботу, за заповіддю, спочивали.
LUKE|24|1|А дня першого в тижні прийшли вони рано вранці до гробу, несучи наготовані пахощі,
LUKE|24|2|та й застали, що камінь від гробу відвалений був.
LUKE|24|3|А ввійшовши, вони не знайшли тіла Господа Ісуса.
LUKE|24|4|І сталось, як безрадні були вони в цім, ось два мужі в одежах блискучих з'явились при них.
LUKE|24|5|А коли налякались вони й посхиляли обличчя додолу, ті сказали до них: Чого ви шукаєте Живого між мертвими?
LUKE|24|6|Нема Його тут, бо воскрес! Пригадайте собі, як Він вам говорив, коли ще перебував в Галілеї.
LUKE|24|7|Він казав: Сину Людському треба бути виданому до рук грішних людей, і розп'ятому бути, і воскреснути третього дня.
LUKE|24|8|І згадали вони ті слова Його!
LUKE|24|9|А вернувшись від гробу, про все те сповістили Одинадцятьох та всіх інших.
LUKE|24|10|То були: Марія Магдалина, і Іванна, і Марія, мати Яковова, і інші з ними, і вони розповіли апостолам це.
LUKE|24|11|Та слова їхні здалися їм вигадкою, і не повірено їм.
LUKE|24|12|Петро ж устав та до гробу побіг, і, нахилившися, бачить лежать самі тільки покривала... І вернувсь він до себе, і дивувався, що сталось...
LUKE|24|13|І ото, двоє з них того ж дня йшли в село, на ім'я Еммаус, що від Єрусалиму лежало на стадій із шістдесят.
LUKE|24|14|І розмовляли вони між собою про все те, що сталося.
LUKE|24|15|І ото, як вони розмовляли, і розпитували один одного, підійшов Сам Ісус, і пішов разом із ними.
LUKE|24|16|Очі ж їхні були стримані, щоб Його не пізнали.
LUKE|24|17|І спитався Він їх: Що за речі такі, що про них між собою в дорозі міркуєте, і чого ви сумні?
LUKE|24|18|І озвався один, йому ймення Клеопа, та й промовив до Нього: Ти хіба тут у Єрусалимі єдиний захожий, що не знає, що сталося в нім цими днями?
LUKE|24|19|І спитався Він їх: Що таке? А вони розповіли Йому: Про Ісуса Назарянина, що Пророк був, могутній у ділі й у слові перед Богом і всім народом.
LUKE|24|20|Як первосвященики й наша старшина Його віддали на суд смертний, і Його розп'яли...
LUKE|24|21|А ми сподівались були, що Це Той, що має Ізраїля визволити. І до того, оце третій день вже сьогодні, як усе оте сталося...
LUKE|24|22|А дехто з наших жінок, що рано були коло гробу, нас здивували:
LUKE|24|23|вони тіла Його не знайшли, та й вернулися й оповідали, що бачили й з'явлення Анголів, які кажуть, що живий Він...
LUKE|24|24|І пішли дехто з наших до гробу, і знайшли так, як казали й жінки; та Його не побачили...
LUKE|24|25|Тоді Він сказав їм: О, безумні й запеклого серця, щоб повірити всьому, про що сповіщали Пророки!
LUKE|24|26|Чи ж Христові не це перетерпіти треба було, і ввійти в Свою славу?
LUKE|24|27|І Він почав від Мойсея, і від Пророків усіх, і виясняв їм зо всього Писання, що про Нього було.
LUKE|24|28|І наблизились вони до села, куди йшли. А Він удавав, ніби хоче йти далі.
LUKE|24|29|А вони не пускали Його й намовляли: Зостанься з нами, бо вже вечоріє, і кінчається день. І Він увійшов, щоб із ними побути.
LUKE|24|30|І ото, коли сів Він із ними до столу, то взяв хліб, поблагословив, і, ламаючи, їм подавав...
LUKE|24|31|Тоді очі відкрилися їм, і пізнали Його. Але Він став для них невидимий...
LUKE|24|32|І говорили вони один одному: Чи не палало нам серце обом, коли промовляв Він до нас по дорозі, і коли виясняв нам Писання?...
LUKE|24|33|І зараз устали вони, і повернулись до Єрусалиму, і знайшли там у зборі Одинадцятьох, і тих, що з ними були,
LUKE|24|34|які розповідали, що Господь дійсно воскрес, і з'явився був Симонові.
LUKE|24|35|А вони розповіли, що сталось було на дорозі, і як пізнали Його в ламанні хліба.
LUKE|24|36|І, як вони говорили оце, Сам Ісус став між ними, і промовив до них: Мир вам!
LUKE|24|37|А вони налякалися та перестрашились, і думали, що бачать духа.
LUKE|24|38|Він же промовив до них: Чого ви стривожились? І пощо ті думки до сердець ваших входять?
LUKE|24|39|Погляньте на руки Мої та на ноги Мої, це ж Я Сам! Доторкніться до Мене й дізнайтесь, бо не має дух тіла й костей, а Я, бачите, маю.
LUKE|24|40|І, промовивши це, показав Він їм руки та ноги.
LUKE|24|41|І, як ще не йняли вони віри з радощів та дивувались, Він сказав їм: Чи не маєте тут чогось їсти?
LUKE|24|42|Вони ж подали Йому кусника риби печеної та стільника медового.
LUKE|24|43|І, взявши, Він їв перед ними.
LUKE|24|44|І промовив до них: Це слова, що казав Я до вас, коли був іще з вами: Потрібно, щоб виконалось усе, що про Мене в Законі Мойсеєвім, та в Пророків, і в Псалмах написане.
LUKE|24|45|Тоді розум розкрив їм, щоб вони розуміли Писання.
LUKE|24|46|І сказав Він до них: Так написано є, і так потрібно було постраждати Христові, і воскреснути з мертвих дня третього,
LUKE|24|47|і щоб у Ймення Його проповідувалось покаяння, і прощення гріхів між народів усіх, від Єрусалиму почавши.
LUKE|24|48|А ви свідки того.
LUKE|24|49|І ось Я посилаю на вас обітницю Мого Отця; а ви позостаньтеся в місті, аж поки зодягнетесь силою з висоти.
LUKE|24|50|І Він вивів за місто їх аж до Віфанії; і, знявши руки Свої, поблагословив їх.
LUKE|24|51|І сталось, як Він благословляв їх, то зачав відступати від них, і на небо возноситись.
LUKE|24|52|А вони поклонились Йому, і повернулись до Єрусалиму з великою радістю.
LUKE|24|53|І постійно вони перебували в храмі, переславляючи й хвалячи Бога. Амінь.
