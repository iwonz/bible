GAL|1|1|Paulus apostolus non ab hominibus neque per hominem sed per Iesum Christum et Deum Patrem qui suscitavit eum a mortuis
GAL|1|2|et qui mecum sunt omnes fratres ecclesiis Galatiae
GAL|1|3|gratia vobis et pax a Deo Patre et Domino nostro Iesu Christo
GAL|1|4|qui dedit semet ipsum pro peccatis nostris ut eriperet nos de praesenti saeculo nequam secundum voluntatem Dei et Patris nostri
GAL|1|5|cui est gloria in saecula saeculorum amen
GAL|1|6|miror quod sic tam cito transferimini ab eo qui vos vocavit in gratiam Christi in aliud evangelium
GAL|1|7|quod non est aliud nisi sunt aliqui qui vos conturbant et volunt convertere evangelium Christi
GAL|1|8|sed licet nos aut angelus de caelo evangelizet vobis praeterquam quod evangelizavimus vobis anathema sit
GAL|1|9|sicut praediximus et nunc iterum dico si quis vobis evangelizaverit praeter id quod accepistis anathema sit
GAL|1|10|modo enim hominibus suadeo aut Deo aut quaero hominibus placere si adhuc hominibus placerem Christi servus non essem
GAL|1|11|notum enim vobis facio fratres evangelium quod evangelizatum est a me quia non est secundum hominem
GAL|1|12|neque enim ego ab homine accepi illud neque didici sed per revelationem Iesu Christi
GAL|1|13|audistis enim conversationem meam aliquando in iudaismo quoniam supra modum persequebar ecclesiam Dei et expugnabam illam
GAL|1|14|et proficiebam in iudaismo supra multos coetaneos in genere meo abundantius aemulator existens paternarum mearum traditionum
GAL|1|15|cum autem placuit ei qui me segregavit de utero matris meae et vocavit per gratiam suam
GAL|1|16|ut revelaret Filium suum in me ut evangelizarem illum in gentibus continuo non adquievi carni et sanguini
GAL|1|17|neque veni Hierosolyma ad antecessores meos apostolos sed abii in Arabiam et iterum reversus sum Damascum
GAL|1|18|deinde post annos tres veni Hierosolyma videre Petrum et mansi apud eum diebus quindecim
GAL|1|19|alium autem apostolorum vidi neminem nisi Iacobum fratrem Domini
GAL|1|20|quae autem scribo vobis ecce coram Deo quia non mentior
GAL|1|21|deinde veni in partes Syriae et Ciliciae
GAL|1|22|eram autem ignotus facie ecclesiis Iudaeae quae erant in Christo
GAL|1|23|tantum autem auditum habebant quoniam qui persequebatur nos aliquando nunc evangelizat fidem quam aliquando expugnabat
GAL|1|24|et in me clarificabant Deum
GAL|2|1|deinde post annos quattuordecim iterum ascendi Hierosolyma cum Barnaba adsumpto et Tito
GAL|2|2|ascendi autem secundum revelationem et contuli cum illis evangelium quod praedico in gentibus seorsum autem his qui videbantur ne forte in vacuum currerem aut cucurrissem
GAL|2|3|sed neque Titus qui mecum erat cum esset gentilis conpulsus est circumcidi
GAL|2|4|sed propter subintroductos falsos fratres qui subintroierunt explorare libertatem nostram quam habemus in Christo Iesu ut nos in servitutem redigerent
GAL|2|5|quibus neque ad horam cessimus subiectioni ut veritas evangelii permaneat apud vos
GAL|2|6|ab his autem qui videbantur esse aliquid quales aliquando fuerint nihil mea interest Deus personam hominis non accipit mihi enim qui videbantur nihil contulerunt
GAL|2|7|sed e contra cum vidissent quod creditum est mihi evangelium praeputii sicut Petro circumcisionis
GAL|2|8|qui enim operatus est Petro in apostolatum circumcisionis operatus est et mihi inter gentes
GAL|2|9|et cum cognovissent gratiam quae data est mihi Iacobus et Cephas et Iohannes qui videbantur columnae esse dextras dederunt mihi et Barnabae societatis ut nos in gentes ipsi autem in circumcisionem
GAL|2|10|tantum ut pauperum memores essemus quod etiam sollicitus fui hoc ipsum facere
GAL|2|11|cum autem venisset Cephas Antiochiam in faciem ei restiti quia reprehensibilis erat
GAL|2|12|prius enim quam venirent quidam ab Iacobo cum gentibus edebat cum autem venissent subtrahebat et segregabat se timens eos qui ex circumcisione erant
GAL|2|13|et simulationi eius consenserunt ceteri Iudaei ita ut et Barnabas duceretur ab eis in illa simulatione
GAL|2|14|sed cum vidissem quod non recte ambularent ad veritatem evangelii dixi Cephae coram omnibus si tu cum Iudaeus sis gentiliter et non iudaice vivis quomodo gentes cogis iudaizare
GAL|2|15|nos natura Iudaei et non ex gentibus peccatores
GAL|2|16|scientes autem quod non iustificatur homo ex operibus legis nisi per fidem Iesu Christi et nos in Christo Iesu credidimus ut iustificemur ex fide Christi et non ex operibus legis propter quod ex operibus legis non iustificabitur omnis caro
GAL|2|17|quod si quaerentes iustificari in Christo inventi sumus et ipsi peccatores numquid Christus peccati minister est absit
GAL|2|18|si enim quae destruxi haec iterum aedifico praevaricatorem me constituo
GAL|2|19|ego enim per legem legi mortuus sum ut Deo vivam Christo confixus sum cruci
GAL|2|20|vivo autem iam non ego vivit vero in me Christus quod autem nunc vivo in carne in fide vivo Filii Dei qui dilexit me et tradidit se ipsum pro me
GAL|2|21|non abicio gratiam Dei si enim per legem iustitia ergo Christus gratis mortuus est
GAL|3|1|o insensati Galatae quis vos fascinavit ante quorum oculos Iesus Christus proscriptus est crucifixus
GAL|3|2|hoc solum volo a vobis discere ex operibus legis Spiritum accepistis an ex auditu fidei
GAL|3|3|sic stulti estis cum Spiritu coeperitis nunc carne consummamini
GAL|3|4|tanta passi estis sine causa si tamen sine causa
GAL|3|5|qui ergo tribuit vobis Spiritum et operatur virtutes in vobis ex operibus legis an ex auditu fidei
GAL|3|6|sicut Abraham credidit Deo et reputatum est ei ad iustitiam
GAL|3|7|cognoscitis ergo quia qui ex fide sunt hii sunt filii Abrahae
GAL|3|8|providens autem scriptura quia ex fide iustificat gentes Deus praenuntiavit Abrahae quia benedicentur in te omnes gentes
GAL|3|9|igitur qui ex fide sunt benedicentur cum fideli Abraham
GAL|3|10|quicumque enim ex operibus legis sunt sub maledicto sunt scriptum est enim maledictus omnis qui non permanserit in omnibus quae scripta sunt in libro legis ut faciat ea
GAL|3|11|quoniam autem in lege nemo iustificatur apud Deum manifestum est quia iustus ex fide vivit
GAL|3|12|lex autem non est ex fide sed qui fecerit ea vivet in illis
GAL|3|13|Christus nos redemit de maledicto legis factus pro nobis maledictum quia scriptum est maledictus omnis qui pendet in ligno
GAL|3|14|ut in gentibus benedictio Abrahae fieret in Christo Iesu ut pollicitationem Spiritus accipiamus per fidem
GAL|3|15|fratres secundum hominem dico tamen hominis confirmatum testamentum nemo spernit aut superordinat
GAL|3|16|Abrahae dictae sunt promissiones et semini eius non dicit et seminibus quasi in multis sed quasi in uno et semini tuo qui est Christus
GAL|3|17|hoc autem dico testamentum confirmatum a Deo quae post quadringentos et triginta annos facta est lex non irritam facit ad evacuandam promissionem
GAL|3|18|nam si ex lege hereditas iam non ex repromissione Abrahae autem per promissionem donavit Deus
GAL|3|19|quid igitur lex propter transgressiones posita est donec veniret semen cui promiserat ordinata per angelos in manu mediatoris
GAL|3|20|mediator autem unius non est Deus autem unus est
GAL|3|21|lex ergo adversus promissa Dei absit si enim data esset lex quae posset vivificare vere ex lege esset iustitia
GAL|3|22|sed conclusit scriptura omnia sub peccato ut promissio ex fide Iesu Christi daretur credentibus
GAL|3|23|prius autem quam veniret fides sub lege custodiebamur conclusi in eam fidem quae revelanda erat
GAL|3|24|itaque lex pedagogus noster fuit in Christo ut ex fide iustificemur
GAL|3|25|at ubi venit fides iam non sumus sub pedagogo
GAL|3|26|omnes enim filii Dei estis per fidem in Christo Iesu
GAL|3|27|quicumque enim in Christo baptizati estis Christum induistis
GAL|3|28|non est Iudaeus neque Graecus non est servus neque liber non est masculus neque femina omnes enim vos unum estis in Christo Iesu
GAL|3|29|si autem vos Christi ergo Abrahae semen estis secundum promissionem heredes
GAL|4|1|dico autem quanto tempore heres parvulus est nihil differt servo cum sit dominus omnium
GAL|4|2|sed sub tutoribus est et actoribus usque ad praefinitum tempus a patre
GAL|4|3|ita et nos cum essemus parvuli sub elementis mundi eramus servientes
GAL|4|4|at ubi venit plenitudo temporis misit Deus Filium suum factum ex muliere factum sub lege
GAL|4|5|ut eos qui sub lege erant redimeret ut adoptionem filiorum reciperemus
GAL|4|6|quoniam autem estis filii misit Deus Spiritum Filii sui in corda nostra clamantem Abba Pater
GAL|4|7|itaque iam non es servus sed filius quod si filius et heres per Deum
GAL|4|8|sed tunc quidem ignorantes Deum his qui natura non sunt dii serviebatis
GAL|4|9|nunc autem cum cognoveritis Deum immo cogniti sitis a Deo quomodo convertimini iterum ad infirma et egena elementa quibus denuo servire vultis
GAL|4|10|dies observatis et menses et tempora et annos
GAL|4|11|timeo vos ne forte sine causa laboraverim in vobis
GAL|4|12|estote sicut et ego quia et ego sicut vos fratres obsecro vos nihil me laesistis
GAL|4|13|scitis autem quia per infirmitatem carnis evangelizavi vobis iam pridem
GAL|4|14|et temptationem vestram in carne mea non sprevistis neque respuistis sed sicut angelum Dei excepistis me sicut Christum Iesum
GAL|4|15|ubi est ergo beatitudo vestra testimonium enim perhibeo vobis quia si fieri posset oculos vestros eruissetis et dedissetis mihi
GAL|4|16|ergo inimicus vobis factus sum verum dicens vobis
GAL|4|17|aemulantur vos non bene sed excludere vos volunt ut illos aemulemini
GAL|4|18|bonum autem aemulamini in bono semper et non tantum cum praesens sum apud vos
GAL|4|19|filioli mei quos iterum parturio donec formetur Christus in vobis
GAL|4|20|vellem autem esse apud vos modo et mutare vocem meam quoniam confundor in vobis
GAL|4|21|dicite mihi qui sub lege vultis esse legem non legistis
GAL|4|22|scriptum est enim quoniam Abraham duos filios habuit unum de ancilla et unum de libera
GAL|4|23|sed qui de ancilla secundum carnem natus est qui autem de libera per repromissionem
GAL|4|24|quae sunt per allegoriam dicta haec enim sunt duo testamenta unum quidem a monte Sina in servitutem generans quae est Agar
GAL|4|25|Sina enim mons est in Arabia qui coniunctus est ei quae nunc est Hierusalem et servit cum filiis eius
GAL|4|26|illa autem quae sursum est Hierusalem libera est quae est mater nostra
GAL|4|27|scriptum est enim laetare sterilis quae non paris erumpe et exclama quae non parturis quia multi filii desertae magis quam eius quae habet virum
GAL|4|28|nos autem fratres secundum Isaac promissionis filii sumus
GAL|4|29|sed quomodo tunc qui secundum carnem natus fuerat persequebatur eum qui secundum spiritum ita et nunc
GAL|4|30|sed quid dicit scriptura eice ancillam et filium eius non enim heres erit filius ancillae cum filio liberae
GAL|4|31|itaque fratres non sumus ancillae filii sed liberae qua libertate nos Christus liberavit
GAL|5|1|state et nolite iterum iugo servitutis contineri
GAL|5|2|ecce ego Paulus dico vobis quoniam si circumcidamini Christus vobis nihil proderit
GAL|5|3|testificor autem rursum omni homini circumcidenti se quoniam debitor est universae legis faciendae
GAL|5|4|evacuati estis a Christo qui in lege iustificamini a gratia excidistis
GAL|5|5|nos enim spiritu ex fide spem iustitiae expectamus
GAL|5|6|nam in Christo Iesu neque circumcisio aliquid valet neque praeputium sed fides quae per caritatem operatur
GAL|5|7|currebatis bene quis vos inpedivit veritati non oboedire
GAL|5|8|persuasio non est ex eo qui vocat vos
GAL|5|9|modicum fermentum totam massam corrumpit
GAL|5|10|ego confido in vobis in Domino quod nihil aliud sapietis qui autem conturbat vos portabit iudicium quicumque est ille
GAL|5|11|ego autem fratres si circumcisionem adhuc praedico quid adhuc persecutionem patior ergo evacuatum est scandalum crucis
GAL|5|12|utinam et abscidantur qui vos conturbant
GAL|5|13|vos enim in libertatem vocati estis fratres tantum ne libertatem in occasionem detis carnis sed per caritatem servite invicem
GAL|5|14|omnis enim lex in uno sermone impletur diliges proximum tuum sicut te ipsum
GAL|5|15|quod si invicem mordetis et comeditis videte ne ab invicem consumamini
GAL|5|16|dico autem spiritu ambulate et desiderium carnis non perficietis
GAL|5|17|caro enim concupiscit adversus spiritum spiritus autem adversus carnem haec enim invicem adversantur ut non quaecumque vultis illa faciatis
GAL|5|18|quod si spiritu ducimini non estis sub lege
GAL|5|19|manifesta autem sunt opera carnis quae sunt fornicatio inmunditia luxuria
GAL|5|20|idolorum servitus veneficia inimicitiae contentiones aemulationes irae rixae dissensiones sectae
GAL|5|21|invidiae homicidia ebrietates comesationes et his similia quae praedico vobis sicut praedixi quoniam qui talia agunt regnum Dei non consequentur
GAL|5|22|fructus autem Spiritus est caritas gaudium pax longanimitas bonitas benignitas
GAL|5|23|fides modestia continentia adversus huiusmodi non est lex
GAL|5|24|qui autem sunt Christi carnem crucifixerunt cum vitiis et concupiscentiis
GAL|5|25|si vivimus spiritu spiritu et ambulemus
GAL|5|26|non efficiamur inanis gloriae cupidi invicem provocantes invicem invidentes
GAL|6|1|fratres et si praeoccupatus fuerit homo in aliquo delicto vos qui spiritales estis huiusmodi instruite in spiritu lenitatis considerans te ipsum ne et tu tempteris
GAL|6|2|alter alterius onera portate et sic adimplebitis legem Christi
GAL|6|3|nam si quis existimat se aliquid esse cum sit nihil ipse se seducit
GAL|6|4|opus autem suum probet unusquisque et sic in semet ipso tantum gloriam habebit et non in altero
GAL|6|5|unusquisque enim onus suum portabit
GAL|6|6|communicet autem is qui catecizatur verbum ei qui se catecizat in omnibus bonis
GAL|6|7|nolite errare Deus non inridetur
GAL|6|8|quae enim seminaverit homo haec et metet quoniam qui seminat in carne sua de carne et metet corruptionem qui autem seminat in spiritu de spiritu metet vitam aeternam
GAL|6|9|bonum autem facientes non deficiamus tempore enim suo metemus non deficientes
GAL|6|10|ergo dum tempus habemus operemur bonum ad omnes maxime autem ad domesticos fidei
GAL|6|11|videte qualibus litteris scripsi vobis mea manu
GAL|6|12|quicumque volunt placere in carne hii cogunt vos circumcidi tantum ut crucis Christi persecutionem non patiantur
GAL|6|13|neque enim qui circumciduntur legem custodiunt sed volunt vos circumcidi ut in carne vestra glorientur
GAL|6|14|mihi autem absit gloriari nisi in cruce Domini nostri Iesu Christi per quem mihi mundus crucifixus est et ego mundo
GAL|6|15|in Christo enim Iesu neque circumcisio aliquid valet neque praeputium sed nova creatura
GAL|6|16|et quicumque hanc regulam secuti fuerint pax super illos et misericordia et super Israhel Dei
GAL|6|17|de cetero nemo mihi molestus sit ego enim stigmata Iesu in corpore meo porto
GAL|6|18|gratia Domini nostri Iesu Christi cum spiritu vestro fratres amen
