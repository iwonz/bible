COL|1|1|Павел, волею Божиею Апостол Иисуса Христа, и Тимофей брат,
COL|1|2|находящимся в Колоссах святым и верным братиям во Христе Иисусе:
COL|1|3|благодать вам и мир от Бога Отца нашего и Господа Иисуса Христа. Благодарим Бога и Отца Господа нашего Иисуса Христа, всегда молясь о вас,
COL|1|4|услышав о вере вашей во Христа Иисуса и о любви ко всем святым,
COL|1|5|в надежде на уготованное вам на небесах, о чем вы прежде слышали в истинном слове благовествования,
COL|1|6|которое пребывает у вас, как и во всем мире, и приносит плод, и возрастает, как и между вами, с того дня, как вы услышали и познали благодать Божию в истине,
COL|1|7|как и научились от Епафраса, возлюбленного сотрудника нашего, верного для вас служителя Христова,
COL|1|8|который и известил нас о вашей любви в духе.
COL|1|9|Посему и мы с того дня, как [о сем] услышали, не перестаем молиться о вас и просить, чтобы вы исполнялись познанием воли Его, во всякой премудрости и разумении духовном,
COL|1|10|чтобы поступали достойно Бога, во всем угождая [Ему], принося плод во всяком деле благом и возрастая в познании Бога,
COL|1|11|укрепляясь всякою силою по могуществу славы Его, во всяком терпении и великодушии с радостью,
COL|1|12|благодаря Бога и Отца, призвавшего нас к участию в наследии святых во свете,
COL|1|13|избавившего нас от власти тьмы и введшего в Царство возлюбленного Сына Своего,
COL|1|14|в Котором мы имеем искупление Кровию Его и прощение грехов,
COL|1|15|Который есть образ Бога невидимого, рожденный прежде всякой твари;
COL|1|16|ибо Им создано все, что на небесах и что на земле, видимое и невидимое: престолы ли, господства ли, начальства ли, власти ли, – все Им и для Него создано;
COL|1|17|и Он есть прежде всего, и все Им стоит.
COL|1|18|И Он есть глава тела Церкви; Он – начаток, первенец из мертвых, дабы иметь Ему во всем первенство,
COL|1|19|ибо благоугодно было [Отцу], чтобы в Нем обитала всякая полнота,
COL|1|20|и чтобы посредством Его примирить с Собою все, умиротворив через Него, Кровию креста Его, и земное и небесное.
COL|1|21|И вас, бывших некогда отчужденными и врагами, по расположению к злым делам,
COL|1|22|ныне примирил в теле Плоти Его, смертью Его, [чтобы] представить вас святыми и непорочными и неповинными пред Собою,
COL|1|23|если только пребываете тверды и непоколебимы в вере и не отпадаете от надежды благовествования, которое вы слышали, которое возвещено всей твари поднебесной, которого я, Павел, сделался служителем.
COL|1|24|Ныне радуюсь в страданиях моих за вас и восполняю недостаток в плоти моей скорбей Христовых за Тело Его, которое есть Церковь,
COL|1|25|которой сделался я служителем по домостроительству Божию, вверенному мне для вас, [чтобы] исполнить слово Божие,
COL|1|26|тайну, сокрытую от веков и родов, ныне же открытую святым Его,
COL|1|27|Которым благоволил Бог показать, какое богатство славы в тайне сей для язычников, которая есть Христос в вас, упование славы,
COL|1|28|Которого мы проповедуем, вразумляя всякого человека и научая всякой премудрости, чтобы представить всякого человека совершенным во Христе Иисусе;
COL|1|29|для чего я и тружусь и подвизаюсь силою Его, действующею во мне могущественно.
COL|2|1|Желаю, чтобы вы знали, какой подвиг имею я ради вас и ради тех, которые в Лаодикии и Иераполе, и ради всех, кто не видел лица моего в плоти,
COL|2|2|дабы утешились сердца их, соединенные в любви для всякого богатства совершенного разумения, для познания тайны Бога и Отца и Христа,
COL|2|3|в Котором сокрыты все сокровища премудрости и ведения.
COL|2|4|Это говорю я для того, чтобы кто–нибудь не прельстил вас вкрадчивыми словами;
COL|2|5|ибо хотя я и отсутствую телом, но духом нахожусь с вами, радуясь и видя ваше благоустройство и твердость веры вашей во Христа.
COL|2|6|Посему, как вы приняли Христа Иисуса Господа, [так] и ходите в Нем,
COL|2|7|будучи укоренены и утверждены в Нем и укреплены в вере, как вы научены, преуспевая в ней с благодарением.
COL|2|8|Смотрите, братия, чтобы кто не увлек вас философиею и пустым обольщением, по преданию человеческому, по стихиям мира, а не по Христу;
COL|2|9|ибо в Нем обитает вся полнота Божества телесно,
COL|2|10|и вы имеете полноту в Нем, Который есть глава всякого начальства и власти.
COL|2|11|В Нем вы и обрезаны обрезанием нерукотворенным, совлечением греховного тела плоти, обрезанием Христовым;
COL|2|12|быв погребены с Ним в крещении, в Нем вы и совоскресли верою в силу Бога, Который воскресил Его из мертвых,
COL|2|13|и вас, которые были мертвы во грехах и в необрезании плоти вашей, оживил вместе с Ним, простив нам все грехи,
COL|2|14|истребив учением бывшее о нас рукописание, которое было против нас, и Он взял его от среды и пригвоздил ко кресту;
COL|2|15|отняв силы у начальств и властей, властно подверг их позору, восторжествовав над ними Собою.
COL|2|16|Итак никто да не осуждает вас за пищу, или питие, или за какой–нибудь праздник, или новомесячие, или субботу:
COL|2|17|это есть тень будущего, а тело – во Христе.
COL|2|18|Никто да не обольщает вас самовольным смиренномудрием и служением Ангелов, вторгаясь в то, чего не видел, безрассудно надмеваясь плотским своим умом
COL|2|19|и не держась главы, от которой все тело, составами и связями будучи соединяемо и скрепляемо, растет возрастом Божиим.
COL|2|20|Итак, если вы со Христом умерли для стихий мира, то для чего вы, как живущие в мире, держитесь постановлений:
COL|2|21|"не прикасайся", "не вкушай", "не дотрагивайся" –
COL|2|22|что все истлевает от употребления, – по заповедям и учению человеческому?
COL|2|23|Это имеет только вид мудрости в самовольном служении, смиренномудрии и изнурении тела, в некотором небрежении о насыщении плоти.
COL|3|1|Итак, если вы воскресли со Христом, то ищите горнего, где Христос сидит одесную Бога;
COL|3|2|о горнем помышляйте, а не о земном.
COL|3|3|Ибо вы умерли, и жизнь ваша сокрыта со Христом в Боге.
COL|3|4|Когда же явится Христос, жизнь ваша, тогда и вы явитесь с Ним во славе.
COL|3|5|Итак, умертвите земные члены ваши: блуд, нечистоту, страсть, злую похоть и любостяжание, которое есть идолослужение,
COL|3|6|за которые гнев Божий грядет на сынов противления,
COL|3|7|в которых и вы некогда обращались, когда жили между ними.
COL|3|8|А теперь вы отложите все: гнев, ярость, злобу, злоречие, сквернословие уст ваших;
COL|3|9|не говорите лжи друг другу, совлекшись ветхого человека с делами его
COL|3|10|и облекшись в нового, который обновляется в познании по образу Создавшего его,
COL|3|11|где нет ни Еллина, ни Иудея, ни обрезания, ни необрезания, варвара, Скифа, раба, свободного, но все и во всем Христос.
COL|3|12|Итак облекитесь, как избранные Божии, святые и возлюбленные, в милосердие, благость, смиренномудрие, кротость, долготерпение,
COL|3|13|снисходя друг другу и прощая взаимно, если кто на кого имеет жалобу: как Христос простил вас, так и вы.
COL|3|14|Более же всего [облекитесь] в любовь, которая есть совокупность совершенства.
COL|3|15|И да владычествует в сердцах ваших мир Божий, к которому вы и призваны в одном теле, и будьте дружелюбны.
COL|3|16|Слово Христово да вселяется в вас обильно, со всякою премудростью; научайте и вразумляйте друг друга псалмами, славословием и духовными песнями, во благодати воспевая в сердцах ваших Господу.
COL|3|17|И все, что вы делаете, словом или делом, все [делайте] во имя Господа Иисуса Христа, благодаря через Него Бога и Отца.
COL|3|18|Жены, повинуйтесь мужьям своим, как прилично в Господе.
COL|3|19|Мужья, любите своих жен и не будьте к ним суровы.
COL|3|20|Дети, будьте послушны родителям вашим во всем, ибо это благоугодно Господу.
COL|3|21|Отцы, не раздражайте детей ваших, дабы они не унывали.
COL|3|22|Рабы, во всем повинуйтесь господам вашим по плоти, не в глазах только служа [им], как человекоугодники, но в простоте сердца, боясь Бога.
COL|3|23|И все, что делаете, делайте от души, как для Господа, а не для человеков,
COL|3|24|зная, что в воздаяние от Господа получите наследие, ибо вы служите Господу Христу.
COL|3|25|А кто неправо поступит, тот получит по своей неправде, [у Него] нет лицеприятия.
COL|4|1|Господа, оказывайте рабам должное и справедливое, зная, что и вы имеете Господа на небесах.
COL|4|2|Будьте постоянны в молитве, бодрствуя в ней с благодарением.
COL|4|3|Молитесь также и о нас, чтобы Бог отверз нам дверь для слова, возвещать тайну Христову, за которую я и в узах,
COL|4|4|дабы я открыл ее, как должно мне возвещать.
COL|4|5|Со внешними обходитесь благоразумно, пользуясь временем.
COL|4|6|Слово ваше [да будет] всегда с благодатию, приправлено солью, дабы вы знали, как отвечать каждому.
COL|4|7|О мне все скажет вам Тихик, возлюбленный брат и верный служитель и сотрудник в Господе,
COL|4|8|которого я для того послал к вам, чтобы он узнал о ваших [обстоятельствах] и утешил сердца ваши,
COL|4|9|с Онисимом, верным и возлюбленным братом нашим, который от вас. Они расскажут вам о всем здешнем.
COL|4|10|Приветствует вас Аристарх, заключенный вместе со мною, и Марк, племянник Варнавы – о котором вы получили приказания: если придет к вам, примите его, –
COL|4|11|также Иисус, прозываемый Иустом, оба из обрезанных. Они – единственные сотрудники для Царствия Божия, бывшие мне отрадою.
COL|4|12|Приветствует вас Епафрас ваш, раб Иисуса Христа, всегда подвизающийся за вас в молитвах, чтобы вы пребыли совершенны и исполнены всем, что угодно Богу.
COL|4|13|Свидетельствую о нем, что он имеет великую ревность и заботу о вас и о находящихся в Лаодикии и Иераполе.
COL|4|14|Приветствует вас Лука, врач возлюбленный, и Димас.
COL|4|15|Приветствуйте братьев в Лаодикии, и Нимфана, и домашнюю церковь его.
COL|4|16|Когда это послание прочитано будет у вас, то распорядитесь, чтобы оно было прочитано и в Лаодикийской церкви; а то, которое из Лаодикии, прочитайте и вы.
COL|4|17|Скажите Архиппу: смотри, чтобы тебе исполнить служение, которое ты принял в Господе.
COL|4|18|Приветствие моею рукою, Павловою. Помните мои узы. Благодать со всеми вами. Аминь.
