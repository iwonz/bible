GEN|1|1|起初，上帝创造天地。
GEN|1|2|地是空虚混沌，深渊上面一片黑暗；上帝的灵 运行在水面上。
GEN|1|3|上帝说：“要有光”，就有了光。
GEN|1|4|上帝看光是好的，于是上帝就把光和暗分开。
GEN|1|5|上帝称光为“昼”，称暗为“夜”。有晚上，有早晨，这是第一日。
GEN|1|6|上帝说：“众水之间要有穹苍，把水和水分开。”
GEN|1|7|上帝就造了穹苍，把穹苍以下的水和穹苍以上的水分开。事就这样成了。
GEN|1|8|上帝称穹苍为“天”。有晚上，有早晨，这是第二日。
GEN|1|9|上帝说：“天下面的水要聚集在一处，使干地露出来。”事就这样成了。
GEN|1|10|上帝称干地为“地”，称聚集在一起的水为“海”。上帝看为好的。
GEN|1|11|上帝说：“地要长出植物，就是含种子的五谷菜蔬，和会结果子、果子里有种子的树，在地上各从其类。”事就这样成了。
GEN|1|12|于是地长出了植物：含种子的五谷菜蔬，各从其类；会结果子、果子里有种子的树，各从其类。上帝看为好的。
GEN|1|13|有晚上，有早晨，这是第三日。
GEN|1|14|上帝说：“天上要有光体来分昼夜，让它们作记号，定季节、日子、年份，
GEN|1|15|它们要在天空发光，照在地上。”事就这样成了。
GEN|1|16|于是上帝造了两个大光体，大的管昼，小的管夜，又造了星辰。
GEN|1|17|上帝把这些光体摆列在天空，照在地上，
GEN|1|18|管理昼夜，分别光暗。上帝看为好的。
GEN|1|19|有晚上，有早晨，这是第四日。
GEN|1|20|上帝说：“水要滋生众多有生命之物；要有鸟飞在地面以上，天空之中。”
GEN|1|21|上帝就创造了大鱼和在水里滋生的各样活动的生物，各从其类，以及各样有翅膀的鸟，各从其类。上帝看为好的。
GEN|1|22|上帝就赐福给这一切，说：“要繁殖增多，充满在海的水里；飞鸟也要在地上增多。”
GEN|1|23|有晚上，有早晨，这是第五日。
GEN|1|24|上帝说：“地要生出有生命之物，各从其类，就是牲畜、爬行动物、地上的走兽，各从其类。”事就这样成了。
GEN|1|25|于是上帝造了地上的走兽，各从其类；牲畜，各从其类；和地上一切的爬行动物，各从其类。上帝看为好的。
GEN|1|26|上帝说：“我们要照着我们的形像，按着我们的样式造人，使他们管理海里的鱼、天空的鸟、地上的牲畜和全地，以及地上爬的一切爬行动物。”
GEN|1|27|上帝就照着他的形像创造人，照着上帝的形像创造他们 ；他创造了他们，有男有女。
GEN|1|28|上帝赐福给他们，上帝对他们说：“要生养众多，遍满这地，治理它；要管理海里的鱼、天空的鸟和地上各样活动的生物。”
GEN|1|29|上帝说：“看哪，我把全地一切含种子的五谷菜蔬和一切会结果子、果子里有种子的树，都赐给你们；这些都可作食物。
GEN|1|30|至于地上一切的走兽、天空一切的飞鸟，并一切在地上爬行的，有生命的动物，我把绿色植物赐给它们作食物。”事就这样成了。
GEN|1|31|上帝看一切所造的，看哪，都非常好。有晚上，有早晨，这是第六日。
GEN|2|1|天和地，以及万象都完成了。
GEN|2|2|到第七日，上帝已经完成了造物之工，就在第七日安息了，歇了他所做一切的工。
GEN|2|3|上帝赐福给第七日，将它分别为圣，因为在这日，上帝安息了，歇了他所做一切创造的工。
GEN|2|4|这就是天地创造的来历。 在耶和华上帝造地和天的时候，
GEN|2|5|地上还没有田野的草木，田间的菜蔬还没有长出来，因为耶和华上帝还没有降雨在地上，也没有人耕种土地。
GEN|2|6|但是，有雾气从地上腾，滋润整个土地的表面。
GEN|2|7|耶和华上帝用地上的尘土造人，将生命之气吹进他的鼻孔，这人就成了有灵的活人 。
GEN|2|8|耶和华上帝在东方的 伊甸 栽了一个园子，把所造的人安置在那里。
GEN|2|9|耶和华上帝使各样的树从土地里长出来，可以悦人的眼目，好作食物。园子当中有生命树和知善恶的树 。
GEN|2|10|有一条河从 伊甸 流出来，滋润那园子，从那里分成四个源头：
GEN|2|11|第一条名叫 比逊 ，它环绕 哈腓拉 全地，在那里有金子。
GEN|2|12|那地的金子很好，在那里也有珍珠 和红玛瑙。
GEN|2|13|第二条河名叫 基训 ，它环绕 古实 全地。
GEN|2|14|第三条河名叫 底格里斯 ，它流到 亚述 的东边。第四条河就是 幼发拉底 。
GEN|2|15|耶和华上帝把那人安置在 伊甸园 ，让他耕耘看管。
GEN|2|16|耶和华上帝吩咐那人说：“园中各样树上所出的，你可以随意吃，
GEN|2|17|只是知善恶的树所出的，你不可吃，因为你吃它的日子必定死！”
GEN|2|18|耶和华上帝说：“那人单独一个不好，我要为他造一个配偶帮助他。”
GEN|2|19|耶和华上帝用泥土造了野地各样的走兽和天空各样的飞鸟，都带到那人面前，看他叫什么。那人怎样叫各样的动物，那就是它的名字。
GEN|2|20|那人就给一切牲畜、天空的飞鸟和野地各样的走兽都起了名。只是 亚当 没有找到配偶帮助他。
GEN|2|21|耶和华上帝使他沉睡，他就睡了；于是取下他的一根肋骨，又在原处把肉合起来。
GEN|2|22|耶和华上帝就用那人身上所取的肋骨造了一个女人，带她到那人面前。
GEN|2|23|那人说： “这正是我骨中的骨， 肉中的肉， 可以称她为女人， 因为她是从男人身上取出来的。”
GEN|2|24|因此，人要离开父母，与妻子结合，二人成为一体。
GEN|2|25|当时夫妻二人赤身露体，并不觉得羞耻。
GEN|3|1|耶和华上帝所造的，惟有蛇比田野一切的走兽更狡猾。蛇对女人说：“上帝岂是真说，你们不可吃园中任何树上所出的吗？”
GEN|3|2|女人对蛇说：“园中树上的果子，我们都可以吃；
GEN|3|3|只是园子中间那棵树的果子，上帝曾说：‘你们不可吃，也不可摸，免得你们死。’”
GEN|3|4|蛇对女人说：“你们不一定死；
GEN|3|5|因为上帝知道，你们吃的日子眼睛就开了，你们就像上帝一样知道善恶。”
GEN|3|6|于是女人见那棵树好作食物，又悦人的眼目，那树令人喜爱，能使人有智慧，她就摘下果子吃了，又给了与她一起的丈夫，他也吃了。
GEN|3|7|他们二人的眼睛就开了，知道自己赤身露体，就编织无花果树的叶子，为自己做成裙子。
GEN|3|8|天起了凉风，那人和他妻子听见耶和华上帝在园中来回行走的声音，就藏在园里的树木中，躲避耶和华上帝的面。
GEN|3|9|耶和华上帝呼唤那人，对他说：“你在哪里？”
GEN|3|10|他说：“我在园中听见你的声音，我就害怕；因为我赤身露体，我就藏了起来。”
GEN|3|11|耶和华上帝说：“谁告诉你，你是赤身露体呢？莫非你吃了那树上所出的，就是我吩咐你不可吃的吗？”
GEN|3|12|那人说：“你赐给我、与我一起的女人，是她把那树上所出的给我，我就吃了。”
GEN|3|13|耶和华上帝对女人说：“你怎么会做这种事呢？”女人说：“那蛇引诱我，我就吃了。”
GEN|3|14|耶和华上帝对蛇说： “你既做了这事，就必受诅咒， 比一切的牲畜和野兽更重。 你必用肚子行走， 终生吃土。
GEN|3|15|我要使你和女人彼此为仇， 你的后裔和女人的后裔也彼此为仇。 他要伤你的头， 你要伤他的脚跟。 ”
GEN|3|16|又对女人说： “我必多多加增你怀胎的痛苦， 你生儿女时必多受痛苦。 你必恋慕你丈夫， 他必管辖你。”
GEN|3|17|又对 亚当 说： “你既听从你妻子的话， 吃了那树上所出的， 就是我吩咐你不可吃的， 土地必因你的缘故受诅咒； 你必终生劳苦才能从土地得吃的。
GEN|3|18|土地必给你长出荆棘和蒺藜来； 你也要吃田间的五谷菜蔬。
GEN|3|19|你必汗流满面才有食物可吃， 直到你归了土地， 因为你是从土地而出的。 你本是尘土，仍要归回尘土。”
GEN|3|20|那人给他妻子起名叫 夏娃 ，因为她是众生之母 。
GEN|3|21|耶和华上帝用兽皮做衣服给 亚当 和他的妻子穿。
GEN|3|22|耶和华上帝说：“看哪，那人已经像我们中间的一个，知道善恶，现在恐怕他又伸手摘生命树所出的来吃，就永远活着。”
GEN|3|23|耶和华上帝就驱逐他出 伊甸园 ，使他耕种土地，他原是从土地里被取出来的。
GEN|3|24|耶和华上帝把那人赶出去，就在 伊甸园 东边安设基路伯和发出火焰转动的剑，把守生命树的道路。
GEN|4|1|那人和他妻子 夏娃 同房， 夏娃 就怀孕，生了 该隐 ，她说：“我靠耶和华得了一个男的。”
GEN|4|2|她又生了 该隐 的弟弟 亚伯 。 亚伯 是牧羊的； 该隐 是耕地的。
GEN|4|3|过了一些日子， 该隐 拿地里的出产为供物献给耶和华；
GEN|4|4|亚伯 也把他羊群中头生的和羊的脂肪献上。耶和华看中了 亚伯 和他的供物，
GEN|4|5|却看不中 该隐 和他的供物。 该隐 就非常生气，沉下脸来。
GEN|4|6|耶和华对 该隐 说：“你为什么生气呢？你为什么沉下脸来呢？
GEN|4|7|你若做得对，岂不仰起头来吗？你若做得不对，罪就伏在门前。它想要控制你，你却要制伏它。”
GEN|4|8|该隐 与他弟弟 亚伯 说话 。 二人正在田间时， 该隐 起来攻击他弟弟 亚伯 ，把他杀了。
GEN|4|9|耶和华对 该隐 说：“你弟弟 亚伯 在哪里？”他说：“我不知道！我岂是看守我弟弟的吗？”
GEN|4|10|耶和华说：“你做了什么事呢？你弟弟血的声音从地里向我哀号。
GEN|4|11|现在你必从这地受诅咒，这地开了口，从你手里接受你弟弟的血。
GEN|4|12|你耕种土地，它不再给你效力；你必流离飘荡在地上。”
GEN|4|13|该隐 对耶和华说：“我的惩罚太重，过于我所能承当的。
GEN|4|14|看哪，今日你赶我离开这块土地，不能见你的面；我必流离飘荡在地上，凡遇见我的必杀我。”
GEN|4|15|耶和华对他说：“既然如此 ，凡杀 该隐 的，必遭报七倍。”耶和华就给 该隐 立一个记号，免得人遇见他就杀他。
GEN|4|16|于是 该隐 离开了耶和华的面，去住在 伊甸 东边 挪得 之地。
GEN|4|17|该隐 与妻子同房，她就怀孕，生了 以诺 。 该隐 建造一座城，就照他儿子的名字称那城为 以诺 。
GEN|4|18|以诺 生 以拿 ， 以拿 生 米户雅利 ， 米户雅利 生 玛土撒利 ， 玛土撒利 生 拉麦 。
GEN|4|19|拉麦 娶了两个妻子：一个名叫 亚大 ，一个名叫 洗拉 。
GEN|4|20|亚大 生 雅八 ； 雅八 是住帐棚、牧养牲畜之人的祖师。
GEN|4|21|雅八 的兄弟名叫 犹八 ；他是所有弹琴吹箫之人的祖师。
GEN|4|22|洗拉 又生了 土八．该隐 ；他是打造各样铜器铁器的工匠。 土八．该隐 的妹妹是 拿玛 。
GEN|4|23|拉麦 对他两个妻子说： 亚大 、 洗拉 啊，听我的声音； 拉麦 的妻子啊，侧耳听我的言语： 大人伤我，我把他杀了； 小孩损我，我把他害了 。
GEN|4|24|若杀 该隐 ，遭报七倍， 杀 拉麦 的，必遭报七十七倍。
GEN|4|25|亚当 又与妻子同房，她就生了一个儿子，给他起名叫 塞特 ，说：“上帝给我立了另一个子嗣代替 亚伯 ，因为 该隐 杀了他。”
GEN|4|26|塞特 也生了一个儿子，起名叫 以挪士 。那时候，人开始求告耶和华的名。
GEN|5|1|这是 亚当 后代的家谱。当上帝造人的日子，他照着自己的样式造人。
GEN|5|2|他造男造女。在他们被造的日子，上帝赐福给他们，称他们为人。
GEN|5|3|亚当 活到一百三十岁，生了一个儿子，形像样式和自己相似，就给他起名叫 塞特 。
GEN|5|4|亚当 生 塞特 之后，又活了八百年，并且生儿育女。
GEN|5|5|亚当 共活了九百三十年，就死了。
GEN|5|6|塞特 活到一百零五岁，生了 以挪士 。
GEN|5|7|塞特 生 以挪士 之后，又活了八百零七年，并且生儿育女。
GEN|5|8|塞特 共活了九百一十二年，就死了。
GEN|5|9|以挪士 活到九十岁，生了 该南 。
GEN|5|10|以挪士 生 该南 之后，又活了八百一十五年，并且生儿育女。
GEN|5|11|以挪士 共活了九百零五年，就死了。
GEN|5|12|该南 活到七十岁，生了 玛勒列 。
GEN|5|13|该南 生 玛勒列 之后，又活了八百四十年，并且生儿育女。
GEN|5|14|该南 共活了九百一十年，就死了。
GEN|5|15|玛勒列 活到六十五岁，生了 雅列 。
GEN|5|16|玛勒列 生 雅列 之后，又活了八百三十年，并且生儿育女。
GEN|5|17|玛勒列 共活了八百九十五年，就死了。
GEN|5|18|雅列 活到一百六十二岁，生了 以诺 。
GEN|5|19|雅列 生 以诺 之后，又活了八百年，并且生儿育女。
GEN|5|20|雅列 共活了九百六十二年，就死了。
GEN|5|21|以诺 活到六十五岁，生了 玛土撒拉 。
GEN|5|22|以诺 生 玛土撒拉 之后，与上帝同行三百年，并且生儿育女。
GEN|5|23|以诺 共活了三百六十五年。
GEN|5|24|以诺 与上帝同行，上帝把他接去，他就不在了。
GEN|5|25|玛土撒拉 活到一百八十七岁，生了 拉麦 。
GEN|5|26|玛土撒拉 生 拉麦 之后，又活了七百八十二年，并且生儿育女。
GEN|5|27|玛土撒拉 共活了九百六十九年，就死了。
GEN|5|28|拉麦 活到一百八十二岁，生了一个儿子，
GEN|5|29|给他起名叫 挪亚 ，说：“在耶和华所诅咒的地上，这个儿子必使我们从工作和手中的劳苦得到安慰。”
GEN|5|30|拉麦 生 挪亚 之后，又活了五百九十五年，并且生儿育女。
GEN|5|31|拉麦 共活了七百七十七年，就死了。
GEN|5|32|挪亚 活到五百岁，生了 闪 、 含 和 雅弗 。
GEN|6|1|当人开始在地面上增多、又生女儿的时候，
GEN|6|2|上帝的儿子们看见人的女子美貌，就随意挑选，娶来为妻。
GEN|6|3|耶和华说：“人既属乎血气，我的灵就不永远住在他里面；然而他的年岁还可到一百二十年。”
GEN|6|4|那时候有巨人在地上，后来也有；上帝的儿子们和人的女子们交合，生了孩子。那些人就是古代的勇士，有名的人物。
GEN|6|5|耶和华见人在地上罪大恶极，终日心里所想的尽都是恶事，
GEN|6|6|耶和华就因造人在地上感到遗憾，心中忧伤。
GEN|6|7|耶和华说：“我要把所造的人和走兽，爬行动物，以及天空的飞鸟，都从地面上除灭，因为我造了他们感到遗憾。”
GEN|6|8|只有 挪亚 在耶和华眼前蒙恩。
GEN|6|9|这是 挪亚 的后代。 挪亚 是个义人，在他的世代中是个完全人。 挪亚 与上帝同行。
GEN|6|10|挪亚 生了三个儿子，就是 闪 、 含 和 雅弗 。
GEN|6|11|这地在上帝面前败坏了，地上充满了暴力。
GEN|6|12|上帝观看这地，看哪，它败坏了，因为凡血肉之躯在地上的行为都败坏了。
GEN|6|13|上帝对 挪亚 说：“在我面前，凡血肉之躯的结局已经临到，因着他们，地上充满了暴力。看哪，我要把他们和这地一起毁灭。
GEN|6|14|你要为自己用歌斐木造一艘方舟，并在方舟内造房间，内外都要抹上沥青。
GEN|6|15|方舟的造法是这样：要长三百肘，宽五十肘，高三十肘。
GEN|6|16|方舟上面要造天窗，向上一肘。方舟的门要开在旁边。方舟要分上、中、下三层。
GEN|6|17|看哪，我要使洪水泛滥在地上，毁灭天下凡有生命气息的血肉之躯，地上的一切都要灭亡。
GEN|6|18|但我要与你立约；你同你的儿子、妻子和媳妇都要进入方舟。
GEN|6|19|凡有血肉的动物，每样一对，一公一母，你要带进方舟，好跟你一起保全生命。
GEN|6|20|飞鸟各从其类，牲畜各从其类，地上的爬行动物各从其类，每样一对，都要到你那里，好保全生命。
GEN|6|21|你要拿各样可吃的食物，储存在你那里，作你和它们的粮食。”
GEN|6|22|挪亚 就去做了；凡上帝吩咐他的，他都照样去做。
GEN|7|1|耶和华对 挪亚 说：“你和你的全家都要进入方舟，因为在这世代中，我看你在我面前是个义人。
GEN|7|2|凡洁净的牲畜，你要各取七公七母；不洁净的牲畜，你要各取一公一母；
GEN|7|3|天空的飞鸟也要各取七公七母，为了要留种，活在全地面上。
GEN|7|4|因为再过七天，我要降雨在地上四十昼夜，把我所造的一切生物从地面上除灭。”
GEN|7|5|挪亚 就遵照耶和华吩咐他的去做。
GEN|7|6|当洪水 在地上泛滥的时候， 挪亚 已六百岁。
GEN|7|7|挪亚 同他的儿子、妻子和媳妇都进入方舟，躲避洪水。
GEN|7|8|洁净的牲畜和不洁净的牲畜，飞鸟及所有爬行在土地上的，
GEN|7|9|都一对一对，有公有母，到 挪亚 那里，进入方舟，正如上帝所吩咐 挪亚 的。
GEN|7|10|过了七天，洪水泛滥在地上。
GEN|7|11|挪亚 六百岁那一年的二月十七日，就在那一天，大深渊的泉源都裂开，天上的窗户也敞开了，
GEN|7|12|四十昼夜有大雨降在地上。
GEN|7|13|正在那日， 挪亚 和他的儿子 闪 、 含 、 雅弗 ，以及 挪亚 的妻子和三个媳妇，都一同进入方舟。
GEN|7|14|他们和一切走兽，各从其类；一切牲畜，各从其类；地上爬的一切爬行动物，各从其类；一切的鸟，就是一切有翅膀的飞禽，各从其类；
GEN|7|15|凡有生命气息的血肉之躯，都一对一对到 挪亚 那里，进入方舟。
GEN|7|16|凡有血肉的，都一公一母进入方舟，正如上帝所吩咐 挪亚 的。耶和华就把他关在方舟里。
GEN|7|17|洪水在地上泛滥四十天，水往上涨，使方舟浮起，方舟就从地上漂起来。
GEN|7|18|水势汹涌，在地上大大上涨，方舟在水面上漂荡。
GEN|7|19|水势在地上极其浩大，普天下所有的高山都淹没了。
GEN|7|20|水势汹涌，比山高出十五肘 ，山岭都淹没了。
GEN|7|21|凡有血肉在地上行动的，就是飞鸟、牲畜、走兽和地上成群的群聚动物，以及所有的人，都死了。
GEN|7|22|在干地上凡鼻孔里有生命气息的都死了。
GEN|7|23|耶和华除灭了地面上各类的生物，包括人和牲畜、爬行动物，以及天空的飞鸟；他们就都从地上除灭了，只剩下 挪亚 和那些与他同在方舟里的。
GEN|7|24|水势汹涌，在地上共一百五十天。
GEN|8|1|上帝记念 挪亚 和 挪亚 方舟里的一切走兽牲畜。上帝使风吹地，水势渐落。
GEN|8|2|深渊的泉源和天上的窗户都关闭了，雨不再从天降下。
GEN|8|3|水从地上逐渐消退。过了一百五十天，水就退了。
GEN|8|4|七月十七日，方舟停在 亚拉腊山 上。
GEN|8|5|水继续退去，直到十月；十月初一，山顶都露出来了。
GEN|8|6|过了四十天， 挪亚 打开他所造的方舟的窗户，
GEN|8|7|放出一只乌鸦。那乌鸦飞来飞去，直到地上的水都干了。
GEN|8|8|他又从他那里放出一只鸽子，要看水从地面上退了没有。
GEN|8|9|但全地面都是水，鸽子找不到落脚之地，就回到方舟 挪亚 那里。 挪亚 伸手接了鸽子，把它带进方舟。
GEN|8|10|挪亚 又另外等了七天，再把鸽子从方舟放出去。
GEN|8|11|到了晚上，鸽子回到他那里，看哪，嘴里有一片刚啄下来的橄榄叶， 挪亚 就知道水已经从地上退了。
GEN|8|12|他又另外等了七天，再放出鸽子，这次鸽子不再回到他那里了。
GEN|8|13|当 挪亚 六百零一岁，正月初一的时候，地上的水都干了。 挪亚 打开方舟的盖观看，看哪，地面干了。
GEN|8|14|到了二月二十七日，地就都干了。
GEN|8|15|上帝对 挪亚 说：
GEN|8|16|“你同你的妻子、儿子、媳妇都要出方舟。
GEN|8|17|凡与你一起有血肉的生物，就是飞鸟、牲畜和地上爬的一切爬行动物，都要带出来。 它们要在地上滋生，繁殖增多。”
GEN|8|18|于是 挪亚 同他的儿子、妻子、媳妇都出来了。
GEN|8|19|一切走兽、爬行动物和飞鸟，地上所有的动物，各从其类，也都出了方舟。
GEN|8|20|挪亚 为耶和华筑了一座坛，拿各种洁净的牲畜和各种洁净的飞鸟，献在坛上为燔祭。
GEN|8|21|耶和华闻了那馨香之气，耶和华心里说：“我不再因人的缘故诅咒土地，因为人从幼年就心里怀着恶念；我也不再照我曾做的毁灭一切生物了。
GEN|8|22|地还存在的时候，撒种、收割、寒暑、冬夏、昼夜都永不止息。”
GEN|9|1|上帝赐福给 挪亚 和他的儿子，对他们说：“你们要生养众多，遍满这地。
GEN|9|2|地上一切的走兽、天空一切的飞鸟、所有爬行在土地上的和海里一切的鱼都必怕你们，畏惧你们，它们都要交在你们手里。
GEN|9|3|凡活的动物都可作你们的食物。这一切我都赐给你们，如同绿色的菜蔬一样。
GEN|9|4|只是带着生命的肉，就是带着血的，你们不可吃。
GEN|9|5|流你们血、害你们命的，我必向他追讨；我要向一切走兽追讨，向人和向人的弟兄追讨人命。
GEN|9|6|凡流人血的，他的血也必被人所流，因为上帝造人，是照自己的形像造的。
GEN|9|7|你们要生养众多，在地上繁衍昌盛。”
GEN|9|8|上帝对 挪亚 和同他一起的儿子说：
GEN|9|9|“看哪，我要与你们和你们后裔立我的约，
GEN|9|10|包括和你们一起所有的生物，就是飞鸟、牲畜、地上一切的走兽，凡从方舟里出来地上一切的生物。
GEN|9|11|我与你们立我的约：凡有血肉的，不再被洪水灭绝，也不再有洪水毁坏这地了。”
GEN|9|12|上帝说：“这是我与你们，以及和你们一起的一切生物所立之约的记号，直到万代：
GEN|9|13|我把彩虹放在云中，这就是我与地立约的记号了。
GEN|9|14|我使云遮地的时候，会有彩虹出现在云中，
GEN|9|15|我就记念我与你们，以及各样有血肉的生物所立的约：不再有洪水泛滥去毁灭一切有血肉的了。
GEN|9|16|彩虹出现在云中，我看见了，就要记念上帝与地上一切有血肉的生物所立的永约。”
GEN|9|17|上帝对 挪亚 说：“这就是我与地上一切有血肉的立约的记号。”
GEN|9|18|挪亚 的儿子，从方舟出来的，有 闪 、 含 和 雅弗 。 含 是 迦南 的父亲。
GEN|9|19|这是 挪亚 的三个儿子，他们的后裔散布全地。
GEN|9|20|挪亚 是农夫，是他开始栽葡萄园的。
GEN|9|21|他喝了一些酒就醉了，在他的帐棚里赤着身子。
GEN|9|22|迦南 的父亲 含 看见他父亲赤身，就到外面告诉他的两个兄弟。
GEN|9|23|于是 闪 和 雅弗 拿了外衣搭在二人肩上，倒退着进去，遮盖父亲的赤身；他们背着脸，看不见父亲的赤身。
GEN|9|24|挪亚 酒醒以后，知道小儿子向他所做的事，
GEN|9|25|就说： “ 迦南 当受诅咒， 必给他弟兄作奴仆的奴仆。”
GEN|9|26|又说： “耶和华— 闪 的上帝是应当称颂的！ 愿 迦南 作 闪 的奴仆。
GEN|9|27|愿上帝使 雅弗 扩张， 愿他住在 闪 的帐棚里； 愿 迦南 作他的奴仆。”
GEN|9|28|洪水以后， 挪亚 又活了三百五十年。
GEN|9|29|挪亚 共活了九百五十年，就死了。
GEN|10|1|这是 挪亚 的儿子 闪 、 含 、 雅弗 的后代。洪水以后，他们都生了儿子。
GEN|10|2|雅弗 的儿子是 歌篾 、 玛各 、 玛代 、 雅完 、 土巴 、 米设 、 提拉 。
GEN|10|3|歌篾 的儿子是 亚实基拿 、 利法 、 陀迦玛 。
GEN|10|4|雅完 的儿子是 以利沙 、 他施 、 基提 、 罗单 人 。
GEN|10|5|从这些人中有沿海国家的人散居各处，有自己的土地，各有各的语言、宗族、国家。
GEN|10|6|含 的儿子是 古实 、 麦西 、 弗 、 迦南 。
GEN|10|7|古实 的儿子是 西巴 、 哈腓拉 、 撒弗他 、 拉玛 、 撒弗提迦 。 拉玛 的儿子是 示巴 、 底但 。
GEN|10|8|古实 又生 宁录 ，他是地上第一个勇士。
GEN|10|9|他在耶和华面前是个英勇的猎人，所以有话说：“像 宁录 在耶和华面前是个英勇的猎人。”
GEN|10|10|他王国的开始是在 巴别 、 以力 、 亚甲 、 甲尼 ，都在 示拿 地。
GEN|10|11|他从那地出来往 亚述 去，建造了 尼尼微 、 利河伯 、 迦拉 ，
GEN|10|12|以及 尼尼微 和 迦拉 之间的 利鲜 ，那是座大城。
GEN|10|13|麦西 生 路低 人、 亚拿米 人、 利哈比 人、 拿弗土希 人、
GEN|10|14|帕斯鲁细 人、 迦斯路希 人、 迦斐托 人； 非利士 人是从 迦斐托 人 出来的。
GEN|10|15|迦南 生了长子 西顿 ，又生 赫
GEN|10|16|和 耶布斯 人、 亚摩利 人、 革迦撒 人、
GEN|10|17|希未 人、 亚基 人、 西尼 人、
GEN|10|18|亚瓦底 人、 洗玛利 人、 哈马 人，后来 迦南 的家族散开了。
GEN|10|19|迦南 的疆界是从 西顿 到 基拉耳 ，直到 迦萨 ，又到 所多玛 、 蛾摩拉 、 押玛 、 洗扁 ，直到 拉沙 。
GEN|10|20|这就是 含 的后裔，各有自己的宗族、语言、土地和国家。
GEN|10|21|闪 也生了儿子，他是 雅弗 的哥哥 ，是 希伯 人的祖先。
GEN|10|22|闪 的儿子是 以拦 、 亚述 、 亚法撒 、 路德 、 亚兰 。
GEN|10|23|亚兰 的儿子是 乌斯 、 户勒 、 基帖 、 玛施 。
GEN|10|24|亚法撒 生 沙拉 ， 沙拉 生 希伯 。
GEN|10|25|希伯 生了两个儿子，一个名叫 法勒 ，因为那时人分地居住； 法勒 的兄弟名叫 约坍 。
GEN|10|26|约坍 生 亚摩答 、 沙列 、 哈萨玛非 、 耶拉 、
GEN|10|27|哈多兰 、 乌萨 、 德拉 、
GEN|10|28|俄巴路 、 亚比玛利 、 示巴 、
GEN|10|29|阿斐 、 哈腓拉 、 约巴 ，这些都是 约坍 的儿子。
GEN|10|30|他们所住的地方是从 米沙 直到 西发 ，到东边的山。
GEN|10|31|这就是 闪 的后裔，各有自己的宗族、语言、土地和国家。
GEN|10|32|这些是 挪亚 儿子的宗族，按着他们的后代立国。洪水以后，邦国就从他们散布在地上。
GEN|11|1|那时，全地只有一种语言，都说一样的话。
GEN|11|2|他们向东迁移的时候，在 示拿 地找到一片平原，就住在那里。
GEN|11|3|他们彼此商量说：“来，让我们来做砖，把砖烧透了。”他们就拿砖当石头，又拿柏油当泥浆。
GEN|11|4|他们说：“来，让我们建造一座城和一座塔，塔顶通天。我们要为自己立名，免得我们分散在全地面上。”
GEN|11|5|耶和华降临，要看世人所建造的城和塔。
GEN|11|6|耶和华说：“看哪，他们成了同一个民族，都有一样的语言。这只是他们开始做的事，现在他们想要做的任何事，就没有什么可拦阻他们了。
GEN|11|7|来，我们下去，在那里变乱他们的语言，使他们彼此语言不通。”
GEN|11|8|于是耶和华使他们从那里分散在全地面上；他们就停止建造那城了。
GEN|11|9|因为耶和华在那里变乱了全地的语言，把人从那里分散在全地面上，所以那城名叫 巴别 。
GEN|11|10|这是 闪 的后代。洪水以后二年， 闪 一百岁生了 亚法撒 。
GEN|11|11|闪 生 亚法撒 之后又活了五百年，并且生儿育女。
GEN|11|12|亚法撒 活到三十五岁，生了 沙拉 。
GEN|11|13|亚法撒 生 沙拉 之后又活了四百零三年，并且生儿育女。
GEN|11|14|沙拉 活到三十岁，生了 希伯 。
GEN|11|15|沙拉 生 希伯 之后又活了四百零三年，并且生儿育女。
GEN|11|16|希伯 活到三十四岁，生了 法勒 。
GEN|11|17|希伯 生 法勒 之后又活了四百三十年，并且生儿育女。
GEN|11|18|法勒 活到三十岁，生了 拉吴 。
GEN|11|19|法勒 生 拉吴 之后又活了二百零九年，并且生儿育女。
GEN|11|20|拉吴 活到三十二岁，生了 西鹿 。
GEN|11|21|拉吴 生 西鹿 之后又活了二百零七年，并且生儿育女。
GEN|11|22|西鹿 活到三十岁，生了 拿鹤 。
GEN|11|23|西鹿 生 拿鹤 之后又活了二百年，并且生儿育女。
GEN|11|24|拿鹤 活到二十九岁，生了 他拉 。
GEN|11|25|拿鹤 生 他拉 之后又活了一百一十九年，并且生儿育女。
GEN|11|26|他拉 活到七十岁，生了 亚伯兰 、 拿鹤 和 哈兰 。
GEN|11|27|这是 他拉 的后代。 他拉 生 亚伯兰 、 拿鹤 和 哈兰 ； 哈兰 生 罗得 。
GEN|11|28|哈兰 死在他父亲 他拉 的面前，死在他的出生地 迦勒底 的 吾珥 。
GEN|11|29|亚伯兰 、 拿鹤 各娶了妻。 亚伯兰 的妻子名叫 撒莱 ， 拿鹤 的妻子名叫 密迦 ，是 哈兰 的女儿。 哈兰 是 密迦 和 亦迦 的父亲。
GEN|11|30|撒莱 不生育，没有孩子。
GEN|11|31|他拉 带着他儿子 亚伯兰 和他孙子， 哈兰 的儿子 罗得 ，以及他的媳妇， 亚伯兰 的妻子 撒莱 ，一同出了 迦勒底 的 吾珥 ，要往 迦南 地去；他们来到 哈兰 ，就住在那里。
GEN|11|32|他拉 共活了二百零五年，就死在 哈兰 。
GEN|12|1|耶和华对 亚伯兰 说：“你要离开本地、本族、父家，往我所要指示你的地去。
GEN|12|2|我必使你成为大国，我必赐福给你，使你的名为大；你要使别人得福 。
GEN|12|3|为你祝福的，我必赐福给他；诅咒你的，我必诅咒他。地上的万族都必因你得福。”
GEN|12|4|亚伯兰 就遵照耶和华的吩咐去了； 罗得 也和他同去。 亚伯兰 离开 哈兰 的时候年七十五岁。
GEN|12|5|亚伯兰 带着他妻子 撒莱 和侄儿 罗得 ，以及他们在 哈兰 积蓄的财物、获得的人口，往 迦南 地去。他们就来到了 迦南 地。
GEN|12|6|亚伯兰 经过那地，直到 示剑 地方， 摩利 橡树那里；当时 迦南 人住在那地。
GEN|12|7|耶和华向 亚伯兰 显现，说：“我要把这地赐给你的后裔。” 亚伯兰 就在那里为向他显现的耶和华筑了一座坛。
GEN|12|8|从那里他又迁到 伯特利 东边的山，支搭帐棚；西边是 伯特利 ，东边是 艾 。他在那里又为耶和华筑了一座坛，求告耶和华的名。
GEN|12|9|后来 亚伯兰 渐渐迁往 尼革夫 去。
GEN|12|10|那地遭遇饥荒。 亚伯兰 因那地的饥荒严重，就下到 埃及 ，要在那里寄居。
GEN|12|11|将近 埃及 ，他对妻子 撒莱 说：“看哪，我知道你是美貌的女人。
GEN|12|12|埃及 人看见你会说：‘这是他的妻子’，他们就会杀我，却让你活着。
GEN|12|13|所以，请你说你是我的妹妹，使我可以因你得平安，我的性命也因你存活。”
GEN|12|14|亚伯兰 到达 埃及 时， 埃及 人看见那女人极其美貌。
GEN|12|15|法老的臣仆看见了她，就在法老面前称赞她。那女人就被带进法老的宫中。
GEN|12|16|法老就因她厚待 亚伯兰 ，给了 亚伯兰 许多牛、羊、公驴、奴仆、婢女、母驴、骆驼。
GEN|12|17|耶和华因 亚伯兰 妻子 撒莱 的缘故，降大灾击打法老和他的全家。
GEN|12|18|法老召了 亚伯兰 来，说：“你向我做的是什么事呢？为什么没有告诉我她是你的妻子？
GEN|12|19|为什么说‘她是我的妹妹’，以致我把她接来要作我的妻子呢？现在 ，看哪，你的妻子在这里，带她走吧！”
GEN|12|20|于是法老吩咐人把 亚伯兰 和他妻子，以及他一切所有的都送走了。
GEN|13|1|亚伯兰 带着他的妻子与 罗得 ，以及一切所有的，从 埃及 上 尼革夫 去。
GEN|13|2|亚伯兰 的牲畜和金银极多。
GEN|13|3|他从 尼革夫 渐渐往 伯特利 去，到了 伯特利 和 艾 的中间，当初他支搭帐棚的地方，
GEN|13|4|也是他起先筑坛的地方。 亚伯兰 在那里求告耶和华的名。
GEN|13|5|与 亚伯兰 同行的 罗得 也有牛群、羊群、帐棚。
GEN|13|6|那地容不下他们住在一起；因为他们的财物非常多，使他们不能同住一起。
GEN|13|7|当时， 迦南 人与 比利洗 人在那地居住。 亚伯兰 的牧人和 罗得 的牧人之间起了争端。
GEN|13|8|亚伯兰 就对 罗得 说：“你我不可以相争，你的牧人和我的牧人也不可以相争，因为我们是一家人。
GEN|13|9|遍地不都在你眼前吗？请你离开我吧！你向左，我就向右；你向右，我就向左。”
GEN|13|10|罗得 举目，看见 约旦河 整个平原，直到 琐珥 ，都是水源充足之地。在耶和华未毁灭 所多玛 、 蛾摩拉 以前，那地好像耶和华的园子，又像 埃及 地。
GEN|13|11|于是 罗得 选择了 约旦河 整个平原。 罗得 往东迁移，他们就彼此分开了。
GEN|13|12|亚伯兰 住在 迦南 地； 罗得 住在平原的城镇，他渐渐迁移帐棚，直到 所多玛 。
GEN|13|13|所多玛 人在耶和华面前罪大恶极。
GEN|13|14|罗得 离开 亚伯兰 以后，耶和华对 亚伯兰 说：“你要从你所在的地方，举目向东西南北观看；
GEN|13|15|你所看见一切的地，我都要把它赐给你和你的后裔，直到永远。
GEN|13|16|我要使你的后裔好像地上的尘沙，人若能数地上的尘沙，才能数你的后裔。
GEN|13|17|你起来，纵横走遍这地，因为我必把这地赐给你。”
GEN|13|18|亚伯兰 就迁移帐棚，来到 希伯仑 ， 幔利 的橡树那里居住，在那里为耶和华筑了一座坛。
GEN|14|1|当 暗拉非 作 示拿 王， 亚略 作 以拉撒 王， 基大老玛 作 以拦 王， 提达 作 戈印 王的时候，
GEN|14|2|他们攻打 所多玛 王 比拉 、 蛾摩拉 王 比沙 、 押玛 王 示纳 、 洗扁 王 善以别 和 比拉 王， 比拉 就是 琐珥 。
GEN|14|3|这些王都会合在 西订谷 ， 西订谷 就是 盐海 。
GEN|14|4|他们已经服事 基大老玛 十二年，第十三年就背叛了。
GEN|14|5|第十四年， 基大老玛 和与他结盟的王都来了，在 亚特律．加宁 击败 利乏音 人，在 哈麦 击败 苏西 人，在 沙微．基列亭 击败 以米 人，
GEN|14|6|在 何利 人的 西珥山 击败 何利 人，一直到靠近旷野的 伊勒．巴兰 。
GEN|14|7|他们转回，来到 安．密巴 ，就是 加低斯 ，击败了 亚玛力 全地的人，以及住在 哈洗逊．他玛 的 亚摩利 人。
GEN|14|8|于是 所多玛 王、 蛾摩拉 王、 押玛 王、 洗扁 王和 比拉 王， 比拉 就是 琐珥 ，都出来，在 西订谷 摆阵，与他们交战，
GEN|14|9|就是与 以拦 王 基大老玛 、 戈印 王 提达 、 示拿 王 暗拉非 、 以拉撒 王 亚略 交战；这就是四王对五王之战。
GEN|14|10|西订谷 有许多柏油坑。 所多玛 王和 蛾摩拉 王逃跑，掉在坑里，其余的人都往山上逃跑。
GEN|14|11|四王就把 所多玛 和 蛾摩拉 所有的财物和所有的粮食都掳掠去了；
GEN|14|12|他们也把 亚伯兰 的侄儿 罗得 和 罗得 的财物都掳掠去了。当时 罗得 住在 所多玛 。
GEN|14|13|有一个逃脱的人来告诉 希伯来 人 亚伯兰 ； 亚伯兰 正住在 亚摩利 人 幔利 的橡树那里。 幔利 、 以实各 和 亚乃 都是弟兄，曾与 亚伯兰 结盟。
GEN|14|14|亚伯兰 听见他侄儿 被掳去，就把三百一十八个生在他家中、受过训练的壮丁全都出动 去追，一直到 但 。
GEN|14|15|在夜间，他和他的仆人分队击败了敌人，并且追杀他们，直到 大马士革 北边的 何把 。
GEN|14|16|他把一切被掳掠的财物夺回，也把他侄儿 罗得 和他的财物，以及人和妇女都夺回来。
GEN|14|17|亚伯兰 击败 基大老玛 和与他结盟的王回来的时候， 所多玛 王出来，在 沙微谷 迎接他， 沙微谷 就是 王的谷 。
GEN|14|18|又有 撒冷 王 麦基洗德 带着饼和酒出来；他是至高上帝的祭司。
GEN|14|19|他为 亚伯兰 祝福，说： “愿至高的上帝、 天地的主赐福给 亚伯兰 ！
GEN|14|20|至高的上帝把敌人交在你手里， 他是应当称颂的！” 亚伯兰 就把所有的拿出十分之一给他。
GEN|14|21|所多玛 王对 亚伯兰 说：“你把人还给我，财物你自己拿去吧！”
GEN|14|22|亚伯兰 对 所多玛 王说：“我指着耶和华—至高的上帝、天地的主起誓：
GEN|14|23|凡是你的东西，就是一根线、一条鞋带，我都不拿，免得你说：‘是我使 亚伯兰 富足！’
GEN|14|24|我什么都不要，只是仆人所吃的，以及与我同去的 亚乃 、 以实各 、 幔利 所应得的份，让他们拿去吧！”
GEN|15|1|这些事以后，耶和华的话在异象中临到 亚伯兰 ，说：“ 亚伯兰 哪，不要惧怕！我是你的盾牌，你必得丰富的赏赐。”
GEN|15|2|亚伯兰 说：“主耶和华啊，我还没有儿子，你能赐我什么呢？承受我家业的是 大马士革 人 以利以谢 。”
GEN|15|3|亚伯兰 又说：“看哪，你没有给我后嗣。你看，那生在我家中的人要继承我。”
GEN|15|4|看哪，耶和华的话又临到他，说：“这人不会继承你，你本身所生的才会继承你。”
GEN|15|5|于是耶和华带他到外面，说：“你向天观看，去数星星，你能数得清吗？”又对他说：“你的后裔将要如此。”
GEN|15|6|亚伯兰 信耶和华，耶和华就以此算他为义。
GEN|15|7|耶和华又对他说：“我是耶和华，曾领你出 迦勒底 的 吾珥 ，为要把这地赐你为业。”
GEN|15|8|亚伯兰 说：“主耶和华啊，我怎能知道我必得这地为业呢？”
GEN|15|9|耶和华对他说：“你为我取一头三岁的母牛犊，一只三岁的母山羊，一只三岁的公绵羊，一只斑鸠和一只雏鸽。”
GEN|15|10|亚伯兰 就把这些都取来，每样从中间劈成两半，一半对着另一半排列，只有鸟没有劈开。
GEN|15|11|当鸷鸟下来，落在这些尸体上时， 亚伯兰 就把它们赶走了。
GEN|15|12|日落的时候， 亚伯兰 沉睡了。看哪，有大而可怕的黑暗落在他身上。
GEN|15|13|耶和华对 亚伯兰 说：“你要确实知道，你的后裔必寄居在别人的地，服事那地的人；那地的人要虐待他们四百年。
GEN|15|14|但我要惩罚他们所服事的那国，以后他们必带着许多财物从那里出来。
GEN|15|15|至于你，你要平平安安归到你祖先那里，必享长寿，被人埋葬。
GEN|15|16|到了第四代，他们必回到这里，因为 亚摩利 人的罪恶到现在还没有满盈。”
GEN|15|17|日落天黑的时候，看哪，有冒烟的炉和烧着的火把从那些肉块中经过。
GEN|15|18|在那日，耶和华与 亚伯兰 立约，说：“我已赐给你的后裔这一片地，从 埃及河 直到 大河 ， 幼发拉底河 ，
GEN|15|19|就是 基尼 人、 基尼洗 人、 甲摩尼 人、
GEN|15|20|赫 人、 比利洗 人、 利乏音 人、
GEN|15|21|亚摩利 人、 迦南 人、 革迦撒 人、 耶布斯 人的地。”
GEN|16|1|亚伯兰 的妻子 撒莱 没有为他生孩子。 撒莱 有一个婢女，是 埃及 人，名叫 夏甲 。
GEN|16|2|撒莱 对 亚伯兰 说：“看哪，耶和华使我不能生育。你来和我的婢女同房，也许我可以从她得孩子 。” 亚伯兰 听从了 撒莱 的话。
GEN|16|3|于是 亚伯兰 的妻子 撒莱 把她的婢女， 埃及 人 夏甲 ，给了丈夫为妾；那时 亚伯兰 在 迦南 已经住了十年。
GEN|16|4|亚伯兰 与 夏甲 同房， 夏甲 就怀了孕。她看见自己有孕，就轻视她的女主人。
GEN|16|5|撒莱 对 亚伯兰 说：“我因你受了委屈。我把我的婢女放在你怀中，她见自己怀了孕，就轻视我。愿耶和华在你我之间判断。”
GEN|16|6|亚伯兰 对 撒莱 说：“看哪，婢女在你手里，你可以照你看为好的对待她。”于是， 撒莱 虐待她，她就从 撒莱 面前逃走了。
GEN|16|7|耶和华的使者在旷野的水泉旁，在 书珥 路上的水泉旁遇见 夏甲 ，
GEN|16|8|对她说：“ 撒莱 的婢女 夏甲 ，你从哪里来？要到哪里去？”她说：“我从我的女主人 撒莱 面前逃出来。”
GEN|16|9|耶和华的使者对她说：“你要回到你的女主人那里，屈服在她手下。”
GEN|16|10|耶和华的使者对她说： “我必使你的后裔极其繁多， 多到不可胜数。”
GEN|16|11|耶和华的使者又对她说： “看哪，你已怀孕， 要生一个儿子。 你要给他起名叫 以实玛利 ， 因为耶和华听见了你的苦楚。
GEN|16|12|他为人必像野驴。 他的手要攻打人， 人的手也要攻打他； 他必常与他的众弟兄作对 。”
GEN|16|13|夏甲 就称那向她说话的耶和华为“你是看见 的上帝”，因为她说：“他看见了我之后，我还能在这里看见他吗？”
GEN|16|14|所以这井名叫 庇耳．拉海．莱 ，看哪，它位于 加低斯 和 巴列 的中间。
GEN|16|15|后来 夏甲 为 亚伯兰 生了一个儿子； 亚伯兰 给 夏甲 生的儿子起名叫 以实玛利 。
GEN|16|16|夏甲 为 亚伯兰 生 以实玛利 的时候， 亚伯兰 年八十六岁。
GEN|17|1|亚伯兰 九十九岁时，耶和华向他显现，对他说：“我是全能的上帝。你当在我面前行走，作完全的人，
GEN|17|2|我要与你立约，使你的后裔极其繁多。”
GEN|17|3|亚伯兰 脸伏于地；上帝又对他说：
GEN|17|4|“看哪，这就是我与你立的约，你要成为多国的父。
GEN|17|5|从今以后，你的名字不再叫 亚伯兰 ，要叫 亚伯拉罕 ，因为我已经立你作多国之父。
GEN|17|6|我必使你生养极其繁多；国度要从你而立，君王要从你而出。
GEN|17|7|我要与你，以及你世世代代的后裔坚立我的约，成为永远的约，是要作你和你后裔的上帝。
GEN|17|8|我要把你现在寄居的地，就是 迦南 全地，赐给你和你的后裔永远为业；我也必作他们的上帝。”
GEN|17|9|上帝又对 亚伯拉罕 说：“你和你的后裔一定要世世代代遵守我的约。
GEN|17|10|这就是我与你，以及你的后裔所立的约，是你们所当遵守的，你们所有的男子都要受割礼。
GEN|17|11|你们要割去肉体的包皮，这是我与你们立约的记号。
GEN|17|12|你们世世代代的男子，无论是在家里生的，或是用银子从外人买来而不是你后裔生的，都要在生下来的第八日受割礼。
GEN|17|13|你家里生的和你用银子买的，都必须受割礼。这样，我的约就在你们肉体上成为永远的约。
GEN|17|14|不受割礼的男子都必从民中剪除，因他违背了我的约。”
GEN|17|15|上帝又对 亚伯拉罕 说：“至于你的妻子 撒莱 ，不可再叫她 撒莱 ，她的名要叫 撒拉 。
GEN|17|16|我必赐福给她，也要从她赐一个儿子给你。我必赐福给 撒拉 ，她要兴起多国；必有百姓的君王从她而出。”
GEN|17|17|亚伯拉罕 就脸伏于地窃笑，心里想：“一百岁的人还能有孩子吗？ 撒拉 已经九十岁了，还能生育吗？”
GEN|17|18|亚伯拉罕 对上帝说：“但愿 以实玛利 活在你面前。”
GEN|17|19|上帝说：“不！你妻子 撒拉 必为你生一个儿子，你要给他起名叫 以撒 。我要与他坚立我的约，成为他后裔永远的约。
GEN|17|20|至于 以实玛利 ，我已听见你了：看哪，我必赐福给他，使他兴旺，极其繁多。他必生十二个族长，我要使他成为大国。
GEN|17|21|到明年所定的时候， 撒拉 必为你生 以撒 ，我要与他坚立我的约。”
GEN|17|22|上帝和 亚伯拉罕 说完了话，就离开他上升去了。
GEN|17|23|在那一天， 亚伯拉罕 遵照上帝所说的，给他的儿子 以实玛利 和家里所有的男丁，无论是在家里生的，或是用银子买来的，都行了割礼 。
GEN|17|24|亚伯拉罕 受割礼时，年九十九岁。
GEN|17|25|他儿子 以实玛利 受割礼时，年十三岁。
GEN|17|26|在那一天， 亚伯拉罕 和他儿子 以实玛利 一同受了割礼。
GEN|17|27|家里所有的男人，无论是在家里生的，或是用银子从外人买来的，也都一同受了割礼。
GEN|18|1|耶和华在 幔利 橡树那里向 亚伯拉罕 显现。天正热的时候， 亚伯拉罕 坐在帐棚门口。
GEN|18|2|他举目观看，看哪，有三个人站在他附近。他一看见，就从帐棚门口跑去迎接他们，俯伏在地，
GEN|18|3|说：“我主，我若在你眼前蒙恩，请不要离开你的仆人走过去。
GEN|18|4|容我拿点水来，请你们洗脚，在树下休息。
GEN|18|5|既然你们来到仆人这里了，我再拿点饼来，让你们恢复心力，然后再走。”他们说：“就照你说的去做吧。”
GEN|18|6|亚伯拉罕 急忙进帐棚到 撒拉 那里，说：“你赶快拿三细亚细面，揉面做饼。”
GEN|18|7|亚伯拉罕 又跑到牛群里，牵了一头又嫩又好的牛犊来，交给仆人，仆人就急忙去预备。
GEN|18|8|亚伯拉罕 取了乳酪和奶，以及预备好了的牛犊来，摆在他们面前，自己在树下站在旁边，他们就吃了。
GEN|18|9|他们对 亚伯拉罕 说：“你妻子 撒拉 在哪里？”他说：“看哪，在帐棚里。”
GEN|18|10|有一位说：“明年这时候 ，我一定会回到你这里。看哪，你的妻子 撒拉 会生一个儿子。” 撒拉 在那人后面的帐棚门口也听见了。
GEN|18|11|亚伯拉罕 和 撒拉 都年纪老迈， 撒拉 的月经已停了。
GEN|18|12|撒拉 心里窃笑，说：“我已衰老，我的主也老了，怎能有这喜事呢？”
GEN|18|13|耶和华对 亚伯拉罕 说：“ 撒拉 为什么窃笑，说：‘我已年老，果真能生育吗？’
GEN|18|14|耶和华岂有难成的事吗？到了所定的时候，我必回到你这里。明年这时候， 撒拉 会生一个儿子。”
GEN|18|15|撒拉 因为害怕，就不承认，说：“我没有笑。”那人说：“不，你的确笑了。”
GEN|18|16|三人从那里起程，面向 所多玛 观望， 亚伯拉罕 与他们同行，要送他们一程。
GEN|18|17|耶和华说：“我所要做的事岂可瞒着 亚伯拉罕 呢？
GEN|18|18|亚伯拉罕 必要成为强大的国；地上的万国都必因他得福。
GEN|18|19|我拣选他 ，为要叫他命令他的子孙和后代家属遵行耶和华的道，秉公行义，使耶和华所应许 亚伯拉罕 的话都实现了。”
GEN|18|20|耶和华说：“ 所多玛 和 蛾摩拉 罪恶极其严重，控告他们的声音很大。
GEN|18|21|我要下去察看他们所做的，是否真的像那达到我这里的声音一样；如果不是，我也要知道。”
GEN|18|22|二人转身离开那里，往 所多玛 去；但 亚伯拉罕 仍然站在耶和华面前。
GEN|18|23|亚伯拉罕 近前来，说：“你真的要把义人和恶人一同剿灭吗？
GEN|18|24|假若那城里有五十个义人，你真的还要剿灭，不因城里这五十个义人饶了那地方吗？
GEN|18|25|你绝不会做这样的事，把义人与恶人一同杀了，使义人与恶人一样。你绝不会这样！审判全地的主岂不做公平的事吗？”
GEN|18|26|耶和华说：“我若在 所多玛城 里找到五十个义人，我就为他们的缘故饶恕那整个地方。”
GEN|18|27|亚伯拉罕 回答说：“看哪，我虽只是尘土灰烬，还敢向主说话。
GEN|18|28|假若这五十个义人少了五个，你就因为少了五个而毁灭全城吗？”他说：“我在那里若找到四十五个，就不毁灭。”
GEN|18|29|亚伯拉罕 又对他说：“假若在那里找到四十个呢？”他说：“为这四十个的缘故，我也不做。”
GEN|18|30|亚伯拉罕 说：“求主不要生气，容我说，假若在那里找到三十个呢？”他说：“我在那里若找到三十个，我也不做。”
GEN|18|31|亚伯拉罕 说：“看哪，我还敢向主说，假若在那里找到二十个呢？”他说：“为这二十个的缘故，我也不毁灭。”
GEN|18|32|亚伯拉罕 说：“求主不要生气，我再说一次，假若在那里找到十个呢？”他说：“为这十个的缘故，我也不毁灭。”
GEN|18|33|耶和华与 亚伯拉罕 说完了话就走了； 亚伯拉罕 也回到自己的地方去了。
GEN|19|1|两个天使在傍晚到了 所多玛 ， 罗得 正坐在 所多玛 的城门口。 罗得 一看见，就起身迎接他们，脸伏于地下拜，
GEN|19|2|说：“看哪，我主，请你们转到仆人家里过夜，洗你们的脚，清早起来再上路。”他们说：“不！我们要在广场上过夜。”
GEN|19|3|罗得 恳切地请他们，他们就转向他，进到他屋里。 罗得 为他们预备宴席，烤无酵饼，他们就吃了。
GEN|19|4|他们还没有躺下， 所多玛城 的人，连老带少所有的人，个个都来围住那屋子。
GEN|19|5|他们呼叫 罗得 ，对他说：“今天晚上到你这里来的人在哪里？把他们带出来，让我们亲近他们。”
GEN|19|6|罗得 出了门，把身后的门关上，到众人那里，
GEN|19|7|说：“我的弟兄们，请你们不要做这恶事。
GEN|19|8|看哪，我有两个女儿，还没有亲近过男人，让我领她们出来给你们，就照你们看为好的对待她们吧！只是这两个人既然到我舍下，请不要向他们做这事。”
GEN|19|9|众人说：“站到一边去吧！”又说：“这个人来寄居，还想扮审判官呢！现在我们要害你比害他们更厉害。”众人就往前冲向 罗得 ，要攻破大门。
GEN|19|10|那两个人伸出手来，把 罗得 拉进屋子他们那里，就关上门。
GEN|19|11|他们击打门外的人，无论老少，都眼睛迷糊，找门找得很烦躁。
GEN|19|12|那两个人对 罗得 说：“你这里还有什么人吗？无论是女婿，是儿女，这城中所有属你的人，你都要把他们从这地方带出去。
GEN|19|13|我们要毁灭这地方，因为控告城内百姓的声音在耶和华面前非常大，耶和华派我们来毁灭这城。”
GEN|19|14|罗得 出去，告诉娶了 他女儿的女婿们说：“起来，离开这地方，因为耶和华要毁灭这城。”他的女婿们却以为他说的是笑话。
GEN|19|15|天亮了，天使催逼 罗得 说：“起来！带着你的妻子和你这里的两个女儿出去，免得你因这城的罪孽同被剿灭。”
GEN|19|16|但 罗得 迟延不走。二人因为耶和华怜悯 罗得 ，就拉着他的手和他妻子的手，以及他两个女儿的手，把他们领出来，安置在城外；
GEN|19|17|领他们出来以后，就说：“逃命吧！不可回头看，也不可在平原站住。要往山上逃跑，免得你被剿灭。”
GEN|19|18|罗得 对他们说：“我主啊，不要这样！
GEN|19|19|看哪，你仆人已经在你眼前蒙恩，你又向我大施慈爱，救我的性命。但是我不能逃到山上去，恐怕这灾祸追上我，我就死了。
GEN|19|20|看哪，这城又近又小，比较容易逃到那里。这不是一座小城吗？求你容我逃到那里，使我的性命可以存活。”
GEN|19|21|天使对他说：“看哪，这事我也应允你，不倾覆你所说的这城。
GEN|19|22|你要赶快逃到那城，因为你还没有到那里，我不能做什么。”因此那城名叫 琐珥 。
GEN|19|23|罗得 到了 琐珥 ，太阳已经升出地面。
GEN|19|24|当时，耶和华把硫磺与火，从天上耶和华那里降与 所多玛 和 蛾摩拉 ，
GEN|19|25|把那些城和全平原，城里所有的居民和土地上生长的，都毁灭了。
GEN|19|26|罗得 的妻子在他后边回头一看，就变成了一根盐柱。
GEN|19|27|亚伯拉罕 清早起来，到了他先前站在耶和华面前的地方，
GEN|19|28|面向 所多玛 和 蛾摩拉 ，以及平原全地观望。他观看，看哪，那地有浓烟上腾，好像烧窑的浓烟。
GEN|19|29|当上帝毁灭平原诸城的时候，他记念 亚伯拉罕 ；在倾覆 罗得 所住之城的时候，就把 罗得 从倾覆中带出来。
GEN|19|30|罗得 因为怕住在 琐珥 ，就同他两个女儿从 琐珥 上去，住在山上。他和两个女儿住在一个洞里。
GEN|19|31|大女儿对小女儿说：“我们的父亲老了，这地又没有男人可以照世上的礼俗来与我们结合。
GEN|19|32|来！我们叫父亲喝酒，然后与他同寝。这样，我们可以从我们的父亲存留后裔。”
GEN|19|33|于是，那晚她们叫父亲喝酒，大女儿就进去和她父亲同寝；她几时躺下，几时起来，父亲都不知道。
GEN|19|34|第二天，大女儿对小女儿说：“看哪，我昨夜与父亲同寝。今晚我们再叫他喝酒，你进去与他同寝。这样，我们可以从父亲存留后裔。”
GEN|19|35|于是，那晚她们又叫父亲喝酒，小女儿起来与她父亲同寝；她几时躺下，几时起来，父亲都不知道。
GEN|19|36|这样， 罗得 的两个女儿都从她们的父亲怀了孕。
GEN|19|37|大女儿生了儿子，给他起名叫 摩押 ，就是现今 摩押 人的始祖。
GEN|19|38|小女儿也生了儿子，给他起名叫 便．亚米 ，就是现今 亚扪 人的始祖。
GEN|20|1|亚伯拉罕 从那里往 尼革夫 迁移，寄居在 加低斯 和 书珥 之间的 基拉耳 。
GEN|20|2|亚伯拉罕 称他的妻子 撒拉 为妹妹。 基拉耳 王 亚比米勒 派人把 撒拉 带走。
GEN|20|3|夜间，上帝在梦中来到 亚比米勒 那里，对他说：“看哪，你要死了，因为你带来的女人，她是有丈夫的女子！”
GEN|20|4|亚比米勒 还未亲近 撒拉 ；他说：“主啊，连公义的国，你也要毁灭吗？
GEN|20|5|那人岂不是自己对我说‘她是我妹妹’吗？连这女人自己也说：‘他是我哥哥。’我做这事是心正手洁的。”
GEN|20|6|上帝在梦中对他说：“我也知道你做这事是心中正直的；是我拦阻了你，免得你得罪我。所以我不让你侵犯她。
GEN|20|7|现在你当把这人的妻子归还给他；因为他是先知，他要为你祷告，使你存活。你若不归还，你当知道，你和你所有的人都必定死。”
GEN|20|8|亚比米勒 清早起来，叫了他的众臣仆来，把这一切事说给他们听，他们就很害怕。
GEN|20|9|亚比米勒 召了 亚伯拉罕 来，对他说：“你怎么向我这样做呢？我什么事得罪你，你竟使我和我的国陷在大罪中呢？你对我做了不该做的事了！”
GEN|20|10|亚比米勒 对 亚伯拉罕 说：“你看见什么才做这事呢？”
GEN|20|11|亚伯拉罕 说：“我以为这地方的人根本不敬畏上帝，必为我妻子的缘故杀我。
GEN|20|12|况且她也真是我的妹妹；她与我是同父异母的，后来作了我的妻子。
GEN|20|13|当上帝叫我离开父家、飘流在外的时候，我对她说：我们无论走到什么地方，你要对人说：‘他是我哥哥’，这就是你以慈爱待我了。”
GEN|20|14|亚比米勒 把牛、羊、奴仆、婢女送给 亚伯拉罕 ，也把他的妻子 撒拉 归还给他。
GEN|20|15|亚比米勒 说：“看哪，我的地都在你面前，你看为好的地方就居住吧。”
GEN|20|16|他对 撒拉 说：“看哪，我给你哥哥一千银子。看哪，这要在你全家人面前遮羞 ，向众人证实你是清白的。”
GEN|20|17|亚伯拉罕 向上帝祷告，上帝就医好 亚比米勒 和他的妻子，以及他的使女们，他们就能生育。
GEN|20|18|因耶和华为 亚伯拉罕 的妻子 撒拉 的缘故，已经使 亚比米勒 家中的妇人不能怀孕。
GEN|21|1|耶和华照着他所说的眷顾 撒拉 ，耶和华实现了他对 撒拉 的应许。
GEN|21|2|亚伯拉罕 年老，到上帝对他说的那所定的时候， 撒拉 怀了孕，给他生了一个儿子。
GEN|21|3|亚伯拉罕 给 撒拉 所生的儿子起名叫 以撒 。
GEN|21|4|以撒 出生后第八日， 亚伯拉罕 遵照上帝所吩咐的，为 以撒 行割礼。
GEN|21|5|他儿子 以撒 出生的时候， 亚伯拉罕 年一百岁。
GEN|21|6|撒拉 说：“上帝使我欢笑，凡听见的人必与我一同欢笑”，
GEN|21|7|又说：“谁能预先对 亚伯拉罕 说， 撒拉 要乳养孩子呢？因为在他年老的时候，我为他生了一个儿子。”
GEN|21|8|孩子渐渐长大，就断了奶。 以撒 断奶的那一天， 亚伯拉罕 摆设丰盛的宴席。
GEN|21|9|那时， 撒拉 看见 埃及 人 夏甲 为 亚伯拉罕 所生的儿子戏笑，
GEN|21|10|就对 亚伯拉罕 说：“你把这使女和她儿子赶出去！因为这使女的儿子不可与我的儿子 以撒 一同承受产业。”
GEN|21|11|亚伯拉罕 为这事非常忧愁，因为关乎他的儿子。
GEN|21|12|上帝对 亚伯拉罕 说：“你不必为这孩子和你的使女忧愁。 撒拉 对你说的话，你都要听从；因为从 以撒 生的，才要称为你的后裔。
GEN|21|13|至于使女的儿子，我也必使他成为一国，因为他是你的后裔。”
GEN|21|14|亚伯拉罕 清早起来，拿饼和一皮袋水，给了 夏甲 ，搭在她肩上，把她和孩子一起送走。 夏甲 就走了，但她却在 别是巴 的旷野流浪。
GEN|21|15|皮袋的水用完了， 夏甲 就把孩子放在一棵小树下，
GEN|21|16|自己走开约有一箭之远，相对而坐，说：“我不忍心看见孩子死”。她就坐在对面，放声大哭。
GEN|21|17|上帝听见孩子的声音，上帝的使者就从天上呼叫 夏甲 说：“ 夏甲 ，你为何这样呢？不要害怕，上帝已经听见孩子在那里的声音了。
GEN|21|18|起来！把孩子扶起来，用你的手握住他，因我必使他成为大国。”
GEN|21|19|上帝开了 夏甲 的眼睛，她就看见一口水井。她就去，把皮袋装满了水，给孩子喝。
GEN|21|20|上帝与这孩子同在，他就渐渐长大，住在旷野，成了一个弓箭手。
GEN|21|21|他住在 巴兰 的旷野；他母亲从 埃及 地为他娶了一个妻子。
GEN|21|22|那时候， 亚比米勒 和他的将军 非各 对 亚伯拉罕 说：“凡你所做的事，上帝都与你同在。
GEN|21|23|我愿你如今在这里指着上帝对我起誓，不要亏待我和我的儿子，以及我的子孙。我怎样忠诚待你，你也要照样忠诚待我和你所寄居的这地。”
GEN|21|24|亚伯拉罕 说：“我愿意起誓。”
GEN|21|25|先前， 亚比米勒 的仆人霸占了一口水井， 亚伯拉罕 为这事责备 亚比米勒 。
GEN|21|26|亚比米勒 说：“我不知道谁做了这事，你也没有告诉我，我到今日才听到。”
GEN|21|27|亚伯拉罕 把羊和牛给了 亚比米勒 ，二人就彼此立约。
GEN|21|28|亚伯拉罕 把七只小母羊另放在一处。
GEN|21|29|亚比米勒 对 亚伯拉罕 说：“你把这七只小母羊另放一处是什么意思呢？”
GEN|21|30|他说：“你要从我手里接受这七只小母羊，作我挖了这口井的证据。”
GEN|21|31|所以他给那地方起名叫 别是巴 ，因为他们二人在那里起了誓。
GEN|21|32|他们在 别是巴 立了约， 亚比米勒 就和他的将军 非各 起身回 非利士 人的地去了。
GEN|21|33|亚伯拉罕 就在 别是巴 种了一棵柳树，在那里求告耶和华—永恒上帝的名。
GEN|21|34|亚伯拉罕 在 非利士 人的地寄居了许多日子。
GEN|22|1|这些事以后，上帝考验 亚伯拉罕 ，对他说：“ 亚伯拉罕 ！”他说：“我在这里。”
GEN|22|2|上帝说：“你要带你的儿子，就是你所爱的独子 以撒 ，往 摩利亚 地去，在我指示你的一座山上，把他献为燔祭。”
GEN|22|3|亚伯拉罕 清早起来，预备了驴，带着跟他一起的两个仆人和他儿子 以撒 ，劈好了燔祭的柴，就起身往上帝指示他的地方去了。
GEN|22|4|到了第三日， 亚伯拉罕 举目遥望那地方。
GEN|22|5|亚伯拉罕 对他的仆人说：“你们和驴留在这里，我和孩子要去那里敬拜，然后回到你们这里来。”
GEN|22|6|亚伯拉罕 把燔祭的柴放在他儿子 以撒 身上，自己手里拿着火与刀；于是二人同行。
GEN|22|7|以撒 对他父亲 亚伯拉罕 说：“我父啊！” 亚伯拉罕 说：“我儿，我在这里。” 以撒 说：“看哪，火与柴都有了，但燔祭的羔羊在哪里呢？”
GEN|22|8|亚伯拉罕 说：“我儿，上帝必自己预备燔祭的羔羊。”于是二人同行。
GEN|22|9|他们到了上帝指示他的地方， 亚伯拉罕 在那里筑坛，把柴摆好，绑了他儿子 以撒 ，放在坛的柴上。
GEN|22|10|亚伯拉罕 就伸手拿刀，要杀他的儿子。
GEN|22|11|耶和华的使者从天上呼唤他说：“ 亚伯拉罕 ！ 亚伯拉罕 ！”他说：“我在这里。”
GEN|22|12|天使说：“不可在这孩子身上下手！一点也不可伤害他！现在我知道你是敬畏上帝的人了，因为你没有把你的儿子，就是你的独子，留下不给我。”
GEN|22|13|亚伯拉罕 举目观看，看哪，一只公绵羊两角缠在灌木丛中。 亚伯拉罕 就去牵了那只公绵羊，献为燔祭，代替他的儿子。
GEN|22|14|亚伯拉罕 给那地方起名叫“耶和华以勒” 。直到今日人还说：“在耶和华的山上必有预备。”
GEN|22|15|耶和华的使者第二次从天上呼唤 亚伯拉罕 ，
GEN|22|16|说：“耶和华说：‘你既行了这事，没有留下你的儿子，就是你的独子，我指着自己起誓：
GEN|22|17|我必多多赐福给你，我必使你的后裔大大增多，如同天上的星、海边的沙。你的后裔必得仇敌的城门，
GEN|22|18|并且地上的万国都必因你的后裔得福，因为你听从了我的话。’”
GEN|22|19|于是 亚伯拉罕 回到他仆人那里。他们一同起身，往 别是巴 去， 亚伯拉罕 就住在 别是巴 。
GEN|22|20|这些事以后，有人告诉 亚伯拉罕 说：“看哪， 密迦 也为你兄弟 拿鹤 生了几个儿子：
GEN|22|21|长子 乌斯 、他的兄弟 布斯 、 亚兰 的父亲 基摩利 、
GEN|22|22|基薛 、 哈琐 、 必达 、 益拉 和 彼土利 。”
GEN|22|23|彼土利 生 利百加 。这八个人都是 密迦 为 亚伯拉罕 的兄弟 拿鹤 生的。
GEN|22|24|拿鹤 的妾名叫 流玛 ，她也生了 提八 、 迦含 、 他辖 和 玛迦 。
GEN|23|1|撒拉 享寿一百二十七岁，这是 撒拉 一生的岁数 。
GEN|23|2|撒拉 死在 迦南 地的 基列．亚巴 ，就是 希伯仑 。 亚伯拉罕 来哀悼 撒拉 ，为她哭泣。
GEN|23|3|然后， 亚伯拉罕 起来，离开死人面前，对 赫 人说：
GEN|23|4|“我在你们中间是外人，是寄居的。请给我你们那里的一块坟地，我好埋葬我的亡妻，使她不在我的面前。”
GEN|23|5|赫 人回答 亚伯拉罕 说：
GEN|23|6|“我主请听。你在我们中间是一位尊贵的王子，只管在我们最好的坟地里埋葬你的死人；我们没有一人会拒绝你在他的坟地里埋葬你的死人。”
GEN|23|7|于是， 亚伯拉罕 起来，向当地的百姓 赫 人下拜，
GEN|23|8|对他们说：“你们若愿意让我埋葬我的亡妻，使她不在我面前，就请听我，为我求 琐辖 的儿子 以弗仑 ，
GEN|23|9|把他田地尽头的 麦比拉洞 卖给我。他可以按照足价卖给我，作为我在你们中间的坟地。”
GEN|23|10|那时， 以弗仑 正坐在 赫 人中间。 赫 人 以弗仑 就回答 亚伯拉罕 ，说给所有出入城门的 赫 人听：
GEN|23|11|“不，我主请听。我要把这块田送给你，连田间的洞也送给你，在我同族的人眼前都给你，让你埋葬你的死人。”
GEN|23|12|亚伯拉罕 就在当地的百姓面前下拜，
GEN|23|13|对 以弗仑 说，也给当地百姓听：“你若应允，请你听我。我要把田的价钱给你，请你收下，我就在那里埋葬我的死人。”
GEN|23|14|以弗仑 回答 亚伯拉罕 说：
GEN|23|15|“我主请听。四百舍客勒银子的地，在你我中间算什么呢？只管埋葬你的死人吧！”
GEN|23|16|亚伯拉罕 听从了 以弗仑 。 亚伯拉罕 就照着他说给 赫 人听的，把买卖通用的银子，秤了四百舍客勒银子给 以弗仑 。
GEN|23|17|于是， 以弗仑 把那块位于 幔利 对面的 麦比拉 田，和其中的洞，以及田间周围的树木都成交了，
GEN|23|18|在所有出入城门的 赫 人眼前，卖给 亚伯拉罕 作为他的产业。
GEN|23|19|后来， 亚伯拉罕 把他妻子 撒拉 安葬在 迦南 地 幔利 对面的 麦比拉 田间的洞里， 幔利 就是 希伯仑 。
GEN|23|20|从此，那块田和田间的洞就从 赫 人移交给 亚伯拉罕 作坟地的产业。
GEN|24|1|亚伯拉罕 年纪老迈，耶和华在一切事上都赐福给他。
GEN|24|2|亚伯拉罕 对他家中管理他一切产业最老的仆人说：“把你的手放在我大腿底下。
GEN|24|3|我要叫你指着耶和华—天和地的上帝起誓，不要为我儿子娶我所居住的 迦南 地的女子为妻。
GEN|24|4|你要往我的本地本族去，为我的儿子 以撒 娶妻。”
GEN|24|5|仆人对他说：“如果那女子不肯跟我来到这地，我必须把你的儿子带回到你出来的地方吗？”
GEN|24|6|亚伯拉罕 对他说：“你要谨慎，不可带我儿子回那里去。
GEN|24|7|耶和华—天上的上帝曾带领我离开父家和本族的地，对我说话，向我起誓说：‘我要将这地赐给你的后裔。’他要差遣使者在你面前，你就可以从那里为我儿子娶妻。
GEN|24|8|倘若那女子不肯跟你来，我叫你起的誓就与你无关了，只是你不可带我的儿子回到那里去。”
GEN|24|9|仆人就把手放在他主人 亚伯拉罕 的大腿底下，为这事向他起誓。
GEN|24|10|那仆人从他主人的骆驼中取了十匹骆驼，他手中也带着他主人各样的贵重物品离开 ，起身往 美索不达米亚 去，到了 拿鹤 的城。
GEN|24|11|傍晚时，众女子出来打水，他就让骆驼跪在城外的水井旁。
GEN|24|12|他说：“耶和华—我主人 亚伯拉罕 的上帝啊，求你施恩给我的主人 亚伯拉罕 ，让我今日就遇见吧！
GEN|24|13|看哪，我站在井旁，城内居民的女子们正出来打水。
GEN|24|14|我向哪一个少女说：‘请你放下水瓶来，给我水喝’，她若说：‘请喝！我也给你的骆驼喝’，愿她作你所选定给你仆人 以撒 的妻。这样，我就知道你施恩给我的主人了。”
GEN|24|15|话还没说完，看哪， 利百加 肩头上扛着水瓶出来。 利百加 是 彼土利 所生的； 彼土利 是 亚伯拉罕 的兄弟 拿鹤 妻子 密迦 的儿子。
GEN|24|16|那少女容貌极其美丽，是未曾与人亲近的童女。她下到井旁，打满了瓶子的水，就上来。
GEN|24|17|仆人跑上前去迎着她，说：“请你让我喝你瓶子里的一点水。”
GEN|24|18|少女说：“我主请喝！”就急忙拿下瓶子托在手上，给他喝水。
GEN|24|19|那少女给他喝足了，又说：“我也为你的骆驼打水，直到骆驼喝足了。”
GEN|24|20|她就急忙把瓶子里的水倒在槽里，又跑到井旁打水，为所有的骆驼打了水。
GEN|24|21|那人定睛看着少女，一句话也不说，要知道耶和华是否使他的道路亨通。
GEN|24|22|骆驼喝足了，那人就拿出一个比加 重的金环，一对十舍客勒重的金手镯，
GEN|24|23|说：“请告诉我，你是谁的女儿？你父亲家里有没有地方可以让我们过夜？”
GEN|24|24|少女说：“我是 密迦 为 拿鹤 生的儿子 彼土利 的女儿。”
GEN|24|25|又说：“我们家里有充足的干草和饲料，也有住宿的地方。”
GEN|24|26|那人就低头向耶和华敬拜，
GEN|24|27|说：“耶和华—我主人 亚伯拉罕 的上帝是应当称颂的，因他不断以慈爱信实待我主人。至于我，耶和华一路引领我，直到我主人的兄弟家里。”
GEN|24|28|那少女跑去，把这些话告诉她母亲家里的人。
GEN|24|29|利百加 有一个哥哥，名叫 拉班 ， 拉班 就跑到外面井旁那人那里。
GEN|24|30|当他看见金环和戴在他妹妹手上的金镯，又听见他妹妹 利百加 说的话：“那人如此对我说”，他就来到那人面前，看哪，他还站在井旁的骆驼旁边，
GEN|24|31|就对他说：“你这蒙耶和华赐福的人，请进来吧！为什么站在外面？我已经收拾了房屋，也为骆驼预备了地方。”
GEN|24|32|那人就进了 拉班 的家。 拉班 卸了骆驼，用饲料喂它们，拿水给那人和随从他的人洗脚，
GEN|24|33|把食物摆在他面前，请他吃。他却说：“我不吃，等我把我的事情说完了再吃。” 拉班 说：“请说。”
GEN|24|34|他说：“我是 亚伯拉罕 的仆人。
GEN|24|35|耶和华大大地赐福给我主人，使他发达，赐给他羊群、牛群、金银、奴仆、婢女、骆驼和驴。
GEN|24|36|我主人的妻子 撒拉 年老的时候为我主人生了一个儿子；我主人把他一切所有的都给了他。
GEN|24|37|我主人叫我起誓说：‘不要为我儿子娶我所居住的 迦南 地的女子为妻。
GEN|24|38|你要往我父家、我本族那里去，为我的儿子娶妻。’
GEN|24|39|我对我主人说：‘恐怕那女子不肯跟我来。’
GEN|24|40|他就说：‘我所事奉的耶和华必要差遣他的使者与你同去，使你的道路亨通，你就可以在我父家、我本族那里，为我的儿子娶妻。
GEN|24|41|只要你到了我本族那里，我叫你起的誓就与你无关。他们若不把女子交给你，我叫你起的誓也与你无关。’
GEN|24|42|“我今日到了井旁，就说：‘耶和华—我主人 亚伯拉罕 的上帝啊，愿你使我所行的道路亨通。
GEN|24|43|看哪，我站在井旁，对哪一个出来打水的女子说：请你让我喝你瓶子里的一点水，
GEN|24|44|她若说：你只管喝，我也为你的骆驼打水；愿那女子作耶和华给我主人儿子所选定的妻子。’
GEN|24|45|“我心里的话还没有说完，看哪， 利百加 肩头上扛着水瓶出来，下到井旁打水。我对她说：‘请你给我水喝。’
GEN|24|46|她就急忙从肩头上拿下瓶子来，说：‘请喝！我也给你的骆驼喝。’我就喝了；她也给我的骆驼喝了。
GEN|24|47|我问她说：‘你是谁的女儿？’她说：‘我是 彼土利 的女儿， 彼土利 是 密迦 和 拿鹤 生的儿子。’我就把环子戴在她鼻子上，把镯子戴在她双手上。
GEN|24|48|然后我低头向耶和华敬拜，称颂耶和华—我主人 亚伯拉罕 的上帝，因为他引导我走合适的道路，使我得着我主人兄弟的孙女，给我主人的儿子为妻。
GEN|24|49|现在你们若愿以慈爱诚信待我主人，就告诉我；若不然，也告诉我，使我可以或向左，或向右。”
GEN|24|50|拉班 和 彼土利 回答说：“这事既然出于耶和华，我们不能向你说好说歹。
GEN|24|51|看哪， 利百加 就在你面前，可以将她带去，遵照耶和华所说的，给你主人的儿子为妻。”
GEN|24|52|亚伯拉罕 的仆人听见他们这些话，就向耶和华俯伏在地。
GEN|24|53|仆人拿出金器、银器和衣服送给 利百加 ，又将贵重的物品送给她哥哥和她母亲。
GEN|24|54|然后，仆人和随从的人才吃喝，并且住了一夜。早晨起来，仆人说：“请让我回我主人那里去吧。”
GEN|24|55|利百加 的哥哥和母亲说：“让她同我们再住几天，也许十天，然后她可以去。”
GEN|24|56|仆人对他们说：“耶和华既然使我道路亨通，你们就不要耽误我，请让我走，回我主人那里去吧！”
GEN|24|57|他们说：“我们把她叫来问问她 。”
GEN|24|58|他们就叫了 利百加 来，对她说：“你和这人同去吗？”她说：“我去。”
GEN|24|59|于是他们送他们的妹妹 利百加 和她的奶妈，同 亚伯拉罕 的仆人，以及随从他的人走了。
GEN|24|60|他们就为 利百加 祝福，对她说： “我们的妹妹啊， 愿你作千万人的母亲！ 愿你的后裔得着仇敌的城门！”
GEN|24|61|利百加 和她的女仆们起来，骑上骆驼，跟着那人去。仆人就带着 利百加 走了。
GEN|24|62|那时， 以撒 住在 尼革夫 。他刚从 庇耳．拉海．莱 回来。
GEN|24|63|傍晚时， 以撒 出来，到田间默想。他举目一看，看哪，来了一队骆驼。
GEN|24|64|利百加 举目看见 以撒 ，就急忙下了骆驼，
GEN|24|65|对那仆人说：“这从田间走来迎接我们的人是谁？”仆人说：“他是我的主人。” 利百加 就拿面纱盖住自己。
GEN|24|66|仆人把他所做的一切事都告诉 以撒 。
GEN|24|67|以撒 就领 利百加 进了母亲 撒拉 的帐棚，娶了她为妻，并且爱她。 以撒 自从母亲离世以后，这才得了安慰。
GEN|25|1|亚伯拉罕 再娶了一个妻子，名叫 基土拉 。
GEN|25|2|她为他生了 心兰 、 约珊 、 米但 、 米甸 、 伊施巴 和 书亚 。
GEN|25|3|约珊 生了 示巴 和 底但 。 底但 的子孙是 亚书利 族、 利都是 族和 利乌米 族。
GEN|25|4|米甸 的儿子是 以法 、 以弗 、 哈诺 、 亚比大 和 以勒大 。这些都是 基土拉 的子孙。
GEN|25|5|亚伯拉罕 把他一切所有的都给了 以撒 。
GEN|25|6|至于 亚伯拉罕 妾的儿子， 亚伯拉罕 趁着自己还活着的时候把财物分给他们，打发他们离开他的儿子 以撒 ，往东方去，直到东方之地。
GEN|25|7|这是 亚伯拉罕 一生的年日，他活了一百七十五年。
GEN|25|8|亚伯拉罕 寿高年迈，安享天年，息劳而终，归到他祖先 那里。
GEN|25|9|他两个儿子 以撒 、 以实玛利 把他安葬在 麦比拉 洞里。这洞在 幔利 的对面、 赫 人 琐辖 的儿子 以弗仑 的田中，
GEN|25|10|就是 亚伯拉罕 向 赫 人买的那块田。 亚伯拉罕 和他妻子 撒拉 都葬在那里。
GEN|25|11|亚伯拉罕 死了以后，上帝赐福给他的儿子 以撒 。 以撒 住在 庇耳．拉海．莱 附近。
GEN|25|12|这是 撒拉 的婢女、 埃及 人 夏甲 为 亚伯拉罕 生的儿子 以实玛利 的后代。
GEN|25|13|以实玛利 儿子们的名字，按着他们后代的名字如下： 以实玛利 的长子 尼拜约 ，又有 基达 、 亚德别 、 米比衫 、
GEN|25|14|米施玛 、 度玛 、 玛撒 、
GEN|25|15|哈大 、 提玛 、 伊突 、 拿非施 ，和 基底玛 。
GEN|25|16|这些都是 以实玛利 的儿子们。他们的村庄和营寨按着他们命名；他们作了十二族的族长。
GEN|25|17|以实玛利 一生的岁数是一百三十七岁，断气而死，归到他祖先那里。
GEN|25|18|他的子孙住在 哈腓拉 ，直到 埃及 东边的 书珥 ，向着 亚述 ，在他众弟兄的对面安顿下来 。
GEN|25|19|这是 亚伯拉罕 的儿子 以撒 的后代。 亚伯拉罕 生 以撒 。
GEN|25|20|以撒 四十岁时娶 利百加 为妻。 利百加 是 巴旦．亚兰 地的 亚兰 人 彼土利 的女儿，是 亚兰 人 拉班 的妹妹。
GEN|25|21|以撒 因他妻子不生育，就为她祈求耶和华。耶和华应允他的祈求，他的妻子 利百加 就怀了孕。
GEN|25|22|胎儿们在她腹中彼此相争，她就说：“若是如此，我为什么会这样呢 ？”她就去求问耶和华。
GEN|25|23|耶和华对她说： 两国在你腹中； 两族要从你身上分立。 这族必强于那族； 将来大的要服侍小的。
GEN|25|24|到了生产的日期，看哪，腹中是对双胞胎。
GEN|25|25|先出生的身体带红，浑身有毛，好像皮衣；他们就给他起名叫 以扫 。
GEN|25|26|随后， 以扫 的弟弟也出生，他的手抓住 以扫 的脚跟，因此给他起名叫 雅各 。两个儿子出生时， 以撒 六十岁。
GEN|25|27|两个孩子渐渐长大， 以扫 善于打猎，常在田野； 雅各 为人安静，常住在帐棚里。
GEN|25|28|以撒 爱 以扫 ，因为常吃他的野味； 利百加 却爱 雅各 。
GEN|25|29|有一天， 雅各 熬了汤， 以扫 从田野回来，疲惫不堪。
GEN|25|30|以扫 对 雅各 说：“我累死了，请你让我吃这红的，这红的汤吧！”因此 以扫 又叫 以东 。
GEN|25|31|雅各 说：“你今日把长子的名分卖给我吧。”
GEN|25|32|以扫 说：“看哪，我快要死了，这长子的名分对我有什么用呢？”
GEN|25|33|雅各 说：“你今日对我起誓吧。” 以扫 就向他起誓，把长子的名分卖给了 雅各 。
GEN|25|34|于是 雅各 把饼和豆汤给了 以扫 ， 以扫 吃喝以后，起来走了。这样， 以扫 轻看他长子的名分。
GEN|26|1|那地有了饥荒，不是 亚伯拉罕 的时候曾有过的那次饥荒， 以撒 就到 基拉耳 ， 非利士 人的王 亚比米勒 那里去。
GEN|26|2|耶和华向 以撒 显现，说：“你不要下 埃及 去，要住在我所指示你的地。
GEN|26|3|你要寄居在这地，我必与你同在，赐福给你，因为我要将这一切的地都赐给你和你的后裔。我必坚定我向你父亲 亚伯拉罕 所起的誓。
GEN|26|4|我要使你的后裔增多，好像天上的星，又要将这一切的地赐给你的后裔，并且地上的万国都必因你的后裔得福，
GEN|26|5|因为 亚伯拉罕 听从我的话，遵守我的吩咐、诫令、律例和教导。”
GEN|26|6|于是， 以撒 住在 基拉耳 。
GEN|26|7|那地方的人问起他的妻子，他就说：“她是我的妹妹。”原来他害怕说“我的妻子”。他想：“或许这地方的人会因 利百加 杀我，因为她容貌美丽。”
GEN|26|8|他在那里住了一段很长的日子。有一天， 非利士 人的王 亚比米勒 从窗户往外观看，看哪， 以撒 在抚爱他的妻子 利百加 。
GEN|26|9|亚比米勒 召 以撒 来，说：“看哪，她实在是你的妻子，你怎么说‘她是我的妹妹’呢？” 以撒 对他说：“因为我想，恐怕我会因她而死。”
GEN|26|10|亚比米勒 说：“你向我们做的是什么事呢？百姓中有一个人几乎要和你的妻子同寝，你就把我们陷在罪中了。”
GEN|26|11|于是 亚比米勒 命令众百姓说：“凡侵犯这个人，或他妻子的，必要把他处死。”
GEN|26|12|以撒 在那地耕种，那一年有百倍的收成。耶和华赐福给他，
GEN|26|13|他就发达，日渐昌盛，成了大富翁。
GEN|26|14|他有羊群牛群，又有许多仆人， 非利士 人就嫉妒他。
GEN|26|15|他父亲 亚伯拉罕 在世的时候，他父亲的仆人所挖的井， 非利士 人全都塞住，填满了土。
GEN|26|16|亚比米勒 对 以撒 说：“你离开我们去吧，因为你比我们强盛得多。”
GEN|26|17|以撒 就离开那里，在 基拉耳谷 支搭帐棚，住在那里。
GEN|26|18|他父亲 亚伯拉罕 在世的时候所挖的水井，在 亚伯拉罕 死后，都被 非利士 人塞住了， 以撒 就重新把井挖出来，仍照他父亲所取的名为它们命名。
GEN|26|19|以撒 的仆人在谷中挖井，就在那里得了一口活水井。
GEN|26|20|基拉耳 的牧人与 以撒 的牧人相争，说：“这水是我们的。” 以撒 就给那井起名叫 埃色 ，因为他们和他相争。
GEN|26|21|以撒 的仆人又挖了一口井，他们又为这井相争， 以撒 就给这井起名叫 西提拿 。
GEN|26|22|以撒 离开那里，又挖了一口井，他们不再为这井相争了，他就给那井起名叫 利河伯 。他说：“耶和华现在给我们宽阔之地，我们必在这地兴旺。”
GEN|26|23|以撒 从那里上 别是巴 去。
GEN|26|24|当夜耶和华向他显现，说：“我是你父亲 亚伯拉罕 的上帝。不要惧怕，因为我与你同在，要赐福给你，也要为我仆人 亚伯拉罕 的缘故，使你的后裔增多。”
GEN|26|25|以撒 就在那里筑了一座坛，求告耶和华的名，并且在那里支搭帐棚；他的仆人就在那里挖了一口井。
GEN|26|26|亚比米勒 同他的顾问 亚户撒 和他军队的元帅 非各 ，从 基拉耳 来到 以撒 那里。
GEN|26|27|以撒 对他们说：“你们既然恨我，赶我离开你们，为什么又到我这里来呢？”
GEN|26|28|他们说：“我们明明看见耶和华与你同在；因此就说，让我们双方彼此起誓，我们跟你立约，
GEN|26|29|使你不加害我们，正如我们未曾侵犯你，素来善待你，并且送你平平安安地走。你是蒙耶和华赐福的！”
GEN|26|30|以撒 为他们摆设宴席，他们就一起吃喝。
GEN|26|31|他们清早起来，彼此起誓。 以撒 送他们走，他们就平平安安地离开他去了。
GEN|26|32|那一天， 以撒 的仆人来，把挖井的消息告诉他，说：“我们得到水了。”
GEN|26|33|他就给那井起名叫 示巴 ，因此那城名叫 别是巴 ，直到今日。
GEN|26|34|以扫 四十岁的时候娶了 赫 人 比利 的女儿 犹滴 ，和 赫 人 以伦 的女儿 巴实抹 为妻。
GEN|26|35|她们使 以撒 和 利百加 心里愁烦。
GEN|27|1|以撒 年老，眼睛昏花，不能看见，就叫他大儿子 以扫 来，对他说：“我儿。” 以扫 对他说：“我在这里。”
GEN|27|2|他说：“看哪，我老了，不知道哪一天死。
GEN|27|3|现在拿你打猎的工具，就是箭囊和弓，到田野去为我打猎，
GEN|27|4|照我所爱的做成美味，拿来给我吃，好让我在未死之前为你祝福。”
GEN|27|5|以撒 对他儿子 以扫 说话的时候， 利百加 听见了。 以扫 往田野去打猎，要把猎物带回来。
GEN|27|6|利百加 就对她儿子 雅各 说：“看哪，我听见你父亲对你哥哥 以扫 说：
GEN|27|7|‘你去把猎物带回来，做成美味给我吃，让我在未死之前，在耶和华面前为你祝福。’
GEN|27|8|现在，我儿，你要听我的话，照我所吩咐你的，
GEN|27|9|到羊群里去，从那里牵两只肥美的小山羊来给我，我就照你父亲所爱的，把它们做成美味给他。
GEN|27|10|然后，你拿到你父亲那里给他吃，好让他在未死之前为你祝福。”
GEN|27|11|雅各 对他母亲 利百加 说：“看哪，我哥哥 以扫 浑身都有毛，我身上却是光滑的；
GEN|27|12|倘若父亲摸着我，我在他眼中就是骗子了。这样，我就自招诅咒，而不是祝福。”
GEN|27|13|他母亲对他说：“我儿，你所受的诅咒临到我身上吧！你只管听我的话，去牵小山羊来给我。”
GEN|27|14|他就去牵来，交给他母亲。他母亲就照他父亲所爱的，做成美味。
GEN|27|15|利百加 把大儿子 以扫 在家里最好的衣服给她小儿子 雅各 穿，
GEN|27|16|又用小山羊的皮包在 雅各 的手上和颈项光滑的地方，
GEN|27|17|就把所做的美味和饼交在她儿子 雅各 的手里。
GEN|27|18|雅各 来到他父亲那里，说：“我的父亲！”他说：“我在这里。我儿，你是谁？”
GEN|27|19|雅各 对他父亲说：“我是你的长子 以扫 。我已照你吩咐我的做了。请起来坐着，吃我的野味，你好为我祝福。”
GEN|27|20|以撒 对他儿子说：“我儿，你怎么这样快就找到了呢？”他说：“因为这是耶和华—你的上帝使我遇见的。”
GEN|27|21|以撒 对 雅各 说：“我儿，靠近一点，让我摸摸你，你真的是我的儿子 以扫 吗？”
GEN|27|22|雅各 就靠近他父亲 以撒 。 以撒 摸着他，说：“声音是 雅各 的声音，手却是 以扫 的手。”
GEN|27|23|以撒 认不出他来，因为他手上有毛，像他哥哥 以扫 的手一样。于是， 以撒 就为他祝福。
GEN|27|24|以撒 说：“你真的是我儿子 以扫 吗？”他说：“我是。”
GEN|27|25|以撒 说：“拿给我，让我吃我儿子的野味，我好为你祝福。” 雅各 拿给他，他就吃了，又拿酒给他，他也喝了。
GEN|27|26|他父亲 以撒 对他说：“我儿，靠近一点来亲我！”
GEN|27|27|他就近前亲吻父亲。他父亲一闻他衣服上的香气，就为他祝福，说： “看，我儿的香气 好像耶和华赐福之田地的香气。
GEN|27|28|愿上帝赐你天上的甘露， 地上的肥土， 和丰富的五谷新酒。
GEN|27|29|愿万民事奉你， 万族向你下拜。 愿你作你弟兄的主， 你母亲的儿子向你下拜。 诅咒你的，愿他受诅咒； 祝福你的，愿他蒙祝福。”
GEN|27|30|以撒 为 雅各 祝福完毕， 雅各 才从他父亲那里出来，他哥哥 以扫 正打猎回来。
GEN|27|31|以扫 也做了美味，拿来给他父亲，对他父亲说：“父亲，请起来，吃你儿子的野味，你好为我祝福。”
GEN|27|32|他父亲 以撒 对他说：“你是谁？”他说：“我是你的儿子，你的长子 以扫 。”
GEN|27|33|以撒 就大大战兢，说：“那么，是谁打了猎物拿来给我呢？你未来之前我已经吃了，也为他祝福了，他将来就必蒙福。”
GEN|27|34|以扫 听了他父亲的话，就大声痛哭，对他父亲说：“我父啊，求你也为我祝福！”
GEN|27|35|以撒 说：“你弟弟已经用诡计来把你的福分夺去了。”
GEN|27|36|以扫 说：“他名叫 雅各 ，岂不是这样吗？他欺骗了我两次：他先前夺了我长子的名分，看哪，他现在又夺了我的福分。” 以扫 又说：“你没有留下给我的祝福吗？”
GEN|27|37|以撒 回答 以扫 说：“看哪，我已立他作你的主，使他的弟兄都给他作仆人，并赐他五谷新酒可以养生。我儿，那么，现在我还能为你做什么呢？”
GEN|27|38|以扫 对他父亲说：“我父啊，你只有一个祝福吗？我父啊，求你也为我祝福！” 以扫 就放声而哭。
GEN|27|39|他父亲 以撒 回答说： “看哪，你所住的地方必缺乏肥沃的土地， 缺乏天上的甘露 。
GEN|27|40|你必倚靠刀剑度日， 又必服侍你的兄弟； 到你强盛的时候， 必从你颈项上挣开他的轭。
GEN|27|41|以扫 因他父亲给 雅各 的祝福，就怨恨 雅各 ，心里说：“为我父亲居丧的时候近了，到那时候，我要杀我的弟弟 雅各 。”
GEN|27|42|有人把 利百加 大儿子 以扫 的话告诉 利百加 ，她就派人去，叫了她小儿子 雅各 来，对他说：“看哪，你哥哥 以扫 想要杀你来泄恨。
GEN|27|43|现在，我儿，听我的话，起来，逃往 哈兰 ，到我哥哥 拉班 那里去，
GEN|27|44|同他住一段日子，直等到你哥哥的怒气消了。
GEN|27|45|等到你哥哥向你消了怒气，忘了你向他所做的事，我就派人去，把你从那里带回来。我何必在一天之内丧失你们二人呢？”
GEN|27|46|利百加 对 以撒 说：“我因这 赫 人的女子活得不耐烦了；倘若 雅各 也从本地女子中娶像这样的 赫 人女子为妻，我为什么要活着呢？”
GEN|28|1|以撒 叫了 雅各 来，为他祝福，并吩咐他说：“你不要娶 迦南 的女子为妻。
GEN|28|2|你起身往 巴旦．亚兰 去，到你外祖父 彼土利 的家，从你舅父 拉班 的女儿中娶一位作你的妻子。
GEN|28|3|愿全能的上帝赐福给你，使你生养众多，成为许多民族，
GEN|28|4|将应许 亚伯拉罕 的福赐给你和你的后裔，使你承受你所寄居的地为业，就是上帝赐给 亚伯拉罕 的地。”
GEN|28|5|以撒 送 雅各 走了， 雅各 就往 巴旦．亚兰 去，到 亚兰 人 彼土利 的儿子 拉班 那里， 拉班 是 利百加 的哥哥， 利百加 是 雅各 和 以扫 的母亲。
GEN|28|6|以扫 见 以撒 已经为 雅各 祝福，而且送他往 巴旦．亚兰 去，在那里娶妻，并且见 以撒 祝福 雅各 的时候吩咐他说：“不要娶 迦南 的女子为妻”，
GEN|28|7|又见 雅各 听从父母的话往 巴旦．亚兰 去了，
GEN|28|8|以扫 就看出他父亲 以撒 看 迦南 女子不顺眼。
GEN|28|9|于是他往 以实玛利 那里去，在两个妻子之外， 又娶了 玛哈拉 为妻，她是 亚伯拉罕 儿子 以实玛利 的女儿，是 尼拜约 的妹妹。
GEN|28|10|雅各 离开 别是巴 ，往 哈兰 去。
GEN|28|11|到了一个地方，因为已经日落，就在那里过夜。他拾起那地方的一块石头枕在头下，就躺在那地方。
GEN|28|12|他做梦，看哪，一个梯子立在地上，梯子的顶端直伸到天；看哪，上帝的使者在梯子上，上去下来。
GEN|28|13|看哪，耶和华站在梯子上面 ，说：“我是耶和华—你祖父 亚伯拉罕 的上帝， 以撒 的上帝。你现在躺卧之地，我要将它赐给你和你的后裔。
GEN|28|14|你的后裔必像地上的尘沙，必向东西南北开展；地上万族必因你和你的后裔得福。
GEN|28|15|看哪，我必与你同在，无论你往哪里去，我必保佑你，领你归回这地。我总不离弃你，直到我实现了对你所说的话。”
GEN|28|16|雅各 睡醒了，说：“耶和华真的在这里，我竟不知道！”
GEN|28|17|他就惧怕，说：“这地方何等可畏！这不是别的，是上帝的殿，是天的门。”
GEN|28|18|雅各 清早起来，拿起枕在头下的石头，立作柱子，浇油在上面。
GEN|28|19|他给那地方起名叫 伯特利 ；那地方原先名叫 路斯 。
GEN|28|20|雅各 许愿说：“上帝若与我同在，在我所行的路上保佑我，给我食物吃，衣服穿，
GEN|28|21|使我平平安安回到我父亲的家，我就必以耶和华为我的上帝。
GEN|28|22|我所立为柱子的这块石头必作上帝的殿；凡你所赐给我的，我必将十分之一献给你。”
GEN|29|1|雅各 起行，到了东方人之地。
GEN|29|2|他观看，看哪，田间有一口井，看哪，有三群羊卧在井旁；因为人都取那井里的水给羊喝。井口上的那块石头很大。
GEN|29|3|羊群都在那里聚集，人就把石头移开井口，取水给羊喝，然后又把石头放回井口原处。
GEN|29|4|雅各 对他们说：“弟兄们，你们从哪里来？”他们说：“我们是从 哈兰 来的。”
GEN|29|5|他对他们说：“你们认识 拿鹤 的孙子 拉班 吗？”他们说：“我们认识。”
GEN|29|6|雅各 对他们说：“他平安吗？”他们说：“平安。看哪，他女儿 拉结 和羊一起来了。”
GEN|29|7|雅各 说：“看哪，日正当中，不是牲畜聚集的时候。你们取水给羊喝，再去牧放吧！”
GEN|29|8|他们说：“我们不能这样，必须等所有的羊群聚集，人把石头移开井口，我们才可以取水给羊喝。”
GEN|29|9|雅各 正和他们说话的时候， 拉结 和她父亲的羊来了，因为她是牧羊的。
GEN|29|10|雅各 看见他舅父 拉班 的女儿 拉结 和舅父 拉班 的羊群，就上前把石头移开井口，取水给舅父 拉班 的羊喝。
GEN|29|11|雅各 亲了 拉结 ，就放声大哭。
GEN|29|12|雅各 告诉 拉结 ，自己是她父亲的亲戚 ，是 利百加 的儿子。 拉结 就跑去告诉她父亲。
GEN|29|13|拉班 听见外甥 雅各 的消息，就跑去迎接他，抱着他，亲他，带他到自己的家。 雅各 把这一切的事告诉 拉班 。
GEN|29|14|拉班 对他说：“你实在是我的骨肉。” 雅各 就和他同住了一个月。
GEN|29|15|拉班 对 雅各 说：“虽然你是我的亲戚，怎么可以让你白白服事我呢？告诉我，你要什么作工资呢？”
GEN|29|16|拉班 有两个女儿，大的名叫 利亚 ，小的名叫 拉结 。
GEN|29|17|利亚 的双眼无神， 拉结 却长得美貌秀丽。
GEN|29|18|雅各 爱 拉结 ，就说：“我愿为你的小女儿 拉结 服事你七年。”
GEN|29|19|拉班 说：“我把她给你，胜过给别人，你与我同住吧！”
GEN|29|20|雅各 就为 拉结 服事了七年；他因为爱 拉结 ，就看这七年如同几天。
GEN|29|21|雅各 对 拉班 说：“日期已经满了，请把我的妻子给我，我好与她同房。”
GEN|29|22|拉班 就摆设宴席，请了当地所有的人。
GEN|29|23|到了晚上， 拉班 带女儿 利亚 来送给 雅各 ， 雅各 就与她同房。
GEN|29|24|拉班 也把自己的婢女 悉帕 给女儿 利亚 作婢女。
GEN|29|25|到了早晨，看哪，她是 利亚 ， 雅各 对 拉班 说：“你向我做的是什么事呢？我服事你，不是为 拉结 吗？你为什么欺骗我呢？”
GEN|29|26|拉班 说：“大女儿还没有给人就先把小女儿给人，我们这地方没有这样的规矩。
GEN|29|27|你先为这个满了七日，我们就把那个也给你，不过你要另外再服事我七年。”
GEN|29|28|雅各 就这样做了。满了 利亚 的七日， 拉班 就把女儿 拉结 给 雅各 为妻。
GEN|29|29|拉班 又把自己的婢女 辟拉 给女儿 拉结 作婢女。
GEN|29|30|雅各 也与 拉结 同房，并且爱 拉结 胜过爱 利亚 ，于是他又服事了 拉班 七年。
GEN|29|31|耶和华见 利亚 失宠 ，就使她生育， 拉结 却不生育。
GEN|29|32|利亚 怀孕生子，给他起名叫 吕便 ，因为她说：“耶和华看见我的苦情，如今我的丈夫必爱我。”
GEN|29|33|她又怀孕生子，给他起名叫 西缅 ，说：“耶和华因为听见我失宠，所以又赐给我这个儿子。”
GEN|29|34|她又怀孕生子，说：“我给丈夫生了三个儿子，现在，这次他必亲近我了。”因此， 雅各 给他起名叫 利未 。
GEN|29|35|她又怀孕生子，说：“这次我要赞美耶和华。”因此给他起名叫 犹大 。于是她停了生育。
GEN|30|1|拉结 见自己不给 雅各 生孩子，就嫉妒她姊姊，对 雅各 说：“你给我孩子，不然，让我死了吧。”
GEN|30|2|雅各 对 拉结 生气，说：“是我代替上帝使你生不出孩子的吗？”
GEN|30|3|拉结 说：“看哪，我的使女 辟拉 在这里，你可以与她同房，使她生子归在我膝下，我也可以藉着她得孩子 。”
GEN|30|4|拉结 就把她的婢女 辟拉 给丈夫为妾， 雅各 与她同房。
GEN|30|5|辟拉 怀孕，为 雅各 生了一个儿子。
GEN|30|6|拉结 给他起名叫 但 ，说：“上帝为我伸冤，也听了我的声音，赐给我一个儿子。”
GEN|30|7|拉结 的婢女 辟拉 又怀孕，为 雅各 生了第二个儿子。
GEN|30|8|拉结 给他起名叫 拿弗他利 ，说：“我与我姊姊大大较力，并且得胜了。”
GEN|30|9|利亚 见自己停了生育，就把她的婢女 悉帕 给 雅各 为妾。
GEN|30|10|利亚 的婢女 悉帕 为 雅各 生了一个儿子。
GEN|30|11|利亚 给他起名叫 迦得 ，说：“真是幸运！”
GEN|30|12|利亚 的婢女 悉帕 又为 雅各 生了第二个儿子。
GEN|30|13|利亚 给他起名叫 亚设 ，说：“我真有福啊，众女子都要称我有福。”
GEN|30|14|收割麦子的时候， 吕便 到田里去，找到曼陀罗草 ，就拿给他的母亲 利亚 。 拉结 对 利亚 说：“请你给我一些你儿子的曼陀罗草吧。”
GEN|30|15|利亚 对她说：“你夺走了我的丈夫还是小事吗？你还要夺取我儿子的曼陀罗草吗？” 拉结 说：“今夜他可以与你同寝，来交换你儿子的曼陀罗草。”
GEN|30|16|到了晚上， 雅各 从田里回来， 利亚 出来迎接他，说：“你要与我同寝，因为我真的用我儿子的曼陀罗草把你雇下了。”那一夜， 雅各 就与她同寝。
GEN|30|17|上帝应允了 利亚 ，她就怀孕，为 雅各 生了第五个儿子。
GEN|30|18|利亚 给他起名叫 以萨迦 ，说：“上帝给了我工价，因为我把婢女给了我的丈夫。”
GEN|30|19|利亚 又怀孕，为 雅各 生了第六个儿子。
GEN|30|20|利亚 给他起名叫 西布伦 ，说：“上帝赐给我厚礼了；这次，我丈夫必看重我，因为我为他生了六个儿子。”
GEN|30|21|后来她又生了一个女儿，给她起名叫 底拿 。
GEN|30|22|上帝顾念 拉结 ，应允她，使她能生育。
GEN|30|23|拉结 怀孕生子，说：“上帝除去了我的羞耻。”
GEN|30|24|拉结 就给他起名叫 约瑟 ，说：“愿耶和华再增添一个儿子给我。”
GEN|30|25|拉结 生 约瑟 之后， 雅各 对 拉班 说：“请让我走，回到我的本乡本土去。
GEN|30|26|请你把我服事你所得的妻子和孩子给我，让我走吧！我怎样服事你，你都知道。”
GEN|30|27|拉班 对他说：“愿你看得起我，因我占卜得知，耶和华赐福给我是因你的缘故。”
GEN|30|28|又说：“请为我定你的工资，我就给你。”
GEN|30|29|雅各 对他说：“我怎样服事你，你的牲畜在我这里变得怎样，你都知道。
GEN|30|30|我未来以前，你拥有的很少，现在却已大量增加，因为耶和华随着我的脚步赐福给你。现在，我到什么时候才可以成家立业呢？”
GEN|30|31|拉班 说：“我该给你什么呢？” 雅各 说：“你什么也不必给我，只要你为我做这件事，我就继续牧放你的羊群。
GEN|30|32|今天我要走遍你的羊群，把绵羊中凡有点的、有斑的，和小绵羊中凡是黑色的羊；以及山羊中凡有斑的、有点的，都从那里挑出来，作为我的工资。
GEN|30|33|以后你来当面查看我的工资，任何我这里的山羊不是有点有斑的，小绵羊不是黑色的，就算是我偷的。这就可以证明我是正直的。”
GEN|30|34|拉班 说：“看哪，就照你所说的做吧。”
GEN|30|35|当日， 拉班 把有纹的、有斑的公山羊，一切有点的、有斑的、有少许白色 的母山羊，以及小绵羊中所有黑色的 ，都挑出来，交在他儿子们的手里，
GEN|30|36|又使自己和 雅各 相隔三天的路程。 雅各 就牧放 拉班 其余的羊。
GEN|30|37|雅各 拿杨树、杏树、枫树的嫩枝，把皮剥出白色的条纹，使枝子露出白色来。
GEN|30|38|他把剥了皮的枝子对着羊群，插在羊喝水的水沟和水槽里。羊来喝水的时候，它们彼此交配。
GEN|30|39|羊对着枝子交配，就生下有纹的、有点的、有斑的来。
GEN|30|40|雅各 把小绵羊分出来，让羊对着 拉班 羊群中有纹的和所有黑色的。于是他把自己的羊群分开，不叫它们和 拉班 的羊混在一起。
GEN|30|41|当肥壮的羊交配的时候， 雅各 就把枝子插在水沟里，使羊对着枝子交配。
GEN|30|42|可是当瘦弱的羊交配的时候，他就不插枝子。这样，瘦弱的就归 拉班 ，肥壮的就归 雅各 。
GEN|30|43|于是这人极其发达，拥有许多的羊群、奴仆、婢女、骆驼和驴。
GEN|31|1|雅各 听见 拉班 儿子们的话，说：“ 雅各 把我们父亲所有的都夺去了！他从我们父亲所拥有的获得这一切的财富。”
GEN|31|2|雅各 见 拉班 的脸色，看哪，待他不如从前了。
GEN|31|3|耶和华对 雅各 说：“你要回你祖先之地，到你本族那里去，我必与你同在。”
GEN|31|4|雅各 就派人叫 拉结 和 利亚 到田野他的羊群那里去，
GEN|31|5|对她们说：“我看你们父亲待我的脸色不如从前了，但我父亲的上帝向来与我同在。
GEN|31|6|你们也知道，我尽了全力服事你们的父亲。
GEN|31|7|可是你们的父亲欺骗我，十次更改我的工资，但上帝不容许他害我。
GEN|31|8|他若说：‘有点的归给你作工资’，羊群所生的都是有点的；他若说：‘有纹的归给你作工资’，羊群所生的都是有纹的。
GEN|31|9|这样，上帝把你们父亲的牲畜拿来赐给我了。
GEN|31|10|“羊群交配的时候，我在梦中举目一看，看哪，跳母羊的公羊都是有纹的、有点的、有花斑的。
GEN|31|11|上帝的使者在梦中呼叫我说：‘ 雅各 。’我说：‘我在这里。’
GEN|31|12|他说：‘你举目观看，跳母羊的公羊都是有纹的、有点的、有花斑的。 拉班 向你所做的一切，我都看见了。
GEN|31|13|我是 伯特利 的上帝；你曾在那里用油膏过柱子，向我许过愿。现在你起来，离开这地，回你本族之地去吧！’”
GEN|31|14|拉结 和 利亚 回答 雅各 说：“在我们父亲家里还有我们可分得的产业吗？
GEN|31|15|我们不是被他看作外人吗？因为他卖了我们，还吞吃了我们的银钱。
GEN|31|16|上帝从我们父亲所拿走的一切财物，都是我们和我们孩子的。现在，凡上帝所吩咐你的，你只管去做吧！”
GEN|31|17|雅各 起来，叫他的孩子和妻子都骑上骆驼，
GEN|31|18|又赶着他一切的牲畜和他所得的一切财物，就是他在 巴旦．亚兰 所得的，他拥有的牲畜 ，往 迦南 地他父亲 以撒 那里去了。
GEN|31|19|当时 拉班 去剪羊毛， 拉结 偷了他父亲家中的神像。
GEN|31|20|雅各 瞒住 亚兰 人 拉班 ，不通知他就逃走了。
GEN|31|21|雅各 带着他所有的逃走了；他起程，渡过 大河 ，面向着 基列山 。
GEN|31|22|到第三天，有人告诉 拉班 ， 雅各 逃跑了。
GEN|31|23|拉班 带着他的弟兄们去追他，追了七天，就在 基列山 追上了。
GEN|31|24|夜间，上帝来到 亚兰 人 拉班 那里，在梦中对他说：“你要小心，不可对 雅各 说好说歹。”
GEN|31|25|拉班 追上 雅各 。 雅各 在山上支搭帐棚； 拉班 和他的弟兄们也在 基列山 上支搭帐棚。
GEN|31|26|拉班 对 雅各 说：“你做的是什么事呢？你瞒着我把我的女儿们带走，好像用刀剑掳去一般。
GEN|31|27|你为什么暗暗地逃跑，瞒着我，不通知我一声，叫我可以欢乐、唱歌、击鼓、弹琴送你回去呢？
GEN|31|28|为什么不容许我与外孙和女儿吻别呢？你现在所做的真是愚蠢！
GEN|31|29|我的手本有能力害你，只是你父亲的上帝昨夜对我说：‘你要小心，不可对 雅各 说好说歹。’
GEN|31|30|现在你既然这么想念你的父家，不得不去，为什么又偷了我的神明呢？”
GEN|31|31|雅各 回答 拉班 说：“因为我害怕，我想，恐怕你把你的女儿从我这里夺走。
GEN|31|32|至于你的神明，你若在谁那里搜出来，就不让谁活。当着我们弟兄面前，你认一认在我这里有什么东西是你的，你就拿去吧。”原来 雅各 并不知道 拉结 偷了神明。
GEN|31|33|拉班 进了 雅各 、 利亚 ，以及两个使女的帐棚，却没有找到，就从 利亚 的帐棚出来，进入 拉结 的帐棚。
GEN|31|34|拉结 拿了神像，藏在骆驼的鞍子里，自己坐在上面。 拉班 搜遍了那帐棚，并没有找到。
GEN|31|35|拉结 对她父亲说：“请我主不要生气，因为我恰有月事，不能在你面前起来。” 拉班 搜寻，却找不到神像。
GEN|31|36|于是 雅各 发怒，斥责 拉班 。 雅各 对 拉班 说：“我有什么过犯，有什么罪恶，你竟这样火速地追我？
GEN|31|37|你搜遍了我一切的物件，你找到什么呢？可以放在你我弟兄面前，叫他们在我们两个之间评评理。
GEN|31|38|我在你那里这二十年，你的母绵羊、母山羊没有掉过胎。你羊群中的公绵羊，我没有吃过；
GEN|31|39|被野兽撕裂的，我没有带来给你，是我自己赔偿的。无论是白日被偷的，或是黑夜被偷的，你都从我手中索取。
GEN|31|40|我常常白日受尽炎热，黑夜受尽寒霜，不得合眼入睡。
GEN|31|41|我这二十年在你家里，为你两个女儿服事了你十四年，为你的羊群服事了你六年，你却十次更改我的工资。
GEN|31|42|若不是我父亲 以撒 所敬畏的上帝，就是 亚伯拉罕 的上帝与我同在，你如今必定打发我空手而去。上帝看见我的苦情和我手的辛劳，就在昨夜责备了你。”
GEN|31|43|拉班 回答 雅各 说：“这两个女儿是我的女儿，这些孩子是我的孩子，这些羊群也都是我的羊群；凡你所看见的都是我的。我的女儿和她们所生的孩子，我今日还能对他们做什么呢？
GEN|31|44|现在，来吧！让我和你立约，作你我之间的证据。”
GEN|31|45|雅各 就拿一块石头立作柱子，
GEN|31|46|对弟兄们说：“大家来堆积石头。”他们拿石头堆成一堆，于是在那里，在石堆旁边吃喝。
GEN|31|47|拉班 称那石堆为 伊迦尔．撒哈杜他 ， 雅各 却称那石堆为 迦累得 。
GEN|31|48|拉班 说：“今日这石堆成为你我之间的证据。”因此这地方名叫 迦累得 ，
GEN|31|49|又叫 米斯巴 ，因为他说：“我们彼此离别以后，愿耶和华在你我中间鉴察 。
GEN|31|50|你若苦待我的女儿，或在我的女儿以外另娶妻，虽没有人在场，你看，有上帝在你我中间作证。”
GEN|31|51|拉班 又对 雅各 说：“看哪，这石堆，看哪，这柱子，是我在你我中间所立的。
GEN|31|52|这石堆是证据，这柱子也是证据。我必不越过这石堆去害你；你也不可越过这石堆和柱子来害我。
GEN|31|53|愿 亚伯拉罕 的上帝和 拿鹤 的上帝，就是他们父亲的上帝 ，在你我中间判断。” 雅各 就指着他父亲 以撒 所敬畏的上帝起誓，
GEN|31|54|又在山上献祭，请弟兄们来吃饭。他们吃了饭，就在山上过夜。
GEN|31|55|拉班 清早起来，与他外孙和女儿亲吻，为他们祝福，就回到自己的地方去了。
GEN|32|1|雅各 继续行路，上帝的使者遇见他。
GEN|32|2|雅各 看见他们就说：“这是上帝的军营。”于是给那地方起名叫 玛哈念 。
GEN|32|3|雅各 派使者在他前面到 西珥 地，就是 以东 地他哥哥 以扫 那里。
GEN|32|4|他吩咐他们说：“你们要对我主 以扫 说：‘你的仆人 雅各 这样说：我在 拉班 那里寄居，延迟到如今。
GEN|32|5|我有牛、驴、羊群、奴仆、婢女，现在派人来报告我主，为了要在你眼前蒙恩。’”
GEN|32|6|使者回到 雅各 那里，说：“我们到了你哥哥 以扫 那里。他正迎着你来，并且有四百人和他一起。”
GEN|32|7|雅各 就很惧怕，而且愁烦。他把跟他同行的人和羊群、牛群、骆驼分成两队，
GEN|32|8|说：“ 以扫 若来击杀其中一队，剩下的另一队还可以逃脱。”
GEN|32|9|雅各 说：“耶和华—我祖父 亚伯拉罕 的上帝，我父亲 以撒 的上帝啊，你曾对我说：‘回你本地本族去，我要厚待你。’
GEN|32|10|你向仆人所施的一切慈爱和信实，我一点也不配得。我先前只用我的一根杖过这 约旦河 ，如今我却成了两队。
GEN|32|11|求你救我脱离我哥哥的手，脱离 以扫 的手，因为我怕他来杀我，连母亲和儿女都不放过。
GEN|32|12|你曾说：‘我必定厚待你，使你的后裔如同海边的沙，多得不可胜数。’”
GEN|32|13|当夜， 雅各 在那里住宿，就从他手中所拥有的拿礼物要送给他哥哥 以扫 ，
GEN|32|14|就是二百只母山羊、二十只公山羊、二百只母绵羊、二十只公绵羊、
GEN|32|15|三十匹哺乳的母骆驼和它们的小骆驼、四十头母牛、十头公牛、二十匹母驴和十匹公驴。
GEN|32|16|他把每种牲畜各分一群，交在仆人手中，对仆人说：“你们要在我的前头过去，使群和群之间保持一段距离”。
GEN|32|17|他又吩咐领头的人说：“我哥哥 以扫 遇见你的时候，问你说：‘你是谁的人？要往哪里去？你前面这些是谁的？’
GEN|32|18|你就说：‘是你仆人 雅各 的，是送给我主 以扫 的礼物。看哪，他自己也在我们后面。’”
GEN|32|19|他又吩咐第二、第三和所有赶畜群的人说：“你们遇见 以扫 的时候要照这样的话对他说，
GEN|32|20|你们还要说：‘看哪，你仆人 雅各 在我们后面。’”因 雅各 说：“我藉着在我前面送去的礼物给他面子，然后再见他的面，或许他会宽容我。”
GEN|32|21|于是礼物在他前面过去了；那夜， 雅各 在营中住宿。
GEN|32|22|他夜间起来，带着两个妻子，两个婢女和十一个孩子，过了 雅博 渡口。
GEN|32|23|他带着他们，送他们过河，他所有的一切也都过去，
GEN|32|24|只剩下 雅各 一人。有一个人来和他摔跤，直到黎明。
GEN|32|25|那人见自己胜不过他，就摸了他的大腿窝一下。 雅各 的大腿窝就在和那人摔跤的时候扭了。
GEN|32|26|那人说：“天快亮了，让我走吧！” 雅各 说：“你不给我祝福，我就不让你走。”
GEN|32|27|那人说：“你叫什么名字？”他说：“ 雅各 。”
GEN|32|28|那人说：“你的名字不要再叫 雅各 ，要叫 以色列 ，因为你与上帝和人较力，都得胜了。”
GEN|32|29|雅各 问他说：“请告诉我你的名字。”那人说：“何必问我的名字呢？”于是他在那里为 雅各 祝福。
GEN|32|30|雅各 就给那地方起名叫 毗努伊勒 ，说：“我面对面见了上帝，我的性命仍得保全。”
GEN|32|31|太阳刚出来的时候， 雅各 经过 毗努伊勒 ，他的大腿就瘸了。
GEN|32|32|因此， 以色列 人不吃大腿窝的筋，直到今日，因为那人摸了 雅各 大腿窝的筋。
GEN|33|1|雅各 举目观看，看哪， 以扫 来了，有四百人和他一起。 雅各 就把孩子们分开交给 利亚 、 拉结 和两个婢女。
GEN|33|2|他叫两个婢女和她们的孩子走在前头， 利亚 和她的孩子跟在后面，而 拉结 和 约瑟 在最后。
GEN|33|3|他自己却走到他们前面，一连七次俯伏在地才挨近他哥哥。
GEN|33|4|以扫 跑来迎接他，将他抱住，伏在他的颈项上亲他，他们都哭了。
GEN|33|5|以扫 举目看见妇人和孩子，就说：“这些和你一起的是谁呢？” 雅各 说：“这些孩子是上帝施恩给你仆人的。”
GEN|33|6|于是两个婢女和她们的孩子前来下拜，
GEN|33|7|利亚 和她的孩子也前来下拜，随后 约瑟 和 拉结 也前来下拜。
GEN|33|8|以扫 说：“我所遇见的这些畜群是什么意思呢？” 雅各 说：“是为了要在我主眼前蒙恩。”
GEN|33|9|以扫 说：“弟弟啊，我的已经够了，你的你自己留着吧！”
GEN|33|10|雅各 说：“不，我若在你眼前蒙恩，就请你从我手里收下这礼物；因为我见了你的面，如同见了上帝的面，并且你也宽容了我。
GEN|33|11|请你收下我带来给你的礼物，因为上帝恩待我，使我一切都充足。” 雅各 再三求他，他才收下。
GEN|33|12|以扫 说：“让我们起身前行，我和你一起走吧。”
GEN|33|13|雅各 对他说：“我主知道孩子们还年幼娇嫩，我的牛羊也正在哺乳中，只要催赶一天，群羊都会死了。
GEN|33|14|请我主在仆人前面先走，我要按着在我面前的牲畜和孩子的步伐慢慢前进，直走到 西珥 我主那里。”
GEN|33|15|以扫 说：“让我把跟随我的人留几个在你这里。” 雅各 说：“何必这样呢？只要能在我主眼前蒙恩就够了。”
GEN|33|16|于是， 以扫 当日起行，回 西珥 去了。
GEN|33|17|雅各 就往 疏割 去，在那里为自己盖房屋，又为牲畜搭棚，因此那地方叫 疏割 。
GEN|33|18|雅各 从 巴旦．亚兰 平安地回到 迦南 地的 示剑城 ，他在城的前面支搭帐棚。
GEN|33|19|他用一百可锡塔 从 示剑 的父亲 哈抹 的众子手中买了搭帐棚的那块地。
GEN|33|20|雅各 在那里筑了一座坛，起名叫 伊利．伊罗伊．以色列 。
GEN|34|1|利亚 给 雅各 所生的女儿 底拿 出去，要探望那地的女子们。
GEN|34|2|那地的族长 希未 人 哈抹 的儿子 示剑 看见她，就拉住她，与她同寝，玷辱了她。
GEN|34|3|示剑 的心喜欢 雅各 的女儿 底拿 ，爱上这少女，甜言蜜语地安慰她。
GEN|34|4|示剑 对他父亲 哈抹 说：“求你为我聘这女孩为妻。”
GEN|34|5|雅各 听见 示剑 污辱了他的女儿 底拿 。那时他的儿子们正和牲畜在田野， 雅各 就沉默，等他们回来。
GEN|34|6|示剑 的父亲 哈抹 出来，到 雅各 那里，要和他讲话。
GEN|34|7|雅各 的儿子们听见这事，就从田野回来，人人悲愤，十分恼怒，因 示剑 在 以色列 中做了丑事，与 雅各 的女儿同寝，这本是不该做的事。
GEN|34|8|哈抹 和他们谈话，说：“我儿子 示剑 的心喜欢你们家的女儿，请你们把她嫁给我的儿子。
GEN|34|9|你们与我们彼此结亲；你们可以把你们家的女儿嫁给我们，也可以娶我们家的女儿。
GEN|34|10|你们与我们同住吧！这地都在你们面前，只管在这里居住，做买卖，置产业。”
GEN|34|11|示剑 对女子的父亲和兄弟们说：“愿你们看得起我，你们向我要什么，我必给你们，
GEN|34|12|无论向我要多贵重的聘金和礼物，我必照你们所说的给你们，只要你们将这少女嫁给我。”
GEN|34|13|雅各 的儿子们因 示剑 污辱了他们的妹妹 底拿 ，就用诡诈的话回答 示剑 和他父亲 哈抹 ，
GEN|34|14|对他们说：“我们不能做这样的事，把我们的妹妹嫁给没有受割礼的人为妻，因为那是我们的羞耻。
GEN|34|15|惟有一个条件，我们才答应你们，就是你们所有的男丁都要受割礼，和我们一样，
GEN|34|16|我们就把我们家的女儿嫁给你们，也娶你们家的女儿；我们就与你们同住，大家成为一族人。
GEN|34|17|倘若你们不听从我们受割礼，我们就带我们家的女儿走了。”
GEN|34|18|这些话在 哈抹 和他儿子 示剑 的眼中看为美。
GEN|34|19|那年轻人毫不迟延做这事，因为他爱上了 雅各 的女儿；他在他父亲家中也是最受人尊重的。
GEN|34|20|哈抹 和他儿子 示剑 到他们的城门口，对城里的人讲说：
GEN|34|21|“这些人对我们友善，不如允许他们在这地居住，做买卖；看哪，这地宽阔，足以容纳他们。我们可以娶他们家的女儿，也可以把我们家的女儿嫁给他们。
GEN|34|22|惟有一个条件，这些人才答应和我们同住，成为一族人，就是我们中间所有的男丁都要受割礼，和他们一样。
GEN|34|23|他们的牲畜、财物和一切的牲口岂不都归给我们吗？只要答应他们，他们就与我们同住。”
GEN|34|24|凡从城门出入的人都听从了 哈抹 和他儿子 示剑 的话。于是，凡从城门出入的男丁都受了割礼。
GEN|34|25|到第三天，他们正疼痛的时候， 雅各 的两个儿子，就是 底拿 的哥哥 西缅 和 利未 ，各拿刀剑，不动声色地来到城中，把所有的男丁都杀了，
GEN|34|26|又用刀杀了 哈抹 和他儿子 示剑 ，把 底拿 从 示剑 家里带走，就离开了。
GEN|34|27|雅各 的儿子们因为他们的妹妹受污辱，就来到被杀的人那里，洗劫那城，
GEN|34|28|夺走了他们的羊群、牛群和驴，以及城里和田间所有的；
GEN|34|29|又俘掳抢劫他们一切的财物、孩童、妇女，以及房屋中所有的。
GEN|34|30|雅各 对 西缅 和 利未 说：“你们连累了我，使我在这地的居民中，就是在 迦南 人和 比利洗 人中坏了名声。我的人丁稀少，他们必聚集来击杀我，我和全家的人都要被灭绝。”
GEN|34|31|他们却说：“他岂可待我们的妹妹如同妓女呢？”
GEN|35|1|上帝对 雅各 说：“起来！上 伯特利 去，住在那里。在那里筑一座坛给上帝，就是你逃避你哥哥 以扫 的时候向你显现的上帝。”
GEN|35|2|雅各 就对他家中的人，以及所有和他一起的人说：“除掉你们中间外邦的神明，要自洁，更换衣服。
GEN|35|3|我们要起来，上 伯特利 去，在那里我要筑一座坛给上帝，就是在我遭难的日子应允我，在我行走的路上与我同在的上帝。”
GEN|35|4|他们就把手中所有外邦的神明和自己耳朵上的环子交给 雅各 ； 雅各 把它们埋在 示剑 那里的橡树下。
GEN|35|5|他们起行。上帝使周围城镇的人都惊恐，就不追赶 雅各 的儿子们了。
GEN|35|6|于是 雅各 和所有与他一起的人到了 迦南 地的 路斯 ，就是 伯特利 。
GEN|35|7|他在那里筑了一座坛，给那地方起名叫 伊勒．伯特利 ，因为他逃避他哥哥的时候，上帝曾在那里向他显现。
GEN|35|8|利百加 的奶妈 底波拉 死了，葬在 伯特利 下边的橡树下；那棵树名叫 亚伦．巴古 。
GEN|35|9|雅各 从 巴旦．亚兰 回来，上帝又向他显现，赐福给他。
GEN|35|10|上帝对他说：“你的名原是 雅各 ，从今以后不要再叫 雅各 ，你的名要叫 以色列 。”于是，上帝就叫他的名为 以色列 。
GEN|35|11|上帝又对他说：“我是全能的上帝；你要生养众多，将来有一国和许多的国从你而来，又有许多君王从你生出 。
GEN|35|12|至于我赐给 亚伯拉罕 和 以撒 的地，我必赐给你；我必赐这地给你的后裔。”
GEN|35|13|上帝就从与 雅各 说话的那地方升上去了。
GEN|35|14|雅各 就在上帝与他说话的地方立了一根柱子，就是石柱，在它上面献浇酒祭，又浇油。
GEN|35|15|雅各 就给上帝与他说话的那地方起名叫 伯特利 。
GEN|35|16|他们从 伯特利 起行，到 以法他 还有一段路程， 拉结 生产，生得十分艰难。
GEN|35|17|她生得十分艰难的时候，接生婆对她说：“不要怕，你又要有一个儿子了。”
GEN|35|18|她快要死，还有一口气的时候，就给她儿子起名叫 便．俄尼 ；他父亲却给他起名叫 便雅悯 。
GEN|35|19|拉结 死了，葬在往 以法他 的路旁； 以法他 就是 伯利恒 。
GEN|35|20|雅各 在她的坟上立了一块碑，就是 拉结 的墓碑，到今日还在。
GEN|35|21|以色列 起行，在 以得台 的那一边支搭帐棚。
GEN|35|22|以色列 住在那地的时候， 吕便 去与他父亲的妾 辟拉 同寝， 以色列 也听见了这件事 。 雅各 共有十二个儿子。
GEN|35|23|利亚 的儿子是 雅各 的长子 吕便 ，还有 西缅 、 利未 、 犹大 、 以萨迦 、 西布伦 。
GEN|35|24|拉结 的儿子是 约瑟 、 便雅悯 。
GEN|35|25|拉结 的婢女 辟拉 的儿子是 但 、 拿弗他利 。
GEN|35|26|利亚 的婢女 悉帕 的儿子是 迦得 、 亚设 。这是 雅各 在 巴旦．亚兰 所生的儿子。
GEN|35|27|雅各 来到他父亲 以撒 那里，到了 幔利 ， 基列．亚巴 ，就是 希伯仑 ，是 亚伯拉罕 和 以撒 寄居的地方。
GEN|35|28|以撒 共活了一百八十年。
GEN|35|29|以撒 年纪老迈，安享天年，息劳而终，归到他祖先 那里。他两个儿子 以扫 和 雅各 把他安葬了。
GEN|36|1|这是 以扫 的后代， 以扫 就是 以东 。
GEN|36|2|以扫 娶 迦南 的女子为妻，就是 赫 人 以伦 的女儿 亚大 和 希未 人 祭便 的孙女， 亚拿 的女儿 阿何利巴玛 ，
GEN|36|3|又娶了 以实玛利 的女儿， 尼拜约 的妹妹 巴实抹 。
GEN|36|4|亚大 为 以扫 生了 以利法 ； 巴实抹 生了 流珥 ；
GEN|36|5|阿何利巴玛 生了 耶乌施 、 雅兰 、 可拉 。这些都是 以扫 的儿子，是在 迦南 地生的。
GEN|36|6|以扫 带着他的妻子、儿女和家中所有的人，以及他的牛羊、牲畜和一切财物，就是他在 迦南 地所得的，往别处去，离开了他的兄弟 雅各 。
GEN|36|7|因为他们拥有的很多，不能住在一起。因为牲畜的缘故，寄居的地方容不下他们。
GEN|36|8|于是 以扫 住在 西珥山 ； 以扫 就是 以东 。
GEN|36|9|这是 以扫 的后代，他是 西珥山 里 以东 人的始祖。
GEN|36|10|以扫 子孙的名字如下： 以扫 的妻子 亚大 生 以利法 ； 以扫 的妻子 巴实抹 生 流珥 。
GEN|36|11|以利法 的儿子是 提幔 、 阿抹 、 洗玻 、 迦坦 、 基纳斯 。
GEN|36|12|亭纳 是 以扫 儿子 以利法 的妾，她为 以利法 生了 亚玛力 。这是 以扫 的妻子 亚大 的子孙。
GEN|36|13|流珥 的儿子是 拿哈 、 谢拉 、 沙玛 、 米撒 。这是 以扫 妻子 巴实抹 的子孙。
GEN|36|14|以扫 的妻子 阿何利巴玛 是 祭便 的孙女， 亚拿 的女儿。她为 以扫 生了 耶乌施 、 雅兰 、 可拉 。
GEN|36|15|这是 以扫 子孙中作族长的： 以扫 的长子 以利法 的子孙中，有 提幔 族长、 阿抹 族长、 洗玻 族长、 基纳斯 族长、
GEN|36|16|可拉 族长、 迦坦 族长、 亚玛力 族长。这是在 以东 地，从 以利法 所出的族长，是 亚大 的子孙。
GEN|36|17|以扫 的儿子 流珥 的子孙中，有 拿哈 族长、 谢拉 族长、 沙玛 族长、 米撒 族长。这是在 以东 地，从 流珥 所出的族长，是 以扫 妻子 巴实抹 的子孙。
GEN|36|18|以扫 的妻子 阿何利巴玛 的子孙中，有 耶乌施 族长、 雅兰 族长、 可拉 族长。这是从 以扫 的妻子， 亚拿 的女儿 阿何利巴玛 的子孙中所出的族长。
GEN|36|19|以上的族长都是 以扫 的子孙； 以扫 就是 以东 。
GEN|36|20|这是那地原来的居民， 何利 人 西珥 的子孙： 罗坍 、 朔巴 、 祭便 、 亚拿 、
GEN|36|21|底顺 、 以察 、 底珊 。这是在 以东 地，从 何利 人 西珥 子孙中所出的族长。
GEN|36|22|罗坍 的儿子是 何利 、 希幔 ， 罗坍 的妹妹是 亭纳 。
GEN|36|23|朔巴 的儿子是 亚勒文 、 玛拿辖 、 以巴录 、 示玻 、 阿南 。
GEN|36|24|祭便 的儿子是 爱亚 、 亚拿 ，当时在旷野牧放他父亲 祭便 的驴，发现温泉的就是这 亚拿 。
GEN|36|25|亚拿 的儿子是 底顺 ， 亚拿 的女儿是 阿何利巴玛 。
GEN|36|26|底顺 的儿子是 欣但 、 伊是班 、 益兰 、 基兰 。
GEN|36|27|以察 的儿子是 辟罕 、 撒番 、 亚干 。
GEN|36|28|底珊 的儿子是 乌斯 、 亚兰 。
GEN|36|29|这是从 何利 人所出的族长： 罗坍 族长、 朔巴 族长、 祭便 族长、 亚拿 族长、
GEN|36|30|底顺 族长、 以察 族长、 底珊 族长。这是从 何利 人所出的族长，都在 西珥 地，按着族长 来分。
GEN|36|31|以色列 未有君王治理之前，这些是在 以东 地作王的。
GEN|36|32|比珥 的儿子 比拉 在 以东 作王，他的城名叫 亭哈巴 。
GEN|36|33|比拉 死了， 波斯拉 人 谢拉 的儿子 约巴 接续他作王。
GEN|36|34|约巴 死了， 提幔 人之地的 户珊 接续他作王。
GEN|36|35|户珊 死了， 比达 的儿子 哈达 接续他作王， 哈达 曾在 摩押 地击败 米甸 人，他的城名叫 亚未得 。
GEN|36|36|哈达 死了， 玛士利加 人 桑拉 接续他作王。
GEN|36|37|桑拉 死了， 大河 边的 利河伯 人 扫罗 接续他作王。
GEN|36|38|扫罗 死了， 亚革波 的儿子 巴勒．哈南 接续他作王。
GEN|36|39|亚革波 的儿子 巴勒．哈南 死了， 哈达尔 接续他作王，他的城名叫 巴乌 。他的妻子名叫 米希她别 ，是 米．萨合 的孙女， 玛特列 的女儿。
GEN|36|40|这些是 以扫 的族长，按着他们的宗族、住处和名字： 亭纳 族长、 亚勒瓦 族长、 耶帖 族长、
GEN|36|41|阿何利巴玛 族长、 以拉 族长、 比嫩 族长、
GEN|36|42|基纳斯 族长、 提幔 族长、 米比萨 族长、
GEN|36|43|玛基叠 族长、 以兰 族长。这些是 以东 人在所得为业的地上，按着他们住处的族长。 以扫 是 以东 人的始祖。
GEN|37|1|雅各 住在 迦南 地，就是他父亲寄居的地。
GEN|37|2|这是 雅各 的事迹。 约瑟 十七岁与他哥哥们一同牧羊。他是个少年，与他父亲的妾 辟拉 和 悉帕 的儿子们常在一起。 约瑟 把他们的恶行报给父亲。
GEN|37|3|以色列 爱 约瑟 过于其他的儿子，因为 约瑟 是他年老生的；他给 约瑟 做了一件长袍 。
GEN|37|4|哥哥们见父亲爱 约瑟 过于他们，就恨 约瑟 ，不与他说友善的话。
GEN|37|5|约瑟 做了一个梦，告诉他哥哥们，他们就更加恨他。
GEN|37|6|约瑟 对他们说：“请听我做的这个梦：
GEN|37|7|看哪，我们在田里捆禾稼；看哪，我的捆起来站着；看哪，你们的捆围着我的捆下拜。”
GEN|37|8|他的哥哥们对他说：“难道你真的要作我们的王吗？难道你真的要统治我们吗？”他们就因他的梦和他的话更加恨他。
GEN|37|9|后来他又做了另一个梦，告诉他哥哥们说：“看哪，我又做了一个梦；看哪，太阳、月亮和十一颗星都向我下拜。”
GEN|37|10|约瑟 告诉他父亲和哥哥们，他父亲就责备他说：“你做的这是什么梦！难道我和你母亲、你的兄弟真的要俯伏在地，来向你下拜吗？”
GEN|37|11|他的哥哥们都嫉妒他，他父亲却把这事存在心里。
GEN|37|12|约瑟 的哥哥们到 示剑 去放他们父亲的羊。
GEN|37|13|以色列 对 约瑟 说：“你哥哥们不是在 示剑 放羊吗？来，我派你到他们那里去。” 约瑟 对他说：“我在这里。”
GEN|37|14|以色列 对他说：“你去看看你哥哥们是否平安，羊群是否平安，再回来告诉我。”于是他派 约瑟 出 希伯仑谷 ， 约瑟 就往 示剑 去了。
GEN|37|15|有人遇见他，看哪，他在田野走迷了路。那人问他说：“你找什么？”
GEN|37|16|他说：“我找我的哥哥们，请告诉我，他们在哪里放羊。”
GEN|37|17|那人说：“他们已经离开这里走了，我听见他们说：‘我们往 多坍 去。’” 约瑟 就去追哥哥们，在 多坍 找到了他们。
GEN|37|18|他们远远看见他，趁他还没有走近他们，就图谋要杀死他。
GEN|37|19|他们彼此说：“看哪！那做梦的来了。
GEN|37|20|现在，来吧！我们把他杀了，丢在一个坑里，就说有恶兽把他吃了。我们且看他的梦将来怎么样。”
GEN|37|21|吕便 听见了，要救 约瑟 脱离他们的手，说：“我们不可害他的性命”；
GEN|37|22|吕便 又对他们说：“不可流他的血，可以把他丢在这旷野的坑里，不可下手害他。” 吕便 要救他脱离他们的手，把他还给他父亲。
GEN|37|23|约瑟 到了他哥哥们那里，他们就剥去他的外衣，就是他身上那件长袍。
GEN|37|24|他们抓住他，把他丢在坑里。那坑是空的，里头没有水。
GEN|37|25|他们坐下吃饭，举目观看，看哪，有一群 以实玛利 人从 基列 来，用骆驼驮着香料、乳香、没药，要带下 埃及 去。
GEN|37|26|犹大 对他的兄弟们说：“我们杀我们的弟弟，遮掩他的血有什么好处呢？
GEN|37|27|来，我们把他卖给 以实玛利 人，不要下手害他，因为他是我们的弟弟，我们的骨肉。”他的兄弟们就听从了他。
GEN|37|28|那时，有些 米甸 的商人从那里经过，就把 约瑟 从坑里拉上来。他们以二十块银子把 约瑟 卖给 以实玛利 人，他们就把 约瑟 带到 埃及 去了。
GEN|37|29|吕便 回到坑旁，看哪， 约瑟 不在坑里，就撕裂自己的衣服，
GEN|37|30|回到他兄弟们那里，说：“孩子不在了。我往哪里去才好呢？”
GEN|37|31|于是，他们宰了一只公山羊，拿了 约瑟 的那件外衣染上了血，
GEN|37|32|派人把长袍送到他们的父亲那里，说：“我们发现这个， 请认一认，是不是你儿子的外衣？”
GEN|37|33|他认出来，就说：“这是我儿子的外衣，恶兽把他吃了， 约瑟 一定被撕碎了！”
GEN|37|34|雅各 就撕裂衣服，腰间围上麻布，为他儿子哀伤了多日。
GEN|37|35|他的儿女都起来安慰他，他却不肯受安慰，说：“我必哀伤着下阴间，到我儿子那里。” 约瑟 的父亲就为他哀哭。
GEN|37|36|米甸 人把 约瑟 卖到 埃及 ，给法老的官员，就是护卫长 波提乏 。
GEN|38|1|那时， 犹大 离开他兄弟们下去，到一个名叫 希拉 的 亚杜兰 人的家附近支搭帐棚。
GEN|38|2|犹大 在那里看见一个名叫 拔．书亚 的 迦南 女子，就娶她为妻，与她同房，
GEN|38|3|她就怀孕生了儿子， 犹大 给他起名叫 珥 。
GEN|38|4|她又怀孕生了儿子，给他起名叫 俄南 。
GEN|38|5|她又再生了儿子，给他起名叫 示拉 。她生 示拉 的时候， 犹大 正在 基悉 。
GEN|38|6|犹大 为长子 珥 娶妻，名叫 她玛 。
GEN|38|7|犹大 的长子 珥 在耶和华眼中看为恶，耶和华就杀死了他。
GEN|38|8|犹大 对 俄南 说：“你当与你哥哥的妻子同房，向她尽你的本分，为你哥哥生子立后。”
GEN|38|9|俄南 知道如果与嫂嫂同房，所生的孩子不属于自己，就泄在地上，不为哥哥生子立后。
GEN|38|10|俄南 所做的在耶和华眼中看为恶，耶和华也杀死了他。
GEN|38|11|犹大 对他媳妇 她玛 说：“你去住在你父亲家里守寡，等我儿子 示拉 长大。”因为他说：“恐怕 示拉 也像两个哥哥一样死去。” 她玛 就去，住在她父亲家里。
GEN|38|12|过了一段很长的日子， 犹大 的妻子， 书亚 的女儿死了。 犹大 受到了安慰，就和他朋友 亚杜兰 人 希拉 上 亭拿 去，到他的剪羊毛的人那里。
GEN|38|13|有人告诉 她玛 说：“看哪，你的公公上 亭拿 剪羊毛去了。”
GEN|38|14|她玛 见 示拉 已经长大，却还没有娶她为妻，就脱去她寡妇的衣裳，用面纱蒙着，盖住自己，坐在往 亭拿 的路上， 伊拿印 城门口。
GEN|38|15|犹大 看见她，以为是妓女，因为她蒙着脸。
GEN|38|16|犹大 就转到路边她那里，说：“来吧！让我与你同寝。”他并不知道她就是他的媳妇。 她玛 说：“你要与我同寝，把什么给我呢？”
GEN|38|17|犹大 说：“我从羊群里取一只小山羊，派人送来给你。” 她玛 说：“在未送之前，你能给我一个信物吗？”
GEN|38|18|他说：“我给你什么信物呢？” 她玛 说：“你的印、你的带子 和你手里的杖。”于是 犹大 给了她，与她同寝，她就从 犹大 怀了孕。
GEN|38|19|她玛 起来走了，除去面纱，照常穿上寡妇的衣裳。
GEN|38|20|犹大 托他朋友 亚杜兰 人送一只小山羊去，要从那女人手里取回信物，却找不到她。
GEN|38|21|他问那地方的人说：“ 伊拿印 路旁的神庙娼妓在哪里？”他们说：“这里没有神庙娼妓。”
GEN|38|22|他回到 犹大 那里说：“我找不到她，并且那地方的人说：‘这里没有神庙娼妓。’”
GEN|38|23|犹大 说：“让她拿去吧，免得我们被人讥笑。看哪，我把这小山羊送去了，可是你找不到她。”
GEN|38|24|大约过了三个月，有人告诉 犹大 说：“你的媳妇 她玛 行淫，并且，看哪，她因行淫而怀了孕。” 犹大 说：“拉她出来，把她烧了！”
GEN|38|25|她玛 被拉出来的时候，就派人到她公公那里，对他说：“这些东西是谁的，我就是从谁怀了孕。”她又说：“请你认一认，这印、这带子和这杖是谁的？”
GEN|38|26|犹大 承认说：“她比我更有理，因为我没有把她给我的儿子 示拉 。” 犹大 再也不跟她同寝。
GEN|38|27|她玛 生产的时候到了，看哪，腹里怀的是双胞胎。
GEN|38|28|生产的时候，一个孩子伸出手来；接生婆拿红线绑在他手上，说：“这是头生的。”
GEN|38|29|这孩子把手收回去，看哪，他哥哥生出来了；接生婆说：“你竟然为自己冲出一个裂缝！”于是，他的名字叫 法勒斯 。
GEN|38|30|后来，那手上有红线的兄弟也生出来，他的名字叫 谢拉 。
GEN|39|1|约瑟 被带下 埃及 去。有一个 埃及 人 波提乏 ，是法老的官员，是护卫长，他从那些带 约瑟 下来的 以实玛利 人手中把 约瑟 买了去。
GEN|39|2|约瑟 在他 埃及 主人的家中，耶和华与他同在，他是一个通达的人。
GEN|39|3|他主人见耶和华与他同在，又见耶和华使他手里所办的事都顺利，
GEN|39|4|约瑟 就在主人眼前蒙恩，伺候他主人，主人派他管理家务，把一切所有的都交在他手里。
GEN|39|5|自从主人派 约瑟 管理家务和他一切所有的，耶和华就因 约瑟 的缘故赐福给那 埃及 人的家；凡家里和田间一切所有的，都蒙耶和华赐福。
GEN|39|6|波提乏 把他一切所有的都交在 约瑟 手中，除了自己所吃的食物，其他的事一概不知。 约瑟 英俊健美。
GEN|39|7|这些事以后， 约瑟 主人的妻子以目送情给 约瑟 ，说：“你与我同寝吧！”
GEN|39|8|约瑟 拒绝，对他主人的妻子说：“看哪，一切家务我主人一概不知，他把所有的都交在我手里。
GEN|39|9|在这家里没有人比我更大，除你以外，他也没有留下一样不交给我，因为你是他的妻子。我怎能行这么大的恶，得罪上帝呢？”
GEN|39|10|她天天这样对 约瑟 说， 约瑟 却不听从她，不与她同寝，也不和她在一起。
GEN|39|11|有一天， 约瑟 进屋里去办事，家里没有一个人在那屋子里，
GEN|39|12|妇人就拉住他的衣服，说：“你与我同寝吧！” 约瑟 把衣服留在她手里，逃出外面去了。
GEN|39|13|妇人看见 约瑟 把衣服留在她手里逃到外面，
GEN|39|14|就叫了家里的人来，对他们说：“看，他带了一个 希伯来 人到我们这里戏弄我们。他到我这里来，要与我同寝，我就大声喊叫。
GEN|39|15|他听见我放声大喊，就把他的衣服留在我这里，逃出外面去了。”
GEN|39|16|妇人把 约瑟 的衣服放在身边，直到他主人回家，
GEN|39|17|就用这样的话对他说：“你带到我们这里来的那 希伯来 仆人进来要调戏我，
GEN|39|18|我放声大喊，他就把衣服留在我身边，逃到外面。”
GEN|39|19|主人听见他妻子对他说的话，说：“你的仆人就是这样对待我”，就非常生气。
GEN|39|20|约瑟 的主人把他抓起来，关在监狱里，就是王的囚犯被关的地方。于是 约瑟 在那里坐牢。
GEN|39|21|但耶和华与 约瑟 同在，向他施恩，使他在监狱长的眼前蒙恩。
GEN|39|22|监狱长就把监狱里所有的囚犯都交在 约瑟 手下；在那里的一切事都由他处理。
GEN|39|23|任何交在 约瑟 手中的事，监狱长一概不察，因为耶和华与 约瑟 同在，耶和华使他所做的都顺利。
GEN|40|1|这些事以后， 埃及 王的司酒长和司膳长得罪了他们的主 埃及 王。
GEN|40|2|法老就对司酒长和司膳长两个官员发怒，
GEN|40|3|把他们关在护卫长府内的监狱里，就是 约瑟 被囚的地方。
GEN|40|4|护卫长把他们交给 约瑟 ， 约瑟 就伺候他们。他们被关了一段日子。
GEN|40|5|关在监狱里的这两个人，就是 埃及 王的司酒长和司膳长，在同一个晚上各自做了一个梦，每个梦都有自己的解释。
GEN|40|6|到了早晨， 约瑟 来到他们那里看他们，看哪，他们很忧愁。
GEN|40|7|他就问一同关在他主人府内法老的官员，说：“你们今日为什么面带愁容呢？”
GEN|40|8|他们对他说：“我们各自做了一个梦，却没有人能讲解。” 约瑟 对他们说：“解梦不是出于上帝吗？请你们把梦告诉我。”
GEN|40|9|司酒长就把梦告诉 约瑟 ，对他说：“在我的梦中，看哪，有一棵葡萄树在我面前，
GEN|40|10|树上有三根枝子。枝子发了芽，开了花，结出串串成熟的葡萄。
GEN|40|11|法老的杯在我手中，我就拿葡萄挤在法老的杯里，把杯递到他手中。”
GEN|40|12|约瑟 对他说：“梦的解释是这样：三根枝子就是三天；
GEN|40|13|三天之内，法老要让你抬起头来，叫你官复原职。你仍要递杯在法老的手中，像先前作他的司酒长一样。
GEN|40|14|但你得福的时候，请你记得我，向我施慈爱，在法老面前提起我，救我出这监牢。
GEN|40|15|我实在是从 希伯来 人之地被拐来的，我在这里也没有做过什么，好叫他们把我关在牢里。”
GEN|40|16|司膳长见梦解得好，就对 约瑟 说：“在我梦中，看哪，我头上顶着三个装饼的篮子；
GEN|40|17|最上面的篮子里有为法老烤的各样食物，有飞鸟来吃我头上篮子里的食物。”
GEN|40|18|约瑟 说：“梦的解释是这样：三个篮子就是三天；
GEN|40|19|三天之内，法老要让你抬起头来，身首异处，把你挂在木架上，必有飞鸟来吃你身上的肉。”
GEN|40|20|到了第三天，正是法老的生日，他为众臣仆摆设宴席，使司酒长和司膳长从众臣仆中抬起头来，
GEN|40|21|让司酒长官复原职，仍旧递杯在法老手中，
GEN|40|22|却把司膳长挂起来，正如 约瑟 向他们所讲解的。
GEN|40|23|然而，司酒长不记得 约瑟 ，竟忘了他。
GEN|41|1|过了两年，法老做梦，看哪，自己站在 尼罗河 边，
GEN|41|2|看哪，有七头母牛从 尼罗河 里上来，长相俊美，肌肉肥壮，在芦苇中吃草。
GEN|41|3|看哪，随后又有七头母牛从 尼罗河 里上来，长相丑陋，肌肉干瘦，与那七头母牛一同站在河边。
GEN|41|4|这长相丑陋，肌肉干瘦的七头母牛吃了那长相俊美又肥壮的七头母牛。法老就醒了。
GEN|41|5|他又睡着，第二次做梦，看哪，一株麦杆长了七个穗子，又肥大又佳美，
GEN|41|6|看哪，随后又长出七个穗子，又细弱又被东风吹焦了。
GEN|41|7|这细弱的穗子吞了那七个又肥大又饱满的穗子。法老醒了，看哪，是个梦。
GEN|41|8|到了早晨，法老心里不安，就派人把 埃及 所有的术士和智慧人都召来。法老把所做的梦告诉他们，但是没有人能为法老解梦。
GEN|41|9|那时司酒长对法老说：“我今日想起我的罪来。
GEN|41|10|从前法老对臣仆发怒，把我和司膳长关在护卫长府内的监牢里。
GEN|41|11|我们两人在同一晚上各做一梦，每个梦都有各自的解释。
GEN|41|12|同我们在一起有一个 希伯来 的年轻人，是护卫长的仆人。我们告诉他，他就为我们解梦，照着各人的梦讲解。
GEN|41|13|后来事情正如他给我们讲解的实现了，我官复原职，司膳长被挂起来了。”
GEN|41|14|于是法老派人去召 约瑟 ，他们就急忙把他从牢里提出来。他就剃头刮脸，换衣服，进到法老面前。
GEN|41|15|法老对 约瑟 说：“我做了一个梦，没有人能讲解。我听人说，你听了梦就能讲解。”
GEN|41|16|约瑟 回答法老说：“这不在乎我。上帝必应允法老平安。”
GEN|41|17|法老对 约瑟 说：“在我的梦中，看哪，我站在 尼罗河 边，
GEN|41|18|看哪，有七头母牛从 尼罗河 里上来，肌肉肥壮，外形俊美，在芦苇中吃草。
GEN|41|19|看哪，随后又有七头母牛上来，虚弱，外形很丑陋，肌肉又干瘦，在 埃及 全地，我没有见过这样丑陋的牛。
GEN|41|20|这干瘦又丑陋的母牛吃了那先前的七头肥母牛，
GEN|41|21|进了肚子以后却看不出已经进了肚子，那丑陋的长相仍旧和先前一样。我就醒了。
GEN|41|22|我又在梦中观看，看哪，一株麦杆长了七个穗子，又饱满又佳美，
GEN|41|23|看哪，随后又长出七个穗子，枯槁，细弱，又被东风吹焦了。
GEN|41|24|这些细弱的穗子吞了那七个佳美的穗子。我告诉术士，却没有人能为我讲解。”
GEN|41|25|约瑟 对法老说：“法老的梦是同一个。上帝已把要做的事指示法老了。
GEN|41|26|七头好母牛是七年，七个佳美的穗子也是七年，这是同一个梦。
GEN|41|27|那随后上来的七头干瘦又丑陋的母牛是七年；那七个空心，被东风吹焦的穗子也一样，都是七个荒年。
GEN|41|28|这就是我对法老所说，上帝已把要做的事显明给法老了。
GEN|41|29|看哪，必有七个大丰年来到 埃及 全地，
GEN|41|30|随后又有七个荒年，甚至 埃及 地的人都忘了先前的丰收，这地必被饥荒所灭。
GEN|41|31|因为那后来的饥荒非常严重，就不觉得这地先前有丰收。
GEN|41|32|至于法老两次做梦，是因为上帝已经确定这事，上帝必速速成就。
GEN|41|33|现在，请法老选一个聪明又有智慧的人，委派他治理 埃及 地。
GEN|41|34|请法老这样做，委派官员治理这地，在七个丰年的期间，征收 埃及 地出产的五分之一，
GEN|41|35|叫他们聚集未来丰年一切的粮食，积存五谷归在法老的手下作粮食，储藏在各城里。
GEN|41|36|这粮食可以为这地作储备，为了 埃及 地要来的七个荒年，免得这地被饥荒所灭。”
GEN|41|37|这事在法老和他众臣仆眼中都觉得好。
GEN|41|38|法老对臣仆说：“像这样的人，有上帝的灵在他里面，我们岂能找得着呢？”
GEN|41|39|法老对 约瑟 说：“上帝既指示你这一切事，就没有人像你这样聪明又有智慧。
GEN|41|40|你可以治理我的家；我的百姓都必服从你口中的命令。惟独在宝座上，我比你大。”
GEN|41|41|法老又对 约瑟 说：“看，我委派你治理 埃及 全地。”
GEN|41|42|法老就脱下手上带印的戒指，戴在 约瑟 的手上，给他穿上细麻衣，把金链戴在他的颈项上，
GEN|41|43|又给 约瑟 坐他的副座车，在他前面有人呼叫说：“跪下 。”于是，法老委派他治理 埃及 全地。
GEN|41|44|法老对 约瑟 说：“我是法老，若没有你的命令， 埃及 全地的人都不可擅自办事 。”
GEN|41|45|法老给 约瑟 起名叫 撒发那特．巴内亚 ，又将 安城 的祭司 波提．非拉 的女儿 亚西纳 给他为妻。 约瑟 就出去治理 埃及 地。
GEN|41|46|约瑟 在 埃及 王法老面前侍立的时候年三十岁。 约瑟 从法老面前出去，巡行 埃及 全地。
GEN|41|47|七个丰年之内，地的出产极其丰盛 ，
GEN|41|48|约瑟 聚集 埃及 地七年一切的粮食，把粮食积存在各城里，就是把各城周围田地的粮食都积存在该城里。
GEN|41|49|约瑟 积存的五谷很多，如同海边的沙，无法计算，数也数不清。
GEN|41|50|荒年未到以前， 安城 的祭司 波提．非拉 的女儿 亚西纳 为 约瑟 生了两个儿子。
GEN|41|51|约瑟 给长子起名叫 玛拿西 ，因为他说：“上帝使我忘了一切的困苦和我父的全家。”
GEN|41|52|他给次子起名叫 以法莲 ，因为他说：“上帝使我在受苦的地方兴盛。”
GEN|41|53|埃及 地的七个丰年一过，
GEN|41|54|七个荒年就来了，正如 约瑟 所说的。各地都有饥荒，惟独 埃及 全地有粮食。
GEN|41|55|等到 埃及 全地也有了饥荒，众百姓就向法老哀求粮食。法老对所有的 埃及 人说：“你们到 约瑟 那里去，凡他所说的，你们都要做。”
GEN|41|56|当时饥荒遍满了全地， 约瑟 就开了各处的粮仓 ，卖粮食给 埃及 人。 埃及 地的饥荒非常严重。
GEN|41|57|各地的人都去 埃及 ，到 约瑟 那里买粮食，因为全地的饥荒非常严重。
GEN|42|1|雅各 见 埃及 有粮，就对儿子们说：“你们为什么彼此对看呢？”
GEN|42|2|他又说：“看哪，我听见 埃及 有粮，你们可以下到那里，从那里为我们买些粮来，我们就可以存活，不至于死。”
GEN|42|3|于是， 约瑟 的十个哥哥都下去，到 埃及 买粮食。
GEN|42|4|至于 约瑟 的弟弟 便雅悯 ， 雅各 没有派他和哥哥们同去，因为 雅各 说：“恐怕他遭难。”
GEN|42|5|以色列 的儿子们来了，在前来的人当中，为要买粮食，因为 迦南 地也有饥荒。
GEN|42|6|当时在 埃及 地掌权的人是 约瑟 ，卖粮给各地众百姓的就是他。 约瑟 的哥哥们来了，脸伏于地，向他下拜。
GEN|42|7|约瑟 看见他哥哥们，就认出他们，却对他们装作陌生人，向他们说严厉的话，对他们说：“你们从哪里来？”他们说：“我们从 迦南 地来买粮。”
GEN|42|8|约瑟 认得他哥哥们，他们却不认得他。
GEN|42|9|约瑟 想起从前所做的那两个梦，就对他们说：“你们是奸细，你们来是要窥探这地的虚实。”
GEN|42|10|他们对他说：“我主啊，不是的，仆人们是来买粮的。
GEN|42|11|我们都是同一个人的儿子，我们是诚实的人。仆人们并不是奸细。”
GEN|42|12|约瑟 对他们说：“不，你们一定是窥探这地的虚实来的。”
GEN|42|13|他们说：“仆人们本是兄弟十二人，我们都是 迦南 地同一个人的儿子。看哪，最小的今日在我们父亲那里，有一个不在了。”
GEN|42|14|约瑟 对他们说：“我刚才对你们说过了，你们是奸细！
GEN|42|15|我指着法老的性命起誓，若是你们最小的弟弟不到这里来，你们就不可以离开这里；这样你们就可以证实自己了。
GEN|42|16|要派你们当中的一个人去，把你们的弟弟带来。至于你们，都要关在这里，好证实你们的话是不是真的。若不是，我指着法老的性命起誓，你们一定是奸细。”
GEN|42|17|于是 约瑟 把他们一起都关在监里三天。
GEN|42|18|第三天， 约瑟 对他们说：“我是敬畏上帝的，你们这么做就可以活。
GEN|42|19|如果你们是诚实的人，留你们兄弟中的一个关在监牢里，你们带粮食回去，救你们家的饥荒，
GEN|42|20|再把你们最小的弟弟带到我这里来。如此，你们的话就是真的了，你们也不至于死。”他们就照样做了。
GEN|42|21|他们彼此说：“我们在弟弟身上实在犯了罪。他哀求我们的时候，我们看见他的痛苦，却不肯听，所以这场苦难临到我们。”
GEN|42|22|吕便 回答他们说：“我不是对你们说过，不可伤害那孩子吗？只是你们不肯听，看哪，他的血在追讨了。”
GEN|42|23|他们不知道 约瑟 在听，因为在他们之间有传译官。
GEN|42|24|约瑟 转身离开他们，哭了一场，又回来对他们说话，就从他们中间抓了 西缅 ，在他们眼前捆绑他。
GEN|42|25|约瑟 吩咐人把他们的器皿装满粮食，把各人的银子退还在各人的袋里，又给他们路上需用的食物。人就为他们这样做了。
GEN|42|26|他们把粮食驮在驴上，离开那里去了。
GEN|42|27|到了住宿的地方，有一个人打开袋子，要拿饲料喂驴，就看见自己的银子，看哪，仍在袋口上。
GEN|42|28|他对兄弟们说：“我的银子退回来了，看哪，还在我袋子里！”他们战战兢兢，心都快跳出来了，彼此说：“上帝向我们做的是什么呢？”
GEN|42|29|他们来到 迦南 地他们的父亲 雅各 那里，把所遭遇的事都告诉他，说：
GEN|42|30|“那地的主对我们说严厉的话，把我们当作窥探那地的奸细。
GEN|42|31|我们对他说：‘我们是诚实的人，并不是奸细。
GEN|42|32|我们本是兄弟十二人，都是同一个父亲的儿子，有一个不在了，最小的今日和我们父亲在 迦南 地。’
GEN|42|33|那地的主对我们说：‘只有这样我才知道你们是诚实的人：留你们兄弟中的一个在我这里，你们带粮食回去，救你们家的饥荒，
GEN|42|34|再把你们最小的弟弟带到我这里来，我就知道你们不是奸细，是诚实的人。然后，我就把你们的兄弟交还你们，你们也可以在此地做买卖。’”
GEN|42|35|后来他们倒空袋子，看哪，各人的银囊都在袋子里。他们和父亲看见银囊就都害怕。
GEN|42|36|他们的父亲 雅各 对他们说：“你们害我丧失了我的儿子： 约瑟 不在了， 西缅 也不在了，你们还要带走 便雅悯 ！这些事都临到我身上了。”
GEN|42|37|吕便 对他父亲说：“我若不带他回来给你，你可以杀我的两个儿子。只管把他交在我手里，我必带他回来给你。”
GEN|42|38|雅各 说：“我的儿子不可与你们一同下去。他哥哥死了，只剩下他。他若在你们行走的路上遭难，你们就害我白发苍苍、悲悲惨惨下阴间去了。”
GEN|43|1|那地的饥荒非常严重。
GEN|43|2|他们从 埃及 带来的粮食吃完了，父亲对他们说：“你们再去给我们买些粮来。”
GEN|43|3|犹大 对他说：“那人严厉地警告我们说：‘你们的弟弟若不和你们同来，你们就不要来见我的面。’
GEN|43|4|你若派我们的弟弟跟我们同去，我们就下去给你买粮；
GEN|43|5|你若不派他去，我们就不下去，因为那人对我们说：‘你们的弟弟若不和你们同来，你们就不要来见我的面。’”
GEN|43|6|以色列 说：“你们为什么这样害我，告诉那人你们还有弟弟呢？”
GEN|43|7|他们说：“那人详细问到我们和我们的家人，说：‘你们的父亲还在吗？你们还有兄弟吗？’我们就按着他的这些话告诉他，我们怎么知道他会说：‘把你们的弟弟带下来’呢？”
GEN|43|8|犹大 又对他父亲 以色列 说：“请派这年轻人和我同去，我们就动身前去，好叫我们和你，以及我们的孩子都得存活，不至于死。
GEN|43|9|我为他担保，你可以从我手中要人，我若不带他回来交在你面前，我就对你永远担当这罪。
GEN|43|10|我们若没有耽搁，现在第二趟都回来了。”
GEN|43|11|父亲 以色列 对他们说：“如果必须如此，你们要这样做：把本地土产中最好的乳香、蜂蜜、香料、没药、坚果、杏仁各取一点，放在器皿里，带下去送给那人作礼物。
GEN|43|12|手里要带双倍的银子，把退还在你们袋口的银子亲手带回去；或许那是个失误。
GEN|43|13|带着你们的弟弟，动身再去见那人。
GEN|43|14|愿全能的上帝使你们在那人面前蒙怜悯，放你们另一个兄弟和 便雅悯 回来。我若要失丧儿子，就丧了吧！”
GEN|43|15|于是，他们拿着那些礼物，手里也带双倍的银子，并且带着 便雅悯 ，动身下到 埃及 ，站在 约瑟 面前。
GEN|43|16|约瑟 见 便雅悯 和他们同来，就对管家说：“把这些人领到屋里。要宰杀牲畜，预备宴席，因为中午这些人要跟我吃饭。”
GEN|43|17|那人就照 约瑟 所说的去做，领他们进 约瑟 的屋里。
GEN|43|18|这些人因为被领到 约瑟 的屋里，就害怕，说：“领我们到这里来，必是因为当初退还在我们袋里的银子，要设计害我们，抓我们去当奴隶，抢夺我们的驴。”
GEN|43|19|他们就挨近 约瑟 的管家，在屋子门口和他说话，
GEN|43|20|说：“我主啊，求求你，我们当初下来，真的是要买粮食。
GEN|43|21|后来到了住宿的地方，我们打开袋子，看哪，各人的银子还在自己的袋口上，银子的分量一点不少。现在我们亲手把它带回来，
GEN|43|22|我们手里又带了另外的银子来买粮食。我们不知道是谁把银子放在我们袋里的。”
GEN|43|23|他说：“你们平安！不要害怕，是你们的上帝和你们父亲的上帝把财宝放在你们的袋里。你们的银子，我已经收了。”他就把 西缅 带出来，交给他们。
GEN|43|24|那人领这些人进 约瑟 的屋里，给他们水洗脚，又给他们饲料喂驴。
GEN|43|25|他们预备好礼物，等候 约瑟 中午来，因为他们听说他们要在那里吃饭。
GEN|43|26|约瑟 来到家里，他们就把手中的礼物拿进屋里给他，俯伏在地，向他下拜。
GEN|43|27|约瑟 问他们安，又说：“你们的父亲，就是你们所说的那位老人家平安吗？他还在吗？”
GEN|43|28|他们说：“你仆人，我们的父亲平安，他还在。”于是他们低头下拜。
GEN|43|29|约瑟 举目看见他同母的弟弟 便雅悯 ，就说：“你们向我所说那最小的弟弟就是这位吗？”又说：“我儿啊，愿上帝赐恩给你！”
GEN|43|30|约瑟 爱弟之情激动，就急忙找个地方去哭。他进入自己的房间，哭了一场。
GEN|43|31|他洗了脸出来，勉强忍住，就说：“开饭吧！”
GEN|43|32|他们为 约瑟 单独摆了一席，为那些人又摆了一席，也为和 约瑟 同吃饭的 埃及 人另摆了一席，因为 埃及 人不和 希伯来 人一同吃饭；那是 埃及 人所厌恶的。
GEN|43|33|兄弟们被安排在 约瑟 面前坐席，都按着长幼的次序，这些人彼此感到诧异。
GEN|43|34|约瑟 把他面前的食物分给他们，但 便雅悯 所得的比别人多五倍。他们就喝酒，和 约瑟 一同畅饮。
GEN|44|1|约瑟 吩咐管家说：“按照他们的驴子所能驮的，把这些人的袋子装满粮食，再把各人的银子放在各人的袋口上，
GEN|44|2|我的杯，就是那个银杯，要和买粮的银子一同放在最年轻的那个人的袋口上。”管家就照 约瑟 所说的话去做了。
GEN|44|3|天一亮，这些人和他们的驴子就被送走了。
GEN|44|4|他们出城走了不远， 约瑟 对管家说：“起来，去追那些人，追上了就对他们说：‘你们为什么以恶报善呢？
GEN|44|5|这不是我主人用来饮酒，确实用它来占卜的吗？你们这么做是不对的！’”
GEN|44|6|管家追上他们，把这些话对他们说了。
GEN|44|7|他们对他说：“我主为什么说这样的话呢？你仆人们绝不会做这样的事。
GEN|44|8|看哪，我们从前在袋口上发现的银子，尚且从 迦南 地带来还你，我们又怎么会从你主人家里偷窃金银呢？
GEN|44|9|你仆人中无论在谁那里找到杯子，就叫他死，我们也要作我主的奴隶。”
GEN|44|10|管家说：“现在就照你们的话做吧！在谁那里找到杯子，谁就作我的奴隶，其余的人都没有罪。”
GEN|44|11|于是他们各人急忙把袋子卸在地上，各人打开自己的袋子。
GEN|44|12|管家就搜查，从年长的开始到年幼的为止，那杯竟在 便雅悯 的袋子里找到了。
GEN|44|13|他们就撕裂衣服，各人把驮子抬在驴上，回城去了。
GEN|44|14|犹大 和他兄弟们来到 约瑟 的屋里， 约瑟 还在那里，他们就在他面前俯伏于地。
GEN|44|15|约瑟 对他们说：“你们做的是什么事呢？你们岂不知像我这样的人必懂得占卜吗？”
GEN|44|16|犹大 说：“我们对我主能说什么呢？还有什么话可说呢？我们还能为自己表白吗？上帝已经查出你仆人的罪孽了。看哪，我们与那在他手中找到杯子的人都是我主的奴隶。”
GEN|44|17|约瑟 说：“我绝不能做这样的事！谁的手中找到杯子，谁就作我的奴隶。至于你们，可以平平安安上到你们父亲那里去。”
GEN|44|18|犹大 挨近他，说：“我主啊，求求你，让仆人说一句话给我主听，不要向仆人发烈怒，因为你如同法老一样。
GEN|44|19|我主曾问仆人们说：‘你们有父亲、兄弟没有？’
GEN|44|20|我们对我主说：‘我们有父亲，他已经年老，还有他老年所生的一个小儿子。他哥哥死了，他的母亲只剩下他一个孩子，父亲也疼爱他。’
GEN|44|21|你对仆人说：‘把他带下到我这里来，让我亲眼看看他。’
GEN|44|22|我们对我主说：‘这年轻人不能离开他父亲，若是离开，父亲就会死。’
GEN|44|23|你对仆人说：‘你们最小的弟弟若不和你们一同下来，你们就不要来见我的面。’
GEN|44|24|我们上到你仆人，我们父亲那里，就把我主的话告诉了他。
GEN|44|25|后来，我们的父亲说：‘你们再去给我买些粮来。’
GEN|44|26|我们说：‘我们不能下去。最小的弟弟若和我们同去，我们就可以下去。因为，最小的弟弟若不和我们同去，我们必不能见那人的面。’
GEN|44|27|你仆人，我父亲对我们说：‘你们知道我的妻子给我生了两个儿子。
GEN|44|28|一个离开我走了，我说他必是被野兽撕碎了，直到如今我再没有见过他；
GEN|44|29|现在你们又要把这个从我面前带走。倘若他遭难，那么你们就害我白发苍苍、悲悲惨惨下阴间去了。’
GEN|44|30|如今我回到你仆人，我父亲那里，若没有这年轻人和我们同去，我父亲的命是与这年轻人的命相连的，
GEN|44|31|当我们的父亲看见没有了这年轻人，他就会死。这样，我们就害你仆人，我们的父亲白发苍苍、悲悲惨惨下阴间去了。
GEN|44|32|仆人曾向我父亲为这年轻人担保，说：‘我若不带他回来交给父亲，我就在父亲面前永远担当这罪。’
GEN|44|33|现在，求你把仆人留下，代替这年轻人作我主的奴隶，让这年轻人和他哥哥们一同上去。
GEN|44|34|若这年轻人不和我一起，我怎能上到我父亲那里呢？恐怕我要看到灾祸临到我父亲了。”
GEN|45|1|约瑟 在所有侍立在他旁边的人面前情不自禁，就喊叫说：“每一个人都离开我，出去吧！” 约瑟 和兄弟相认的时候没有一人站在他那里。
GEN|45|2|他放声大哭， 埃及 人听见了，法老家中的人也听见了。
GEN|45|3|约瑟 对他兄弟们说：“我就是 约瑟 。我的父亲还在吗？”他兄弟们不敢回答他，因为他们在他面前都很惊惶。
GEN|45|4|约瑟 又对他兄弟们说：“靠近我一点。”他们就近前来。他说：“我是被你们卖到 埃及 的兄弟 约瑟 。
GEN|45|5|现在，不要因为把我卖到这里而忧伤，对自己生气，因为上帝差我在你们以先来，为要保全性命。
GEN|45|6|现在这地的饥荒已经二年了，还有五年不能耕种，没有收成。
GEN|45|7|上帝差我在你们以先来，为要给你们在世上存留余种，大施拯救，保全你们的性命。
GEN|45|8|这样看来，差我到这里来的不是你们，而是上帝。他又使我如同法老之父，作他全家之主，和 埃及 全地掌权的人。
GEN|45|9|你们要赶紧上到我父亲那里，对他说：‘你儿子 约瑟 这样说：上帝已立我作全 埃及 之主，请你下到我这里来，不要耽搁。
GEN|45|10|你和你的儿子孙子，羊群牛群，以及一切所有的，都可以住在 歌珊 地，与我相近。
GEN|45|11|我要在那里奉养你，因为还有五年的饥荒，免得你和你的家属，以及一切所有的，都陷入穷困中。’
GEN|45|12|看哪，你们的眼睛和我弟弟 便雅悯 的眼睛都看见，是我亲口对你们说话。
GEN|45|13|你们要把我在 埃及 一切的尊荣和你们所有看见的事情都告诉我父亲，也要赶紧请我父亲下到这里来。”
GEN|45|14|于是 约瑟 伏在他弟弟 便雅悯 的颈项上哭， 便雅悯 也在他的颈项上哭。
GEN|45|15|他又亲众兄弟，伏着他们哭。过后，他的兄弟就和他说话。
GEN|45|16|这消息传到法老的宫里，说：“ 约瑟 的兄弟们来了。”法老和他的臣仆眼中都看为好。
GEN|45|17|法老对 约瑟 说：“你要吩咐你的兄弟们说：‘你们要这样做：把驮子抬在牲口上，动身到 迦南 地去，
GEN|45|18|请你们的父亲和你们的家属都到我这里来，我要把 埃及 地的美物赐给你们，你们也要吃这地肥美的出产。’
GEN|45|19|你要吩咐他们：‘要这样做：从 埃及 地带着车辆去，把你们的孩子和妻子，以及你们的父亲都接来。
GEN|45|20|你们的眼不要顾惜你们的家具，因为 埃及 全地的美物都是你们的。’”
GEN|45|21|以色列 的儿子们就照样做了。 约瑟 遵照法老的吩咐，给他们车辆和路上需用的食物。
GEN|45|22|他又给所有哥哥每人一套衣服， 却给 便雅悯 三百银子，五套衣服。
GEN|45|23|他也送给父亲十匹公驴，驮着 埃及 的美物，以及十匹母驴，驮着给他父亲在路上需用的谷物、饼和粮食。
GEN|45|24|于是 约瑟 送他的兄弟们回去，对他们说：“你们不要在路上争吵。”
GEN|45|25|他们从 埃及 上去，来到 迦南 地他们的父亲 雅各 那里，
GEN|45|26|告诉他说：“ 约瑟 还活着，并且作了 埃及 全地掌权的人。” 雅各 心里冰凉，因为不信他们。
GEN|45|27|他们就把 约瑟 对他们所说一切的话都告诉了他。他看见 约瑟 派来接他的车辆，他们父亲 雅各 的灵就苏醒了。
GEN|45|28|以色列 说：“够了！我的儿子 约瑟 还活着，我要趁我未死之前去见他。”
GEN|46|1|以色列 带着一切所有的，起程到 别是巴 去，献祭给他父亲 以撒 的上帝。
GEN|46|2|夜间，上帝在异象中对 以色列 说：“ 雅各 ！ 雅各 ！”他说：“我在这里。”
GEN|46|3|上帝说：“我是上帝，你父亲的上帝。不要害怕下 埃及 去，因为我必使你在那里成为大国。
GEN|46|4|我要和你同下 埃及 去，也必定带你上来； 约瑟 要亲手合上你的眼睛。”
GEN|46|5|雅各 就从 别是巴 起行。 以色列 的儿子让他们的父亲 雅各 和他们的孩子、妻子都坐在法老为 雅各 派来的车上。
GEN|46|6|他们也带着 迦南 地所得的牲畜和财物来到 埃及 。 雅各 和他所有的子孙都一同来了。
GEN|46|7|他把他的儿子、孙子、女儿、孙女，他所有的子孙一同带到 埃及 。
GEN|46|8|这些是来到 埃及 的 以色列 人， 雅各 和他子孙的名字： 雅各 的长子是 吕便 。
GEN|46|9|吕便 的儿子是 哈诺 、 法路 、 希斯伦 、 迦米 。
GEN|46|10|西缅 的儿子是 耶母利 、 雅悯 、 阿辖 、 雅斤 、 琐辖 ，还有 迦南 女子生的儿子 扫罗 。
GEN|46|11|利未 的儿子是 革顺 、 哥辖 、 米拉利 。
GEN|46|12|犹大 的儿子是 珥 、 俄南 、 示拉 、 法勒斯 、 谢拉 ； 珥 与 俄南 死在 迦南 地。 法勒斯 的儿子是 希斯仑 、 哈母勒 。
GEN|46|13|以萨迦 的儿子是 陀拉 、 普瓦 、 约伯 、 伸仑 。
GEN|46|14|西布伦 的儿子是 西烈 、 以伦 、 雅利 。
GEN|46|15|这是 利亚 在 巴旦．亚兰 为 雅各 所生的儿孙，还有女儿 底拿 ，儿孙共三十三人。
GEN|46|16|迦得 的儿子是 洗非芸 、 哈基 、 书尼 、 以斯本 、 以利 、 亚罗底 、 亚列利 。
GEN|46|17|亚设 的儿子是 音拿 、 亦施瓦 、 亦施韦 、 比利亚 ，还有他们的妹妹 西拉 。 比利亚 的儿子是 希别 、 玛结 。
GEN|46|18|这是 拉班 给他女儿 利亚 的婢女 悉帕 的儿孙，她为 雅各 所生的共有十六人。
GEN|46|19|雅各 之妻 拉结 的儿子是 约瑟 和 便雅悯 。
GEN|46|20|约瑟 在 埃及 地生了 玛拿西 和 以法莲 ，是 安城 的祭司 波提非拉 的女儿 亚西纳 为 约瑟 生的。
GEN|46|21|便雅悯 的儿子是 比拉 、 比结 、 亚实别 、 基拉 、 乃幔 、 以希 、 罗实 、 母平 、 户平 、 亚勒 。
GEN|46|22|这是 拉结 为 雅各 所生的儿孙，共有十四人。
GEN|46|23|但 的儿子是 户伸 。
GEN|46|24|拿弗他利 的儿子是 雅薛 、 沽尼 、 耶色 、 示冷 。
GEN|46|25|这是 拉班 给他女儿 拉结 的婢女 辟拉 的儿孙，她为 雅各 所生的共有七人。
GEN|46|26|那与 雅各 同到 埃及 的，除了他媳妇之外，凡从他生的共有六十六人。
GEN|46|27|还有 约瑟 在 埃及 所生的两个儿子。到 埃及 的 雅各 全家共有七十人。
GEN|46|28|雅各 派 犹大 先到 约瑟 那里，请他先指示到 歌珊 去的路；于是他们来到了 歌珊 地。
GEN|46|29|约瑟 备好座车，上 歌珊 去迎接他的父亲 以色列 。他见到父亲，就伏在父亲的颈项上，在父亲的颈项上哭了许久。
GEN|46|30|以色列 对 约瑟 说：“我见了你的面，知道你还活着，现在我可以死了。”
GEN|46|31|约瑟 对他兄弟和他父亲的全家说：“我要上去告诉法老，对他说：‘我在 迦南 地的兄弟和我父亲的全家，都到我这里来了。
GEN|46|32|他们是牧羊人，是牧放牲畜的人；他们把羊群牛群和一切所有的都带来了。’
GEN|46|33|等到法老召见你们，说：‘你们是做什么的？’
GEN|46|34|你们就说：‘你的仆人，从幼年直到现在，都是牧放牲畜的人，我们和我们的祖宗都是这样。’如此，你们就可以住在 歌珊 地，因为凡牧羊的都被 埃及 人厌恶。”
GEN|47|1|约瑟 进去告诉法老说：“我的父亲和我的兄弟带着羊群牛群，以及他们一切所有的，从 迦南 地来了。看哪，他们正在 歌珊 地。”
GEN|47|2|约瑟 从他所有兄弟中挑选五个人，引他们到法老面前。
GEN|47|3|法老对 约瑟 的兄弟说：“你们是做什么的？”他们对法老说：“你仆人是牧羊的，我们和我们的祖宗都是这样。”
GEN|47|4|他们又对法老说：“ 迦南 地的饥荒非常严重，仆人的羊群没有牧草，所以我们来到这地寄居。现在求你准许仆人住在 歌珊 地。”
GEN|47|5|法老对 约瑟 说：“你的父亲和你的兄弟到你这里来了，
GEN|47|6|埃及 地都在你面前，只管让你父亲和你兄弟住在最好的地，他们可以住在 歌珊 地。你若知道他们中间有能干的人，就派他们看管我的牲畜。”
GEN|47|7|约瑟 带他父亲 雅各 来，站在法老面前， 雅各 就为法老祝福。
GEN|47|8|法老对 雅各 说：“你平生的年日是多少呢？”
GEN|47|9|雅各 对法老说：“我在世寄居的年日是一百三十年，我一生的岁月又短又苦，比不上我祖先在世寄居的年日。”
GEN|47|10|雅各 又为法老祝福，就从法老面前退出去了。
GEN|47|11|约瑟 安顿他的父亲和兄弟，遵照法老的命令，把 埃及 境内最好的地，就是 兰塞 地，给他们作为产业。
GEN|47|12|约瑟 用粮食供给他父亲和兄弟们，以及他父亲全家的人，照扶养亲属的人口供给。
GEN|47|13|饥荒非常严重，全地都绝了粮， 埃及 地和 迦南 地都因饥荒耗损了。
GEN|47|14|约瑟 收集了 埃及 地和 迦南 地所有的银子，就是众人买粮的银子， 约瑟 就把那些银子都带到法老的宫里。
GEN|47|15|埃及 地和 迦南 地的银子都花光了， 埃及 众人到 约瑟 那里，说：“我们的银子都用完了，求你给我们粮食吧！我们为什么要死在你面前呢？”
GEN|47|16|约瑟 说：“银子若是用完了，可以把你们的牲畜卖给我，我就以你们的牲畜换粮食给你们。”
GEN|47|17|于是他们把牲畜带到 约瑟 那里， 约瑟 就拿粮食换了他们的马、羊、牛、驴；那一年他因换他们一切的牲畜，用粮食养活他们。
GEN|47|18|那一年过去，第二年他们又来到 约瑟 那里，对他说：“不瞒我主，我们的银子都花光了，牲畜也都归于我主了。我们在我主面前，除了自己的身体和土地以外，一无所剩。
GEN|47|19|你为什么要眼看着我们人死地荒呢？求你用粮食买我们和我们的地，我们和我们的地就要为法老效力。求你给我们种子，使我们可以存活，不致死亡，土地也不致荒芜。”
GEN|47|20|于是， 约瑟 为法老买了 埃及 所有的土地， 埃及 人因饥荒所迫，都卖了自己的田地；那些地都归给法老了。
GEN|47|21|至于百姓，从 埃及 边界的一端到另一端， 约瑟 使他们作奴隶。
GEN|47|22|只有祭司的土地， 约瑟 没有买，因为祭司从法老领取薪俸，靠法老的薪俸过活，所以没有卖自己的土地。
GEN|47|23|约瑟 对百姓说：“看哪，我今日为法老买了你们和你们的土地。看，这些种子是给你们的，你们可以耕种土地。
GEN|47|24|将来收割的时候，你们要把五分之一纳给法老，另外四分可以给你们作田地的种子，作你们和你们全家大小的食物。”
GEN|47|25|他们说：“你救了我们的性命，愿我们在我主眼前蒙恩，我们情愿作法老的奴隶。”
GEN|47|26|于是 约瑟 为 埃及 的土地立下定例，直到今日，就是收成的五分之一要归法老。惟独祭司的土地例外，不归于法老。
GEN|47|27|以色列 人住在 埃及 境内的 歌珊 地。他们在那里得了产业，并且生养众多。
GEN|47|28|雅各 住在 埃及 地十七年。 雅各 一生的年日是一百四十七年。
GEN|47|29|以色列 的死期快到了，就叫了他儿子 约瑟 来，对他说：“我若在你眼前蒙恩，把你的手放在我大腿底下，以慈爱和诚实向我承诺，必不将我葬在 埃及 。
GEN|47|30|我与我祖先同睡的时候，你要将我带出 埃及 ，把我葬在他们所葬的地方。” 约瑟 说：“我必遵照你的吩咐去做。”
GEN|47|31|雅各 说：“你向我起誓吧！” 约瑟 就向他起了誓。于是 以色列 在床头 敬拜。
GEN|48|1|这些事以后，有人告诉 约瑟 说：“看哪，你的父亲病了。”他就带着两个儿子 玛拿西 和 以法莲 同去。
GEN|48|2|有人告诉 雅各 说：“看哪，你的儿子 约瑟 到你这里来了。” 以色列 就勉强在床上坐起来。
GEN|48|3|雅各 对 约瑟 说：“全能的上帝曾在 迦南 地的 路斯 向我显现，赐福给我，
GEN|48|4|对我说：‘看哪，我必使你生养众多，成为许多民族，又要将这地赐给你的后裔，永远为业。’
GEN|48|5|我未到 埃及 你那里之前，你在 埃及 地所生的 以法莲 和 玛拿西 这两个儿子，现在他们是我的，正如 吕便 和 西缅 是我的一样。
GEN|48|6|你在他们以后所生的后裔就是你的，这些后裔可以在自己兄弟的名下得产业。
GEN|48|7|至于我，我从 巴旦 回来的时候， 拉结 在我身旁死了，就是在往 迦南 地的路上，离 以法他 还有一段路程。我就把她葬在往 以法他 的路旁； 以法他 就是 伯利恒 。”
GEN|48|8|以色列 看见 约瑟 的儿子，就说：“这些是谁？”
GEN|48|9|约瑟 对他父亲说：“这是上帝在这里赐给我的儿子。” 以色列 说：“领他们到我跟前，我要为他们祝福。”
GEN|48|10|以色列 年纪老迈，眼睛昏花，不能看见。 约瑟 领他们到他跟前，他就和他们亲吻，抱着他们。
GEN|48|11|以色列 对 约瑟 说：“我没有想到能够见你的面。看哪，上帝还让我看见你的儿子。”
GEN|48|12|约瑟 把他们从 以色列 两膝中间领出来，自己脸伏于地下拜。
GEN|48|13|然后， 约瑟 牵着他们两个，带到父亲跟前，右手牵 以法莲 到 以色列 的左边，左手牵 玛拿西 到 以色列 的右边。
GEN|48|14|以色列 却伸出右手来，按在次子 以法莲 的头上，又交叉伸出左手来，按在长子 玛拿西 的头上。
GEN|48|15|他就为 约瑟 祝福说： “愿我祖父 亚伯拉罕 和我父亲 以撒 所事奉的上帝， 就是一生牧养我直到今日的上帝，
GEN|48|16|救赎我脱离一切患难的那位使者，赐福给这两个孩子。 愿我的名，我祖父 亚伯拉罕 和我父亲 以撒 的名藉着他们得以流传。 又愿他们在全地上多多繁衍。”
GEN|48|17|约瑟 见父亲把右手按在 以法莲 的头上，他看为不好，就提起他父亲的手，要从 以法莲 的头上移到 玛拿西 的头上。
GEN|48|18|约瑟 对父亲说：“我父，不是这样。这个才是长子，请你把右手按在他头上。”
GEN|48|19|他父亲却不肯，说：“我知道，我儿，我知道。他也要成为一族，也要强大。可是他的弟弟将来比他还要强大；他弟弟的后裔要成为许多国家。”
GEN|48|20|以色列 就在当日为他们祝福，说：“ 以色列 人要指着你们祝福，说：‘愿上帝使你如 以法莲 、 玛拿西 一样。’”于是他立 以法莲 在 玛拿西 之上。
GEN|48|21|以色列 又对 约瑟 说：“看哪，我快要死了，但上帝必与你们同在，领你们回到你们祖先之地。
GEN|48|22|从前我用刀用弓从 亚摩利 人手下夺取的那一份，我要把它赐给你，使你比你的兄弟多得一份 。”
GEN|49|1|雅各 叫了他的儿子来，说：“你们都来聚集，让我把你们日后要遇到的事告诉你们。
GEN|49|2|雅各 的儿子们，你们要聚集，要聆听， 听你们父亲 以色列 的话。
GEN|49|3|吕便 啊，你是我的长子，我的力量， 我壮年头生之子， 极有尊荣，权力超群。
GEN|49|4|你却放纵如水，必不得居首位； 因为你上了你父亲的床， 你 上了我的榻，污辱了它！
GEN|49|5|西缅 和 利未 是兄弟； 他们的刀剑是残暴的兵器。
GEN|49|6|愿我的心不与他们同谋， 愿我的灵 不与他们合伙； 因为他们在烈怒中杀人， 任意割断牛腿的筋。
GEN|49|7|他们火爆的烈怒可诅， 他们凶残的愤恨可咒！ 我要把他们分散在 雅各 中， 使他们散居在 以色列 。
GEN|49|8|犹大 啊，你的兄弟必赞美你， 你的手必掐住仇敌的颈项， 你父亲的儿子要向你下拜。
GEN|49|9|犹大 是只小狮子； 我儿啊，你捕获了猎物就上去。 他蹲伏，他躺卧，如公狮， 又如母狮，谁敢惹他呢？
GEN|49|10|权杖必不离 犹大 ， 统治者的杖必不离他两脚之间， 直等细罗 来到， 万民都要归顺他。
GEN|49|11|犹大 把小驴拴在葡萄树上， 把驴驹拴在佳美的葡萄树上。 他在葡萄酒中洗衣服， 在葡萄汁 中洗长袍。
GEN|49|12|他的眼睛比 酒红润， 他的牙齿比奶洁白。
GEN|49|13|西布伦 必住在海边， 必成为停船的港口； 他的疆界必延到 西顿 。
GEN|49|14|以萨迦 是匹强壮的驴， 卧在羊圈之中。
GEN|49|15|他看见居所安舒， 土地肥美， 就屈肩负重， 成为服劳役的仆人。
GEN|49|16|但 必为他的百姓伸冤 ， 作为 以色列 支派之一。
GEN|49|17|但 必作道旁的蛇， 路边的毒蛇， 咬伤马蹄， 使骑马的人向后坠落。
GEN|49|18|耶和华啊，我等候你的救恩。
GEN|49|19|迦得 必被袭击者袭击 ， 他却要袭击他们的脚跟。
GEN|49|20|亚设 必出丰盛的粮食， 要供应君王的佳肴。
GEN|49|21|拿弗他利 是被释放的母鹿， 他要生出可爱的小鹿 。
GEN|49|22|约瑟 是多结果子的树枝， 是泉旁多结果的枝子； 他的枝条伸出墙外。
GEN|49|23|弓箭手恶意攻击他， 敌对他，向他射箭。
GEN|49|24|但他的弓仍旧坚硬， 他的手臂灵活敏捷， 这是因 雅各 的大能者的手， 从那里，他是 以色列 的牧者， 以色列 的磐石 。
GEN|49|25|你父亲的上帝必帮助你； 全能者必赐福给你： 天上的福， 深渊下面蕴藏的福， 以及生育哺养的福。
GEN|49|26|你父亲的福 胜过我祖先的福， 直到永世山岭的极限。 这些福必降在 约瑟 的头上， 临到那与兄弟有分别之人的头顶上。
GEN|49|27|便雅悯 是只抓撕掠物的狼， 早晨要吃他的猎物， 晚上要分他的掳物。”
GEN|49|28|这一切是 以色列 的十二个支派。这是他们的父亲对他们所说的话，他按照各人的福分为他们祝福。
GEN|49|29|他又吩咐他们说：“我快要归到我祖先 那里。你们要将我葬在 赫 人 以弗仑 田间的洞里，与我的祖先在一处，
GEN|49|30|就是在 迦南 地 幔利 对面的 麦比拉 田间的洞里，那田是 亚伯拉罕 向 赫 人 以弗仑 买来作坟地的产业。
GEN|49|31|亚伯拉罕 和他的妻子 撒拉 葬在那里； 以撒 和他的妻子 利百加 也葬在那里。我也在那里葬了 利亚 。
GEN|49|32|那块田和田间的洞是向 赫 人买的。”
GEN|49|33|雅各 嘱咐众子完毕后，就把脚收在床上断了气，归到他祖先 那里去了。
GEN|50|1|约瑟 伏在他父亲的脸上，在他脸上哭，又亲他。
GEN|50|2|约瑟 吩咐伺候他的医生们用香料涂他父亲，医生就用香料涂了 以色列 。
GEN|50|3|四十天满了，就是涂香料所规定的日子满了。 埃及 人为他哀哭了七十天。
GEN|50|4|过了哀悼的日子， 约瑟 对法老家中的人说：“我若在你们眼前蒙恩，请你们对法老说：
GEN|50|5|‘我父亲曾叫我起誓说：看哪，我快要死了，你要将我葬在 迦南 地，在我为自己所掘的坟墓里。’现在求你准我上去葬我父亲，然后我必回来。”
GEN|50|6|法老说：“你可以上去，照你父亲叫你起的誓，将他安葬。”
GEN|50|7|于是 约瑟 上去葬他父亲。与他一同上去的有法老的众臣仆和法老家中的长老，以及 埃及 地所有的长老，
GEN|50|8|还有 约瑟 的全家和他的兄弟们，以及他父亲的家属；只留下他们的孩子和羊群牛群在 歌珊 地。
GEN|50|9|又有车辆和驾驶兵和他一同上去，队伍非常庞大。
GEN|50|10|他们到了 约旦河 东 亚达 的禾场，就在那里大大地号啕痛哭。 约瑟 为他父亲哀哭了七天。
GEN|50|11|迦南 的居民看见 亚达 禾场上的哀哭，就说：“这是 埃及 人一场极大的哀哭。”因此那地方名叫 亚伯．麦西 ，是在 约旦河 东。
GEN|50|12|雅各 的儿子们遵照父亲的吩咐去办了，
GEN|50|13|他们把他送到 迦南 地，葬在 幔利 对面的 麦比拉 田间的洞里；那田是 亚伯拉罕 向 赫 人 以弗仑 买来作坟地的产业。
GEN|50|14|约瑟 葬了他父亲以后，就和他的兄弟，以及所有同他上去葬他父亲的人，都回 埃及 去了。
GEN|50|15|约瑟 的哥哥们见父亲死了，就说：“也许 约瑟 仍然怀恨我们，会照我们从前待他一切的恶，重重报复我们。”
GEN|50|16|他们就传口信给 约瑟 说：“你父亲未死之前曾吩咐说：
GEN|50|17|‘你们要对 约瑟 这样说：从前你哥哥们恶待你，你要饶恕他们的过犯和罪恶。’现在求你饶恕你父亲的上帝之仆人们的过犯。”他们对 约瑟 说了这话， 约瑟 就哭了。
GEN|50|18|他的哥哥们又来俯伏在他面前，说：“看哪，我们是你的奴隶。”
GEN|50|19|约瑟 对他们说：“不要怕，我岂能代替上帝呢？
GEN|50|20|从前你们的意思是要害我，但上帝的意思原是好的，要使许多百姓得以存活，成就今日的光景。
GEN|50|21|现在你们不要害怕，我必养活你们和你们的孩子。”于是 约瑟 安慰他们，讲了使他们安心的话。
GEN|50|22|约瑟 和他父亲的家属都住在 埃及 。 约瑟 活了一百一十年。
GEN|50|23|约瑟 看到 以法莲 第三代的子孙。 玛拿西 的孙子， 玛吉 的儿子，出生时都放在 约瑟 的膝上。
GEN|50|24|约瑟 对他的兄弟说：“我快要死了，但上帝必定看顾你们，领你们从这地上去，到他起誓应许给 亚伯拉罕 、 以撒 、 雅各 之地。”
GEN|50|25|约瑟 叫 以色列 的子孙起誓：“上帝必定眷顾你们，你们要把我的骸骨从这里带上去。”
GEN|50|26|约瑟 死了，那时他一百一十岁。人用香料涂了他，把他收殓在棺材里，停放在 埃及 。
EXOD|1|1|以色列 的众儿子各带着家眷，和 雅各 一同来到 埃及 ，他们的名字如下：
EXOD|1|2|吕便 、 西缅 、 利未 、 犹大 、
EXOD|1|3|以萨迦 、 西布伦 、 便雅悯 、
EXOD|1|4|但 、 拿弗他利 、 迦得 、 亚设 。
EXOD|1|5|凡从 雅各 生的，共有七十人。那时， 约瑟 已经在 埃及 。
EXOD|1|6|约瑟 和他所有的兄弟，以及那一代的人都死了。
EXOD|1|7|然而， 以色列 人生养众多，繁衍昌盛，极其强盛，遍满了那地。
EXOD|1|8|有一位不认识 约瑟 的新王兴起，统治 埃及 。
EXOD|1|9|他对自己的百姓说：“看哪， 以色列 人的百姓比我们还多，又比我们强盛。
EXOD|1|10|来吧，让我们机巧地待他们，恐怕他们增多起来，将来若有战争，他们就联合我们的仇敌来攻击我们，然后离开这地去了。”
EXOD|1|11|于是 埃及 人派监工管辖他们，用劳役苦待他们。他们为法老建造储货城，就是 比东 和 兰塞 。
EXOD|1|12|可是越苦待他们，他们就越发增多，更加繁衍， 埃及 人就因 以色列 人愁烦。
EXOD|1|13|埃及 人严厉地强迫 以色列 人做工，
EXOD|1|14|使他们因苦工而生活痛苦；无论是和泥，是做砖，是做田间各样的工，一切的工 埃及 人都严厉地对待他们。
EXOD|1|15|埃及 王又对 希伯来 的接生婆，一个名叫 施弗拉 ，另一个名叫 普阿 的说：
EXOD|1|16|“你们为 希伯来 妇人接生，临盆的时候要注意 ，若是男的，就把他杀了，若是女的，就让她活。”
EXOD|1|17|但是接生婆敬畏上帝，不照 埃及 王的吩咐去做，却让男孩活着。
EXOD|1|18|埃及 王召了接生婆来，对她们说：“你们为什么做这事，让男孩活着呢？”
EXOD|1|19|接生婆对法老说：“因为 希伯来 妇人与 埃及 妇人不同； 希伯来 妇人健壮，接生婆还没有到，她们已经生产了。”
EXOD|1|20|上帝恩待接生婆； 以色列 人增多起来，极其强盛。
EXOD|1|21|接生婆因为敬畏上帝，上帝就叫她们成立家室。
EXOD|1|22|法老吩咐他的众百姓说：“把所生的 每一个男孩都丢到 尼罗河 里去，让所有的女孩存活。”
EXOD|2|1|有一个 利未 家的人娶了一个 利未 女子为妻。
EXOD|2|2|那女人怀孕，生了一个儿子，见他俊美，就把他藏了三个月，
EXOD|2|3|后来不能再藏，就取了一个蒲草箱，抹上柏油和树脂，将孩子放在里面，把箱子搁在 尼罗河 边的芦苇中。
EXOD|2|4|孩子的姊姊远远站着，要知道他究竟会怎样。
EXOD|2|5|法老的女儿来到 尼罗河 边洗澡，她的女仆们在河边行走。她看见在芦苇中的箱子，就派一个使女把它拿来。
EXOD|2|6|她打开箱子，看见那孩子。看哪，男孩在哭，她就可怜他，说：“这是 希伯来 人的一个孩子。”
EXOD|2|7|孩子的姊姊对法老的女儿说：“我去叫一个 希伯来 妇人来作奶妈，替你乳养这孩子，好吗？”
EXOD|2|8|法老的女儿对她说：“去吧！”那女孩就去叫了孩子的母亲来。
EXOD|2|9|法老的女儿对她说：“你把这孩子抱去，替我乳养这孩子，我必给你工钱。”那妇人就把孩子接过来，乳养他。
EXOD|2|10|孩子长大了，妇人把他带到法老的女儿那里，就作了她的儿子。她给孩子起名叫 摩西 ，说：“因我把他从水里拉出来。”
EXOD|2|11|过了一段日子， 摩西 长大了，他出去到他同胞那里，看见他们的劳役。他看见一个 埃及 人打他的同胞，一个 希伯来 人。
EXOD|2|12|他左右观看，见没有人，就把 埃及 人打死了，藏在沙土里。
EXOD|2|13|第二天他出去，看哪，有两个 希伯来 人在打架，他就对那凶恶的人说：“你为什么打你同族的人呢？”
EXOD|2|14|那人说：“谁立你作我们的领袖和审判官呢？难道你要杀我，像杀那 埃及 人一样吗？” 摩西 就惧怕，说：“这事一定是让人知道了。”
EXOD|2|15|法老听见这事，就设法要杀 摩西 。于是 摩西 逃走，躲避法老，到了 米甸 地，坐在井旁。
EXOD|2|16|米甸 的祭司有七个女儿；她们来打水，打满了槽，要给父亲的羊群喝水。
EXOD|2|17|有一些牧羊人来，把她们赶走， 摩西 却起来帮助她们，取水给她们的羊群喝。
EXOD|2|18|她们回到父亲 流珥 那里；他说：“今日你们为何这么快就回来了呢？”
EXOD|2|19|她们说：“有一个 埃及 人来救我们脱离牧羊人的手，他甚至打水给我们的羊群喝。”
EXOD|2|20|他对女儿们说：“那人在哪里？你们为什么撇下他呢？去请他来吃饭吧！”
EXOD|2|21|摩西 愿意和那人同住， 那人就把女儿 西坡拉 给 摩西 为妻。
EXOD|2|22|西坡拉 生了一个儿子， 摩西 给他起名叫 革舜 ，因他说：“我在外地作了寄居者。”
EXOD|2|23|过了许多年， 埃及 王死了。 以色列 人因做苦工，就叹息哀求；他们因苦工所发出的哀声达于上帝。
EXOD|2|24|上帝听见他们的哀声，就记念他与 亚伯拉罕 、 以撒 、 雅各 所立的约。
EXOD|2|25|上帝看顾 以色列 人，上帝是知道的 。
EXOD|3|1|摩西 牧放他岳父 米甸 祭司 叶特罗 的羊群，他领羊群往旷野的那一边去，到了上帝的山，就是 何烈山 。
EXOD|3|2|耶和华的使者在荆棘的火焰中向他显现。 摩西 观看，看哪，荆棘在火中焚烧，却没有烧毁。
EXOD|3|3|摩西 说：“我要转过去看这大异象，这荆棘为何没有烧毁呢？”
EXOD|3|4|耶和华见 摩西 转过去看，上帝就从荆棘里呼叫他说：“ 摩西 ！ 摩西 ！”他说：“我在这里。”
EXOD|3|5|上帝说：“不要靠近这里。把你脚上的鞋脱下来，因为你所站的地方是圣地”。
EXOD|3|6|他又说：“我是你父亲的上帝，是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。” 摩西 蒙上脸，因为怕看上帝。
EXOD|3|7|耶和华说：“我确实看见了我百姓在 埃及 所受的困苦，我也听见了他们因受监工苦待所发的哀声；我确实知道他们的痛苦。
EXOD|3|8|我下来是要救他们脱离 埃及 人的手，领他们从那地上来，到美好与宽阔之地，到流奶与蜜之地，就是 迦南 人、 赫 人、 亚摩利 人、 比利洗 人、 希未 人、 耶布斯 人之地。
EXOD|3|9|现在，看哪， 以色列 人的哀声达到我这里，我也看见 埃及 人怎样欺压他们。
EXOD|3|10|现在，你去，我要差派你到法老那里，把我的百姓 以色列 人从 埃及 领出来。”
EXOD|3|11|摩西 对上帝说：“我是什么人，竟能去见法老，把 以色列 人从 埃及 领出来呢？”
EXOD|3|12|上帝说：“我必与你同在。这就是我差派你去，给你的凭据：你把百姓从 埃及 领出来之后，你们必在这山上事奉上帝。”
EXOD|3|13|摩西 对上帝说：“看哪，我到 以色列 人那里，对他们说：‘你们祖宗的上帝差派我到你们这里来。’他们若对我说：‘他叫什么名字？’我要对他们说什么呢？”
EXOD|3|14|上帝对 摩西 说：“我是自有永有的”；又说：“你要对 以色列 人这样说：‘那自有永有的差派我到你们这里来。’”
EXOD|3|15|上帝又对 摩西 说：“你要对 以色列 人这样说：‘耶和华－你们祖宗的上帝，就是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝差派我到你们这里来。’这是我的名，直到永远；这也是我的称号 ，直到万代。
EXOD|3|16|你去召集 以色列 的长老，对他们说：‘耶和华－你们祖宗的上帝，就是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝向我显现，说：我实在眷顾了你们，眷顾你们在 埃及 的遭遇。
EXOD|3|17|我也曾说：要把你们从 埃及 的困苦中领出来，往 迦南 人、 赫 人、 亚摩利 人、 比利洗 人、 希未 人、 耶布斯 人的地去，就是到流奶与蜜之地。’
EXOD|3|18|他们必听你的话。你和 以色列 的长老要到 埃及 王那里，对他说：‘耶和华－ 希伯来 人的上帝向我们显现，现在求你让我们往旷野去，走三天的路程，为要向耶和华我们的上帝献祭。’
EXOD|3|19|我知道若不用大能的手， 埃及 王不会放你们走。
EXOD|3|20|因此，我必伸出我的手，在 埃及 施行我一切的神迹，击打这地，然后，他才放你们走。
EXOD|3|21|我必使 埃及 人看得起你们，你们离开的时候就不至于空手而去。
EXOD|3|22|每一个妇女必向她的邻舍，以及寄居在她家里的女人，索取金器、银器和衣裳，给你们的儿女穿戴。这样你们就掠夺了 埃及 人。”
EXOD|4|1|摩西 回答说：“看哪！他们不会信我，也不会听我的话，因为他们必说：‘耶和华并没有向你显现。’”
EXOD|4|2|耶和华对 摩西 说：“你手里的是什么？”他说：“是杖。”
EXOD|4|3|耶和华说：“把它丢在地上！”他一丢在地上，杖就变成一条蛇； 摩西 逃走避开它。
EXOD|4|4|耶和华对 摩西 说：“伸出手来，拿住它的尾巴─ 摩西 就伸出手，抓住它，它就在 摩西 的手掌中变为杖─
EXOD|4|5|为了要使他们信耶和华他们祖宗的上帝，就是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝，曾向你显现了。”
EXOD|4|6|耶和华又对他说：“把手放进怀里。”他就把手放进怀里。当他把手抽出来，看哪，手竟然长了痲疯 ，像雪一样白。
EXOD|4|7|耶和华说：“把手放回怀里─他就把手放回怀里。当他把手从怀里再抽出来，看哪，手复原了，与全身的肉一样─
EXOD|4|8|倘若他们不信你，也不听第一个神迹的声音，他们会信第二个神迹的声音。
EXOD|4|9|倘若他们不信这两个神迹，不听你的话，你就从 尼罗河 里取些水，倒在干的地上。你从 尼罗河 里所取的水必在干地上变成血。”
EXOD|4|10|摩西 对耶和华说：“主啊，求求你，我并不是一个能言善道的人，以前这样，就是你对仆人说话以后也是这样，因为我是拙口笨舌的。”
EXOD|4|11|耶和华对他说：“谁造人的口呢？谁使人口哑、耳聋、目明、眼瞎呢？岂不是我－耶和华吗？
EXOD|4|12|现在，去吧，我必赐你口才，指教你应当说的。”
EXOD|4|13|摩西 说：“主啊，求求你，你要藉着谁的手，就差派谁去吧！”
EXOD|4|14|耶和华的怒气向 摩西 发作，说：“你不是有一个哥哥 利未 人 亚伦 吗？我知道他是个能言善道的人。看哪，他正出来迎接你。他一见到你，心里就欢喜。
EXOD|4|15|你要跟他说话，把话放在他的口里，我要赐你口才，也要赐他口才，又要教你们做当做的事。
EXOD|4|16|他要替你向百姓说话；他要当你的口，你要当他的上帝。
EXOD|4|17|你手里要拿这杖，用它来行神迹。”
EXOD|4|18|于是， 摩西 回到他岳父 叶特罗 那里，对他说：“请你让我回 埃及 我同胞那里，看他们还在不在。” 叶特罗 对 摩西 说：“平平安安地去吧！”
EXOD|4|19|耶和华在 米甸 对 摩西 说：“你要回 埃及 去，因为那些寻索你命的人都死了。”
EXOD|4|20|摩西 就带着妻子和两个儿子，让他们骑上驴，回 埃及 地去。 摩西 手里拿着上帝的杖。
EXOD|4|21|耶和华对 摩西 说：“你回到 埃及 去的时候，要留意将我交在你手中的一切奇事行在法老面前。但我要任凭他的心刚硬，他必不放百姓走。
EXOD|4|22|你要对法老说：‘耶和华如此说： 以色列 是我的儿子，我的长子。
EXOD|4|23|我对你说过：放我的儿子走，好事奉我。你还是不肯放他走。看哪，我要杀你头生的儿子。’”
EXOD|4|24|在路上住宿的地方，耶和华遇见 摩西 ，想要杀他。
EXOD|4|25|西坡拉 就拿一块火石，割下她儿子的包皮，碰触 摩西 的脚，说：“你真是我血的新郎了。”
EXOD|4|26|这样，耶和华才放了他。那时， 西坡拉 说：“你因割礼就是血的新郎 了”。
EXOD|4|27|耶和华对 亚伦 说：“你往旷野去迎接 摩西 。”他就去，在上帝的山遇见 摩西 ，就亲他。
EXOD|4|28|摩西 将耶和华差派他所说的话和吩咐他所行的神迹都告诉了 亚伦 。
EXOD|4|29|摩西 和 亚伦 就去召集 以色列 的众长老。
EXOD|4|30|亚伦 将耶和华对 摩西 所说的一切话述说了一遍，又在百姓眼前行了那些神迹，
EXOD|4|31|百姓就信了。他们听见耶和华眷顾 以色列 人，鉴察他们的困苦，就低头敬拜。
EXOD|5|1|后来， 摩西 和 亚伦 去对法老说：“耶和华－ 以色列 的上帝这样说：‘放我的百姓走，好让他们在旷野向我守节。’”
EXOD|5|2|法老说：“耶和华是谁，要我听他的话，让 以色列 人去？我不认识耶和华，也不放 以色列 人走！”
EXOD|5|3|他们说：“ 希伯来 人的上帝已向我们显现了。求你让我们往旷野去，走三天的路程，向耶和华我们的上帝献祭，免得他用瘟疫、刀剑攻击我们。”
EXOD|5|4|埃及 王对他们说：“ 摩西 、 亚伦 ！你们为什么叫百姓不做工呢？去，服你们的劳役吧！”
EXOD|5|5|他又说：“看哪，这地的 以色列 人如今这么多，你们竟然叫他们歇下劳役！”
EXOD|5|6|当天，法老吩咐监工和工头说：
EXOD|5|7|“你们不可照以前一样提供草给百姓做砖，要叫他们自己去捡草。
EXOD|5|8|他们平时做砖的数目，你们仍旧向他们要，一点不可减少，因为他们是懒惰的，所以才呼求说：‘让我们去向我们的上帝献祭。’
EXOD|5|9|你们要把更重的工作加在这些人身上，使他们在其中劳碌，不去理会谎言。”
EXOD|5|10|监工和工头出来对百姓说：“法老这样说：‘我不给你们草，
EXOD|5|11|你们自己在哪里能找到草，就往哪里去找吧！但你们的工作一点也不可减少。’”
EXOD|5|12|于是，百姓分散在 埃及 全地，捡碎秸当草用。
EXOD|5|13|监工催逼他们，说：“你们每天要做完一天的工，与先前有草一样。”
EXOD|5|14|法老的监工击打他们所派的 以色列 工头，说：“为什么昨天和今天你们没有按照以前做砖的数目，完成你们的工作呢？”
EXOD|5|15|以色列 人的工头来哀求法老说：“为什么这样待你的仆人呢？
EXOD|5|16|监工不把草给仆人，并且对我们说：‘做砖吧！’看哪，你仆人挨了打，其实是你百姓的错。”
EXOD|5|17|法老却说：“懒惰，你们真是懒惰！所以你们说：‘让我们去向耶和华献祭吧。’
EXOD|5|18|现在，去做工吧！草是不会给你们，砖却要如数交纳。”
EXOD|5|19|以色列 人的工头听见“你们每天做砖的工作一点也不可减少”，就知道惹上祸了。
EXOD|5|20|他们离开法老出来，正遇见 摩西 和 亚伦 站在那里等候他们，
EXOD|5|21|就向他们说：“愿耶和华鉴察你们，施行判断，因为你们使我们在法老和他臣仆面前有了臭名，把刀递在他们手中来杀我们。”
EXOD|5|22|摩西 回到耶和华那里，说：“主啊，你为什么苦待这百姓呢？为什么差派我呢？
EXOD|5|23|自从我到法老那里，奉你的名说话，他就苦待这百姓，你却一点也没有拯救你的百姓。”
EXOD|6|1|耶和华对 摩西 说：“现在你必看见我向法老所行的事，使他因我大能的手放 以色列 人走，因我大能的手把他们赶出他的地。”
EXOD|6|2|上帝吩咐 摩西 ，对他说：“我是耶和华。
EXOD|6|3|我从前向 亚伯拉罕 、 以撒 、 雅各 显现为全能的上帝；至于我的名耶和华，我未曾让他们知道。
EXOD|6|4|我要与他们坚立我的约，要把 迦南 地，他们寄居的地赐给他们。
EXOD|6|5|我听见 以色列 人被 埃及 人奴役的哀声，我就记念我的约。
EXOD|6|6|所以你要对 以色列 人说：‘我是耶和华；我要除去 埃及 人加给你们的劳役，救你们脱离他们的奴役。我要用伸出来的膀臂，藉严厉的惩罚救赎你们。
EXOD|6|7|我要以你们为我的百姓，我也要作你们的上帝。我除去 埃及 人加给你们的劳役，你们就知道我是耶和华你们的上帝。
EXOD|6|8|我起誓应许给 亚伯拉罕 、 以撒 、 雅各 的地，我要领你们进去，将那地赐给你们为业。我是耶和华。’”
EXOD|6|9|摩西 把这话告诉 以色列 人，但是他们因心里愁烦，又因苦工，就不肯听 摩西 的话。
EXOD|6|10|耶和华吩咐 摩西 说：
EXOD|6|11|“你去对 埃及 王法老说，让 以色列 人离开他的地。”
EXOD|6|12|摩西 在耶和华面前说：“看哪， 以色列 人尚且不听我，法老怎么会听我这不会讲话的人呢？”
EXOD|6|13|耶和华吩咐 摩西 和 亚伦 ，命令他们到 以色列 人和 埃及 王法老那里，把 以色列 人从 埃及 地领出来。
EXOD|6|14|以色列 人族长的名字如下： 以色列 长子 吕便 的儿子是 哈诺 、 法路 、 希斯伦 、 迦米 ；这是 吕便 的家族。
EXOD|6|15|西缅 的儿子是 耶母利 、 雅悯 、 阿辖 、 雅斤 、 琐辖 ，和 迦南 女子生的儿子 扫罗 ；这是 西缅 的家族。
EXOD|6|16|以下是 利未 的儿子按着家谱的名字： 革顺 、 哥辖 、 米拉利 。 利未 一生的岁数是一百三十七岁。
EXOD|6|17|革顺 的儿子按着家族是 立尼 、 示每 。
EXOD|6|18|哥辖 的儿子是 暗兰 、 以斯哈 、 希伯伦 、 乌薛 。 哥辖 一生的岁数是一百三十三岁。
EXOD|6|19|米拉利 的儿子是 抹利 和 母示 ；这是 利未 按着家谱的家族。
EXOD|6|20|暗兰 娶了他父亲的妹妹 约基别 为妻，她为他生了 亚伦 和 摩西 。 暗兰 一生的岁数是一百三十七岁。
EXOD|6|21|以斯哈 的儿子是 可拉 、 尼斐 、 细基利 。
EXOD|6|22|乌薛 的儿子是 米沙利 、 以利撒反 、 西提利 。
EXOD|6|23|亚伦 娶了 亚米拿达 的女儿， 拿顺 的妹妹， 以利沙巴 为妻，她为他生了 拿答 、 亚比户 、 以利亚撒 、 以他玛 。
EXOD|6|24|可拉 的儿子是 亚惜 、 以利加拿 、 亚比亚撒 ；这是 可拉 的家族。
EXOD|6|25|亚伦 的儿子 以利亚撒 娶了 普铁 的一个女儿为妻，她为他生了 非尼哈 。这是 利未 人按着家族的族长。
EXOD|6|26|这就是曾听见耶和华说“把 以色列 人按着队伍从 埃及 地领出来”的 亚伦 和 摩西 ，
EXOD|6|27|对 埃及 王法老说要将 以色列 人从 埃及 领出来的，也是这 摩西 和 亚伦 。
EXOD|6|28|当耶和华在 埃及 地对 摩西 说话的时候，
EXOD|6|29|耶和华对 摩西 说：“我是耶和华；我对你所说的一切话，你都要告诉 埃及 王法老。”
EXOD|6|30|摩西 在耶和华面前说：“看哪，我是不会讲话的人，法老怎么会听我呢？”
EXOD|7|1|耶和华对 摩西 说：“我使你在法老面前像上帝一样，你的哥哥 亚伦 是你的代言人 。
EXOD|7|2|凡我所吩咐你的，你都要说。你的哥哥 亚伦 要对法老说，让 以色列 人离开他的地。
EXOD|7|3|我要使法老的心固执，我也要在 埃及 地多行神迹奇事。
EXOD|7|4|法老必不听从你们，因此我要伸手严厉地惩罚 埃及 ，把我的军队，就是我的百姓 以色列 人从 埃及 地领出来。
EXOD|7|5|我伸手攻击 埃及 ，把 以色列 人从他们中间领出来的时候， 埃及 人就知道我是耶和华。”
EXOD|7|6|摩西 和 亚伦 就去做；他们照耶和华吩咐的去做了。
EXOD|7|7|摩西 和 亚伦 与法老说话的时候， 摩西 八十岁， 亚伦 八十三岁。
EXOD|7|8|耶和华对 摩西 和 亚伦 说：
EXOD|7|9|“法老若吩咐你们说：‘你们行一件奇事吧！’你就对 亚伦 说：‘把杖丢在法老面前！杖会变成蛇。’”
EXOD|7|10|摩西 和 亚伦 到法老那里去，照耶和华所吩咐的去做。 亚伦 把杖丢在法老和他臣仆面前，杖就变成蛇。
EXOD|7|11|法老也召了智慧人和行邪术的人来，这些 埃及 术士也用邪术照样做。
EXOD|7|12|他们各人丢下自己的杖，杖就变成蛇；但 亚伦 的杖吞了他们的杖。
EXOD|7|13|法老心里刚硬，不听 摩西 和 亚伦 ，正如耶和华所说的。
EXOD|7|14|耶和华对 摩西 说：“法老心硬，不肯放百姓走。
EXOD|7|15|明天早晨你要到法老那里去，看哪，他出来往水边去，你要到 尼罗河 边去迎见他，手里拿着那根变过蛇的杖。
EXOD|7|16|你要对他说：‘耶和华－ 希伯来 人的上帝差派我到你这里，说：放我的百姓走，到旷野事奉我。看哪，到如今你还是不听。
EXOD|7|17|耶和华如此说：看哪，我要用我手里的杖击打 尼罗河 中的水，水就变成血；这样，你就知道我是耶和华。
EXOD|7|18|河里的鱼必死，河也要发臭， 埃及 人就厌恶喝这河里的水。’”
EXOD|7|19|耶和华对 摩西 说：“你要对 亚伦 说：‘拿你的杖，伸出你的手在 埃及 所有的水上，在他们的江、河、池塘，所有水聚集的地方上，叫水变成血。在 埃及 全地，无论在木器中，石器中，都必有血。’”
EXOD|7|20|摩西 和 亚伦 就照耶和华所吩咐的去做。 亚伦 在法老和他臣仆眼前举杖击打 尼罗河 里的水，河里的水都变成血了。
EXOD|7|21|河里的鱼死了，河也臭了， 埃及 人就不能喝这河里的水； 埃及 遍地都有了血。
EXOD|7|22|但是， 埃及 的术士也用邪术照样做了；法老心里刚硬，不听 摩西 和 亚伦 ，正如耶和华所说的。
EXOD|7|23|法老转身回宫去，并不把这事放在心上。
EXOD|7|24|所有的 埃及 人都沿着 尼罗河 边挖掘，要找水喝，因为他们不能喝河里的水。
EXOD|7|25|耶和华击打 尼罗河 后，过了七天。
EXOD|8|1|耶和华对 摩西 说：“你要到法老那里，对他说：‘耶和华如此说：放我的百姓走，好事奉我。
EXOD|8|2|你若不肯放他们走，看哪，我必以青蛙之灾击打你的疆土。
EXOD|8|3|尼罗河 要滋生青蛙；这青蛙要上来进你的宫殿和你的卧房，上你的床榻，进你臣仆的房屋，上你百姓的身上，进你的炉灶和你的揉面盆。
EXOD|8|4|这些青蛙要跳上你、你百姓和你众臣仆的身上。’”
EXOD|8|5|耶和华对 摩西 说：“你要对 亚伦 说：‘伸出你手里的杖在江、河、池塘上，把青蛙带上 埃及 地来。’”
EXOD|8|6|亚伦 伸手在 埃及 的众水上，青蛙就上来，遮满了 埃及 地。
EXOD|8|7|术士也用他们的邪术照样去做，把青蛙带上 埃及 地。
EXOD|8|8|法老召 摩西 和 亚伦 来，说：“请你们祈求耶和华使这些青蛙离开我和我的百姓，我就让这百姓去向耶和华献祭。”
EXOD|8|9|摩西 对法老说：“悉听尊便，告诉我何时为你、你臣仆和你的百姓祈求，使青蛙被剪除，离开你和你的宫殿，只留在 尼罗河 里。”
EXOD|8|10|他说：“明天。” 摩西 说：“就照你的话吧，为要叫你知道没有像耶和华我们上帝的，
EXOD|8|11|青蛙必会离开你、你宫殿、你臣仆和你的百姓，只留在 尼罗河 里。”
EXOD|8|12|于是 摩西 和 亚伦 离开法老出去。 摩西 为了青蛙的事呼求耶和华，因为他带来青蛙搅扰法老。
EXOD|8|13|耶和华就照 摩西 的请求去做；在屋里、院中、田间的青蛙都死了。
EXOD|8|14|众人把青蛙聚拢成堆，地就发出臭气。
EXOD|8|15|但法老见灾祸舒缓了，就硬着心，不听从他们，正如耶和华所说的。
EXOD|8|16|耶和华对 摩西 说：“你要对 亚伦 说：‘伸出你的杖击打地上的尘土，使尘土在 埃及 全地变成蚊子 。’”
EXOD|8|17|他们就照样做了。 亚伦 伸出他手里的杖，击打地上的尘土，人和牲畜身上就有了蚊子； 埃及 全地的尘土都变成蚊子了。
EXOD|8|18|术士也用邪术要照样产生蚊子，却做不成。于是人和牲畜的身上都有了蚊子。
EXOD|8|19|术士对法老说：“这是上帝的手指。”法老心里刚硬，不听 摩西 和 亚伦 ，正如耶和华所说的。
EXOD|8|20|耶和华对 摩西 说：“你要清早起来，站在法老面前。看哪，法老来到水边，你就对他说：‘耶和华如此说：放我的百姓走，好事奉我。
EXOD|8|21|你若不放我的百姓走，看哪，我要派成群的苍蝇到你、你臣仆和你百姓身上，进你的宫殿； 埃及 人的房屋和他们所住的地都要满了成群的苍蝇。
EXOD|8|22|那一日，我必把我百姓所住的 歌珊 地分别出来，使那里没有成群的苍蝇，好叫你知道我─耶和华是在全地之中。
EXOD|8|23|我要施行救赎，区隔我的百姓和你的百姓。明天必有这神迹。’”
EXOD|8|24|耶和华就这样做了。大群的苍蝇进入法老的宫殿和他臣仆的房屋；在 埃及 全地，地就因这成群的苍蝇毁坏了。
EXOD|8|25|法老召了 摩西 和 亚伦 来，说：“去，在此地向你们的上帝献祭。”
EXOD|8|26|摩西 说：“这样做是不妥的，因为我们要献给耶和华－我们上帝的祭物是 埃及 人所厌恶的；看哪，我们在 埃及 人眼前献他们所厌恶的，他们岂不拿石头打死我们吗？
EXOD|8|27|我们要遵照耶和华－我们上帝所吩咐我们的，往旷野去，走三天路程，向他献祭。”
EXOD|8|28|法老说：“我可以放你们走，在旷野向耶和华－你们的上帝献祭，只是不可走得太远。你们要为我祈祷。”
EXOD|8|29|摩西 说：“看哪，我要从你这里出去祈求耶和华，使成群的苍蝇明天离开法老、法老的臣仆和法老的百姓；法老却不可再欺骗，不让百姓去向耶和华献祭。”
EXOD|8|30|于是 摩西 离开法老，去祈求耶和华。
EXOD|8|31|耶和华就照 摩西 的请求去做，使成群的苍蝇离开法老、他的臣仆和他的百姓，一只也没有留下。
EXOD|8|32|但这一次法老又硬着心，不放百姓走。
EXOD|9|1|耶和华对 摩西 说：“你要到法老那里，对他说：‘耶和华－ 希伯来 人的上帝如此说：放我的百姓走，好事奉我。
EXOD|9|2|你若不肯放他们走，仍要强留他们，
EXOD|9|3|看哪，耶和华的手必以严重的瘟疫加在你田间的牲畜上，就是在马、驴、骆驼、牛群和羊群的身上。
EXOD|9|4|耶和华却要分别 以色列 的牲畜和 埃及 的牲畜，凡属 以色列 人的，一只都不死。’”
EXOD|9|5|耶和华就设定时间，说：“明天耶和华必在此地行这事。”
EXOD|9|6|第二天，耶和华行了这事。 埃及 的牲畜全都死了，只是 以色列 人的牲畜，一只都没有死。
EXOD|9|7|法老派人去，看哪， 以色列 人的牲畜连一只都没有死。可是法老硬着心，不放百姓走。
EXOD|9|8|耶和华对 摩西 和 亚伦 说：“你们从炉里满满捧出炉灰， 摩西 要在法老眼前把它撒在空中。
EXOD|9|9|这灰要在 埃及 全地变成尘土，使 埃及 全地的人和牲畜身上起泡生疮。”
EXOD|9|10|摩西 和 亚伦 取了炉灰，站在法老面前。 摩西 把它撒在空中，人和牲畜的身上就起泡生疮了。
EXOD|9|11|因为这疮，术士在 摩西 面前站立不住，术士和所有 埃及 人的身上都生了疮。
EXOD|9|12|但耶和华任凭法老的心刚硬，不听 摩西 和 亚伦 ，正如耶和华对 摩西 所说的。
EXOD|9|13|耶和华对 摩西 说：“你要清早起来，站在法老面前，对他说：‘耶和华－ 希伯来 人的上帝如此说：放我的百姓走，好事奉我。
EXOD|9|14|因为这一次我要使一切的灾祸临到你自己，你臣仆和你百姓的身上，为要叫你知道在全地没有像我的。
EXOD|9|15|现在，我若伸手用瘟疫攻击你和你的百姓，你就会从地上除灭了。
EXOD|9|16|然而，我让你存活，是为了要使你看见我的大能，并要使我的名传遍全地。
EXOD|9|17|可是你仍然向我的百姓自高自大，不放他们走。
EXOD|9|18|看哪，明天大约这时候，我必使大量的冰雹降下，这是从 埃及 立国直到如今没有出现过的。
EXOD|9|19|现在，你要派人把你的牲畜和你田间一切所有的带去躲避；任何在田间，无论是人是牲畜没有回到屋内的，冰雹必降在他们身上，他们就必死。’”
EXOD|9|20|法老的臣仆中，惧怕耶和华这话的，就让他的奴仆和牲畜逃进屋里。
EXOD|9|21|但那不把耶和华这话放在心上的，就把他的奴仆和牲畜留在田里。
EXOD|9|22|耶和华对 摩西 说：“你向天伸出你的手，使冰雹降在 埃及 全地，降在 埃及 地的人和牲畜身上，以及田间各样菜蔬上。”
EXOD|9|23|摩西 向天伸杖，耶和华就打雷下雹，有火降到地上；耶和华下雹在 埃及 地上。
EXOD|9|24|那时，有雹，也有火在雹中闪烁，极其严重；自从 埃及 立国以来，全地没有像这样的。
EXOD|9|25|在 埃及 全地，冰雹击打田间所有的人和牲畜，击打一切的菜蔬，也打坏了田间一切的树木。
EXOD|9|26|惟独 以色列 人所住的 歌珊 地没有冰雹。
EXOD|9|27|法老差派人去召 摩西 和 亚伦 来，对他们说：“这一次我犯罪了。耶和华是公义的；我和我的百姓是邪恶的。
EXOD|9|28|请你们祈求耶和华，因上帝的雷轰和冰雹已经够了。我要放你们走，你们不用再留下来了。”
EXOD|9|29|摩西 对他说：“我一出城就向耶和华举起双手；雷必止住，也不再有冰雹，叫你知道地是属于耶和华的。
EXOD|9|30|至于你和你的臣仆，我知道你们仍然不敬畏耶和华上帝。”
EXOD|9|31|那时，亚麻和大麦被摧毁了，因为大麦已经吐穗，亚麻也开了花。
EXOD|9|32|只是小麦和粗麦没有被摧毁，因为它们还没有长成。
EXOD|9|33|摩西 离开法老出了城，向耶和华举起双手，雷和雹就止住，雨也不再下在地上了。
EXOD|9|34|法老见雨、雹、雷止住，又再犯罪；他和他的臣仆都硬着心。
EXOD|9|35|法老的心刚硬，不放 以色列 人走，正如耶和华藉着 摩西 所说的。
EXOD|10|1|耶和华对 摩西 说：“你要到法老那里，因我使他硬着心，也使他臣仆硬着心，为要在他们中间 显出我的这些神迹来，
EXOD|10|2|并要叫你将我严厉对付 埃及 的事，和在他们中间所行的神迹，传于儿子和孙子的耳中，好叫你们知道我是耶和华。”
EXOD|10|3|摩西 和 亚伦 就到法老那里，对他说：“耶和华－ 希伯来 人的上帝这样说：‘你在我面前不肯谦卑要到几时呢？放我的百姓走，好事奉我。
EXOD|10|4|你若不肯放我的百姓走，看哪，明天我要使蝗虫进入你的境内，
EXOD|10|5|遮满地面 ，甚至地也看不见了。它们要吃那冰雹后所剩，就是留给你们的；并且要吃那生长在田间的一切树木。
EXOD|10|6|你的宫殿和你众臣仆的房屋，以及一切 埃及 人的房屋，都要被蝗虫占满；你祖宗和你祖宗的祖宗在世以来，直到今日都没有见过。’” 摩西 就转身离开法老出去。
EXOD|10|7|法老的臣仆对法老说：“这家伙成为我们的罗网要到几时呢？让这些人去事奉耶和华－他们的上帝吧！ 埃及 快要灭亡了，你还不知道吗？”
EXOD|10|8|于是 摩西 和 亚伦 被召回来见法老。法老对他们说：“去，事奉耶和华－你们的上帝吧！但要去的是哪些人呢？”
EXOD|10|9|摩西 说：“我们要带着年老的和年少的同去，要带着我们的儿子和女儿，以及我们的羊群牛群一起去，因为我们要向耶和华守节。”
EXOD|10|10|法老对他们说：“愿耶和华与你们同在吧！我若让你们带着你们的孩子同去，看，灾祸就在你们面前 ！
EXOD|10|11|不可都去！你们壮年人去事奉耶和华吧，因为这是你们所求的。”于是法老把他们从自己面前赶出去。
EXOD|10|12|耶和华对 摩西 说：“你向 埃及 地伸出你的手，使蝗虫上到 埃及 地，吃地上冰雹后所剩一切的植物。”
EXOD|10|13|摩西 就向 埃及 地伸杖；整整一昼一夜，耶和华使东风刮在 埃及 地上，到了早晨，东风把蝗虫刮了来。
EXOD|10|14|蝗虫上到 埃及 全地，落在 埃及 全境，非常厉害；蝗虫这么多，是空前绝后的。
EXOD|10|15|蝗虫遮满地面，地上一片黑暗。它们吃尽了地上一切的植物和冰雹过后所剩树上的果子。 埃及 全地，无论是树木，是田间的植物，连一点绿的也没有留下。
EXOD|10|16|于是法老急忙召了 摩西 和 亚伦 来，说：“我得罪了耶和华－你们的上帝，又得罪了你们。
EXOD|10|17|现在求你，就这一次，饶恕我的罪，祈求耶和华－你们的上帝救我脱离这次的死亡。”
EXOD|10|18|摩西 就离开法老，去祈求耶和华。
EXOD|10|19|耶和华转变风向，使强劲的西风吹来，把蝗虫刮起，吹入 红海 ；在 埃及 全境连一只也没有留下。
EXOD|10|20|但耶和华任凭法老的心刚硬，不放 以色列 人走。
EXOD|10|21|耶和华对 摩西 说：“你向天伸出你的手，使黑暗笼罩 埃及 地；这黑暗甚至可以摸得到。”
EXOD|10|22|摩西 向天伸出他的手，浓密的黑暗就笼罩了 埃及 全地三天之久。
EXOD|10|23|三天内，人人彼此看不见，谁也不敢起身离开原地；但所有 以色列 人住的地方却有光。
EXOD|10|24|法老就召 摩西 来，说：“去，事奉耶和华吧！只是你们的羊群牛群要留下来。你们的孩子可以和你们同去。”
EXOD|10|25|摩西 说：“你必须把祭物和燔祭牲交在我们手中，让我们可以向耶和华我们的上帝献祭。
EXOD|10|26|我们的牲畜也要与我们同去，连一蹄也不留下，因为我们要从牲畜中挑选来事奉耶和华－我们的上帝。未到那里之前，我们还不知道要用什么来事奉耶和华。”
EXOD|10|27|但耶和华任凭法老的心刚硬，法老不肯放他们走。
EXOD|10|28|法老对 摩西 说：“离开我去吧！你要小心，不要再见我的面，因为再见我面的那日，你就必死！”
EXOD|10|29|摩西 说：“就照你说的，我也不要再见你的面了！”
EXOD|11|1|耶和华对 摩西 说：“我要再降一个灾祸给法老和 埃及 ，然后他必让你们离开这里。他放你们走的时候，一定会赶你们全都离开这里。
EXOD|11|2|你要传于百姓耳中，叫他们男的女的各向邻舍索取金器银器。”
EXOD|11|3|耶和华使 埃及 人看得起他的百姓 ，并且 摩西 在 埃及 地，在法老臣仆和百姓眼中看为伟大。
EXOD|11|4|摩西 说：“耶和华如此说：‘约到半夜，我必出去走遍 埃及 。
EXOD|11|5|凡在 埃及 地，从坐宝座的法老到推磨 的婢女所生的长子，以及一切头生的牲畜，都必死。
EXOD|11|6|埃及 全地必有大大的哀号，这将是空前绝后的。
EXOD|11|7|至于 以色列 人中，无论是人是牲畜，连狗也不敢向他们吠叫，使你们知道耶和华区别 埃及 和 以色列 。’
EXOD|11|8|你所有的这些臣仆都要下到我这里，向我下拜说：‘请你和跟从你的百姓都离开吧！’然后我才离开。”于是， 摩西 气愤愤地离开法老出去了。
EXOD|11|9|耶和华对 摩西 说：“法老必不听你们，为了要使我在 埃及 地多行奇事。”
EXOD|11|10|摩西 和 亚伦 在法老面前行了这一切奇事，但耶和华任凭法老的心刚硬，不让 以色列 人离开他的地。
EXOD|12|1|耶和华在 埃及 地对 摩西 和 亚伦 说：
EXOD|12|2|“你们要以本月为正月，为一年之首。
EXOD|12|3|你们要吩咐 以色列 全会众说：本月初十，各人要按着家庭 取羔羊，一家一只羔羊。
EXOD|12|4|若一家的人太少，吃不了一只羔羊，就要按照人数和隔壁的邻舍共取一只；你们要按每人的食量来估算羔羊。
EXOD|12|5|你们要从绵羊或山羊中取一只无残疾、一岁的公羔羊，
EXOD|12|6|要把它留到本月十四日；那日黄昏的时候， 以色列 全会众要把羔羊宰了。
EXOD|12|7|他们要取一些血，涂在他们吃羔羊的房屋两边的门框上和门楣上。
EXOD|12|8|当晚要吃羔羊的肉；要用火烤了，与无酵饼和苦菜一起吃。
EXOD|12|9|不可吃生的，或用水煮的，要把羔羊连头带腿和内脏用火烤了吃。
EXOD|12|10|一点也不可留到早晨；若有留到早晨的，要用火烧了。
EXOD|12|11|你们要这样吃羔羊：腰间束带，脚上穿鞋，手中拿杖，快快地吃。这是耶和华的逾越。
EXOD|12|12|因为那夜我要走遍 埃及 地，把 埃及 地一切头生的，无论是人是牲畜，都击杀了；我要对 埃及 所有的神明施行审判。我是耶和华。
EXOD|12|13|这血要在你们所住的房屋上作记号；我一见这血，就逾越你们。我击打 埃及 地的时候，灾殃必不临到你们身上施行毁灭。”
EXOD|12|14|“你们要记念这日，世世代代守这日为耶和华的节日，作为你们永远的定例。
EXOD|12|15|你们要吃无酵饼七日。第一日要把酵从你们各家中除去，因为从第一日到第七日，任何吃有酵之物的，必从 以色列 中剪除。
EXOD|12|16|第一日当有圣会，第七日也当有圣会。在这两日，任何工作都不可做，只能预备各人的食物，这是惟一可做的工作。
EXOD|12|17|你们要守除酵节，因为我在这一日把你们的军队从 埃及 地领出来。所以，你们要世世代代守这日，立为永远的定例。
EXOD|12|18|从正月十四日晚上，直到二十一日晚上，你们要吃无酵饼。
EXOD|12|19|在你们各家中，七日之内不可有酵，因为凡吃有酵之物的，无论是寄居的，是本地的，必从 以色列 的会中剪除。
EXOD|12|20|任何有酵的物，你们都不可吃；在你们一切的住处要吃无酵饼。”
EXOD|12|21|于是， 摩西 召了 以色列 的众长老来，对他们说：“你们要为家人取羔羊，把逾越的羔羊宰了。
EXOD|12|22|要拿一把牛膝草，蘸盆里的血，把盆里的血涂在门楣上和两边的门框上。直到早晨你们谁也不可出自己家里的门。
EXOD|12|23|因为耶和华要走遍 埃及 ，施行击杀，他看见血在门楣上和两边的门框上，耶和华就必逾越那门，不让灭命者进你们的家，施行击杀。
EXOD|12|24|你们要守这命令，作为你们和你们子孙永远的定例。
EXOD|12|25|日后，你们到了耶和华所应许赐给你们的那地，就要守这礼仪。
EXOD|12|26|你们的儿女对你们说：‘这礼仪是什么意思呢？’
EXOD|12|27|你们就说：‘这是献给耶和华逾越节的祭物。当耶和华击杀 埃及 人的时候，他逾越了 以色列 人在 埃及 的房屋，救了我们各家。’”于是百姓低头敬拜。
EXOD|12|28|以色列 人就去做；他们照耶和华吩咐 摩西 和 亚伦 的去做了。
EXOD|12|29|到了半夜，耶和华把 埃及 地所有头生的，就是从坐宝座的法老，到关在牢里的人的长子，以及一切头生的牲畜，尽都杀了。
EXOD|12|30|法老和他众臣仆，以及所有的 埃及 人，都在夜间起来了。在 埃及 有大大的哀号，因为没有一家不死人的。
EXOD|12|31|夜间，法老召了 摩西 和 亚伦 来，说：“起来！你们和 以色列 人，都离开我的百姓出去，照你们所说的，去事奉耶和华吧！
EXOD|12|32|照你们所说的，连羊群牛群也带走，也为我祝福吧！”
EXOD|12|33|埃及 人催促百姓赶快离开那地，因为 埃及 人说：“我们都快死了。”
EXOD|12|34|百姓就拿着没有发酵的生面，把揉面盆包在衣服中，扛在肩上。
EXOD|12|35|以色列 人照 摩西 的话去做，向 埃及 人索取金器、银器和衣裳。
EXOD|12|36|耶和华使 埃及 人看得起他的百姓， 埃及 人就给了他们所要的。他们就掠夺了 埃及 人。
EXOD|12|37|以色列 人从 兰塞 起程，往 疏割 去。除了小孩，步行的男人约有六十万。
EXOD|12|38|又有许多不同族群的人，以及众多的羊群牛群，和他们一同上去。
EXOD|12|39|他们用 埃及 带出来的生面烤成无酵饼。这生面是没有发酵的；因为他们被催促离开 埃及 ，不能耽延，就没有为自己预备食物。
EXOD|12|40|以色列 人住在 埃及 共四百三十年。
EXOD|12|41|正满四百三十年的那一天，耶和华的全军从 埃及 地出来了。
EXOD|12|42|这是向耶和华守的夜，他领他们出 埃及 地；这是 以色列 众人世世代代要向耶和华守的夜。
EXOD|12|43|耶和华对 摩西 和 亚伦 说：“逾越节的条例是这样：外邦人不可吃这羔羊。
EXOD|12|44|但是你们用银子买来，又受过割礼的奴仆可以吃。
EXOD|12|45|寄居的和雇工都不可吃。
EXOD|12|46|应当在一个屋子里吃，不可把肉带到屋外，骨头一根也不可折断。
EXOD|12|47|以色列 全会众都要守这礼仪。
EXOD|12|48|若有外人寄居在你那里，要向耶和华守逾越节，他所有的男子务要先受割礼，然后才可以当他是本地人，容许他守这礼仪。但未受割礼的都不可吃这羔羊。
EXOD|12|49|本地人和寄居在你们中间的外人当守同一个条例。”
EXOD|12|50|以色列 众人就去做，他们照耶和华吩咐 摩西 和 亚伦 的去做了。
EXOD|12|51|正当那日，耶和华将 以色列 人按着他们的队伍从 埃及 地领了出来。
EXOD|13|1|耶和华吩咐 摩西 说：
EXOD|13|2|“头生的要分别为圣归我； 以色列 中凡头生的，无论是人是牲畜，都是我的。”
EXOD|13|3|摩西 对百姓说：“你们要记念从 埃及 为奴之家出来的这日，因为耶和华用大能的手将你们从这地领出来。有酵之物都不可吃。
EXOD|13|4|亚笔月的这一日你们走出来了。
EXOD|13|5|将来耶和华领你进 迦南 人、 赫 人、 亚摩利 人、 希未 人、 耶布斯 人之地，就是他向你祖宗起誓应许给你的那流奶与蜜之地，那时你要在这一个月守这礼仪。
EXOD|13|6|你要吃无酵饼七日，在第七日要向耶和华守节。
EXOD|13|7|这七日之内，要吃无酵饼；在你的全境内不可见有酵之物，也不可见酵母。
EXOD|13|8|当那日，你要告诉你的儿子说：‘这样做是因为耶和华在我出 埃及 的时候为我所做的事。’
EXOD|13|9|这要在你手上作记号，在你额上 作纪念，使耶和华的教导常在你口中，因为耶和华用大能的手将你从 埃及 领出来。
EXOD|13|10|所以你每年要按着日期守这条例。”
EXOD|13|11|“当耶和华照他向你和你祖宗所起的誓将你领进 迦南 人之地，把那地赐给你的时候，
EXOD|13|12|你要将一切头生的献给耶和华；你牲畜中头生的，公的都归耶和华。
EXOD|13|13|然而，凡头生的驴，你要用羔羊赎回；若不赎它，就要打断它的颈项。你儿子中的长子都要赎出来。
EXOD|13|14|日后，你的儿子问你说：‘这是什么意思？’你就说：‘耶和华用大能的手将我们从 埃及 为奴之家领出来。
EXOD|13|15|那时法老固执，不肯放我们走，耶和华就把 埃及 地所有头生的，无论是人是牲畜，都杀了。因此，我把一切头生的公的牲畜献给耶和华为祭，却将所有头生的儿子赎出来。
EXOD|13|16|这要在你手上作记号，在你额上作经匣 ，因为耶和华用大能的手将我们从 埃及 领出来。’”
EXOD|13|17|法老放百姓走的时候， 非利士 人之地的路虽近，上帝却不领他们从那里走，因为上帝说：“恐怕百姓遇见战争就后悔，转回 埃及 去。”
EXOD|13|18|上帝领百姓绕道而行，走旷野的路到 红海 。 以色列 人出 埃及 地，都带着兵器上去 。
EXOD|13|19|摩西 把 约瑟 的骸骨一起带走；因为 约瑟 曾叫 以色列 人郑重地起誓，对他们说：“上帝必定眷顾你们，你们要把我的骸骨从这里一起带上去。”
EXOD|13|20|他们从 疏割 起程，在旷野边上的 以倘 安营。
EXOD|13|21|耶和华走在他们前面，日间用云柱引领他们的路，夜间用火柱照亮他们，使他们日夜都可以行走。
EXOD|13|22|日间的云柱，夜间的火柱，总不离开百姓的面前。
EXOD|14|1|耶和华吩咐 摩西 说：
EXOD|14|2|“你吩咐 以色列 人转回，要在 比．哈希录 前面， 密夺 和海的中间， 巴力．洗分 的前面安营。你们要在对面，靠近海边安营。
EXOD|14|3|以色列 人这样做，法老必说：‘他们在此地迷了路，旷野把他们困住了。’
EXOD|14|4|我要任凭法老的心刚硬，他要追赶他们。我必在法老和他全军身上得荣耀， 埃及 人就知道我是耶和华。”于是 以色列 人照样做了。
EXOD|14|5|有人报告 埃及 王说：“百姓逃跑了！”法老和他的臣仆对百姓改变了心意，说：“我们放 以色列 人走，不再服事我们，我们怎么会做这种事呢？”
EXOD|14|6|法老就预备战车，带领他的军兵同去，
EXOD|14|7|他带了六百辆特选的战车和 埃及 所有的战车，每辆都有军官。
EXOD|14|8|耶和华任凭 埃及 王法老的心刚硬，他就追赶 以色列 人； 以色列 人却抬起头 来出去了。
EXOD|14|9|埃及 人追赶他们，法老一切的马匹、战车、战车长，与军兵就在海边上，靠近 比．哈希录 ，在 巴力．洗分 的前面，在他们安营的地方追上了。
EXOD|14|10|法老逼近的时候， 以色列 人举目，看哪， 埃及 人追来了，就非常惧怕， 以色列 人向耶和华哀求。
EXOD|14|11|他们对 摩西 说：“难道 埃及 没有坟地，你要把我们带来死在旷野吗？你为什么这样待我们，将我们从 埃及 领出来呢？
EXOD|14|12|我们在 埃及 岂没有对你说过，不要搅扰我们，让我们服事 埃及 人吗？因为服事 埃及 人总比死在旷野好。”
EXOD|14|13|摩西 对百姓说：“不要怕，要站稳，看耶和华今天向你们所要施行的拯救，因为你们今天所看见的 埃及 人必永远不再看见了。
EXOD|14|14|耶和华必为你们争战，你们要安静！”
EXOD|14|15|耶和华对 摩西 说：“你为什么向我哀求呢？你吩咐 以色列 人往前走。
EXOD|14|16|你举手向海伸杖，把水分开。 以色列 人要下到海中，走在干地上。
EXOD|14|17|看哪，我要任凭 埃及 人的心刚硬，他们就跟着下去。我要在法老和他的全军、战车、战车长身上得荣耀。
EXOD|14|18|我在法老和他的战车、战车长身上得荣耀的时候， 埃及 人就知道我是耶和华。”
EXOD|14|19|在 以色列 营前行走的上帝的使者移动，走到他们后面；云也从他们的前面移动，站在他们后面。
EXOD|14|20|它来到 埃及 营和 以色列 营的中间：一边有云和黑暗，另一边它照亮夜晚，整夜彼此不得接近。
EXOD|14|21|摩西 向海伸手，耶和华就用强劲的东风，使海水在一夜间退去，海就成了干地；水分开了。
EXOD|14|22|以色列 人下到海中，走在干地上，水在他们左右成了墙壁。
EXOD|14|23|埃及 人追赶他们，法老一切的马匹、战车和战车长都跟着下到海中。
EXOD|14|24|破晓时分，耶和华从云柱、火柱中了望 埃及 的军兵，使 埃及 的军兵混乱。
EXOD|14|25|他使他们的车轮脱落 ，难以前行， 埃及 人说：“我们从 以色列 人面前逃跑吧！因耶和华为他们作战，攻击 埃及 了。”
EXOD|14|26|耶和华对 摩西 说：“你要向海伸手，使水回流到 埃及 人，他们的战车和战车长身上。”
EXOD|14|27|摩西 就向海伸手，到了天亮的时候，海恢复原状。 埃及 人逃避水的时候，耶和华把他们推入海中。
EXOD|14|28|海水回流，淹没了战车和战车长，以及那些跟着 以色列 人下到海中的法老全军，连一个也没有剩下。
EXOD|14|29|以色列 人却在海中走干地，水在他们的左右成了墙壁。
EXOD|14|30|那一日，耶和华拯救 以色列 脱离 埃及 人的手。 以色列 人看见 埃及 人死在海边。
EXOD|14|31|以色列 人看见耶和华向 埃及 人所施展的大能，百姓就敬畏耶和华，并且信服耶和华和他的仆人 摩西 。
EXOD|15|1|那时， 摩西 和 以色列 人向耶和华唱这歌，说： “我要向耶和华歌唱，因他大大得胜， 将马和骑马的投在海中。
EXOD|15|2|耶和华是我的力量，是我的诗歌， 他也成了我的拯救。 这是我的上帝，我要赞美他； 我父亲的上帝，我要尊崇他。
EXOD|15|3|耶和华是战士； 耶和华是他的名。
EXOD|15|4|“法老的战车、军兵，他已抛在海中； 法老精选的军官都沉于 红海 。
EXOD|15|5|深水淹没他们； 他们好像石头坠到深处。
EXOD|15|6|耶和华啊，你的右手施展能力，大显荣耀； 耶和华啊，你的右手摔碎仇敌。
EXOD|15|7|你大发威严，摧毁了你的敌人； 你发出烈怒，吞灭他们如同碎秸。
EXOD|15|8|因你鼻中的气，水就聚成堆， 大水竖立如垒， 海的中心深水凝结。
EXOD|15|9|仇敌说：‘我要追赶，我要追上， 我要分掳物，在他们身上满足我的心愿， 我要拔刀，亲手毁灭他们。’
EXOD|15|10|你用风一吹，海水就淹没他们； 他们像铅沉在大水之中。
EXOD|15|11|“耶和华啊，众神明中，谁能像你？ 谁能像你，至圣至荣， 可颂可畏，施行奇事！
EXOD|15|12|你伸出右手， 地就吞灭他们。
EXOD|15|13|“你以慈爱引领你所救赎的百姓； 你以能力引导他们到你的圣所。
EXOD|15|14|万民听见就战抖； 疼痛抓住 非利士 的居民。
EXOD|15|15|那时， 以东 的族长惊惶， 摩押 的英雄被战兢抓住， 迦南 所有的居民都融化。
EXOD|15|16|惊骇恐惧临到他们； 耶和华啊，因你膀臂的大能， 他们如石头寂静不动， 等候你百姓过去， 等候你所赎的百姓过去。
EXOD|15|17|你要将他们领进去，栽在你产业的山上， 耶和华啊，就是你为自己所造的住处， 主啊，就是你手所建立的圣所。
EXOD|15|18|耶和华必作王，直到永永远远！”
EXOD|15|19|法老的马匹、战车和战车长下到海中，耶和华使海水回流到他们身上； 以色列 人却走在海中的干地上。
EXOD|15|20|那时， 米利暗 女先知， 亚伦 的姊姊，手里拿着铃鼓；众妇女也跟她出去打鼓跳舞。
EXOD|15|21|米利暗 回应他们： “你们要歌颂耶和华，因他大大得胜， 将马和骑马的投在海中。”
EXOD|15|22|摩西 领 以色列 人从 红海 起程，到了 书珥 的旷野，在旷野走了三天，找不到水。
EXOD|15|23|到了 玛拉 ，他们不能喝 玛拉 的水，因为水是苦的；所以那地名叫 玛拉 。
EXOD|15|24|百姓就向 摩西 发怨言，说：“我们喝什么呢？”
EXOD|15|25|摩西 呼求耶和华，耶和华指示他一棵树 。他把树丢在水里，水就变甜了。 耶和华在那里为他们定了律例、典章，在那里考验他们。
EXOD|15|26|他说：“你若留心听从耶和华－你上帝的话，行我眼中看为正的事，侧耳听我的诫令，遵守我一切的律例，我就不将所加于 埃及 人的疾病加在你身上，因为我是医治你的耶和华。”
EXOD|15|27|他们到了 以琳 ，在那里有十二股水泉，七十棵棕树；他们就在那里的水边安营。
EXOD|16|1|以色列 全会众从 以琳 起程，在出 埃及 之后第二个月十五日到了 以琳 和 西奈 中间， 汛 的旷野。
EXOD|16|2|以色列 全会众在旷野向 摩西 和 亚伦 发怨言。
EXOD|16|3|以色列 人对他们说：“我们宁愿在 埃及 地死在耶和华手中！那时我们坐在肉锅旁，吃饼得饱。你们却将我们领出来，到这旷野，要叫这全会众都饿死啊！”
EXOD|16|4|耶和华对 摩西 说：“看哪，我要从天降食物给你们。百姓可以出去，每天收集当天的分量。这样，我就可以考验他们是否遵行我的指示。
EXOD|16|5|到第六天，他们预备食物，所收集的分量要比每天所收的多一倍。”
EXOD|16|6|摩西 和 亚伦 对 以色列 众人说：“到了晚上，你们就知道是耶和华将你们从 埃及 地领出来的。
EXOD|16|7|早晨，你们要看见耶和华的荣耀，因为耶和华听见你们向他所发的怨言了。我们算什么，你们竟然向我们发怨言呢？”
EXOD|16|8|摩西 又说：“耶和华晚上必给你们肉吃，早晨必给你们食物得饱，因为耶和华已经听见你们向他所发的怨言。我们算什么呢？你们的怨言不是向我们发的，而是向耶和华发的。”
EXOD|16|9|摩西 对 亚伦 说：“你对 以色列 全会众说：‘你们来到耶和华面前，因为他已经听见你们的怨言了。’”
EXOD|16|10|亚伦 正对 以色列 全会众说话的时候，他们转向旷野，看哪，耶和华的荣光在云中显现。
EXOD|16|11|耶和华吩咐 摩西 说：
EXOD|16|12|“我已经听见 以色列 人的怨言了。你要对他们说：‘到黄昏的时候 ，你们要吃肉，早晨也必有食物得饱。你们就知道我是耶和华－你们的上帝。’”
EXOD|16|13|到了晚上，有鹌鹑上来，遮满营地；早晨，营地周围有一层露水。
EXOD|16|14|那一层露水蒸发之后，看哪，旷野的表面出现了小圆物，好像地上的薄霜一样。
EXOD|16|15|以色列 人看见了，不知道是什么，就彼此说：“这是什么？ ” 摩西 对他们说：“这是耶和华给你们吃的食物。
EXOD|16|16|耶和华所吩咐的是这样：‘你们每个人要按自己的食量收集，各人要为帐棚里的人收集，按照人口数每个人一俄梅珥。’”
EXOD|16|17|以色列 人就照样去做；有的收多，有的收少。
EXOD|16|18|用俄梅珥量一量，多收的没有余，少收的也没有缺；各人都按着自己的食量收集。
EXOD|16|19|摩西 对他们说：“任何人都不可以把所收的留到早晨。”
EXOD|16|20|然而他们不听从 摩西 ，当中有人把食物留到早晨，食物就生虫发臭了。 摩西 就向他们发怒。
EXOD|16|21|他们每日早晨按着各人的食量收集；太阳一发热，食物就融化了。
EXOD|16|22|到第六天，他们收集了双倍的食物，每个人二俄梅珥。会众的官长来告诉 摩西 ，
EXOD|16|23|摩西 对他们说：“耶和华吩咐：‘明天是安息日，是向耶和华守的圣安息日。你们要烤的就烤，要煮的就煮，所剩下的都留到早晨。’”
EXOD|16|24|他们就照 摩西 的吩咐把剩下的留到早晨，这些食物既不发臭，里头也没有生虫。
EXOD|16|25|摩西 说：“你们今天就吃这些吧！因为今天是向耶和华守的安息日，你们在野外必找不着食物了。
EXOD|16|26|六天可以收集，第七天是安息日，这一天什么也没有了。”
EXOD|16|27|第七天，百姓中有人出去收，什么也找不着。
EXOD|16|28|耶和华对 摩西 说：“你们不肯遵守我的诫令和教导，要到几时呢？
EXOD|16|29|你们看，耶和华既然将安息日赐给你们，所以第六天他就赐给你们两天的食物，第七天各人都要留在自己的地方，不许任何人从这里出去。”
EXOD|16|30|于是百姓在第七天安息了。
EXOD|16|31|以色列 家给这食物取名叫吗哪，它的样子像芫荽子，颜色是白的，吃起来像和蜜的薄饼。
EXOD|16|32|摩西 说：“耶和华所吩咐的是这样：‘要装满一俄梅珥的吗哪留给你们的后代，使他们可以看见我领你们出 埃及 地的时候，在旷野所给你们吃的食物。’”
EXOD|16|33|摩西 对 亚伦 说：“你拿一个罐子，装满一俄梅珥的吗哪，存在耶和华面前，留给你们的后代。”
EXOD|16|34|耶和华怎么吩咐 摩西 ， 亚伦 就照样做，把吗哪存留作见证 。
EXOD|16|35|以色列 人吃吗哪共四十年，直到进入有人居住的地方；他们吃吗哪，直到 迦南 地的边境。
EXOD|16|36|一俄梅珥是一伊法的十分之一。
EXOD|17|1|以色列 全会众遵照耶和华的吩咐，从 汛 的旷野一段一段地往前行。他们在 利非订 安营，但百姓没有水喝。
EXOD|17|2|百姓就与 摩西 争闹，说：“给我们水喝吧！” 摩西 对他们说：“你们为什么与我争闹呢？你们为什么试探耶和华呢？”
EXOD|17|3|百姓在那里口渴要喝水，就向 摩西 发怨言，说：“你为什么把我们从 埃及 领出来，使我们和我们的儿女，以及牲畜都渴死呢？”
EXOD|17|4|摩西 就呼求耶和华说：“我要怎样对待这百姓呢？他们差一点就要拿石头打死我了。”
EXOD|17|5|耶和华对 摩西 说：“你带着 以色列 的几个长老，走在百姓前面，手里拿着你先前击打 尼罗河 的杖，去吧！
EXOD|17|6|看哪，我要在 何烈 的磐石那里，站在你面前。你要击打磐石，水就会从磐石流出来，给百姓喝。” 摩西 就在 以色列 的长老眼前这样做了。
EXOD|17|7|他给那地方起名叫 玛撒 ，又叫 米利巴 ，因为 以色列 人在那里争闹，并且试探耶和华，说：“耶和华是否在我们中间呢？”
EXOD|17|8|那时， 亚玛力 来到 利非订 ，和 以色列 争战。
EXOD|17|9|摩西 对 约书亚 说：“你为我们选出人来，出去和 亚玛力 争战。明天我要站在山顶上，手里拿着上帝的杖。”
EXOD|17|10|于是， 约书亚 照着 摩西 对他所说的话去做，和 亚玛力 争战。 摩西 、 亚伦 和 户珥 都上了山顶。
EXOD|17|11|摩西 何时举手， 以色列 就得胜；何时垂手， 亚玛力 就得胜。
EXOD|17|12|但 摩西 的双手沉重，他们就搬一块石头来放在他下面，他就坐在上面。 亚伦 与 户珥 扶着他的手，一个在这边，一个在那边，他的手就稳住，直到日落。
EXOD|17|13|约书亚 用刀打败了 亚玛力 和他的百姓。
EXOD|17|14|耶和华对 摩西 说：“你要把这事记录在书上作纪念，又念给 约书亚 听：我要把 亚玛力 的名字从天下全然涂去。”
EXOD|17|15|摩西 筑了一座坛，起名叫“耶和华尼西 ”。
EXOD|17|16|他说：“我指着耶和华的宝座发誓 ，耶和华必世世代代和 亚玛力 争战。”
EXOD|18|1|摩西 的岳父， 米甸 祭司 叶特罗 ，听见上帝为 摩西 和为他百姓 以色列 所行的一切事，就是耶和华将 以色列 从 埃及 领了出来。
EXOD|18|2|摩西 的岳父 叶特罗 带着 西坡拉 ，就是 摩西 先前送回家的妻子，
EXOD|18|3|又带着她的两个儿子：一个名叫 革舜 ，因为 摩西 说：“我在外地作了寄居者”；
EXOD|18|4|另一个名叫 以利以谢 ，因为他说：“我父亲的上帝帮助我，救我脱离法老的刀。”
EXOD|18|5|摩西 的岳父 叶特罗 带着 摩西 的妻子和两个儿子来到上帝的山，就是 摩西 在旷野安营的地方。
EXOD|18|6|他对 摩西 说：“我是 你岳父 叶特罗 ，带着你的妻子和两个儿子来到你这里。”
EXOD|18|7|摩西 迎接他的岳父，向他下拜，亲他，彼此问安，然后进入帐棚。
EXOD|18|8|摩西 将耶和华为 以色列 的缘故向法老和 埃及 人所行的一切事，他们在路上遭遇的一切艰难，以及耶和华怎样搭救他们，都述说给他的岳父听。
EXOD|18|9|叶特罗 因耶和华待 以色列 的一切恩惠，就是拯救他们脱离 埃及 人的手，就非常喜乐。
EXOD|18|10|叶特罗 说：“耶和华是应当称颂的，他救了你们脱离 埃及 人和法老的手，将这百姓从 埃及 人的手里救出来 。
EXOD|18|11|现在，从 埃及 人狂傲地对待 以色列 人这件事上，我知道耶和华比万神更大。”
EXOD|18|12|摩西 的岳父 叶特罗 把燔祭和祭物献给上帝。 亚伦 和 以色列 的众长老都来了，与 摩西 的岳父在上帝面前吃饭。
EXOD|18|13|第二天， 摩西 坐着审判百姓，百姓从早到晚站在 摩西 的旁边。
EXOD|18|14|摩西 的岳父看见他为百姓所做的一切事，就说：“你为百姓所做的，这是什么事呢？你为什么独自一人坐着，而众百姓从早到晚都站在你旁边呢？”
EXOD|18|15|摩西 对岳父说：“这是因为百姓到我这里来求问上帝。
EXOD|18|16|他们有事的时候，就到我这里来，我就在双方之间作判决；我又叫他们知道上帝的律例和法度。”
EXOD|18|17|摩西 的岳父对他说：“你这样做不好。
EXOD|18|18|你和这些与你在一起的百姓都必疲惫，因为这事太重，你独自一人做不了。
EXOD|18|19|现在，听我的话，我给你出个主意，愿上帝与你同在。你要代替百姓到上帝面前，将事件带到上帝那里，
EXOD|18|20|又要用律例和法度警戒他们，指示他们当行的道，当做的事。
EXOD|18|21|你也要从百姓中选出有才能的人，敬畏上帝、诚实可靠、恨恶不义之财的人，派他们作千夫长、百夫长、五十夫长、十夫长来管理百姓。
EXOD|18|22|他们要随时审判百姓；重大的事要送到你这里，小事就由他们自行判决。这样，你就可以轻省一些，他们可以与你分担。
EXOD|18|23|你若这样做，上帝也这样吩咐你，你就能承受得住，众百姓也可以和睦地回到自己的地方。”
EXOD|18|24|摩西 听了他岳父的话，照着他所说的一切去做。
EXOD|18|25|摩西 从 以色列 人中选出有才能的人，立他们为百姓的领袖，作千夫长、百夫长、五十夫长、十夫长。
EXOD|18|26|他们随时审判百姓：难断的事就送到 摩西 那里，各样小事就由他们自行判决。
EXOD|18|27|于是， 摩西 给他的岳父送行，他就回到本地去了。
EXOD|19|1|以色列 人出 埃及 地以后，第三个月的初一，就在那一天他们来到了 西奈 的旷野。
EXOD|19|2|他们从 利非订 起程，来到 西奈 的旷野，在那里的山下安营。
EXOD|19|3|摩西 到上帝那里，耶和华从山上呼唤他说：“你要这样告诉 雅各 家，对 以色列 人说：
EXOD|19|4|‘我向 埃及 人所行的事，你们都看见了， 我如鹰将你们背在翅膀上，带你们来归我。
EXOD|19|5|如今你们若真的听从我的话，遵守我的约，就要在万民中作属我的子民 ，因为全地都是我的。
EXOD|19|6|你们要归我作祭司的国度，为神圣的国民。’这些话你要告诉 以色列 人。”
EXOD|19|7|摩西 去召了百姓中的长老来，将耶和华吩咐他的话当面告诉他们。
EXOD|19|8|百姓都同声回答：“凡耶和华所说的，我们一定遵行。” 摩西 就将百姓的话回覆耶和华。
EXOD|19|9|耶和华对 摩西 说：“看哪，我要在密云中临到你那里，叫百姓在我与你说话的时候可以听见，就可以永远相信你了。”于是， 摩西 将百姓的话禀告耶和华。
EXOD|19|10|耶和华对 摩西 说：“你往百姓那里去，使他们今天明天分别为圣，又叫他们洗衣服。
EXOD|19|11|第三天要预备好，因为第三天耶和华要在众百姓眼前降临在 西奈山 。
EXOD|19|12|你要在山的周围给百姓划定界限，说：‘你们当谨慎，不可上山去，也不可摸山的边界。凡摸这山的，必被处死。
EXOD|19|13|不可用手碰他，要用石头打死，或射死；无论是人是牲畜，都不可活。’到角声拉长的时候，他们才可到山脚来。”
EXOD|19|14|摩西 下山到百姓那里去，使他们分别为圣，他们就洗衣服。
EXOD|19|15|他对百姓说：“第三天要预备好；不可亲近女人。”
EXOD|19|16|到了第三天早晨，山上有雷轰、闪电和密云，并且角声非常响亮，营中的百姓尽都战抖。
EXOD|19|17|摩西 率领百姓出营迎见上帝，都站在山下。
EXOD|19|18|西奈山 全山冒烟，因为耶和华在火中降临山上。山的烟雾上腾，仿佛烧窑，整座山剧烈震动。
EXOD|19|19|角声越来越响， 摩西 说话，上帝以声音回答他。
EXOD|19|20|耶和华降临在 西奈山 顶上，耶和华召 摩西 上山顶， 摩西 就上去了。
EXOD|19|21|耶和华对 摩西 说：“你下去警告百姓，免得他们闯过来看耶和华，就会有许多人死亡。
EXOD|19|22|那些亲近耶和华的祭司也要把自己分别为圣，免得耶和华忽然出来击杀他们。”
EXOD|19|23|摩西 对耶和华说：“百姓不能上 西奈山 ，因为你已经警告我们说：‘要在山的周围划定界限，使山成圣。’”
EXOD|19|24|耶和华对他说：“下去吧，你要和 亚伦 一起上来；只是祭司和百姓不可闯上来到耶和华这里，免得耶和华忽然出来击杀他们。”
EXOD|19|25|于是， 摩西 下到百姓那里告诉他们。
EXOD|20|1|上帝吩咐这一切的话，说：
EXOD|20|2|“我是耶和华－你的上帝，曾将你从 埃及 地为奴之家领出来。
EXOD|20|3|“除了我以外，你不可有别的神。
EXOD|20|4|“不可为自己雕刻偶像，也不可做什么形像，仿佛上天、下地和地底下水中的百物。
EXOD|20|5|不可跪拜那些像，也不可事奉它们，因为我耶和华─你的上帝是忌邪 的上帝。恨我的，我必惩罚他们的罪，自父及子，直到三、四代；
EXOD|20|6|爱我，守我诫命的，我必向他们施慈爱，直到千代。
EXOD|20|7|“不可妄称耶和华－你上帝的名，因为妄称耶和华名的，耶和华必不以他为无罪。
EXOD|20|8|“当记念安息日，守为圣日。
EXOD|20|9|六日要劳碌做你一切的工，
EXOD|20|10|但第七日是向耶和华─你的上帝当守的安息日。这一日你和你的儿女、奴仆、婢女、牲畜，以及你城里寄居的客旅，都不可做任何的工。
EXOD|20|11|因为六日之内，耶和华造天、地、海和其中的万物，第七日就安息了；所以耶和华赐福与安息日，定为圣日。
EXOD|20|12|“当孝敬父母，使你的日子在耶和华－你上帝所赐你的地上得以长久。
EXOD|20|13|“不可杀人。
EXOD|20|14|“不可奸淫。
EXOD|20|15|“不可偷盗。
EXOD|20|16|“不可做假见证陷害你的邻舍。
EXOD|20|17|“不可贪恋你邻舍的房屋；不可贪恋你邻舍的妻子、奴仆、婢女、牛驴，以及他一切所有的。”
EXOD|20|18|众百姓见雷轰、闪电、角声、山上冒烟，百姓看见 就都战抖，远远站着。
EXOD|20|19|他们对 摩西 说：“请你向我们说话，我们必听；不要让上帝向我们说话，免得我们死亡。”
EXOD|20|20|摩西 对百姓说：“不要害怕；因为上帝降临是要考验你们，要你们敬畏他，不致犯罪。”
EXOD|20|21|于是百姓远远站着，但 摩西 却挨近上帝所在的幽暗中。
EXOD|20|22|耶和华对 摩西 说：“你要向 以色列 人这样说：‘你们亲自看见我从天上向你们说话了。
EXOD|20|23|你们不可为我制造偶像，不可为自己造任何金银的神像。
EXOD|20|24|你要为我筑一座土坛，在上面献牛羊为燔祭和平安祭。凡在我叫你记念我名的地方，我必到那里赐福给你。
EXOD|20|25|你若为我筑一座石坛，不可用凿过的石头，因为你在石头上动了工具，就使坛污秽了。
EXOD|20|26|你不可用台阶上我的坛，免得露出你的下体来。’”
EXOD|21|1|“你在百姓面前所要立的典章是这样：
EXOD|21|2|“你若买 希伯来 人作奴仆，他服事你六年，第七年他可以自由，白白地离去。
EXOD|21|3|他若单身来就可以单身去；他若是有妻子的，他的妻子可以同他离去。
EXOD|21|4|若他主人给他娶了妻，妻子为他生了儿子或女儿，妻子和儿女要归主人，他要独自离去。
EXOD|21|5|倘若奴仆声明：‘我爱我的主人和我的妻子儿女，不愿意自由离去。’
EXOD|21|6|他的主人就要带他到审判官 前，再带他到门或门框那里，用锥子穿他的耳朵，他就要永远服事主人。
EXOD|21|7|“人若卖女儿作婢女，婢女不可像男的奴仆那样离去。
EXOD|21|8|主人若选定她归自己，后来看不顺眼，就要允许她赎身；主人既然对她失信，就没有权柄把她卖给外邦人。
EXOD|21|9|主人若选定她给自己的儿子，就当照女儿的规矩对待她。
EXOD|21|10|若另娶一个，她的饮食、衣服和房事不可减少。
EXOD|21|11|若不向她行这三样，她就可以白白离去，不必付赎金。”
EXOD|21|12|“打人致死的，必被处死。
EXOD|21|13|他若不是出于预谋 ，而是上帝交在他手中，我就设立一个地方，让他可以逃到那里。
EXOD|21|14|人若蓄意用诡计杀了他的邻舍，就是逃到我的坛那里，也当把他捉去处死。
EXOD|21|15|“打父母的，必被处死。
EXOD|21|16|“诱拐人口的，无论是把人卖了，或是扣留在他手中，必被处死。
EXOD|21|17|“咒骂父母的，必被处死。
EXOD|21|18|“人若彼此争吵，一个用石头或拳头打另一个，被打的人没有死去，却要躺卧在床，
EXOD|21|19|若他还能起来扶杖行走，那打他的可免处刑，却要赔偿他不能工作的损失，并要把他完全医好。
EXOD|21|20|“人若用棍子打奴仆或婢女，当场死在他的手下，他必受报应。
EXOD|21|21|若能撑过一两天，主人就不必受惩罚，因为那是他的财产。
EXOD|21|22|“人若彼此打斗，伤害有孕的妇人，以致胎儿掉了出来，随后却无别的伤害，那伤害她的人，总要按妇人的丈夫所提出的，照审判官所裁定的赔偿。
EXOD|21|23|若有别的伤害，就要以命抵命，
EXOD|21|24|以眼还眼，以牙还牙，以手还手，以脚还脚，
EXOD|21|25|以灼伤还灼伤，以损伤还损伤，以鞭打还鞭打。
EXOD|21|26|“人若打奴仆或婢女的眼睛，毁了一只，就要因他的眼让他自由离去。
EXOD|21|27|若打掉了奴仆或婢女的一颗牙，就要因他的牙让他自由离去。”
EXOD|21|28|“牛若抵死男人或女人，总要用石头打死那牛，却不可吃它的肉；牛的主人可免处刑。
EXOD|21|29|倘若那牛向来是抵人的，牛的主人虽然受过警告，仍不把它拴好，以致把男人或女人抵死，牛要用石头打死，主人也要被处死。
EXOD|21|30|若罚他付赎命的赔款，他就要照所罚的数目赎他的命。
EXOD|21|31|牛若抵了男孩或女孩，也要照这条例处理。
EXOD|21|32|牛若抵了奴仆或婢女，就要把三十舍客勒银子给他的主人，牛要用石头打死。
EXOD|21|33|“人若敞开井口，或挖井不盖住它，有牛或驴掉进井里，
EXOD|21|34|井的主人要拿钱赔偿牲畜的主人，死牲畜要归自己。
EXOD|21|35|“人的牛若抵死邻舍的牛，他们就要卖了那活牛，平分价钱；也要平分死牛。
EXOD|21|36|若这牛向来是以好抵人出名的，主人竟不把牛拴好，他必要以牛赔牛，死牛却归自己。”
EXOD|22|1|“人若偷牛或羊，无论是宰了或卖了，他就要以五牛赔一牛， 四羊赔一羊。
EXOD|22|2|贼挖洞，若被发现而被打死，打的人没有流血的罪。
EXOD|22|3|若太阳已经出来，打的人就有流血的罪。贼总要赔偿，若他一无所有，就要被卖来还他所偷的东西。
EXOD|22|4|若发现他所偷的，无论是牛、驴，或羊，在他手中还活着，他就要加倍赔偿。
EXOD|22|5|“人若在田间或葡萄园里牧放牲畜，任凭牲畜上别人田里去吃 ，他就要拿自己田间和葡萄园里上好的赔偿。
EXOD|22|6|“若火冒出，延烧到荆棘，以致将堆积的禾捆，直立的庄稼，或田地，都烧尽了，那点火的必要赔偿。
EXOD|22|7|“人若将银钱或物件托邻舍保管，东西从这人的家中被偷去，若找到了贼，贼要加倍赔偿；
EXOD|22|8|若找不到贼，这家的主人就要到审判官 那里，声明 自己没有伸手拿邻舍的物件。
EXOD|22|9|“关于任何侵害的案件，无论是为牛、驴、羊、衣服，或任何失物，有一人说：‘这是我的’，双方就要将案件带到审判官面前，审判官定谁有罪，谁就要加倍赔偿给他的邻舍。
EXOD|22|10|“人将驴、牛、羊，或别的牲畜托邻舍看管，若牲畜死亡，受了伤，或被抢走，无人看见，
EXOD|22|11|双方要在耶和华前起誓，受托人要表明自己没有伸手拿邻舍的东西，原主要接受誓言，受托人不必赔偿。
EXOD|22|12|牲畜若从受托人那里被偷去，他就要赔偿原主；
EXOD|22|13|若被野兽撕碎，受托人要带回来作证据，被撕碎的就不必赔偿。
EXOD|22|14|“人若向邻舍借牲畜 ，所借的或伤或死，原主没有在场，借的人总要赔偿。
EXOD|22|15|若原主在场，借的人不必赔偿；若是租用的，只要付租金 。”
EXOD|22|16|“人若引诱没有订婚的处女，与她同寝，他就必须交出聘礼，娶她为妻。
EXOD|22|17|若女子的父亲坚决不将女子给他，他就要按着处女的聘礼交出钱来。
EXOD|22|18|“行邪术的女人，不可让她存活。
EXOD|22|19|“凡与兽交合的，必被处死。
EXOD|22|20|“向别神献祭，不单单献给耶和华的，那人必要灭绝。
EXOD|22|21|“不可亏待寄居的，也不可欺压他，因为你们在 埃及 地也作过寄居的。
EXOD|22|22|不可苛待寡妇和孤儿；
EXOD|22|23|若你确实苛待他，他向我苦苦哀求，我一定会听他的呼求，
EXOD|22|24|并要发烈怒，用刀杀你们，使你们的妻子成为寡妇，儿女成为孤儿。
EXOD|22|25|“我的子民中有困苦人在你那里，你若借钱给他，不可如放债的向他取利息。
EXOD|22|26|你果真拿了邻舍的外衣作抵押，也要在日落前还给他；
EXOD|22|27|因为他只有这一件用来作被子，是他蔽体的衣服。他还可以拿什么睡觉呢？当他哀求我，我就应允，因为我是有恩惠的。
EXOD|22|28|“不可毁谤上帝；也不可诅咒你百姓的领袖。
EXOD|22|29|“不可迟延献你的庄稼、酒和油 。 “要将你头生的儿子归给我。
EXOD|22|30|你的牛羊也要照样做：七天当跟着它母亲，第八天你要把它归给我。
EXOD|22|31|“你们要分别为圣归给我。因此，田间被野兽撕裂的肉，你们不可吃，要把它丢给狗。”
EXOD|23|1|“不可散布谣言；不可与恶人连手作恶意的见证。
EXOD|23|2|不可附和群众作恶；不可在诉讼中附和群众歪曲公正，作歪曲的见证；
EXOD|23|3|也不可在诉讼中偏袒贫寒人。
EXOD|23|4|“若遇见你仇敌的牛或驴迷了路，务必牵回来交给他。
EXOD|23|5|若看见恨你的人的驴被压在重驮之下，不可走开，务要和他一同卸下驴的重驮。
EXOD|23|6|“不可在贫穷人的诉讼中屈枉正直。
EXOD|23|7|当远离诬告的事。不可杀害无辜和义人，因我必不以恶人为义。
EXOD|23|8|不可接受贿赂，因为贿赂能使明眼人变瞎，又能曲解义人的证词。
EXOD|23|9|“不可欺压寄居的，因为你们在 埃及 地作过寄居的，知道寄居者的心情。”
EXOD|23|10|“六年你要耕种田地，收集地的出产。
EXOD|23|11|只是第七年你要让地歇息，不耕不种，使你百姓中的贫穷人有吃的；他们吃剩的，野兽可以吃。你的葡萄园和橄榄园也要照样办理。
EXOD|23|12|“六日你要做工，第七日要安息，使牛、驴可以歇息，也让你使女的儿子和寄居的可以恢复精力。
EXOD|23|13|“凡我对你们说的话，你们都要谨守。别神的名，你不可提，也不可用口说给人听。”
EXOD|23|14|“一年三次，你要向我守节。
EXOD|23|15|你要守除酵节，照我所吩咐你的，在亚笔月内所定的日期吃无酵饼七天，因为你是在这月离开了 埃及 。谁也不可空手来朝见我。
EXOD|23|16|你要守收割节，收田间所种、劳碌所得初熟之物。你年底收藏田间劳碌所得时，要守收藏节。
EXOD|23|17|所有的男丁都要一年三次朝见主耶和华。
EXOD|23|18|“不可将我祭牲的血和有酵之物一同献上，也不可将我节期中祭牲的脂肪留到早晨。
EXOD|23|19|“要把地里最好的初熟之物带到耶和华－你上帝的殿中。 “不可用母山羊的奶来煮它的小山羊。”
EXOD|23|20|“看哪，我要差遣使者在你前面，在路上保护你，领你到我所预备的地方。
EXOD|23|21|你们要在他面前谨慎，听从他的话。不可抗拒 他，否则他必不赦免你们的过犯，因为我的名在他身上。
EXOD|23|22|“你若真的听从他的话，照我一切所说的去做，我就以你的仇敌为仇敌，以你的敌人为敌人。
EXOD|23|23|“我的使者要走在你前面，领你到 亚摩利 人、 赫 人、 比利洗 人、 迦南 人、 希未 人、 耶布斯 人那里，我必将他们除灭。
EXOD|23|24|你不可跪拜事奉他们的神明，也不可随从他们的习俗，却要彻底废除，完全打碎他们的柱像。
EXOD|23|25|你们要事奉耶和华－你们的上帝，他必赐福给你的粮食和水，也必从你中间除去疾病。
EXOD|23|26|你境内必没有流产的、不生育的。我要使你享满你年日的数目。
EXOD|23|27|凡你所到的地方，我要使那里的众百姓在你面前惊慌失措，又要使你所有的仇敌转身逃跑。
EXOD|23|28|我要派瘟疫 在你的前面，把 希未 人、 迦南 人、 赫 人从你面前赶出去。
EXOD|23|29|我不在一年之内把他们从你面前赶出去，恐怕地会荒废，野地的走兽增多危害你。
EXOD|23|30|我要逐渐把他们从你面前赶出去，直到你的人数增多，承受那地为业。
EXOD|23|31|我要定你的疆界，从 红海 直到 非利士海 ，从旷野直到 大河 。我要把那地的居民交在你手中，你要把他们从你面前赶出去。
EXOD|23|32|不可跟他们和他们的神明立约。
EXOD|23|33|他们不可住在你的地上，免得他们使你得罪我。你若事奉他们的神明，必成为你的圈套。”
EXOD|24|1|耶和华对 摩西 说：“你和 亚伦 、 拿答 、 亚比户 ，以及 以色列 长老中的七十人，都要上到耶和华这里来，远远地下拜。
EXOD|24|2|只有 摩西 可以接近耶和华，其他的人却不可接近；百姓也不可和他一同上来。”
EXOD|24|3|摩西 下山，向百姓陈述耶和华一切的命令和典章。众百姓齐声说：“耶和华所吩咐的一切，我们都必遵行。”
EXOD|24|4|摩西 将耶和华一切的命令都写下来。 他清早起来，在山脚筑了一座坛，按着 以色列 十二支派立了十二根石柱。
EXOD|24|5|他差派 以色列 的年轻人去献燔祭，又宰牛献给耶和华为平安祭。
EXOD|24|6|摩西 将血的一半盛在盆中，另一半洒在坛上。
EXOD|24|7|然后，他拿起约书来，念给百姓听。他们说：“耶和华所吩咐的一切，我们都必遵行，也必听从。”
EXOD|24|8|摩西 把血洒在百姓身上，说：“看哪！这是立约的血，是耶和华按照这一切的命令和你们立约的凭据。”
EXOD|24|9|摩西 、 亚伦 、 拿答 、 亚比户 ，以及 以色列 长老中的七十人都上去，
EXOD|24|10|看见了 以色列 的上帝。在他的脚下，仿佛有蓝宝石铺道，明净如天。
EXOD|24|11|他不把手伸在 以色列 领袖的身上。他们瞻仰上帝，又吃又喝。
EXOD|24|12|耶和华对 摩西 说：“你上山到我这里来，就在那里，我要将石版，就是我所写的律法和诫命赐给你，使你可以教导他们。”
EXOD|24|13|摩西 和他的助手 约书亚 站起来； 摩西 上了上帝的山。
EXOD|24|14|摩西 对长老们说：“你们在这里等我们，直到我们再回到你们这里。看哪， 亚伦 和 户珥 与你们同在。谁有诉讼，可以去找他们。”
EXOD|24|15|摩西 上山，有云彩把山遮盖。
EXOD|24|16|耶和华的荣耀驻在 西奈山 ，云彩遮盖了山六天，第七天他从云中呼叫 摩西 。
EXOD|24|17|耶和华的荣耀在山顶上，在 以色列 人眼前，形状如吞噬的火。
EXOD|24|18|摩西 进入云中，登上了山。 摩西 在山上四十昼夜。
EXOD|25|1|耶和华吩咐 摩西 说：
EXOD|25|2|“你要吩咐 以色列 人献礼物给我。凡甘心乐意献给我的礼物，你们都可以收下。
EXOD|25|3|要从他们收的礼物是：金、银、铜，
EXOD|25|4|蓝色、紫色、朱红色纱 ，细麻，山羊毛，
EXOD|25|5|染红的公羊皮、精美的皮料，金合欢木，
EXOD|25|6|点灯的油，做膏油的香料、做香的香料，
EXOD|25|7|红玛瑙与宝石，可以镶嵌在以弗得和胸袋上。
EXOD|25|8|他们要为我造圣所，使我住在他们中间。
EXOD|25|9|你们要按照我指示你的，帐幕和其中一切器具的样式，照样去做。”
EXOD|25|10|“他们要用金合欢木做一个柜子，长二肘半，宽一肘半，高一肘半。
EXOD|25|11|你要把它里里外外包上纯金，四围要镶上金边。
EXOD|25|12|要铸造四个金环，安在柜子的四脚上；这边两个环，那边两个环。
EXOD|25|13|要用金合欢木做两根杠，包上金子。
EXOD|25|14|要把杠穿过柜旁的环，以便抬柜。
EXOD|25|15|这杠要留在柜的环内，不可抽出来。
EXOD|25|16|要把我所要赐给你的法版 放在柜里。
EXOD|25|17|要用纯金做一个柜盖 ，长二肘半，宽一肘半。
EXOD|25|18|要造两个用金子锤出的基路伯，从柜盖的两端锤出它们。
EXOD|25|19|这端锤出一个基路伯，那端锤出一个基路伯；从柜盖的两端锤出两个基路伯。
EXOD|25|20|二基路伯的翅膀要向上张开，用翅膀遮住柜盖，脸要彼此相对；基路伯的脸要朝向柜盖。
EXOD|25|21|要把柜盖安在柜的上边，又要把我所要赐给你的法版放在柜里。
EXOD|25|22|我要在那里与你相会，并要从法版之柜的柜盖上，两个基路伯的中间，将我要吩咐 以色列 人的一切事告诉你。”
EXOD|25|23|“你要用金合欢木做一张供桌，长二肘，宽一肘，高一肘半，
EXOD|25|24|把它包上纯金，四围镶上金边。
EXOD|25|25|供桌的四围各做一掌宽的边缘，边缘周围要镶上金边。
EXOD|25|26|要为供桌做四个金环，把环安在四个桌脚的四角上。
EXOD|25|27|环要靠近边缘，以便穿杠抬供桌。
EXOD|25|28|要用金合欢木做两根杠，包上金子，用来抬供桌。
EXOD|25|29|要用纯金做桌上的盘、碟，以及浇酒祭的壶和杯。
EXOD|25|30|要把供饼摆在桌上，常在我面前。”
EXOD|25|31|“要造一座用纯金锤出的灯台。灯台的座、干、杯、花萼和花瓣，都要和灯台接连一块。
EXOD|25|32|灯台两旁要伸出六根枝子：这边三根，那边三根。
EXOD|25|33|这边枝子上有三个杯，形状像杏花，有花萼有花瓣；那边枝子上也有三个杯，形状像杏花，有花萼有花瓣。从灯台伸出来的六根枝子都是如此。
EXOD|25|34|灯台本身要有四个杯，形状像杏花，有花萼有花瓣。
EXOD|25|35|灯台的第一对枝子下面有花萼，灯台的第二对枝子下面有花萼，灯台的第三对枝子下面也有花萼；灯台伸出的六根枝子都是如此。
EXOD|25|36|花萼和枝子都要和灯台接连一块，全是从一块纯金锤出来的。
EXOD|25|37|要做灯台的七盏灯，灯要点燃，照亮前面。
EXOD|25|38|要用纯金做灯剪和灯盘。
EXOD|25|39|做灯台和这一切的器具要用一他连得纯金。
EXOD|25|40|要谨慎，照着在山上指示你的样式去做。”
EXOD|26|1|“你要用十幅幔子做帐幕。这些幔子要用搓的细麻和蓝色、紫色、朱红色纱织成，并且以刺绣的手艺绣上基路伯。
EXOD|26|2|每幅幔子要长二十八肘，每幅幔子宽四肘，全部的幔子尺寸都要一样。
EXOD|26|3|这五幅幔子要彼此相连；那五幅也彼此相连。
EXOD|26|4|在这一组相连幔子的末幅边上要缝蓝色的钮环；在另一组相连幔子的末幅边上也要照样做。
EXOD|26|5|这幅幔子上要缝五十个钮环，另一组相连幔子的末幅上也缝五十个钮环，环环相对。
EXOD|26|6|要做五十个金钩，用钩子使幔子彼此相连，成为一个帐幕。
EXOD|26|7|“你要用山羊毛织十一幅幔子来作帐幕的罩棚。
EXOD|26|8|每幅幔子要长三十肘，每幅幔子宽四肘；十一幅幔子的尺寸都要一样。
EXOD|26|9|要把五幅幔子连成一幅，又把六幅幔子连成一幅，这第六幅幔子要在罩棚的前面摺上去。
EXOD|26|10|在这一组相连幔子的末幅边上要缝五十个钮环；在另一组相连幔子的末幅边上也缝五十个钮环。
EXOD|26|11|要做五十个铜钩，钩在钮环中，使罩棚相连成为一个。
EXOD|26|12|罩棚幔子余下垂着的，那余下的半幅要垂在帐幕的背面。
EXOD|26|13|罩棚的幔子两旁所余下的，这边一肘，那边一肘，要垂在帐幕的两边，盖住帐幕。
EXOD|26|14|要用染红的公羊皮做罩棚的盖，再用精美皮料做外层的盖。
EXOD|26|15|“你要用金合欢木做竖立帐幕的木板，
EXOD|26|16|木板要长十肘，每块板宽一肘半，
EXOD|26|17|每块板有两个榫头可以彼此衔接。帐幕一切的板都要这样做。
EXOD|26|18|你要做帐幕的木板：南面，就是面向南方的那一边，要做二十块板。
EXOD|26|19|在这二十块板底下要做四十个带卯眼的银座；两个卯眼接连这块板上的两个榫头，另外两个卯眼接连那块板上的两个榫头。
EXOD|26|20|帐幕的第二边，就是北面，也要做二十块板，
EXOD|26|21|和四十个带卯眼的银座；这块板底下有两个卯眼，那块板底下也有两个卯眼。
EXOD|26|22|帐幕的后面，就是西面，要做六块板。
EXOD|26|23|帐幕后面的角落要做两块板。
EXOD|26|24|下端的板是成双的，上端要连在一起，直到顶端的第一个环子；两块板都要这样，做成两个角落。
EXOD|26|25|一共有八块板和十六个带卯眼的银座；这块板底下有两个卯眼，那块板底下也有两个卯眼。
EXOD|26|26|“你要用金合欢木做横木：为帐幕这面的板做五根横木，
EXOD|26|27|为帐幕那面的板做五根横木，又为帐幕后面，就是朝西的板做五根横木。
EXOD|26|28|板腰间的横木，要从一头通到另一头。
EXOD|26|29|板要包上金子，又要做板上的金环来套横木；横木也要包上金子。
EXOD|26|30|要照着在山上所指示你的样式，把帐幕竖立起来。
EXOD|26|31|“你要用蓝色、紫色、朱红色纱，和搓的细麻织幔子，以刺绣的手艺绣上基路伯。
EXOD|26|32|要把幔子挂在四根包金的金合欢木柱子上，柱子有金钩，并且安在四个带卯眼的银座上。
EXOD|26|33|要把幔子垂挂在钩子上，把法柜抬进幔子内；这幔子要将圣所和至圣所隔开。
EXOD|26|34|又要把柜盖安在至圣所内的法柜上，
EXOD|26|35|把供桌安在幔子的外面，供桌在北面，灯台在帐幕的南面，和供桌相对。
EXOD|26|36|“你要用蓝色、紫色、朱红色纱，和搓的细麻，以刺绣的手艺为帐幕织门帘。
EXOD|26|37|要用金合欢木为帘子做五根柱子，包上金子。柱子有金钩，又为柱子铸造五个带卯眼的铜座。”
EXOD|27|1|“你要用金合欢木做祭坛，长五肘，宽五肘，这坛是正方形的，高三肘。
EXOD|27|2|要在坛的四角做四个翘角，与坛接连一块；要把坛包上铜。
EXOD|27|3|要做桶子来盛坛上的灰，又要做铲子、盘子、肉叉和火盆；坛上一切的器具都要用铜做。
EXOD|27|4|要为坛做一个铜网，在网的四角做四个铜环，
EXOD|27|5|把网安在坛四围的边的下面，使网垂到坛的半腰。
EXOD|27|6|又要用金合欢木为坛做杠，包上铜。
EXOD|27|7|这杠要穿过坛两旁的环子，用来抬坛。
EXOD|27|8|要用板做坛，坛的中心是空的，都照着在山上所指示你的样式做。”
EXOD|27|9|“你要做帐幕的院子。南面，就是面向南方的那一边，要用搓的细麻做院子的帷幔，长一百肘，
EXOD|27|10|院子要有二十根柱子，二十个带卯眼的铜座。要用银做柱子的钩和箍。
EXOD|27|11|北面的长度也一样，帷幔长一百肘，要有二十根柱子，二十个带卯眼的铜座。要用银做柱子的钩和箍。
EXOD|27|12|院子的西面有帷幔，宽五十肘，帷幔要有十根柱子，十个带卯眼的座。
EXOD|27|13|院子的东面，就是面向东方的那一边，宽五十肘。
EXOD|27|14|一边的帷幔有十五肘，要有三根柱子，三个带卯眼的座。
EXOD|27|15|另一边的帷幔也有十五肘，要有三根柱子，三个带卯眼的座。
EXOD|27|16|院子的门要有二十肘长的帘子，用蓝色、紫色、朱红色纱，和搓的细麻，以刺绣的手艺织成；要有四根柱子，四个带卯眼的座。
EXOD|27|17|院子四围一切的柱子都要用银子箍着，要用银做柱子的钩子，用铜做带卯眼的座。
EXOD|27|18|院子要长一百肘，宽五十肘 ，高五肘。要用搓的细麻做帷幔，用铜做带卯眼的座。
EXOD|27|19|帐幕中各样用途的器具，以及帐幕一切的橛子和院子里一切的橛子，都要用铜做。”
EXOD|27|20|“你要吩咐 以色列 人，把捣成的纯橄榄油拿来给你，用以点灯，使灯经常点着；
EXOD|27|21|在会幕中法柜前的幔子外， 亚伦 和他的儿子要从晚上到早晨，在耶和华面前照管这灯。这要成为 以色列 人世世代代永远的定例。”
EXOD|28|1|“你要从 以色列 人中，叫你的哥哥 亚伦 和他的儿子 拿答 、 亚比户 、 以利亚撒 、 以他玛 一同亲近你，作事奉我的祭司。
EXOD|28|2|你要为你哥哥 亚伦 做圣衣，以示尊严和华美。
EXOD|28|3|要吩咐一切心中有智慧的，就是我用智慧的灵所充满的人，为 亚伦 做衣服，使他分别为圣，作事奉我的祭司。
EXOD|28|4|所要做的是胸袋、以弗得、外袍、织成的内袍、礼冠和腰带。他们要为你哥哥 亚伦 和他的儿子做圣衣，使他们作祭司事奉我。
EXOD|28|5|要用金色、蓝色、紫色、朱红色纱，和细麻去缝制。
EXOD|28|6|“他们要用金色、蓝色、紫色、朱红色纱，和搓的细麻，以刺绣的手艺做以弗得。
EXOD|28|7|以弗得当有两条肩带，接上两端，使它相连。
EXOD|28|8|以弗得的精致带子，要以一样的手艺，用金色、蓝色、紫色、朱红色纱，和搓的细麻缝制，与以弗得接连在一起。
EXOD|28|9|要取两块红玛瑙，在上面刻 以色列 儿子的名字：
EXOD|28|10|六个名字在一块宝石上，六个名字在另一块宝石上，都按照他们出生的次序。
EXOD|28|11|要以雕刻宝石的手艺，如同刻印章，把 以色列 儿子的名字刻在这两块宝石上，并把宝石镶在金槽里。
EXOD|28|12|要把这两块宝石安在以弗得的两条肩带上，为 以色列 人作纪念石。 亚伦 要在耶和华面前把他们的名字带在两肩上，作为纪念。
EXOD|28|13|要用金子做两个槽，
EXOD|28|14|再用纯金打两条链子，像编成的绳子一样，把这编成的金链扣在槽上。”
EXOD|28|15|“你要以刺绣的手艺做一个决断的胸袋，和做以弗得的方法一样，用金色、蓝色、紫色、朱红色纱，和搓的细麻缝制。
EXOD|28|16|胸袋是正方形的，叠成两层，长一虎口，宽一虎口。
EXOD|28|17|要在上面镶四行宝石：第一行是红宝石、红璧玺、红玉；
EXOD|28|18|第二行是绿宝石、蓝宝石、金刚石；
EXOD|28|19|第三行是紫玛瑙、白玛瑙、紫晶；
EXOD|28|20|第四行是水苍玉、红玛瑙、碧玉。这些都要镶在金槽中。
EXOD|28|21|这些宝石要有 以色列 十二个儿子的名字，如同刻印章，每一颗有自己的名字，代表十二个支派。
EXOD|28|22|要在胸袋上用纯金打链子，像编成的绳子一样。
EXOD|28|23|要为胸袋做两个金环，把这两个环安在胸袋的两端。
EXOD|28|24|要把那两条编成的金链系在胸袋两端的两个环上。
EXOD|28|25|又要把链子的另外两端扣在两个槽上，安在以弗得前面的肩带上。
EXOD|28|26|要做两个金环，安在胸袋的两端，在以弗得里面的边上。
EXOD|28|27|再做两个金环，安在以弗得前面两条肩带的下边，靠近接缝处，在以弗得精致带子的上面。
EXOD|28|28|要用蓝色的带子把胸袋的环与以弗得的环系住，使胸袋绑在以弗得的精致带子上，不致松脱。
EXOD|28|29|亚伦 进圣所的时候，要把刻着 以色列 儿子名字的决断胸袋带着，放在心上，在耶和华面前常作纪念。
EXOD|28|30|又要将乌陵和土明 放在决断胸袋里； 亚伦 进到耶和华面前的时候，要放在心上。这样， 亚伦 在耶和华面前要把 以色列 人的决断胸袋常常带着，放在心上。”
EXOD|28|31|“你要做以弗得的外袍，颜色全是蓝的。
EXOD|28|32|袍上方的中间要留一个领口，领口周围的领边要以手艺编织而成，好像铠甲的领口，免得破裂。
EXOD|28|33|袍子下摆，就是下摆的周围要用蓝色、紫色、朱红色纱做石榴，周围的石榴中间要有金铃铛：
EXOD|28|34|一个金铃铛一个石榴，一个金铃铛一个石榴，在袍子下摆的周围。
EXOD|28|35|亚伦 供职的时候要穿这袍。他进入圣所到耶和华面前，以及出来的时候，袍上的铃声必被听见，使他不至于死。
EXOD|28|36|“你要用纯金做一面牌，如同刻印章，在上面刻‘归耶和华为圣’。
EXOD|28|37|要用蓝色的带子把牌系在礼冠上，在礼冠的正前面。
EXOD|28|38|这牌必在 亚伦 的额上， 亚伦 要担当干犯圣物的罪孽；这圣物是 以色列 人在一切圣礼物上所分别为圣的。这牌要常在他的额上，使他们可以在耶和华面前蒙悦纳。
EXOD|28|39|要用细麻编织内袍，用细麻做礼冠，又以刺绣的手艺做腰带。
EXOD|28|40|“你要为 亚伦 的儿子做内袍、腰带、头巾，以示尊严和华美。
EXOD|28|41|要把这些给你哥哥 亚伦 和他的儿子穿戴，又要膏他们，授予圣职，使他们分别为圣，作事奉我的祭司。
EXOD|28|42|要用细麻布给他们做裤子来遮掩下体，从腰间直到大腿。
EXOD|28|43|亚伦 和他儿子进入会幕，或接近祭坛，在圣所供职的时候要穿上裤子，免得担当罪孽而死。这要成为 亚伦 和他后裔永远的定例。”
EXOD|29|1|“这是你使他们分别为圣，作事奉我的祭司时要做的事：取一头公牛犊，两只无残疾的公绵羊，
EXOD|29|2|无酵饼、用油调和的无酵饼，和抹油的无酵薄饼；这些饼都要用细麦面做成。
EXOD|29|3|这些饼要装在一个篮子里，用篮子带来，又把公牛和两只公绵羊牵来。
EXOD|29|4|要带 亚伦 和他儿子到会幕的门口，用水洗他们。
EXOD|29|5|要拿服装，给 亚伦 穿上内袍和以弗得的外袍，以及以弗得，又带上胸袋，束上以弗得精致的带子。
EXOD|29|6|要把礼冠戴在他头上，将圣冕加在礼冠上，
EXOD|29|7|把膏油倒在他头上膏他。
EXOD|29|8|要带他的儿子来，给他们穿上内袍。
EXOD|29|9|要给 亚伦 和他的儿子束上腰带，裹上头巾，他们就凭永远的定例得祭司的职分。又要授圣职给 亚伦 和他的儿子。
EXOD|29|10|“你要把公牛牵到会幕前， 亚伦 和他的儿子要按手在公牛的头上。
EXOD|29|11|你要在耶和华面前，在会幕的门口宰这公牛。
EXOD|29|12|要取些公牛的血，用指头抹在祭坛的四个翘角上，把其余的血全倒在坛的底座上。
EXOD|29|13|要把所有包着内脏的脂肪、肝上的网油、两个肾和肾上的脂肪，都烧在坛上。
EXOD|29|14|只是公牛的肉、皮、粪都要在营外用火焚烧；这牛是赎罪祭。
EXOD|29|15|“你要牵一只公绵羊来， 亚伦 和他儿子要按手在这羊的头上。
EXOD|29|16|你要宰这羊，把血洒在祭坛的周围。
EXOD|29|17|再把羊切成肉块，洗净内脏和腿，连肉块和头放在一处。
EXOD|29|18|要把全羊烧在坛上。这是献给耶和华的燔祭，是献给耶和华馨香的火祭。”
EXOD|29|19|“你要把第二只公绵羊牵来， 亚伦 和他儿子要按手在这羊的头上。
EXOD|29|20|你要宰这羊，取些血抹在 亚伦 的右耳垂和他儿子的右耳垂上，又抹在他们右手的大拇指和右脚的大脚趾上，然后把其余的血洒在坛的周围。
EXOD|29|21|你要取些膏油和坛上的血，弹在 亚伦 和他的衣服上，以及他儿子和他们的衣服上； 亚伦 和他的衣服，他儿子和他们的衣服都成为圣了。
EXOD|29|22|“你要取这羊的脂肪，肥尾巴、包着内脏的脂肪、肝上的网油、两个肾、肾上的脂肪和右腿，这是圣职礼所献的公绵羊；
EXOD|29|23|再从耶和华面前那装无酵饼的篮子中取一个饼、一个油饼和一个薄饼，
EXOD|29|24|把它们都放在 亚伦 的手和他儿子的手上，在耶和华面前摇一摇，作为摇祭。
EXOD|29|25|然后，你要从他们手中接过来，放在燔祭上，一起烧在坛上，作为耶和华面前馨香之气；这是献给耶和华的火祭。
EXOD|29|26|“你要取 亚伦 圣职礼所献公绵羊的胸，在耶和华面前摇一摇，作为摇祭；这份就是你的。
EXOD|29|27|那摇祭的胸和举祭的腿，就是圣职礼献公绵羊时所摇的、所举的，你要使它们分别为圣，是归给 亚伦 和他儿子的。
EXOD|29|28|这是 亚伦 和他子孙凭永远的定例从 以色列 人中所应得的；因为这是举祭，是从 以色列 人的平安祭中取出，作为献给耶和华的举祭。
EXOD|29|29|“ 亚伦 的圣衣要传给他的子孙，使他们在受膏和承接圣职的时候穿上。
EXOD|29|30|他的子孙接续他当祭司的，每逢进入会幕在圣所供职的时候，要穿这圣衣七天。
EXOD|29|31|“你要拿圣职礼所献的公绵羊，在圣处煮它的肉。
EXOD|29|32|亚伦 和他儿子要在会幕的门口吃这羊的肉和篮子里的饼。
EXOD|29|33|他们要吃那些用来赎罪之物，好承接圣职，使他们分别为圣。外人不可吃，因为这是圣物。
EXOD|29|34|那圣职礼所献的肉或饼，若有剩余留到早晨，就要把剩下的用火烧了，不可再吃，因为这是圣物。
EXOD|29|35|“你要这样照我一切所吩咐的，向 亚伦 和他儿子行授圣职礼七天。
EXOD|29|36|为了赎罪，每天要献一头公牛为赎罪祭。你要为祭坛赎罪，使坛洁净，并要用膏抹坛，使坛成为圣。
EXOD|29|37|要为坛赎罪七天，使坛成为圣，坛就成为至圣。凡触摸坛的都成为圣。”
EXOD|29|38|“这是你要献在坛上的：每天不可间断地献两只一岁的羔羊；
EXOD|29|39|早晨献第一只羔羊，黄昏献第二只羔羊。
EXOD|29|40|献第一只羔羊时，要同时献上十分之一伊法细面，调和四分之一欣捣成的油，再献四分之一欣酒作浇酒祭。
EXOD|29|41|黄昏你献第二只羔羊，要照早晨的素祭和同献的浇酒祭献上，作为献给耶和华馨香的火祭。
EXOD|29|42|这要在耶和华面前，在会幕的门口，作为你们世世代代经常献的燔祭。我要在那里与你们 相会，和你说话。
EXOD|29|43|我要在那里与 以色列 人相会，会幕就要因我的荣耀成为圣。
EXOD|29|44|我要使会幕和祭坛分别为圣，也要使 亚伦 和他的儿子分别为圣，作事奉我的祭司。
EXOD|29|45|我要住在 以色列 人中，作他们的上帝。
EXOD|29|46|他们必知道我是耶和华－他们的上帝，是将他们从 埃及 地领出来的，为要住在他们中间。我是耶和华－他们的上帝 。”
EXOD|30|1|“你要用金合欢木做一座烧香的坛，
EXOD|30|2|长一肘，宽一肘，这坛是正方形的，高二肘。坛的四个翘角与坛接连一块。
EXOD|30|3|要把坛的上面与坛的四围，以及坛的四个翘角包上纯金；又要在坛的四围镶上金边。
EXOD|30|4|要在坛的两个对侧，金边下面做两个金环，用来穿杠抬坛。
EXOD|30|5|要用金合欢木做杠，包上金子。
EXOD|30|6|要把坛放在法柜前的幔子外，对着法柜上的柜盖，就是我与你相会的地方。
EXOD|30|7|亚伦 要在坛上烧芬芳的香；每早晨整理灯的时候，他都要烧这香。
EXOD|30|8|黄昏点灯的时候， 亚伦 也要烧这香。这是你们世世代代在耶和华面前常烧的香。
EXOD|30|9|在这坛上不可烧别样的香，不可献燔祭、素祭，也不可献浇酒祭。
EXOD|30|10|亚伦 每年一次要为坛的四个翘角赎罪。他每年一次要用赎罪祭的血为坛赎罪，作为世世代代的定例。这坛在耶和华面前是至圣的。”
EXOD|30|11|耶和华吩咐 摩西 说：
EXOD|30|12|“你数点 以色列 人，计算人头时，被数的每一个人要把他生命的赎价献给耶和华，免得灾殃在数点中临到他们。
EXOD|30|13|每一个被数的人要按照圣所的舍客勒，付半舍客勒，一舍客勒是二十季拉；这半舍客勒是献给耶和华的礼物。
EXOD|30|14|每一个被数的人，就是二十岁以上的，要将这礼物献给耶和华。
EXOD|30|15|富有的不必多付，贫穷的也不可少出，各人都要献半舍客勒给耶和华，作你们生命的赎价。
EXOD|30|16|你要向 以色列 人收这赎罪的银子，用在会幕的事工。这要在耶和华面前为 以色列 人作纪念，作你们生命的赎价。”
EXOD|30|17|耶和华吩咐 摩西 说：
EXOD|30|18|“你要用铜做洗濯盆和盆座，用来洗濯。要将盆放在会幕和祭坛的中间，盆里盛水。
EXOD|30|19|亚伦 和他的儿子要用这盆洗手洗脚。
EXOD|30|20|他们进会幕，或是走近坛前供职，献火祭给耶和华的时候，必须用水洗濯，免得死亡；
EXOD|30|21|他们要洗手洗脚，免得死亡。这是 亚伦 和他的后裔世世代代永远的定例。”
EXOD|30|22|耶和华吩咐 摩西 说：
EXOD|30|23|“你要取上等的香料，就是五百舍客勒流质的没药、二百五十香肉桂、二百五十香菖蒲，
EXOD|30|24|和五百桂皮，都按照圣所的舍客勒；再取一欣橄榄油，
EXOD|30|25|以做香的方法调和制成圣膏油，它就成为圣膏油。
EXOD|30|26|要用这膏油抹会幕和法柜，
EXOD|30|27|供桌和供桌的一切器具，灯台和灯台的器具 ，以及香坛、
EXOD|30|28|燔祭坛和坛的一切器具，洗濯盆和盆座。
EXOD|30|29|你要使这些分别为圣，成为至圣；凡触摸它们的都成为圣。
EXOD|30|30|要膏 亚伦 和他的儿子，使他们分别为圣，作事奉我的祭司。
EXOD|30|31|你要吩咐 以色列 人说：‘你们要世世代代以这油为我的圣膏油。
EXOD|30|32|不可把这油倒在别人身上，也不可用配制这膏油的方法制成同样的膏油。这膏油是圣的，你们要以它为圣。
EXOD|30|33|凡调和与此类似的膏油，或将它膏在别人身上的，这人要从百姓中剪除。’”
EXOD|30|34|耶和华吩咐 摩西 说：“你要取香料，就是拿他弗、施喜列、喜利比拿，这些香料再加纯乳香，每样都要相同的分量。
EXOD|30|35|你要用这些加上盐，以配制香料的方法，制成纯净又神圣的香。
EXOD|30|36|要取一点这香，捣成细的粉，放在会幕中的法柜前，就是我和你相会的地方。你们要以这香为至圣。
EXOD|30|37|你们不可用这配制的方法为自己做香；要以这香为圣，归于耶和华。
EXOD|30|38|为要闻香味而配制同样的香的，这人要从百姓中剪除。”
EXOD|31|1|耶和华吩咐 摩西 说：
EXOD|31|2|“你看，我已经题名召 犹大 支派中 户珥 的孙子， 乌利 的儿子 比撒列 。
EXOD|31|3|我以上帝的灵充满他，使他有智慧，有聪明，有知识，能做各样的工，
EXOD|31|4|能设计图案，用金、银、铜制造各物，
EXOD|31|5|又能雕刻镶嵌用的宝石，雕刻木头，做各样的工。
EXOD|31|6|看哪，我委派 但 支派中 亚希撒抹 的儿子 亚何利亚伯 与他同工。凡心里有智慧的，我更要赐给他们智慧的心，能做我所吩咐你的一切，
EXOD|31|7|就是会幕、法柜和其上的柜盖、会幕中一切的器具、
EXOD|31|8|供桌和供桌的器具、纯金的灯台和灯台的一切器具、香坛、
EXOD|31|9|燔祭坛和坛的一切器具、洗濯盆与盆座、
EXOD|31|10|供祭司职分用的精致礼服， 亚伦 祭司的圣衣和他儿子的衣服，
EXOD|31|11|以及膏油和圣所用的芬芳的香。他们都要照我所吩咐的一切去做。”
EXOD|31|12|耶和华对 摩西 说：
EXOD|31|13|“你要吩咐 以色列 人说：‘你们务要守我的安息日，因为这是你我之间世世代代的记号，叫你们知道我是耶和华，是使你们分别为圣的。
EXOD|31|14|你们要守安息日，以它为圣日。凡干犯这日的，必被处死；凡在这日做工的，那人必从百姓中剪除。
EXOD|31|15|六日要做工，但第七日是向耶和华守完全安息的安息圣日。凡在安息日做工的，必被处死。’
EXOD|31|16|以色列 人要守安息日，世世代代守安息日为永远的约。
EXOD|31|17|这是我和 以色列 人之间永远的记号，因为六日之内耶和华造天地，第七日就安息舒畅。”
EXOD|31|18|耶和华在 西奈山 和 摩西 说完了话，就把两块法版交给他，是上帝用指头写的石版。
EXOD|32|1|百姓见 摩西 迟迟不下山，就聚集到 亚伦 那里，对他说：“起来！为我们造神明，在我们前面引路，因为领我们出 埃及 地的那个 摩西 ，我们不知道他遭遇了什么事。”
EXOD|32|2|亚伦 对他们说：“你们去摘下你们妻子、儿女耳上的金环，拿来给我。”
EXOD|32|3|众百姓就摘下他们耳上的金环，拿来给 亚伦 。
EXOD|32|4|亚伦 从他们手里接过来，用模子塑造它，把它铸成一头牛犊。他们就说：“ 以色列 啊，这是领你出 埃及 地的神明！”
EXOD|32|5|亚伦 看见，就在牛犊面前筑坛。 亚伦 宣告说：“明日要向耶和华守节。”
EXOD|32|6|次日清早，百姓起来献燔祭和平安祭，就坐下吃喝，起来玩乐。
EXOD|32|7|耶和华吩咐 摩西 ：“下去吧，因为你从 埃及 领上来的百姓已经败坏了。
EXOD|32|8|他们这么快偏离了我所吩咐的道，为自己铸了一头牛犊，向它跪拜，向它献祭，说：‘ 以色列 啊，这就是领你出 埃及 地的神明。’”
EXOD|32|9|耶和华对 摩西 说：“我看这百姓，看哪，他们真是硬着颈项的百姓。
EXOD|32|10|现在，你且由着我，我要向他们发烈怒，灭绝他们，但我要使你成为大国。”
EXOD|32|11|摩西 就恳求耶和华－他的上帝，说：“耶和华啊，你为什么向你的百姓发烈怒呢？这百姓是你用大能大力的手从 埃及 地领出来的！
EXOD|32|12|为什么让 埃及 人说：‘他领他们出去，是要降灾祸给他们，在山中把他们杀了，将他们从地上除灭’呢？求你回心转意，不发你的烈怒，不降灾祸给你的百姓。
EXOD|32|13|求你记念你的仆人 亚伯拉罕 、 以撒 、 以色列 。你曾向他们指着自己起誓说：‘我必使你们的后裔像天上的星那样多，并且我要将所应许的这全地赐给你们的后裔，让他们永远承受为业。’”
EXOD|32|14|于是耶和华改变心意，不把所说的灾祸降给他的百姓。
EXOD|32|15|摩西 转身下山，手里拿着两块法版。这版的两面都写着字，正面背面都有字。
EXOD|32|16|版是上帝的工作，字是上帝写的字，刻在版上。
EXOD|32|17|约书亚 一听见百姓呼喊的声音，就对 摩西 说：“在营里有战争的声音。”
EXOD|32|18|摩西 说：“这不是打胜仗的声音，也不是打败仗的声音，我听见的是歌唱的声音。”
EXOD|32|19|摩西 走近营前，看见牛犊，又看见人在跳舞，就发烈怒，把两块版从手中扔到山下摔碎了。
EXOD|32|20|他将他们所铸的牛犊用火焚烧，磨得粉碎，撒在水面上，叫 以色列 人喝。
EXOD|32|21|摩西 对 亚伦 说：“这百姓向你做了什么呢？你竟使他们陷入大罪中！”
EXOD|32|22|亚伦 说：“求我主不要发烈怒。你知道这百姓，他们是向恶的。
EXOD|32|23|他们对我说：‘你为我们造神明，在我们前面引路，因为领我们出 埃及 地的那个 摩西 ，我们不知道他遭遇了什么事。’
EXOD|32|24|我对他们说：‘凡有金环的可以摘下来’，他们就给了我。我把金环扔在火中，这牛犊就出来了。”
EXOD|32|25|摩西 见百姓放肆，因 亚伦 纵容他们，使这事成了敌人的笑柄，
EXOD|32|26|就站在营门前，说：“凡属耶和华的人，都到我这里来！”于是 利未 人都聚集到他那里。
EXOD|32|27|他对他们说：“耶和华－ 以色列 的上帝这样说：‘你们各人把刀佩在腰间，从这门到那门，来回走遍全营，各人要杀自己的弟兄、邻舍和亲人。’”
EXOD|32|28|利未 人遵照 摩西 的话做了。那一天百姓中倒下的约有三千人。
EXOD|32|29|摩西 说：“今天你们要奉献自己 来事奉耶和华，因为各人牺牲自己的儿子和弟兄，使耶和华今天赐福给你们。”
EXOD|32|30|第二天， 摩西 对百姓说：“你们犯了大罪。我如今要上耶和华那里去，或许可以为你们赎罪。”
EXOD|32|31|摩西 回到耶和华那里，说：“唉！这百姓犯了大罪，为自己造了金的神明。
EXOD|32|32|现在，求你赦免他们的罪；不然，就把我从你所写的册上除名。”
EXOD|32|33|耶和华对 摩西 说：“谁得罪我，我就把他从我的册上除去。
EXOD|32|34|现在你去，领这百姓往我所告诉你的地方去，看哪，我的使者必在你的前面引路。到了该惩罚的时候，我必惩罚他们的罪。”
EXOD|32|35|耶和华降灾与百姓，因为他们和 亚伦 一起造了牛犊。
EXOD|33|1|耶和华吩咐 摩西 说：“去，离开这里，你和你从 埃及 地领出来的百姓要上到我起誓应许给 亚伯拉罕 、 以撒 和 雅各 之地去；我曾对他们说：‘我要将这地赐给你的后裔’。
EXOD|33|2|我要差遣使者在你前面，把 迦南 人、 亚摩利 人、 赫 人、 比利洗 人、 希未 人、 耶布斯 人赶出
EXOD|33|3|那流奶与蜜之地。但我不与你们上去，因为你们是硬着颈项的百姓，免得我在路上把你们灭绝。”
EXOD|33|4|百姓一听见这坏的信息，他们就悲哀，没有人佩戴首饰。
EXOD|33|5|耶和华对 摩西 说：“你对 以色列 人说：‘你们是硬着颈项的百姓，我若在你们中间一起上去，只一瞬间，就必把你们灭绝。现在把你们身上的首饰摘下来，我好知道该怎样处置你们。’”
EXOD|33|6|以色列 人离开 何烈山 以后，就把身上的首饰全都摘下来。
EXOD|33|7|摩西 拿一个帐棚支搭在营外，离营有一段距离，他称这帐棚为会幕。凡求问耶和华的，就到营外的会幕那里去。
EXOD|33|8|当 摩西 出营到会幕去的时候，百姓就都起来，各人站在自己帐棚的门口，望着 摩西 ，直到他进了会幕。
EXOD|33|9|摩西 进会幕的时候，云柱就降下来，停在会幕的门前，耶和华就与 摩西 说话。
EXOD|33|10|众百姓看见云柱停在会幕的门前，就都起来，各人在自己帐棚的门口下拜。
EXOD|33|11|耶和华与 摩西 面对面说话，好像人与朋友说话。 摩西 回到营里去，他的年轻助手 嫩 的儿子 约书亚 却没有离开会幕。
EXOD|33|12|摩西 对耶和华说：“看，你曾对我说：‘将这百姓领上去’；却没有让我知道你要差派谁与我同去。你还说：‘我按你的名认识你，你也在我眼前蒙了恩。’
EXOD|33|13|我如今若在你眼前蒙恩，求你将你的道指示我，使我可以认识你，并在你眼前蒙恩。求你顾念这国是你的子民。”
EXOD|33|14|耶和华说：“我必亲自去，让你安心。”
EXOD|33|15|摩西 说：“你若不亲自去，就不要把我们从这里领上去。
EXOD|33|16|现在，人如何得知我和你的百姓在你眼前蒙恩呢？岂不是因为你与我们同去，使我和你的百姓与地面上的万民有分别吗？”
EXOD|33|17|耶和华对 摩西 说：“你所说的这件事，我也会去做，因为你在我眼前蒙了恩，并且我按你的名认识你。”
EXOD|33|18|摩西 说：“求你显出你的荣耀给我看。”
EXOD|33|19|耶和华说：“我要显示我一切的美善，在你面前经过，并要在你面前宣告耶和华的名。我要恩待谁就恩待谁，要怜悯谁就怜悯谁。”
EXOD|33|20|他又说：“只是你不能看见我的面，因为没有人看见我还可以存活。”
EXOD|33|21|耶和华说：“看哪，靠近我这里有个地方，你可以站在这磐石上。
EXOD|33|22|当我的荣耀经过的时候，我必将你放在磐石缝里，用我的手掌遮掩你，等我过去，
EXOD|33|23|然后我要将我的手掌收回，你就可以看见我的背，却看不到我的面。”
EXOD|34|1|耶和华对 摩西 说：“你要凿出两块石版，和先前的一样；我要把你摔碎的那版上先前所写的字，写在这版上。
EXOD|34|2|明日早晨，你要预备好了，上 西奈山 ，在山顶那里站在我面前。
EXOD|34|3|谁也不可和你上去，整座山都不可见到人，也不可有羊群牛群在山下吃草。”
EXOD|34|4|摩西 就凿出两块石版，和先前的一样。他清晨起来，遵照耶和华吩咐他的，上 西奈山 去，手里拿着两块石版。
EXOD|34|5|耶和华在云中降临，与 摩西 一同站在那里，宣告耶和华的名。
EXOD|34|6|耶和华在他面前经过，宣告： “耶和华，耶和华， 有怜悯，有恩惠的上帝， 不轻易发怒， 且有丰盛的慈爱和信实，
EXOD|34|7|为千代的人存留慈爱， 赦免罪孽、过犯和罪恶， 万不以有罪的为无罪， 必惩罚人的罪， 自父及子，直到三、四代。”
EXOD|34|8|摩西 急忙俯伏在地敬拜，
EXOD|34|9|说：“主啊，我若在你眼前蒙恩，求主在我们中间同行。虽然这是硬着颈项的百姓，求你赦免我们的罪孽和罪恶，接纳我们为你的产业。”
EXOD|34|10|耶和华说：“看哪，我要立约，要在你众百姓面前行奇妙的事，是在全地万国中未曾做过的。你周围的万民要看见我藉着你所行，耶和华可畏惧的作为。
EXOD|34|11|“我今天所吩咐你的，你要谨守。看哪，我要从你面前赶出 亚摩利 人、 迦南 人、 赫 人、 比利洗 人、 希未 人、 耶布斯 人。
EXOD|34|12|你要谨慎，不可与你所要去那地的居民立约，免得他们成为你中间的圈套。
EXOD|34|13|你要拆毁他们的祭坛，打碎他们的柱像，砍断他们的 亚舍拉 。
EXOD|34|14|不可敬拜别神，因为耶和华是忌邪 的上帝，他的名是忌邪者。
EXOD|34|15|你不可与那地的居民立约，因为他们随从自己的神明行淫；祭他们神明的时候，有人邀请你参加，你就会吃他的祭物。
EXOD|34|16|你为你儿子娶他们的女儿为妻，他们的女儿因着随从她们的神明行淫，就引诱你的儿子也随从她们的神明行淫。
EXOD|34|17|“不可为自己铸造神像。
EXOD|34|18|“你要守除酵节，照我所吩咐你的，在亚笔月内所定的日期吃无酵饼七天，因为你是在亚笔月内出了 埃及 。
EXOD|34|19|“凡头生的都是我的；无论是牛是羊，一切头生的公的牲畜都要分别出来 。
EXOD|34|20|头生的驴可以用羔羊代赎。若不赎它，就要打断它的颈项。凡头生的儿子都要赎出来。没有人可以空手来朝见我。
EXOD|34|21|“六日你要做工，第七日要安息，即使在耕种或收割的时候也要安息。
EXOD|34|22|在收割初熟麦子的时候要守七七节，又要在年底守收藏节。
EXOD|34|23|你所有的男丁要一年三次朝见主耶和华－ 以色列 的上帝。
EXOD|34|24|我要从你面前赶走列国，扩张你的疆界。你一年三次上去朝见耶和华－你上帝的时候，必没有人贪图你的地。
EXOD|34|25|“不可将我祭牲的血和有酵之物一同献上。逾越节的祭牲也不可留到早晨。
EXOD|34|26|土地里上好的初熟之物要奉到耶和华－你上帝的殿。不可用母山羊的奶来煮它的小山羊。”
EXOD|34|27|耶和华对 摩西 说：“你要将这些话写上，因为我按这话与你和 以色列 人立约。”
EXOD|34|28|摩西 在耶和华那里四十昼夜，不吃饭不喝水。他把这约的话，那十条诫命 ，写在版上。
EXOD|34|29|摩西 下 西奈山 。 摩西 从山上下来的时候，手里拿着两块法版。 摩西 不知道自己脸上的皮肤因耶和华和他说话而发光。
EXOD|34|30|亚伦 和 以色列 众人看见 摩西 ，看哪，他脸上的皮肤发光，他们就怕靠近他。
EXOD|34|31|摩西 叫他们来， 亚伦 和会众的官长回到他那里， 摩西 就跟他们说话。
EXOD|34|32|随后 以色列 众人都近前来，他就把耶和华在 西奈山 与他所说的一切话都吩咐他们。
EXOD|34|33|摩西 跟他们说完了话，就用面纱蒙上脸。
EXOD|34|34|但 摩西 进到耶和华面前与他说话的时候，就把面纱揭下，直到出来。 摩西 出来，将所吩咐他的话告诉 以色列 人。
EXOD|34|35|以色列 人看见 摩西 的脸，他脸上的皮肤发光。 摩西 就用面纱蒙上脸，直到他进去与耶和华说话才揭下。
EXOD|35|1|摩西 召集 以色列 全会众，对他们说：“这是耶和华吩咐你们遵行的事：
EXOD|35|2|六日要做工，第七日你们要奉为向耶和华守完全安息的安息圣日。凡在这日做工的，要被处死。
EXOD|35|3|在安息日这一天，不可在你们一切的住处生火。”
EXOD|35|4|摩西 对 以色列 全会众说：“这是耶和华所吩咐的话，说：
EXOD|35|5|要从你们当中拿礼物献给耶和华；凡甘心乐意的，可以把耶和华的礼物拿来，就是金、银、铜，
EXOD|35|6|蓝色、紫色、朱红色纱，细麻，山羊毛，
EXOD|35|7|染红的公羊皮，精美的皮料，金合欢木，
EXOD|35|8|点灯的油，做膏油的香料、做香的香料，
EXOD|35|9|红玛瑙与宝石，可以镶嵌在以弗得和胸袋上。”
EXOD|35|10|“你们当中凡心里有智慧的都要来，制造一切耶和华所吩咐的，
EXOD|35|11|就是帐幕、帐幕的罩棚、帐幕的盖、钩子、竖板、横木、柱子和带卯眼的座，
EXOD|35|12|柜子、柜子的杠、柜盖和遮掩的幔子，
EXOD|35|13|供桌、供桌的杠、供桌一切的器具和供饼，
EXOD|35|14|灯台、灯台的器具、灯和点灯的油，
EXOD|35|15|香坛、坛的杠、膏油和芬芳的香，帐幕门口的门帘，
EXOD|35|16|燔祭坛、坛的铜网、坛的杠和坛的一切器具，洗濯盆和盆座，
EXOD|35|17|院子的帷幔、柱子、带卯眼的座和院子的门帘，
EXOD|35|18|帐幕的橛子、院子的橛子和绳子，
EXOD|35|19|以及圣所事奉用的精致礼服， 亚伦 祭司的圣衣和他儿子的衣服，供祭司职分用。”
EXOD|35|20|以色列 全会众从 摩西 的面前出去。
EXOD|35|21|凡心受感动，灵被驱策的，都带耶和华的礼物来，为要造会幕和其中一切的器具，以及缝制圣衣。
EXOD|35|22|凡甘心乐意的，连男带女都来了，各将金器，就是胸针、耳环、打印的戒指，和项链带来，摇着金器的摇祭献给耶和华。
EXOD|35|23|凡有蓝色、紫色、朱红色纱、细麻、山羊毛、染红的公羊皮、精美皮料的，都拿了来；
EXOD|35|24|凡愿意献银和铜作礼物的，都拿礼物来献给耶和华；凡有金合欢木可做各种用途的也都拿了来。
EXOD|35|25|凡心中有智慧，可以亲手纺织的妇女，也把所纺的蓝色、紫色、朱红色纱，和细麻都拿了来。
EXOD|35|26|凡有智慧，心里受感动的妇女都来纺山羊毛。
EXOD|35|27|众官长把红玛瑙和宝石，可以镶嵌在以弗得与胸袋上的，都拿了来，
EXOD|35|28|又拿做香，做膏油，和点灯所需的香料和油来。
EXOD|35|29|以色列 人，无论男女，凡心里受感动的，都带甘心祭来献给耶和华，为要做耶和华藉 摩西 所吩咐的一切工。
EXOD|35|30|摩西 对 以色列 人说：“看， 犹大 支派中 户珥 的孙子， 乌利 的儿子 比撒列 ，耶和华已经题名召他，
EXOD|35|31|又以上帝的灵充满他，使他有智慧、聪明、知识，能做各样的工，
EXOD|35|32|能设计图案，用金、银、铜制造各物，
EXOD|35|33|又能雕刻镶嵌用的宝石，雕刻木头，做各样精巧的工。
EXOD|35|34|耶和华又赐给他和 但 支派中， 亚希撒抹 的儿子 亚何利亚伯 能教导人的心。
EXOD|35|35|耶和华使他们的心满有智慧，能做各样的工，无论是雕刻的工，图案设计的工，用蓝色、紫色、朱红色纱，和细麻作刺绣的工，以及编织的工，他们都能胜任，也能设计图案。”
EXOD|36|1|比撒列 和 亚何利亚伯 ，以及一切心里有智慧，蒙耶和华赐智慧和聪明，懂得做圣所各样用途之工的人，都照耶和华所吩咐的去做。
EXOD|36|2|摩西 把 比撒列 和 亚何利亚伯 ，以及那些蒙耶和华赐他心里有智慧，心受感动愿意前来做工的人都召来。
EXOD|36|3|这些人就从 摩西 收了 以色列 人为建造圣所，以及圣所各用途之工而奉献的礼物。每天早晨，百姓继续把甘心祭拿来。
EXOD|36|4|凡有智慧能做圣所一切工的人，都各自离开他们原本的工作前来，
EXOD|36|5|对 摩西 说：“百姓送来的礼物很多，已经超过耶和华吩咐建造之工所需要的了。”
EXOD|36|6|摩西 吩咐，他们就在营中传令说：“无论男女，不必再为圣所的礼物做任何的工。”这样才使百姓停止，不再拿礼物来，
EXOD|36|7|他们所有的材料已经足够整个工程之用，而且有余。
EXOD|36|8|做工的人当中，凡心里有智慧的，用十幅幔子做帐幕，幔子是用搓的细麻和蓝色、紫色、朱红色纱织成的，并且以刺绣的手艺绣上基路伯。
EXOD|36|9|每幅幔子长二十八肘，每幅幔子宽四肘，全部的幔子都是一样的尺寸。
EXOD|36|10|他使这五幅幔子彼此相连，又使那五幅幔子彼此相连。
EXOD|36|11|他在这一组相连幔子的末幅边上缝了蓝色的钮环；在另一组相连幔子的末幅边上也照样做。
EXOD|36|12|他在这幅幔子上缝五十个钮环，在另一组相连幔子的末幅上也缝五十个钮环，环环相对。
EXOD|36|13|他又做了五十个金钩，用钩子使幔子彼此相连，成为一个帐幕。
EXOD|36|14|他用山羊毛织十一幅幔子，作为帐幕上的罩棚。
EXOD|36|15|每幅幔子长三十肘，每幅幔子宽四肘；十一幅幔子都是一样的尺寸。
EXOD|36|16|他把五幅幔子连成一幅，又把六幅幔子连成一幅。
EXOD|36|17|他在这一组相连幔子的末幅边上缝了五十个钮环；在另一组相连幔子的末幅边上也缝了五十个钮环。
EXOD|36|18|他又做五十个铜钩，使罩棚相连成为一个。
EXOD|36|19|他用染红的公羊皮做罩棚的盖，再用精美皮料做外层的盖。
EXOD|36|20|他用金合欢木做竖立帐幕的木板，
EXOD|36|21|木板长十肘，每块板宽一肘半，
EXOD|36|22|每块板有两个榫头可以彼此衔接。帐幕一切的板都是这样做。
EXOD|36|23|他做帐幕的木板：南面，就是面向南方的那一边，做二十块板，
EXOD|36|24|在这二十块板底下做了四十个带卯眼的银座：两个卯眼接连这块板上的两个榫头，另外两个卯眼接连那块板上的两个榫头。
EXOD|36|25|他在帐幕的第二边，就是北面，也做二十块板，
EXOD|36|26|和四十个带卯眼的银座；这块板底下有两个卯眼，那块板底下也有两个卯眼。
EXOD|36|27|他在帐幕的后面，就是西面，做六块板，
EXOD|36|28|在帐幕后面的角落做两块板。
EXOD|36|29|下端的板是成双的，上端连在一起，直到顶端的第一个环子；两块板都是这样，做成两个角落。
EXOD|36|30|一共有八块板和十六个带卯眼的银座，每块板底下有两个卯眼。
EXOD|36|31|他用金合欢木做横木：为帐幕这面的板做五根横木，
EXOD|36|32|为帐幕那面的板做五根横木，又为帐幕后面，就是朝西的板做五根横木，
EXOD|36|33|他做了板腰间的横木，从一头通到另一头。
EXOD|36|34|他将板包上金子，又做板上的金环来套横木；横木也包上金子。
EXOD|36|35|他用蓝色、紫色、朱红色纱，和搓的细麻织幔子，以刺绣的手艺绣上基路伯。
EXOD|36|36|他又用金合欢木为幔子做四根柱子，包上金子，柱子有金钩，又为柱子铸了四个带卯眼的银座。
EXOD|36|37|他用蓝色、紫色、朱红色纱，和搓的细麻，以刺绣的手艺为帐幕织门帘，
EXOD|36|38|又为帘子做五根柱子和柱子的钩子，把柱顶和柱子的箍包上金子。柱子有五个带卯眼的铜座。
EXOD|37|1|比撒列 用金合欢木做一个柜子，长二肘半，宽一肘半，高一肘半。
EXOD|37|2|里里外外包上金子，四围镶上金边。
EXOD|37|3|他又铸了四个金环，安在柜子的四脚上；这边两个环，那边两个环。
EXOD|37|4|他用金合欢木做了两根杠，包上金子，
EXOD|37|5|又把杠穿过柜旁的环，以便抬柜。
EXOD|37|6|他用纯金做了一个柜盖，长二肘半，宽一肘半，
EXOD|37|7|他造两个用金子锤出的基路伯，从柜盖的两端锤出它们。
EXOD|37|8|这端一个基路伯，那端一个基路伯；从柜盖的两端锤出两个基路伯。
EXOD|37|9|二基路伯的翅膀向上张开，用翅膀遮住柜盖，脸彼此相对；基路伯的脸朝向柜盖。
EXOD|37|10|他用金合欢木做了一张供桌，长二肘，宽一肘，高一肘半，
EXOD|37|11|把它包上纯金，四围镶上金边。
EXOD|37|12|供桌的四围各做了一掌宽的边缘，边缘镶上金边。
EXOD|37|13|他又铸了四个金环，把环安在四个桌脚的四角上。
EXOD|37|14|环靠近边缘，以便穿杠抬供桌。
EXOD|37|15|他用金合欢木做了两根杠，包上金子，用来抬供桌。
EXOD|37|16|他又用纯金做了桌上的器具，就是盘、碟，以及浇酒祭的杯和壶。
EXOD|37|17|他造一座用纯金锤出的灯台；灯台的座、干、杯、花萼和花瓣，都和灯台接连一块。
EXOD|37|18|灯台两旁伸出六根枝子：这边三根，那边三根。
EXOD|37|19|这边的枝子上有三个杯，形状像杏花，有花萼有花瓣；那边的枝子上也有三个杯，形状像杏花，有花萼有花瓣。从灯台伸出来的六根枝子都是如此。
EXOD|37|20|灯台本身有四个杯，形状像杏花，有花萼有花瓣。
EXOD|37|21|灯台的第一对枝子下面有花萼，灯台的第二对枝子下面有花萼，灯台的第三对枝子下面也有花萼；灯台伸出的六根枝子都是如此。
EXOD|37|22|花萼和枝子都和灯台接连一块，全是从一块纯金锤出来的。
EXOD|37|23|他用纯金做灯台的七盏灯，以及灯剪和灯盘。
EXOD|37|24|他用一他连得的纯金做灯台和灯台的一切器具。
EXOD|37|25|他用金合欢木做香坛，长一肘，宽一肘，这坛是正方形的，高二肘。坛的四个翘角与坛接连一块。
EXOD|37|26|他把坛的上面与坛的四围，以及坛的四个翘角包上纯金，又在坛的四围镶上金边。
EXOD|37|27|他在坛的两个对侧，金边下面做了两个金环，用来穿杠抬坛。
EXOD|37|28|他又用金合欢木做杠，包上金子。
EXOD|37|29|他按配制香料的方法制成圣膏油和芬芳的纯香。
EXOD|38|1|他用金合欢木做燔祭坛，长五肘，宽五肘，是正方形的，高三肘。
EXOD|38|2|在坛的四角做四个翘角，与坛接连一块，把坛包上铜。
EXOD|38|3|他做坛的一切器具，就是桶子、铲子、盘子、肉叉和火盆；这一切器具都是用铜做的。
EXOD|38|4|他又为坛做一个铜网，安在坛四围的边的下面，垂到坛的半腰。
EXOD|38|5|他在铜网的四角上铸了四个环，用来穿杠。
EXOD|38|6|他用金合欢木做杠，包上铜，
EXOD|38|7|把杠穿过坛两旁的环子，用来抬坛。他用板做坛，坛的中心是空的。
EXOD|38|8|他用铜做洗濯盆和盆座，是用会幕门前事奉之妇人的铜镜做的。
EXOD|38|9|他又做院子，在南面，就是面向南方的那一边，用搓的细麻做院子的帷幔，一百肘。
EXOD|38|10|帷幔有二十根柱子，二十个带卯眼的铜座；柱子的钩和箍都是银的。
EXOD|38|11|北面的帷幔一百肘。帷幔有二十根柱子，二十个带卯眼的铜座；柱子的钩和箍都是银的。
EXOD|38|12|西面的帷幔五十肘。帷幔有十根柱子，十个带卯眼的座；柱子的钩和箍都是银的。
EXOD|38|13|院子的东面，就是面向东方的那一边，五十肘。
EXOD|38|14|一边的帷幔有十五肘，有三根柱子，三个带卯眼的座。
EXOD|38|15|另一边也一样，院子门口左右的帷幔也有十五肘，有三根柱子，三个带卯眼的座。
EXOD|38|16|院子四面的帷幔都是用搓的细麻做的。
EXOD|38|17|柱子带卯眼的座是铜的，柱子的钩和箍是银的，柱顶是用银包的。院子一切的柱子都是用银子箍着的。
EXOD|38|18|院子的门帘是以刺绣的手艺，用蓝色、紫色、朱红色纱，和搓的细麻织的，长二十肘，宽也就是高五肘，与院子帷幔的高度相同。
EXOD|38|19|门帘有四根柱子，四个带卯眼的铜座；柱子上的钩和箍是银的，柱顶是用银包的。
EXOD|38|20|帐幕一切的橛子和院子四围的橛子都是铜的。
EXOD|38|21|这是帐幕，就是法柜帐幕中物件的总数，是照 摩西 的吩咐， 亚伦 祭司的儿子 以他玛 经手， 利未 人数点的。
EXOD|38|22|凡耶和华吩咐 摩西 的，都是由 犹大 支派中 户珥 的孙子， 乌利 的儿子 比撒列 去做的；
EXOD|38|23|与他同工的有 但 支派中 亚希撒抹 的儿子 亚何利亚伯 ；他是雕刻师，也是设计师，又是用蓝色、紫色、朱红色纱，和细麻的刺绣师。
EXOD|38|24|为圣所一切工作用的金子，就是所奉献的金子，按圣所的舍客勒，一共是二十九他连得，七百三十舍客勒。
EXOD|38|25|会中被数的人所献的银子，按圣所的舍客勒，一共是一百他连得，一千七百七十五舍客勒。
EXOD|38|26|凡曾被数的，就是二十岁以上的人，共有六十万三千五百五十人。按圣所的舍客勒，每人半舍客勒，就是一比加。
EXOD|38|27|一百他连得银子是用来铸造圣所带卯眼的座和幔子下带卯眼的座；用一百他连得铸造一百个带卯眼的座，每个带卯眼的座一他连得。
EXOD|38|28|一千七百七十五舍客勒是用来铸造柱子的钩，包柱顶，以及箍着柱子。
EXOD|38|29|所奉献的铜共有七十他连得，二千四百舍客勒。
EXOD|38|30|这些铜是用来做会幕门口带卯眼的座，铜坛、坛的铜网和坛的一切器具，
EXOD|38|31|院子四围带卯眼的座和院子门口带卯眼的座，以及帐幕一切的橛子和院子四围所有的橛子。
EXOD|39|1|他们用蓝色、紫色、朱红色纱缝制精致的礼服，在圣所用以供职；他们为 亚伦 做圣衣，是照耶和华所吩咐 摩西 的。
EXOD|39|2|以弗得是用金色、蓝色、紫色、朱红色纱，和搓的细麻做的。
EXOD|39|3|他们把金子锤成薄片，剪成细线，与蓝色、紫色、朱红色纱，以刺绣的手艺织在一起。
EXOD|39|4|他们又为以弗得做两条相连的肩带，接连在以弗得的两端。
EXOD|39|5|以弗得的精致带子以一样的手艺，用金色、蓝色、紫色、朱红色纱，和搓的细麻缝制，与以弗得接连在一起，是照耶和华所吩咐 摩西 的。
EXOD|39|6|他们琢出两块红玛瑙，镶在金槽里，如同刻印章，刻上 以色列 众子的名字。
EXOD|39|7|他把这两块宝石安在以弗得的两条肩带上，为 以色列 人作纪念石，是照耶和华所吩咐 摩西 的。
EXOD|39|8|胸袋是以刺绣的手艺，如同以弗得的做法，用金色、蓝色、紫色、朱红色纱，和搓的细麻缝制。
EXOD|39|9|胸袋是正方形的，他们把它做成两层，这两层各长一虎口，宽一虎口。
EXOD|39|10|他们在上面镶四行宝石：第一行是红宝石、红璧玺、红玉；
EXOD|39|11|第二行是绿宝石、蓝宝石、金刚石；
EXOD|39|12|第三行是紫玛瑙、白玛瑙、紫晶；
EXOD|39|13|第四行是水苍玉、红玛瑙、碧玉。这些都镶在金槽中。
EXOD|39|14|这些宝石有 以色列 十二个儿子的名字，如同刻印章，每一颗有自己的名字，代表十二个支派。
EXOD|39|15|他们在胸袋上用纯金打链子，像编成的绳子一样。
EXOD|39|16|他们又做了两个金槽和两个金环，把这两个环安在胸袋的两端。
EXOD|39|17|他们把那两条编成的金链系在胸袋两端的两个环上，
EXOD|39|18|又把链子的另外两端扣在两个槽上，安在以弗得前面的肩带上。
EXOD|39|19|他们做了两个金环，安在胸袋的两端，在以弗得里面的边上，
EXOD|39|20|又做两个金环，安在以弗得前面两条肩带的下边，靠近接缝处，在精致带子的上面。
EXOD|39|21|他们用蓝色的带子把胸袋的环与以弗得的环系住，使胸袋绑在以弗得精致的带子上，不致松脱，是照耶和华所吩咐 摩西 的。
EXOD|39|22|以弗得的外袍是以编织的手艺做的，颜色全是蓝的。
EXOD|39|23|袍上方的中间留了一个领口，领口的周围织出领边，好像铠甲的领口，免得破裂。
EXOD|39|24|他们在袍子下摆用蓝色、紫色、朱红色纱，和搓的细麻 做石榴，
EXOD|39|25|又用纯金铸了铃铛，把铃铛钉在石榴中间，袍子下摆周围的石榴中间：
EXOD|39|26|一个铃铛一个石榴，一个铃铛一个石榴，在袍子下摆的周围，用以供职，是照耶和华所吩咐 摩西 的。
EXOD|39|27|他们用编织的工为 亚伦 和他的儿子做细麻布内袍、
EXOD|39|28|细麻布礼冠、细麻布精致头巾，和搓的细麻布裤子，
EXOD|39|29|又用蓝色、紫色、朱红色纱，和搓的细麻，以刺绣的手艺做腰带，是照耶和华所吩咐 摩西 的。
EXOD|39|30|他们用纯金做一面圣冠上的牌，如同刻印章，在上面写着“归耶和华为圣”，
EXOD|39|31|又用蓝色的带子把牌系在礼冠上，是照耶和华所吩咐 摩西 的。
EXOD|39|32|会幕的帐幕一切的工程就这样做完了。凡耶和华所吩咐 摩西 的， 以色列 人都照样做了。
EXOD|39|33|他们把帐幕运到 摩西 那里，帐幕和帐幕的一切器具，就是钩、板、横木、柱子、带卯眼的座，
EXOD|39|34|染红公羊皮的盖、精美皮料的盖、遮掩的幔子，
EXOD|39|35|法柜、柜的杠、柜盖，
EXOD|39|36|供桌、供桌的一切器具、供饼，
EXOD|39|37|纯金的灯台、摆列的灯、灯台的一切器具、点灯的油，
EXOD|39|38|金坛、膏油、芬芳的香、帐幕的门帘，
EXOD|39|39|铜坛、坛的铜网、坛的杠、坛的一切器具，洗濯盆和盆座，
EXOD|39|40|院子的帷幔、柱子、带卯眼的座、院子的门帘、绳子、橛子，帐幕，就是会幕使用的一切器具，
EXOD|39|41|以及圣所事奉用的精致礼服， 亚伦 祭司的圣衣和他儿子的衣服，供祭司职分用。
EXOD|39|42|这一切工作都是 以色列 人照耶和华所吩咐 摩西 做的。
EXOD|39|43|摩西 看见这一切的工，看哪，耶和华怎样吩咐，他们就照样做了， 摩西 就为他们祝福。
EXOD|40|1|耶和华吩咐 摩西 说：
EXOD|40|2|“正月初一，你要立起会幕的帐幕，
EXOD|40|3|把法柜安放在里面，用幔子将柜遮掩。
EXOD|40|4|把供桌搬进去，摆设桌上的器具。又把灯台搬进去，点上灯。
EXOD|40|5|把金香坛安在法柜前，挂上帐幕的门帘。
EXOD|40|6|把燔祭坛安在会幕的帐幕门前。
EXOD|40|7|把洗濯盆安在会幕和坛的中间，在盆里盛水。
EXOD|40|8|又要在院子周围支起帷幔，把院子的门帘挂上。
EXOD|40|9|你要用膏油抹帐幕和其中所有的，使帐幕和一切器具分别为圣，就都成为圣。
EXOD|40|10|又要抹燔祭坛和坛的一切器具，使坛分别为圣，坛就成为至圣。
EXOD|40|11|要抹洗濯盆和盆座，使盆分别为圣。
EXOD|40|12|你要带 亚伦 和他儿子到会幕门口，用水洗身。
EXOD|40|13|要给 亚伦 穿上圣衣，又膏他，使他分别为圣，作事奉我的祭司。
EXOD|40|14|又要带他的儿子来，给他们穿上内袍。
EXOD|40|15|你怎样膏他们的父亲，也要照样膏他们，使他们成为事奉我的祭司。他们受了膏，就必世世代代永远得祭司的职分。”
EXOD|40|16|摩西 这样做了；耶和华怎样吩咐 摩西 ，他就照样做了。
EXOD|40|17|第二年正月初一，帐幕就立起来。
EXOD|40|18|摩西 支起帐幕，安上带卯眼的座，安上板，穿上横木，立起柱子。
EXOD|40|19|他在帐幕的上面搭上罩棚，把罩棚外层的盖子盖在其上，是照着耶和华所吩咐他的。
EXOD|40|20|他把法版放在柜里，把杠穿在柜的两旁，把柜盖安在柜上。
EXOD|40|21|把柜抬进帐幕，挂上遮掩柜的幔子，把法柜遮盖了，是照耶和华所吩咐 摩西 的。
EXOD|40|22|他把供桌安在会幕内，在帐幕的北边，幔子的外面。
EXOD|40|23|把饼摆设在供桌上，在耶和华面前，是照耶和华所吩咐 摩西 的。
EXOD|40|24|他把灯台安在会幕内，在帐幕的南边，供桌的对面，
EXOD|40|25|并在耶和华面前点灯，是照耶和华所吩咐 摩西 的。
EXOD|40|26|他把金坛安在会幕内，幔子的前面，
EXOD|40|27|又在坛上烧芬芳的香，是照耶和华所吩咐 摩西 的。
EXOD|40|28|他又挂上帐幕的门帘。
EXOD|40|29|在会幕的帐幕门口安设燔祭坛，把燔祭和素祭献在坛上，是照耶和华所吩咐 摩西 的。
EXOD|40|30|他又把洗濯盆安在会幕和祭坛的中间，盆里盛水，以便洗濯。
EXOD|40|31|摩西 和 亚伦 ，以及 亚伦 的儿子用这盆洗手洗脚。
EXOD|40|32|他们进会幕或走近坛的时候，就都洗濯，是照耶和华所吩咐 摩西 的。
EXOD|40|33|他在帐幕和祭坛的四围支起院子的帷幔，把院子的门帘挂上。这样， 摩西 就做完了工。
EXOD|40|34|那时，云彩遮盖会幕，耶和华的荣光充满了帐幕。
EXOD|40|35|摩西 不能进会幕，因为云彩停在其上，耶和华的荣光充满了帐幕。
EXOD|40|36|每逢云彩从帐幕升上去， 以色列 人就起程前行；
EXOD|40|37|云彩若不升上去，他们就不起程，直等到云彩升上去。
EXOD|40|38|在他们所行的路上，在 以色列 全家的眼前，白天，耶和华的云彩在帐幕上，黑夜，有火在云彩中。
LEV|1|1|耶和华从会幕中呼叫 摩西 ，吩咐他说：
LEV|1|2|“你要吩咐 以色列 人，对他们说：你们中间若有人要献供物给耶和华，可以从牛群羊群中献牲畜为供物。
LEV|1|3|“他的供物若以牛为燔祭，要献一头没有残疾的公牛，献在会幕的门口，他就可以在耶和华面前蒙悦纳。
LEV|1|4|他要按手在燔祭牲的头上，为自己赎罪，就蒙悦纳。
LEV|1|5|他要在耶和华面前宰公牛犊； 亚伦 子孙作祭司的要献上血，把血洒在会幕门口坛的周围。
LEV|1|6|他要剥去燔祭牲的皮，把燔祭牲切成块。
LEV|1|7|亚伦 祭司的子孙要在坛上生火，把柴摆在火上。
LEV|1|8|亚伦 子孙作祭司的要把肉块连头和脂肪，摆在坛上烧着火的柴上。
LEV|1|9|燔祭牲的内脏与小腿要用水洗净，祭司要把整只全烧在坛上，当作燔祭，是献给耶和华为馨香的火祭。
LEV|1|10|“人的供物若以绵羊或山羊为燔祭，要献一只没有残疾的公羊。
LEV|1|11|他要在坛的北边，在耶和华面前宰羊； 亚伦 子孙作祭司的要把血洒在坛的周围。
LEV|1|12|他要把燔祭牲切成块，祭司就要把肉块连头和脂肪，摆在坛上烧着火的柴上。
LEV|1|13|内脏与小腿要用水洗净，祭司要把整只献上，全烧在坛上。这是燔祭，是献给耶和华为馨香的火祭。
LEV|1|14|“人献给耶和华的供物若以鸟为燔祭，就要献斑鸠或雏鸽为他的供物。
LEV|1|15|祭司要把鸟拿到坛前，扭断它的头，把鸟烧在坛上，鸟的血要流在坛的旁边；
LEV|1|16|又要把鸟的嗉囊和里面的脏物 除掉，丢在坛东边倒灰的地方。
LEV|1|17|他要拿着鸟的两个翅膀，把鸟撕开，却不可撕断；祭司要把它摆在坛上烧着火的柴上焚烧。这是燔祭，是献给耶和华为馨香的火祭。”
LEV|2|1|“若有人献素祭为供物给耶和华，就要献细面为供物，把油浇在上面，加上乳香，
LEV|2|2|带到 亚伦 子孙作祭司的那里。祭司要从细面中取出满满的一把，又取些油和所有的乳香，把这些作为纪念的烧在坛上，是献给耶和华为馨香的火祭。
LEV|2|3|素祭所剩的要归给 亚伦 和他的子孙；在献给耶和华的火祭中，这是至圣的。
LEV|2|4|“若献炉中烤的素祭为供物，要用调了油的无酵细面饼，或抹了油的无酵薄饼。
LEV|2|5|若以铁盘上的素祭为供物，就要用调了油的无酵细面，
LEV|2|6|分成小块，浇上油；这是素祭。
LEV|2|7|若以煎锅煎的素祭为供物，就要用油与细面做成。
LEV|2|8|要把这样做成的素祭带到耶和华面前，拿给祭司，祭司要带到坛前。
LEV|2|9|祭司要从素祭中取出作为纪念的烧在坛上，是献给耶和华为馨香的火祭。
LEV|2|10|素祭所剩的要归给 亚伦 和他的子孙；在献给耶和华的火祭中，这是至圣的。
LEV|2|11|“凡献给耶和华的素祭都不可以有酵，因为你们不可把任何的酵或蜜烧了，当作火祭献给耶和华。
LEV|2|12|你们可以把这些献给耶和华当作初熟的供物，但是不可献在坛上作为馨香的祭。
LEV|2|13|凡献为素祭的供物都要用盐调和；在素祭中，不可缺少你与上帝立约的盐。一切的供物都要加盐献上。
LEV|2|14|“你若献初熟之物给耶和华为素祭，就要献在火中烘过的新麦穗，就是磨碎的新谷物，当作初熟之物的素祭。
LEV|2|15|你要加上油和乳香；这是素祭。
LEV|2|16|祭司要把供物中作为纪念的，就是一些磨碎的新谷物和一些油，以及所有的乳香，都焚烧，是献给耶和华的火祭。”
LEV|3|1|“人献平安祭为供物，若是从牛群中献，无论是公的母的，要用没有残疾的，献在耶和华面前。
LEV|3|2|他要按手在供物的头上，在会幕的门口宰了它。 亚伦 子孙作祭司的，要把血洒在坛的周围。
LEV|3|3|从平安祭中，他要把火祭献给耶和华，就是包着内脏的脂肪和内脏上所有的脂肪，
LEV|3|4|两个肾和肾上的脂肪，即靠近肾两旁的脂肪，以及肝上的网油，连同肾一起取下。
LEV|3|5|亚伦 的子孙要把这些摆在烧着火的柴上，烧在坛的燔祭上，是献给耶和华为馨香的火祭。
LEV|3|6|“人向耶和华献平安祭为供物，若是从羊群中献，无论是公的母的，要用没有残疾的。
LEV|3|7|若他献一只绵羊为供物，就要把它献在耶和华面前。
LEV|3|8|要按手在供物的头上，在会幕前宰了它。 亚伦 的子孙要把血洒在坛的周围。
LEV|3|9|从平安祭中，他要取脂肪当作火祭献给耶和华，就是靠近脊骨处取下的整条肥尾巴，包着内脏的脂肪和内脏上所有的脂肪，
LEV|3|10|两个肾和肾上的脂肪，即靠近肾两旁的脂肪，以及肝上的网油，连同肾一起取下。
LEV|3|11|祭司要把这些烧在坛上，是献给耶和华为食物的火祭。
LEV|3|12|“人的供物若是山羊，就要把它献在耶和华面前。
LEV|3|13|要按手在它的头上，在会幕前宰了它。 亚伦 的子孙要把血洒在坛的周围，
LEV|3|14|又要从供物中把火祭献给耶和华，就是包着内脏的脂肪和内脏上所有的脂肪，
LEV|3|15|两个肾和肾上的脂肪，即靠近肾两旁的脂肪，以及肝上的网油，连同肾一起取下。
LEV|3|16|祭司要把这些烧在坛上，作为馨香火祭的食物；所有的脂肪都是耶和华的。
LEV|3|17|在你们一切的住处，脂肪和血都不可吃，这要成为你们世世代代永远的定例。”
LEV|4|1|耶和华吩咐 摩西 说：
LEV|4|2|“你要吩咐 以色列 人说：若有人无意中犯罪，在任何事上犯了一条耶和华所吩咐的禁令，
LEV|4|3|或是受膏的祭司犯了罪，使百姓陷在罪里，他就当为自己所犯的罪，把没有残疾的公牛犊献给耶和华为赎罪祭。
LEV|4|4|他要把公牛牵到会幕的门口，在耶和华面前按手在牛的头上，把牛宰于耶和华面前。
LEV|4|5|受膏的祭司要取些公牛的血，带到会幕那里。
LEV|4|6|祭司要把手指蘸在血中，在耶和华面前对着圣所的幔子弹血七次，
LEV|4|7|又要把一些血抹在会幕内，耶和华面前香坛的四个翘角上，再把公牛其余的血全倒在会幕门口燔祭坛的底座上；
LEV|4|8|又要取出这头赎罪祭公牛所有的脂肪，就是包着内脏的脂肪和内脏上所有的脂肪，
LEV|4|9|两个肾和肾上的脂肪，即靠近肾两旁的脂肪，以及肝上的网油，连同肾一起取下，
LEV|4|10|正如从平安祭的牛身上所取的，祭司要把这些烧在燔祭坛上。
LEV|4|11|但公牛的皮和所有的肉，以及头、腿、内脏、粪，
LEV|4|12|就是全公牛，要搬到营外清洁的地方倒灰之处，放在柴上用火焚烧。
LEV|4|13|“ 以色列 全会众若犯了错，在任何事上犯了一条耶和华所吩咐的禁令，而有了罪，会众看不出这隐藏的事；
LEV|4|14|他们一知道犯了罪，就要献一头公牛犊为赎罪祭，牵它到会幕前。
LEV|4|15|会众的长老要在耶和华面前按手在公牛的头上，把牛宰于耶和华面前。
LEV|4|16|受膏的祭司要取些公牛的血，带到会幕那里。
LEV|4|17|祭司要用手指蘸一些血，在耶和华面前对着幔子弹七次，
LEV|4|18|又要把一些血抹在会幕内，耶和华面前坛的四个翘角上，再把其余的血全倒在会幕门口燔祭坛的底座上。
LEV|4|19|他要取出公牛所有的脂肪，烧在坛上。
LEV|4|20|他要处理这牛，正如处理那头赎罪祭的公牛一样，他要如此去做。祭司要为他们赎罪，他们就蒙赦免。
LEV|4|21|他要把牛搬到营外烧了，像烧前一头公牛一样；这是会众的赎罪祭。
LEV|4|22|“官长若犯罪，在任何事上无意中犯了一条耶和华－他的上帝所吩咐的禁令，而有了罪，
LEV|4|23|他一知道自己犯了罪，就要牵一只没有残疾的公山羊为供物。
LEV|4|24|他要按手在羊的头上，在耶和华面前宰燔祭牲的地方把它宰了；这是赎罪祭。
LEV|4|25|祭司要用手指蘸一些赎罪祭牲的血，抹在燔祭坛的四个翘角上，再把其余的血倒在燔祭坛的底座上。
LEV|4|26|祭牲所有的脂肪都要烧在坛上，正如平安祭的脂肪一样。祭司要为他的罪赎了他，他就蒙赦免。
LEV|4|27|“这地的百姓若有人无意中犯罪，在任何事上犯了一条耶和华所吩咐的禁令，而有了罪，
LEV|4|28|他一知道自己犯了罪，就要为所犯的罪牵一只没有残疾的母山羊为供物。
LEV|4|29|他要按手在赎罪祭牲的头上，在燔祭牲的地方把它宰了。
LEV|4|30|祭司要用手指蘸一些祭牲的血，抹在燔祭坛的四个翘角上，再把其余的血全倒在坛的底座上；
LEV|4|31|又要把祭牲所有的脂肪都取下，正如取平安祭牲的脂肪一样。祭司要把脂肪烧在坛上，在耶和华面前作为馨香的祭。祭司要为他赎罪，他就蒙赦免。
LEV|4|32|“人若牵一只绵羊为赎罪祭作供物，就要牵一只没有残疾的母羊。
LEV|4|33|他要按手在赎罪祭牲的头上，在宰燔祭牲的地方宰了它，作为赎罪祭。
LEV|4|34|祭司要用手指蘸一些赎罪祭牲的血，抹在燔祭坛的四个翘角上，再把其余的血全倒在坛的底座上；
LEV|4|35|又要把祭牲所有的脂肪都取下，正如取平安祭的羊的脂肪一样。祭司要按献给耶和华火祭的条例，把脂肪烧在坛上。祭司要为他所犯的罪赎了他，他就蒙赦免。”
LEV|5|1|“若有人犯了罪，就是听见了誓言，他本来可以作证，却不把所看见、所知道的说出来，必须担当他的罪孽。
LEV|5|2|若有人摸了任何不洁之物，无论是野兽的不洁尸体，家畜的不洁尸体，或是群聚动物的不洁尸体，他虽不察觉，也是不洁净，就有罪了。
LEV|5|3|或是他摸了人的不洁之物，就是任何使人成为不洁的不洁之物，他虽不察觉，但一知道，就有罪了。
LEV|5|4|若有人随口发誓，或出于恶意，或出于善意，这人无论在什么事上随意发誓，虽不察觉，但一知道，就在这其中的一件事上有罪了。
LEV|5|5|当他在这其中的一件事上有罪的时候，就要承认所犯的罪，
LEV|5|6|并要为所犯的罪，把他的赎愆祭牲，就是羊群中的一只母绵羊或母山羊，献给耶和华为赎罪祭，祭司要为他的罪赎了他。
LEV|5|7|“若他的力量不够献一只绵羊，就要为所犯的罪，把两只斑鸠或是两只雏鸽献给耶和华为赎愆祭：一只作赎罪祭，一只作燔祭。
LEV|5|8|他要把这些带到祭司那里，祭司就先把赎罪祭献上，从鸟的颈项上扭断它的头，但不把鸟撕断。
LEV|5|9|祭司要把一些赎罪祭牲的血弹在祭坛的边上，其余的血要倒在坛的底座上；这是赎罪祭。
LEV|5|10|他要依照条例献第二只鸟为燔祭。祭司要为他所犯的罪赎了他，他就蒙赦免。
LEV|5|11|“他的力量若不够献两只斑鸠或两只雏鸽，就要为所犯的罪把供物，就是十分之一伊法细面，献上为赎罪祭；不可加上油，也不可加上乳香，因为这是赎罪祭。
LEV|5|12|他要把细面带到祭司那里，祭司要取出满满的一把，作为纪念，按照献火祭给耶和华的条例把它烧在坛上；这是赎罪祭。
LEV|5|13|至于他在这几件事中所犯的任何罪，祭司要为他赎了，他就蒙赦免。剩下的都归给祭司，和素祭一样。”
LEV|5|14|耶和华吩咐 摩西 说：
LEV|5|15|“若有人在耶和华的圣物上无意中犯了罪，有了过犯，就要献羊群中一只没有残疾的公绵羊给耶和华为赎愆祭，或依圣所的舍客勒所估定的银子，作为赎愆祭。
LEV|5|16|他要为在圣物上的疏忽赔偿，另外加五分之一，把这些都交给祭司。祭司要用赎愆祭的公绵羊为他赎罪，他就蒙赦免。
LEV|5|17|“若有人犯罪，在任何事上犯了一条耶和华所吩咐的禁令，他虽不察觉，仍算有罪，必须担当自己的罪孽。
LEV|5|18|他要牵羊群中一只没有残疾的公绵羊，或照你所估定的价值，给祭司作赎愆祭。祭司要为他赎他因不知道而无意中所犯的罪，他就蒙赦免。
LEV|5|19|这是赎愆祭；因他确实得罪了耶和华。”
LEV|6|1|耶和华吩咐 摩西 说：
LEV|6|2|“若有人犯罪，得罪了耶和华，就是在邻舍寄托他的东西或抵押品上行诡诈，或抢夺，或欺压邻舍，
LEV|6|3|或是捡了失物行了诡诈，起了假誓，在人所做的任何事上犯了罪；
LEV|6|4|他既犯了罪，有了过犯，就要归还他所抢夺的，或是因欺压所得的，或是别人寄托他的，或是他所捡到的失物，
LEV|6|5|或是起假誓得来的任何东西，就要全数归还，另外再加五分之一。在查出他有罪的日子，就要立刻赔还给原主。
LEV|6|6|他要献羊群中一只没有残疾的公绵羊，给耶和华为赎愆祭，或照你所估定的价值，给祭司 作赎愆祭。
LEV|6|7|祭司要在耶和华面前为他赎罪；他无论做了什么事，以致有了罪，都必蒙赦免。”
LEV|6|8|耶和华吩咐 摩西 说：
LEV|6|9|“你要吩咐 亚伦 和他的子孙说，燔祭的条例是这样：燔祭要放在坛的底盘上，从晚上到天亮，坛上的火要不断地烧着。
LEV|6|10|祭司要穿上细麻布衣服，又要把细麻布裤子穿在身上，把在坛上烧剩的燔祭灰收起来，放在坛的旁边。
LEV|6|11|然后，他要脱去这衣服，穿上别的衣服，把灰拿到营外洁净之处。
LEV|6|12|坛上的火要不断地烧着，不可熄灭。每日早晨，祭司要在坛上烧柴，把燔祭摆在坛上，并烧平安祭牲的脂肪。
LEV|6|13|坛上的火要不断地烧着，不可熄灭。”
LEV|6|14|“素祭的条例是这样： 亚伦 的子孙要在坛前把这祭献在耶和华面前。
LEV|6|15|祭司要从素祭中的细面取出一把，再取些油和素祭上所有的乳香，把这些作为纪念的烧在坛上，是献给耶和华为馨香的祭。
LEV|6|16|亚伦 和他子孙要吃素祭剩下的；要在圣处吃这无酵饼，在会幕的院子里吃。
LEV|6|17|烤饼不可加酵。这是从献给我的火祭中归给他们的一份；如赎罪祭和赎愆祭一样，这份是至圣的。
LEV|6|18|亚伦 子孙中的男丁都要吃，因为这是你们世世代代从献给耶和华的火祭中，他们永远应得的份。凡摸这些祭物的都要成为圣。”
LEV|6|19|耶和华吩咐 摩西 说：
LEV|6|20|“这是 亚伦 受膏的日子，他和他的子孙所要献给耶和华的供物：十分之一伊法细面，如他们经常献的素祭，早晨一半，晚上一半。
LEV|6|21|要在铁盘上用油调和，调匀后，就拿去烤。素祭烤熟了要分成小块，作为献给耶和华馨香的祭。
LEV|6|22|亚伦 子孙中接续他受膏为祭司的，要把这素祭献上，全烧给耶和华。这是永远的定例。
LEV|6|23|祭司一切的素祭要全部烧了，不可以吃。”
LEV|6|24|耶和华吩咐 摩西 说：
LEV|6|25|“你要吩咐 亚伦 和他的子孙说，赎罪祭的条例是这样：要在耶和华面前宰燔祭牲的地方宰赎罪祭牲；这是至圣的。
LEV|6|26|献赎罪祭的祭司要吃这祭物；要在圣处，就是在会幕的院子里吃。
LEV|6|27|凡摸这祭肉的都要成为圣；这祭牲的血若溅在衣服上，你要在圣处洗净那溅到血的衣服 。
LEV|6|28|煮这祭物的瓦器要打碎；若祭物是在铜器里煮，要把这铜器擦净，用水冲洗。
LEV|6|29|祭司中所有的男丁都可以吃；这是至圣的。
LEV|6|30|若将任何赎罪祭的血带进会幕，为要在圣所赎罪，那肉就不可吃，要用火焚烧。”
LEV|7|1|“赎愆祭的条例是这样：这祭是至圣的。
LEV|7|2|人在哪里宰燔祭牲，也要在哪里宰赎愆祭牲；其血，祭司要洒在坛的周围。
LEV|7|3|祭司要献上它所有的脂肪，把肥尾巴和包着内脏的脂肪，
LEV|7|4|两个肾和肾上的脂肪，即靠近肾两旁的脂肪，以及肝上的网油，连同肾一起取下。
LEV|7|5|祭司要把这些烧在坛上，献给耶和华为火祭，作为赎愆祭。
LEV|7|6|祭司中所有的男丁都可以吃这祭物，要在圣处吃；这是至圣的。
LEV|7|7|赎罪祭怎样，赎愆祭也是怎样，都有一样的条例，用赎愆祭赎罪的祭司要得这祭物。
LEV|7|8|献燔祭的祭司，无论为谁献，所献燔祭牲的皮要归给那祭司，那是他的。
LEV|7|9|任何素祭，无论是在炉中烤的，用煎锅或铁盘做成的，都要归给献祭的祭司。
LEV|7|10|任何素祭，无论是用油调和的，是干的，都要归 亚伦 的子孙，大家均分。”
LEV|7|11|“献给耶和华平安祭的条例是这样：
LEV|7|12|若有人为感谢献祭，就要把用油调和的无酵饼、抹了油的无酵薄饼，和用油调匀细面做成的饼，与感谢祭一同献上。
LEV|7|13|要用有酵的饼，和那为感谢而献的平安祭，与供物一同献上。
LEV|7|14|他要从每一种供物中拿一个饼，献给耶和华为举祭，是要归给那洒平安祭牲血的祭司。
LEV|7|15|为感谢而献的平安祭的肉，要在献祭当天吃，一点也不可留到早晨。
LEV|7|16|若所献的是还愿祭或甘心祭，要在献祭当天吃，剩下的，第二天也可以吃。
LEV|7|17|第三天，所剩下的祭肉要用火焚烧。
LEV|7|18|第三天若吃平安祭的肉，必不蒙悦纳，所献的也不算为祭；这祭物是不洁净的，凡吃这祭物的，必担当自己的罪孽。
LEV|7|19|“沾了不洁净之物的肉就不可吃，要用火焚烧。至于其他的肉，凡洁净的人都可以吃这肉；
LEV|7|20|但不洁净的人若吃了献给耶和华平安祭的肉，这人必从民中剪除。
LEV|7|21|若有人摸了不洁之物，无论是人体的不洁净，或是不洁的牲畜，或是不洁的可憎之物 ，再吃了献给耶和华平安祭的肉，这人必从民中剪除。”
LEV|7|22|耶和华吩咐 摩西 说：
LEV|7|23|“你要吩咐 以色列 人说：牛、绵羊、山羊的脂肪，你们都不可吃。
LEV|7|24|自然死去的或被野兽撕裂的，那脂肪可以作别的用途，你们却万不可吃。
LEV|7|25|任何人吃了献给耶和华作火祭祭牲的脂肪，这人必从民中剪除。
LEV|7|26|在你们一切的住处，无论是鸟或兽的血，你们都不可吃。
LEV|7|27|无论谁吃了血，这人必从民中剪除。”
LEV|7|28|耶和华吩咐 摩西 说：
LEV|7|29|“你要吩咐 以色列 人说：献平安祭给耶和华的，要从他的平安祭中取些供物来献给耶和华。
LEV|7|30|他要亲手把献给耶和华的火祭带来，要把脂肪和胸带来，把胸在耶和华面前摇一摇，作为摇祭。
LEV|7|31|祭司要把脂肪烧在坛上，但胸要归给 亚伦 和他的子孙。
LEV|7|32|你们要从平安祭牲中把右腿作为举祭，送给祭司。
LEV|7|33|亚伦 子孙中献平安祭牲的血和脂肪的，要得这右腿，作为他当得的份。
LEV|7|34|因为我从 以色列 人的平安祭中，把这摇祭的胸和这举祭的腿给 亚伦 祭司和他子孙，作为他们在 以色列 人中永远当得的份。”
LEV|7|35|这是从耶和华的火祭中取出，作为 亚伦 和他子孙受膏的份，就是 摩西 叫他们前来，给耶和华供祭司职分的那一天开始的。
LEV|7|36|这是在 摩西 膏他们的日子，耶和华吩咐给他们的，作为他们在 以色列 人中世世代代永远当得的份。
LEV|7|37|这就是燔祭、素祭、赎罪祭、赎愆祭、圣职礼和平安祭的条例，
LEV|7|38|都是耶和华在 西奈山 上吩咐 摩西 的，也是他在 西奈 旷野吩咐 以色列 人献供物给耶和华的日子所说的。
LEV|8|1|耶和华吩咐 摩西 说：
LEV|8|2|“你领 亚伦 和他儿子前来，并将圣衣、膏油，与赎罪祭的一头公牛、两只公绵羊、一筐无酵饼都一同带来；
LEV|8|3|又要召集全会众到会幕的门口。”
LEV|8|4|摩西 就遵照耶和华的吩咐做了，于是会众聚集在会幕的门口。
LEV|8|5|摩西 对会众说：“这是耶和华所吩咐当做的事。”
LEV|8|6|摩西 领了 亚伦 和他儿子前来，用水洗他们。
LEV|8|7|他给 亚伦 穿上内袍，束上腰带，套上外袍，加上以弗得，再束上精致的带子，把以弗得系在他身上。
LEV|8|8|他又给 亚伦 戴上胸袋，把乌陵和土明放在胸袋内。
LEV|8|9|他把礼冠戴在 亚伦 的头上，礼冠前面安上金牌，成为圣冕，是照耶和华所吩咐 摩西 的。
LEV|8|10|摩西 用膏油抹帐幕和其中所有的，使它们成为圣。
LEV|8|11|他又用膏油在祭坛上弹了七次，抹了坛和坛的一切器皿，以及洗濯盆和盆座，使它们成为圣。
LEV|8|12|他把膏油倒在 亚伦 的头上膏他，使他成为圣。
LEV|8|13|摩西 带了 亚伦 的儿子来，给他们穿上内袍，束上腰带，裹上头巾，是照耶和华所吩咐 摩西 的。
LEV|8|14|他把赎罪祭的公牛牵来， 亚伦 和他儿子按手在赎罪祭公牛的头上，
LEV|8|15|就宰了公牛。 摩西 取了血，用指头抹在祭坛周围的四个翘角上，使坛洁净，再把其余的血倒在坛的底座上，使坛成为圣，为坛赎罪。
LEV|8|16|摩西 把内脏所有的脂肪和肝上的网油，以及两个肾与肾上的脂肪取出，都烧在坛上。
LEV|8|17|至于公牛，连皮带肉和粪，他都用火烧在营外，是照耶和华所吩咐 摩西 的。
LEV|8|18|他把燔祭的公绵羊牵来， 亚伦 和他儿子按手在羊的头上，
LEV|8|19|就宰了公羊。 摩西 把血洒在祭坛的周围，
LEV|8|20|把羊切成块，把头和肉块，以及脂肪拿去烧，
LEV|8|21|他用水洗了内脏和腿之后，就把全羊烧在坛上，作为馨香的燔祭，是献给耶和华的火祭，都是照耶和华所吩咐 摩西 的。
LEV|8|22|他又牵来第二只公绵羊，就是圣职礼的羊， 亚伦 和他儿子按手在羊的头上，
LEV|8|23|就宰了羊。 摩西 把一些血抹在 亚伦 的右耳垂上，右手的大拇指上和右脚的大脚趾上。
LEV|8|24|他领了 亚伦 的儿子来，把一些血抹在他们的右耳垂上，右手的大拇指上和右脚的大脚趾上。 摩西 把其余的血洒在坛的周围。
LEV|8|25|他把脂肪，肥尾巴、内脏所有的脂肪、肝上的网油、两个肾、肾上的脂肪，和右腿取下，
LEV|8|26|再从耶和华面前那装无酵饼的篮子中取一个无酵饼、一个油饼和一个薄饼，把这些放在脂肪和右腿上。
LEV|8|27|他把这一切放在 亚伦 和他儿子的手上，在耶和华面前摇一摇，作为摇祭。
LEV|8|28|摩西 从他们的手上把这些祭物拿来，放在坛的燔祭上烧，这就是圣职礼中献给耶和华馨香的火祭。
LEV|8|29|摩西 拿羊的胸，在耶和华面前摇一摇，作为摇祭，这是圣职礼的羊归给 摩西 的一份，是照耶和华所吩咐 摩西 的。
LEV|8|30|摩西 取些膏油和坛上的血，弹在 亚伦 和他的衣服上，以及他儿子和他们的衣服上，使 亚伦 和他的衣服，他儿子和他们的衣服都成为圣。
LEV|8|31|摩西 对 亚伦 和他儿子说：“你们要在会幕的门口把肉煮了，在那里吃这肉和圣职礼中篮子里的饼，按我所吩咐的说：‘这是 亚伦 和他儿子当吃的。’
LEV|8|32|剩下的肉和饼，你们要用火焚烧。
LEV|8|33|这七天，你们不可走出会幕的门口，直等到你们圣职礼的日子满了，因为授予你们圣职需要七天 。
LEV|8|34|今天所做的，都是耶和华吩咐要做的，好为你们赎罪。
LEV|8|35|这七天，你们要昼夜留在会幕门内，遵守耶和华所吩咐的，免得你们死亡，因为所吩咐我的就是这样。”
LEV|8|36|于是， 亚伦 和他的儿子就做了耶和华藉着 摩西 所吩咐的一切事。
LEV|9|1|到了第八天， 摩西 召 亚伦 和他儿子，以及 以色列 的众长老来，
LEV|9|2|对 亚伦 说：“你当取一头公牛犊作赎罪祭，一只公绵羊作燔祭，都要没有残疾的，献在耶和华面前。
LEV|9|3|你要对 以色列 人说：‘你们当取一只公山羊作赎罪祭，再取一头牛犊和一只小绵羊，都要一岁没有残疾的，作燔祭；
LEV|9|4|又当取一头公牛，一只公绵羊作平安祭，宰杀献在耶和华面前，再加上调油的素祭。因为今天耶和华要向你们显现。’”
LEV|9|5|于是，他们把 摩西 所吩咐的带到会幕前；全会众都近前来，站在耶和华面前。
LEV|9|6|摩西 说：“这是耶和华吩咐你们当做的事，耶和华的荣光要向你们显现。”
LEV|9|7|摩西 对 亚伦 说：“你靠近祭坛前，献你的赎罪祭和燔祭，为自己与百姓赎罪，再献上百姓的供物，为他们赎罪，都是照耶和华所吩咐的。”
LEV|9|8|于是， 亚伦 靠近坛前，宰了那头为自己赎罪的牛犊。
LEV|9|9|亚伦 的儿子把血递给他，他就把指头蘸在血中，抹在坛的四个翘角上，再把其余的血倒在坛的底座上。
LEV|9|10|他把赎罪祭的脂肪和肾，以及肝上的网油，烧在坛上，是照耶和华所吩咐 摩西 的。
LEV|9|11|他用火将肉和皮烧在营外。
LEV|9|12|亚伦 把燔祭牲宰了，他儿子把血递给他，他就把血洒在坛的周围。
LEV|9|13|他们又把燔祭一块一块地，连头递给他，他就烧在坛上。
LEV|9|14|他又洗了内脏和腿，放在坛的燔祭上烧。
LEV|9|15|然后，他奉上百姓的供物。他牵来给百姓作赎罪祭的公山羊，把它宰了，献为赎罪祭，和先前的一样。
LEV|9|16|他也奉上燔祭，按照条例献上。
LEV|9|17|除了早晨的燔祭以外，他又献上素祭，用手取了满满的一把，烧在坛上。
LEV|9|18|亚伦 宰了那给百姓作平安祭的公牛和公绵羊，他儿子把血递给他，他就把血洒在坛的周围；
LEV|9|19|他们把公牛和公绵羊的脂肪、肥尾巴，包着内脏的脂肪，肾和肝上的网油，都递给他。
LEV|9|20|他们把脂肪放在祭牲的胸上，他就把脂肪烧在坛上。
LEV|9|21|亚伦 把祭牲的胸和右腿在耶和华面前摇一摇，作为摇祭，是照 摩西 所吩咐的。
LEV|9|22|亚伦 向百姓举手，为他们祝福。他献了赎罪祭、燔祭、平安祭就下来了。
LEV|9|23|摩西 和 亚伦 进了会幕。他们出来，为百姓祝福；耶和华的荣光向全体百姓显现。
LEV|9|24|有火从耶和华面前出来，焚烧了坛上的燔祭和脂肪；全体百姓一看见，就都欢呼，脸伏于地。
LEV|10|1|亚伦 的儿子 拿答 和 亚比户 各拿着自己的香炉，把火放在炉里，加上香，在耶和华面前献上凡火，是耶和华没有吩咐他们的。
LEV|10|2|有火从耶和华面前出来，把他们吞灭，他们就死在耶和华面前。
LEV|10|3|于是， 摩西 对 亚伦 说：“这就是耶和华所吩咐的，说：‘我在那亲近我的人中要显为圣；在全体百姓面前，我要得着荣耀。’” 亚伦 就默默不言。
LEV|10|4|摩西 召 亚伦 的叔父 乌薛 的儿子 米沙利 和 以利撒反 前来，对他们说：“过来，把你们的亲属从圣所前抬到营外。”
LEV|10|5|于是，二人过来把尸体连袍子一起抬到营外，是照 摩西 所吩咐的。
LEV|10|6|摩西 对 亚伦 和他儿子 以利亚撒 和 以他玛 说：“不可蓬头散发，也不可撕裂衣服，免得你们死亡，免得耶和华向全会众发怒。但你们的弟兄 以色列 全家却要为耶和华发出的火哀哭。
LEV|10|7|你们也不可出会幕的门口，免得你们死亡，因为耶和华的膏油在你们身上。”他们就遵照 摩西 的话去做了。
LEV|10|8|耶和华吩咐 亚伦 说：
LEV|10|9|“你和你儿子进会幕的时候，清酒烈酒都不可喝，免得你们死亡，这要作你们世世代代永远的定例。
LEV|10|10|你们必须分辨圣的俗的，洁净的和不洁净的，
LEV|10|11|也要将耶和华藉 摩西 吩咐 以色列 人的一切律例教导他们。”
LEV|10|12|摩西 对 亚伦 和他剩下的儿子 以利亚撒 和 以他玛 说：“献给耶和华的火祭中所剩下的素祭，你们要拿来，在祭坛旁吃这无酵饼，因为它是至圣的。
LEV|10|13|你们要在圣处吃，因为在献给耶和华的火祭中，这是你和你儿子当得的份；所吩咐我的就是这样。
LEV|10|14|这摇祭的胸和这举祭的腿，你要在洁净的地方和你的儿女一同吃，因为这些是从 以色列 人的平安祭中归给你，作为你和你儿子当得的份。
LEV|10|15|他们要把举祭的腿、摇祭的胸和火祭的脂肪一同带来，在耶和华面前摇一摇，作为摇祭。这些要归给你和你儿子，作永远当得的份，都是照耶和华所吩咐的。”
LEV|10|16|那时， 摩西 急切地寻找那只赎罪祭的公山羊，看哪，它已经烧掉了。他向 亚伦 剩下的儿子 以利亚撒 和 以他玛 发怒，说：
LEV|10|17|“你们为何没有在圣所吃这赎罪祭呢？它是至圣的，是耶和华给你们的，为了除掉会众的罪孽，在耶和华面前为他们赎罪。
LEV|10|18|看哪，这祭牲的血没有拿到圣所里去！你们应当照我所吩咐的，在圣所里吃这祭肉。”
LEV|10|19|亚伦 对 摩西 说：“看哪，他们今天在耶和华面前献上赎罪祭和燔祭，但是我却遭遇这样的灾难。我若今天吃这赎罪祭，耶和华岂能看为美呢？”
LEV|10|20|摩西 听了，就看为美。
LEV|11|1|耶和华吩咐 摩西 和 亚伦 ，对他们说：
LEV|11|2|“你们要吩咐 以色列 人说，地上一切的走兽中可吃的动物是这些：
LEV|11|3|凡蹄分两瓣，分趾蹄而又反刍食物的走兽，你们都可以吃。
LEV|11|4|但那反刍或分蹄之中不可吃的是：骆驼，反刍却不分蹄，对你们是不洁净的；
LEV|11|5|石獾，反刍却不分蹄，对你们是不洁净的；
LEV|11|6|兔子，反刍却不分蹄，对你们是不洁净的；
LEV|11|7|猪，蹄分两瓣，分趾蹄却不反刍，对你们是不洁净的。
LEV|11|8|这些兽的肉，你们不可吃；它们的尸体，你们也不可摸，对你们都是不洁净的。
LEV|11|9|“水中可吃的是这些：凡在水里，无论是海或河，有鳍有鳞的，都可以吃。
LEV|11|10|凡在海里、河里和水里滋生的动物，就是在水里所有的动物，无鳍无鳞的，对你们是可憎的。
LEV|11|11|它们对你们都是可憎的。你们不可吃它们的肉；它们的尸体，也当以为可憎。
LEV|11|12|凡在水里无鳍无鳞的，对你们是可憎的。
LEV|11|13|“飞鸟中你们当以为可憎，不可吃且可憎的是：雕、狗头雕、红头雕，
LEV|11|14|鹞鹰、小鹰的类群，
LEV|11|15|所有乌鸦的类群，
LEV|11|16|鸵鸟、夜鹰、鱼鹰、鹰的类群，
LEV|11|17|鸮鸟、鸬鹚、猫头鹰，
LEV|11|18|角鸱、鹈鹕、秃雕，
LEV|11|19|鹳、鹭鸶的类群，戴鵀与蝙蝠。
LEV|11|20|“凡有翅膀却用四足爬行的群聚动物，对你们是可憎的。
LEV|11|21|只是有翅膀却用四足爬行的群聚动物中，足上有腿在地上跳的，你们还可以吃；
LEV|11|22|其中你们可以吃的有蝗虫的类群，蚂蚱的类群，蟋蟀的类群和蚱蜢的类群。
LEV|11|23|其余有翅膀有四足的群聚动物，对你们都是可憎的。
LEV|11|24|“这些都能使你们不洁净。凡摸它们尸体的，必不洁净到晚上。
LEV|11|25|任何人搬动了它们的尸体，要把衣服洗净，必不洁净到晚上。
LEV|11|26|凡蹄分两瓣却不分趾或不反刍食物的走兽，对你们是不洁净的；谁摸了它们就不洁净。
LEV|11|27|凡用脚掌行走，四足行走的动物，对你们是不洁净的；凡摸它们尸体的，必不洁净到晚上。
LEV|11|28|谁搬动了它们的尸体，要把衣服洗净，必不洁净到晚上。这些对你们是不洁净的。
LEV|11|29|“在地上成群的群聚动物中，对你们不洁净的是这些：鼬鼠、鼫鼠、蜥蜴的类群，
LEV|11|30|壁虎、龙子、守宫、蛇医、蝘蜓。
LEV|11|31|这些群聚动物对你们都是不洁净的。在它们死后，凡摸了它们尸体的，必不洁净到晚上。
LEV|11|32|其中死了的，若掉在任何东西上，这东西就不洁净，无论是木器、衣服、皮革、麻袋，或是任何工作需用的器皿，都要泡在水中，必不洁净到晚上，然后才是洁净的。
LEV|11|33|若有一点掉在瓦器里，里面的任何东西就不洁净了； 你们要把这瓦器打破。
LEV|11|34|其中一切可吃的食物，沾到那水的就不洁净；器皿里可喝的东西，也必不洁净。
LEV|11|35|它们的尸体，只要有一点掉在任何物件上，那物件就不洁净。无论是烤炉或炉灶，都要打碎；它们不洁净，而且对你们也不洁净。
LEV|11|36|但是水泉或池子，就是聚水的地方，仍是洁净的；凡摸这些尸体的才不洁净。
LEV|11|37|若它们的尸体有一点掉在要播的种子上，种子仍是洁净的；
LEV|11|38|若水已经浇在种子上，它们的尸体有一点掉在上面，这种子对你们就是不洁净的了。
LEV|11|39|“你们可吃的走兽中若有死了的，谁摸了它的尸体，就必不洁净到晚上。
LEV|11|40|人若吃了那已死的走兽，要把衣服洗净，必不洁净到晚上。人若搬动了那已死的牲畜，要把衣服洗净，必不洁净到晚上。
LEV|11|41|“凡在地上成群的群聚动物都是可憎的，都不可吃。
LEV|11|42|凡用肚子爬行或用四脚爬行，或是用多足的，地上一切群聚的动物，你们都不可吃，因为是可憎的。
LEV|11|43|你们不可因任何群聚的动物使自己成为可憎的，也不可因它们成为不洁净，染了污秽。
LEV|11|44|我是耶和华－你们的上帝。你们要使自己分别为圣，要成为圣，因为我是神圣的。你们不可因地上爬行的群聚动物使自己不洁净。
LEV|11|45|我是把你们从 埃及 地领出来的耶和华，要作你们的上帝。你们要成为圣，因为我是神圣的。”
LEV|11|46|这是牲畜、飞鸟、水中一切游动的生物和地上一切爬行的动物的条例，
LEV|11|47|为要使你们能分辨洁净的和不洁净的，可吃的和不可吃的动物。
LEV|12|1|耶和华吩咐 摩西 说：
LEV|12|2|“你要吩咐 以色列 人说：妇人若怀孕生男孩，就不洁净七天，像在月经污秽的期间不洁净一样。
LEV|12|3|第八天，要给婴孩行割礼。
LEV|12|4|妇人产后流血的洁净，要家居三十三天。她洁净的日子未满，不可摸圣物，也不可进入圣所。
LEV|12|5|她若生女孩，就不洁净两个七天，像经期中一样。她产后流血的洁净，要家居六十六天。
LEV|12|6|“洁净的日子满了，无论生儿子或女儿，她要把一只一岁的羔羊作燔祭，一只雏鸽或一只斑鸠作赎罪祭，带到会幕的门口交给祭司。
LEV|12|7|祭司要把这祭物献在耶和华面前，为她赎罪。这样，她就从流血中得洁净了。这是为生男或生女之妇人的条例。
LEV|12|8|妇人的能力若不足，无法献一只羔羊，她就要取两只斑鸠或两只雏鸽，一只为燔祭，一只为赎罪祭。祭司要为她赎罪，她就洁净了。”
LEV|13|1|耶和华吩咐 摩西 和 亚伦 说：
LEV|13|2|“人身上的皮肤若肿胀，或发疹，或有斑点，可能成为痲疯 的灾病，就要把他带到 亚伦 祭司或 亚伦 的一个作祭司的子孙那里。
LEV|13|3|祭司要检查他身上皮肤的患处，若患处的毛已经变白，灾病的现象深入身上皮肤内，这就是痲疯的灾病。祭司检查后，要宣布他为不洁净。
LEV|13|4|若这人身上的皮肤有白斑，看起来并没有深入皮肤内，其上的毛也没有变白，祭司就要将这病人隔离七天。
LEV|13|5|第七天，祭司要检查他，看哪，若灾病在祭司眼前止住了，没有在皮肤上扩散，要将他再隔离七天。
LEV|13|6|到了第七天，祭司要再检查他。看哪，若灾病减轻，没有在皮肤上扩散，祭司就要宣布他为洁净，因为他患的不过是疹子。那人要洗自己的衣服，就洁净了。
LEV|13|7|他给祭司检查宣布为洁净后，疹子若在皮肤上大大扩散，他就要再给祭司检查。
LEV|13|8|祭司要检查，看哪，疹子若在皮肤上扩散了，祭司就要宣布他为不洁净，是痲疯病。
LEV|13|9|“人若得了痲疯的灾病，就要把他带到祭司那里。
LEV|13|10|祭司要检查，看哪，若皮肤有白色肿块，使毛变白，肿块里有嫩的新长的肉，
LEV|13|11|这就是他身上皮肤慢性的痲疯病。祭司要宣布他为不洁净，不必将他隔离，因为他已是不洁净了。
LEV|13|12|若痲疯在皮肤四处扩散，长满在患灾病之人的皮肤上，据祭司察看，从头到脚无处不有，
LEV|13|13|祭司就要检查，看哪，若这病人全身已长满了痲疯，就要宣布他为洁净；他全身都变白了，他是洁净的。
LEV|13|14|但他身上一旦出现新长的肉，就不洁净了。
LEV|13|15|祭司一见新长的肉，就要宣布他为不洁净。新长的肉是不洁净的，这就是痲疯病。
LEV|13|16|新长的肉若变白了，他就要到祭司那里。
LEV|13|17|祭司要检查，看哪，患处若变白了，祭司就要宣布那患灾病的人为洁净，他就洁净了。
LEV|13|18|“人身上的皮肤 若长了疮，却已经好了，
LEV|13|19|在长疮之处又发肿变白，或是出现白中带红的斑点，就要给祭司检查。
LEV|13|20|祭司要检查，看哪，若灾病的现象已深入皮肤内，其上的毛也变白了，祭司就要宣布他为不洁净，有痲疯的灾病生在疮中。
LEV|13|21|祭司若检查，看哪，其上没有白毛，也没有深入皮肤内，而且灾病减轻，祭司就要将他隔离七天。
LEV|13|22|若在皮肤上大大扩散，祭司就要宣布他为不洁净，这是灾病。
LEV|13|23|斑点若留在原处，没有扩散，这就是疮的疤痕，祭司就要宣布他为洁净。
LEV|13|24|“人身上的皮肤若被火烧伤，伤口新长的肉有了斑点，无论是白中带红，或是全白，
LEV|13|25|祭司就要检查，看哪，斑点上的毛若变白了，现象又深入皮肤内，这就是痲疯长在烧伤处；祭司就要宣布他为不洁净，是痲疯的灾病。
LEV|13|26|若祭司检查，看哪，斑点上没有白毛，也没有深入皮肤内，而且灾病减轻，祭司就要将他隔离七天。
LEV|13|27|第七天，祭司要检查他。斑点若在皮肤上大大扩散，祭司就要宣布他为不洁净，是患了痲疯的灾病。
LEV|13|28|斑点若留在原处，没有在皮肤上扩散，并减轻了，它只是烧伤的肿块，祭司要宣布他为洁净，这不过是烧伤后的疤痕。
LEV|13|29|“无论男女，若在头上或下巴有灾病，
LEV|13|30|祭司就要检查这灾病，看哪，若灾病的现象深入皮肤内，其上有黄色的细毛，祭司就要宣布他为不洁净，这是疥疮，是头上或下巴的痲疯病。
LEV|13|31|祭司要检查这疥疮的灾病，看哪，现象若未深入皮肤内，其上也没有黑毛，祭司就要将长疥疮的人隔离七天。
LEV|13|32|第七天，祭司要检查这灾病，看哪，若疥疮没有扩散，其上没有黄色的毛，疥疮的现象也没有深入皮肤内，
LEV|13|33|那人就要剃去须发，但不可剃长疥疮之处。祭司要将那长疥疮的人，再隔离七天。
LEV|13|34|第七天，祭司要检查疥疮，看哪，疥疮若没有在皮肤上扩散，现象也未深入在皮肤内，祭司就要宣布他为洁净；那人要洗自己的衣服，就洁净了。
LEV|13|35|但他被宣布为洁净后，疥疮若在皮肤上大大扩散，
LEV|13|36|祭司就要检查他。看哪，疥疮若在皮肤上扩散，祭司就不必找黄色的毛，这人是不洁净了。
LEV|13|37|若疥疮在祭司眼前止住了，其上长了黑毛，疥疮就已痊愈了，那人是洁净的，祭司要宣布他为洁净。
LEV|13|38|“无论男女，身上的皮肤若有斑点，是白色的斑点，
LEV|13|39|祭司就要检查，看哪，若皮肤的斑点是暗白色的，这是皮肤长了斑；那人是洁净的。
LEV|13|40|“人的头发若掉了，变成秃头，他是洁净的。
LEV|13|41|他头顶的前面若掉了头发，以致顶门光秃，他是洁净的。
LEV|13|42|头秃处或顶门秃处，若有白中带红的灾病，这就是痲疯长在他的头秃处或顶门秃处。
LEV|13|43|祭司要检查他，看哪，若头秃处或顶门秃处的灾病肿块白中带红，像身上皮肤痲疯病的现象一样，
LEV|13|44|那人就是患了痲疯病，是不洁净的。祭司要宣布他为不洁净；他的灾病是生在头上。
LEV|13|45|“患有痲疯灾病的人，他的衣服要撕裂，也要蓬头散发，遮住上唇，喊着说：‘不洁净！不洁净！’
LEV|13|46|灾病还在他身上的时候，他就是不洁净的；既然不洁净，他就要独居，住在营外。”
LEV|13|47|“衣服若发霉 了，无论是羊毛衣服、麻布衣服，
LEV|13|48|无论是经线、纬线，是麻布的、羊毛的，是皮革，或是任何皮制的物件；
LEV|13|49|若是衣服、皮革、经线、纬线，或是任何皮制的物件呈现绿色或红色，这就是发霉，必须给祭司检查。
LEV|13|50|祭司要检查这霉，把发霉的物件隔离七天。
LEV|13|51|第七天，他要检查这霉。若霉在衣服上，无论是经线、纬线，或任何用途的皮制物件上扩散，这是侵蚀性的霉，是不洁净的。
LEV|13|52|发霉的衣服，无论在经线、纬线，羊毛的、麻布的，或是任何皮制物件，都要把它烧掉；因为这是侵蚀性的霉，必须用火焚烧。
LEV|13|53|祭司检查，看哪，霉若在衣服上，无论是经线、纬线，或在任何的皮制物件上没有扩散，
LEV|13|54|祭司就要吩咐人把发霉的物件洗了，再隔离七天。
LEV|13|55|洗过之后，祭司要检查，看哪，若那霉在他眼前没有变色，霉虽没有扩散，也是不洁净的。这是侵蚀性的灾病，无论是在正面或反面，都要用火焚烧那物件。
LEV|13|56|祭司若检查，看哪，那霉在洗过之后已经褪色，他就要从衣服，皮革，或经线、纬线，把发霉的部分撕去。
LEV|13|57|若霉再出现在衣服上，无论是经线、纬线、或在任何皮制物件上，这就是旧霉复发，必须用火将那发霉的物件焚烧。
LEV|13|58|洗过的衣服，或是经线，纬线，或是任何皮制的物件，若霉已经消失了，仍要再洗，这衣服就洁净了。”
LEV|13|59|这就是衣服发霉的条例。无论是羊毛衣服，麻布衣服，或是经线、纬线，或任何皮制的物件，都按照这条例宣布为洁净或不洁净。
LEV|14|1|耶和华吩咐 摩西 说：
LEV|14|2|“这是患痲疯病的人得洁净时的条例：要带他到祭司那里，
LEV|14|3|祭司要出到营外，检查那患痲疯病的人，看哪，他的痲疯灾病已经痊愈了，
LEV|14|4|祭司就要吩咐人为那求洁净的人带两只洁净的活鸟和香柏木、朱红色纱，以及牛膝草来。
LEV|14|5|祭司要吩咐用瓦器盛清水，把第一只鸟宰在上面。
LEV|14|6|至于那只活鸟，祭司要把它和香柏木、朱红色纱，以及牛膝草，一同蘸在宰于清水上的鸟血中。
LEV|14|7|他要向那从痲疯病中得洁净的人身上弹血七次，宣布他为洁净，然后把那活鸟在野地里放走。
LEV|14|8|求洁净的人要洗衣服，剃去所有的毛发，用水洗澡，他就洁净了。然后，他可以进营，不过仍要在自己的帐棚外居住七天。
LEV|14|9|到了第七天，他要剃所有的毛发，头发、胡须、眼睛的眉毛，他全身的毛都剃了；然后，他要洗衣服，用水洗身，才洁净了。
LEV|14|10|“第八天，他要取两只没有残疾的小公羊和一只没有残疾、一岁的小母羊，以及作为素祭的十分之三伊法调了油的细面和一罗革的油。
LEV|14|11|宣布洁净的祭司要将那求洁净的人，连同这些东西，安置在耶和华面前，会幕的门口。
LEV|14|12|祭司要取一只小公羊献为赎愆祭，又取一罗革的油，把它们在耶和华面前摇一摇，作为摇祭；
LEV|14|13|再把小公羊宰于圣处，就是宰赎罪祭牲和燔祭牲的地方。赎愆祭要归给祭司，与赎罪祭一样，是至圣的。
LEV|14|14|祭司要取一些赎愆祭牲的血，抹在求洁净的人的右耳垂上、右手的大拇指上和右脚的大脚趾上。
LEV|14|15|祭司要从那一罗革的油中，取一些倒在自己的左手掌里，
LEV|14|16|祭司要用右手指蘸在他左手掌的油里，在耶和华面前用手指弹七次。
LEV|14|17|祭司要把手掌里剩下的油抹在那求洁净的人的右耳垂上、右手的大拇指上和右脚的大脚趾上，在赎愆祭牲之血抹过的上面。
LEV|14|18|祭司手掌里剩下的油要抹在那求洁净的人的头上，祭司就在耶和华面前为他赎罪。
LEV|14|19|祭司要献赎罪祭，为那从不洁净中得洁净的人赎罪，然后要宰燔祭牲，
LEV|14|20|祭司要把燔祭和素祭献在坛上，祭司要为他赎罪，他就洁净了。
LEV|14|21|“他若贫穷，手头财力不及，就要取一只小公羊作赎愆祭，作摇祭为他赎罪。他也要把作为素祭的十分之一伊法调了油的细面，和一罗革的油，一同取来。
LEV|14|22|他又要照手头财力所及，取两只斑鸠或两只雏鸽，一只作赎罪祭，一只作燔祭。
LEV|14|23|第八天，为了使自己洁净，他要把这些祭物带到耶和华面前，在会幕的门口交给祭司。
LEV|14|24|祭司要把赎愆祭的羔羊和那一罗革的油一同在耶和华面前摇一摇，作为摇祭。
LEV|14|25|祭司要宰赎愆祭的羔羊，取一些赎愆祭牲的血，抹在那求洁净的人的右耳垂上、右手的大拇指上和右脚的大脚趾上。
LEV|14|26|祭司要把一些油倒在自己的左手掌里，
LEV|14|27|祭司要用右手指，把他左手掌里的油在耶和华面前弹七次。
LEV|14|28|祭司要把手掌里的油抹一些在那求洁净的人的右耳垂上、右手的大拇指上和右脚的大脚趾上，在赎愆祭牲之血抹过之处的上面。
LEV|14|29|祭司手掌里剩下的油要抹在那求洁净的人的头上，在耶和华面前为他赎罪。
LEV|14|30|那人又要照他手头财力所及，献上斑鸠中的一只或雏鸽中的一只，
LEV|14|31|照他手头财力所及，一只为赎罪祭，一只为燔祭，与素祭一同献上。祭司就在耶和华面前为他赎罪。
LEV|14|32|这是为患痲疯灾病，手头财力不及而求洁净的人所定的条例。”
LEV|14|33|耶和华吩咐 摩西 和 亚伦 说：
LEV|14|34|“你们到了我所赐给你们为业的 迦南 地，我若使你们所得为业之地的房屋发霉 ，
LEV|14|35|屋主就要去告诉祭司说：‘据我看，房屋似乎发霉了。’
LEV|14|36|祭司进去检查这霉之前，要吩咐把屋内的东西全部搬走，免得屋子里所有的东西成为不洁净。然后，祭司要进去检查房屋。
LEV|14|37|他要检查这霉，看哪，若屋子墙上的霉有发绿或发红凹入的斑纹，其现象深入墙内，
LEV|14|38|祭司就要出到屋子的门外，把屋子封锁七天。
LEV|14|39|第七天，祭司要再去检查，看哪，霉若在屋子的墙上扩散，
LEV|14|40|祭司要吩咐把发霉的石头挖出来，扔在城外不洁净之处。
LEV|14|41|他也要叫人刮屋内的四围，把刮出来的灰泥倒在城外不洁净之处。
LEV|14|42|他们要用别的石头取代挖出来的石头，用别的灰泥涂抹屋子。
LEV|14|43|“他挖出石头，刮了屋子，涂抹以后，霉若又在屋子里出现，
LEV|14|44|祭司就要进去检查，看哪，霉若在屋子里扩散，那就是有侵蚀性的霉在屋子里，是不洁净的。
LEV|14|45|他要拆毁屋子，把石头、木料和所有的灰泥都搬到城外不洁净之处。
LEV|14|46|屋子封锁的任何时候，进去的人必不洁净到晚上。
LEV|14|47|在屋子里躺卧的人必须把衣服洗净，在屋子里吃饭的人也必须把衣服洗净。
LEV|14|48|“屋子涂抹了之后，祭司若进去检查，看哪，霉没有在屋内扩散，就要宣布这房屋为洁净，因为霉已经消除了。
LEV|14|49|他要为洁净房屋取两只鸟和香柏木、朱红色纱，以及牛膝草，
LEV|14|50|用瓦器盛清水，把一只鸟宰在上面。
LEV|14|51|他要把香柏木、牛膝草、朱红色纱和那一只活鸟，都蘸在被宰的鸟血和清水中，用来弹屋子七次。
LEV|14|52|他要用鸟血、清水、活鸟、香柏木、牛膝草和朱红色纱洁净那房屋。
LEV|14|53|他要把活鸟在城外野地里放走。他要为房屋赎罪，房屋就洁净了。”
LEV|14|54|这条例是为痲疯灾病和疥疮，
LEV|14|55|衣服和房屋发霉，
LEV|14|56|以及皮肤肿胀、发疹、有斑点等，
LEV|14|57|用以分辨何时洁净，何时不洁净。这是痲疯病的条例。
LEV|15|1|耶和华吩咐 摩西 和 亚伦 说：
LEV|15|2|“你们要吩咐 以色列 人，对他们说：人若身体 患了漏症，他因这症就不洁净了。
LEV|15|3|这就是他因漏症而有的不洁净：无论是身体流出液体，或身体已经止住不再有液体，他都是不洁净的。
LEV|15|4|那患漏症的人所躺的床都不洁净，所坐的任何东西也不洁净。
LEV|15|5|凡摸他床的人，要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|6|人坐了漏症患者坐过的东西，他要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|7|人摸了漏症患者，他要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|8|若漏症患者吐唾沫在洁净的人身上，这人要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|9|漏症患者所骑的任何鞍子也不洁净。
LEV|15|10|凡摸了他坐过的任何东西，必不洁净到晚上；拿了这些东西的，要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|11|漏症患者若没有用水冲洗他的手，无论摸了谁，谁就要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|12|漏症患者所摸的瓦器必要打破；他所摸的一切木器必要用水冲洗。
LEV|15|13|“漏症患者的漏症痊愈了，就要为洁净自己计算七天，也要洗衣服，用清水洗身，就洁净了。
LEV|15|14|第八天，他要带两只斑鸠或两只雏鸽，来到耶和华面前，在会幕门口把鸟交给祭司。
LEV|15|15|祭司要献上一只为赎罪祭，一只为燔祭。祭司要因这人所患的漏症，在耶和华面前为他赎罪。
LEV|15|16|“人若遗精，他要用水洗全身，必不洁净到晚上。
LEV|15|17|无论是衣服或皮革，若沾染了精液，要用水洗净，必不洁净到晚上。
LEV|15|18|女人，若有男人与她同寝，沾染了精液，二人要用水洗澡，必不洁净到晚上。”
LEV|15|19|“女人月经期间，有血从体内流出，她必不洁净七天；凡摸她的，必不洁净到晚上。
LEV|15|20|在不洁净期间，女人所躺的东西都不洁净，所坐的任何东西也不洁净。
LEV|15|21|凡摸她床的，要洗衣服，用水洗澡，必不洁净到晚上；
LEV|15|22|凡摸她坐过的东西的，要洗衣服，用水洗澡，必不洁净到晚上；
LEV|15|23|不论是床，或她坐过的东西，人摸了，必不洁净到晚上。
LEV|15|24|男人若和这女人同寝，沾了她的不洁净，就不洁净七天，所躺的床也都不洁净。
LEV|15|25|“女人若在经期之外仍然流血多日，或是经期过长，她在流血的一切日子都不洁净，和她在经期的日子不洁净一样。
LEV|15|26|在流血的日子，她所躺的床、所坐的任何东西都不洁净，和在月经期间不洁净一样。
LEV|15|27|凡摸这些东西的，就不洁净；他要洗衣服，用水洗澡，必不洁净到晚上。
LEV|15|28|这女人的血漏若痊愈了，就要计算七天，然后才洁净。
LEV|15|29|第八天，她要取两只斑鸠或两只雏鸽，带到会幕门口祭司那里。
LEV|15|30|祭司要献一只为赎罪祭，一只为燔祭。祭司要因这女人血漏的不洁净，在耶和华面前为她赎罪。
LEV|15|31|“你们要使 以色列 人与他们的不洁净隔离，免得他们玷污我在他们中间的帐幕，因自己的不洁净死亡。”
LEV|15|32|这条例是为漏症患者或遗精而不洁净者，
LEV|15|33|女人经期的不洁，男女患漏症，以及男人与不洁净女人同寝而立的。
LEV|16|1|亚伦 的两个儿子靠近耶和华面前，死了。他们死后，耶和华吩咐 摩西 ；
LEV|16|2|耶和华对 摩西 说：“你要吩咐你哥哥 亚伦 ，不可随时进入圣所的幔子内、到柜盖 前，免得他死亡，因为我在柜盖上的云中显现。
LEV|16|3|亚伦 进圣所要带这些：一头公牛犊为赎罪祭，一只公绵羊为燔祭。
LEV|16|4|他要穿上细麻布圣内袍，把细麻布裤子穿在身上，腰束细麻布带子，头戴细麻布礼冠；这些都是圣服。他要用水洗身，然后穿上圣服。
LEV|16|5|他要从 以色列 会众中取两只公山羊为赎罪祭，一只公绵羊为燔祭。
LEV|16|6|“亚伦要把他自己赎罪祭的公牛献上，为自己和家人赎罪；
LEV|16|7|也要把两只公山羊牵到耶和华面前，安置在会幕的门口。
LEV|16|8|亚伦 要为那两只山羊抽签，一签归给耶和华，一签归给 阿撒泻勒 。
LEV|16|9|亚伦 要把那抽中归给耶和华的山羊牵来献为赎罪祭，
LEV|16|10|至于抽中归给 阿撒泻勒 的山羊，却要活着安放在耶和华面前，用以赎罪，然后送到旷野去，归给 阿撒泻勒 。
LEV|16|11|“ 亚伦 要把他自己赎罪祭的公牛献上，为自己和家人赎罪，他要宰作自己赎罪祭的公牛。
LEV|16|12|他要从耶和华面前的坛上取盛满火炭的香炉，再拿一捧捣细的香料，把这些都带入幔子内。
LEV|16|13|在耶和华面前，他要把香放在火上，使香的烟云遮着法柜上的盖子，免得他死亡。
LEV|16|14|他要取一些公牛的血，用手指弹在柜盖的前面，就是东面，又在柜盖的前面用手指弹血七次。
LEV|16|15|“他要宰那只为百姓作赎罪祭的公山羊，把羊的血带入幔子内，把血弹在柜盖的上面和前面，好像弹公牛的血一样。
LEV|16|16|因 以色列 人的不洁净和过犯，就是他们一切的罪，他要为圣所赎罪；因会幕在他们不洁净之中，他也要为会幕照样做。
LEV|16|17|他进圣所赎罪的时候，会幕里都不准有人，直等到他为自己和家人，以及 以色列 全会众赎了罪出来。
LEV|16|18|他出来后，要到耶和华面前的祭坛那里，为坛赎罪。他要取一些公牛的血和公山羊的血，抹在坛周围的四个翘角上。
LEV|16|19|他也要用手指把血弹在坛上七次，使坛从 以色列 人的不洁净中得以洁净，成为圣。”
LEV|16|20|“ 亚伦 为圣所和会幕，以及祭坛赎罪后，就要把那只活的公山羊牵来。
LEV|16|21|他的双手要按在活的山羊的头上，承认 以色列 人所有的罪孽过犯，就是他们一切的罪，把这些罪都归在羊的头上，再指派一个人把它送到旷野去。
LEV|16|22|这羊要担当他们一切的罪孽，带到无人之地；那人要把羊送到旷野去。
LEV|16|23|“ 亚伦 要进入会幕，把他进圣所时所穿的细麻布衣服脱下，放在那里，
LEV|16|24|又要在圣处用水洗身，穿上衣服出来，把自己的燔祭和百姓的燔祭献上，为自己和百姓赎罪。
LEV|16|25|赎罪祭牲的脂肪要烧在坛上。
LEV|16|26|那放走山羊归给 阿撒泻勒 的人要洗衣服，用水洗身，然后才可以回到营里。
LEV|16|27|作赎罪祭的公牛和作赎罪祭的公山羊的血被带入圣所赎罪之后，就要把这牛羊搬到营外，皮、肉、粪都用火焚烧。
LEV|16|28|焚烧的人要洗衣服，用水洗身，然后才可以回到营里。”
LEV|16|29|“这是你们永远的定例：每年七月初十，你们要刻苦己心；无论是本地人，是寄居在你们中间的外人，任何工都不可做。
LEV|16|30|因为这日要为你们赎罪，洁净你们，使你们脱离一切的罪，在耶和华面前得以洁净。
LEV|16|31|这日你们要守完全安息的安息日，刻苦己心；这是永远的定例。
LEV|16|32|那受膏接续他父亲担任圣职的祭司要赎罪，穿上细麻布衣服，就是圣衣，
LEV|16|33|为至圣所和会幕赎罪，为祭坛赎罪，并要为祭司和会众的全体百姓赎罪。
LEV|16|34|这要作你们永远的定例：因 以色列 人一切的罪，要一年一次为他们赎罪。”于是， 亚伦 照耶和华所吩咐 摩西 的做了 。
LEV|17|1|耶和华吩咐 摩西 说：
LEV|17|2|“你要吩咐 亚伦 和他儿子，以及 以色列 众人，对他们说，耶和华所吩咐的话是这样：
LEV|17|3|凡 以色列 家中的人宰公牛，或小绵羊，或山羊，无论是在营内或营外，
LEV|17|4|若不把牲畜牵到会幕门口耶和华的帐幕前，献给耶和华为供物，所流的血必归到那人身上。他既使血流出，就要从百姓中剪除。
LEV|17|5|这是为要使 以色列 人把他们在野地里所宰的祭牲带来，带到耶和华前，会幕门口祭司那里，宰杀这些祭牲，把它们献给耶和华为平安祭。
LEV|17|6|祭司要在会幕门口，把血洒在耶和华的祭坛上，把脂肪焚烧，献给耶和华为馨香的祭。
LEV|17|7|他们不可再宰杀祭牲献给他们行淫所随从的山羊鬼魔。这要作他们世世代代永远的定例。
LEV|17|8|“你要对他们说：凡 以色列 家中的任何人，或寄居在他们中间的外人献燔祭或祭物，
LEV|17|9|若不带到会幕门口献给耶和华，那人必从百姓中剪除。
LEV|17|10|“凡 以色列 家中的任何人，或寄居在他们中间的外人，吃任何的血，我必向那吃血的人变脸，把他从百姓中剪除。
LEV|17|11|因为动物的生命是在血中。我把这血赐给你们，可以在祭坛上为你们的生命赎罪；因为血就是生命，能够赎罪。
LEV|17|12|因此，我对 以色列 人说：你们都不可吃血；寄居在你们中间的外人也不可吃血。
LEV|17|13|凡 以色列 人，或寄居在他们中间的外人，猎取了可吃的飞禽走兽，必须把它的血放出来，用土掩盖。
LEV|17|14|“因一切动物的生命，它的血就是它的生命。所以我对 以色列 人说：无论什么动物的血，你们都不可吃，因为一切动物的生命就是它的血。凡吃血的必被剪除。
LEV|17|15|无论是本地人，是寄居的，若吃了自然死去或被野兽撕裂的动物，要洗衣服，用水洗澡，必不洁净到晚上，晚上就洁净了。
LEV|17|16|但他若不洗衣服，也不洗身，就要担当自己的罪孽。”
LEV|18|1|耶和华吩咐 摩西 说：
LEV|18|2|“你要吩咐 以色列 人，对他们说：我是耶和华－你们的上帝。
LEV|18|3|你们不可做你们从前住 埃及 地的人所做的，也不可做我要领你们去的 迦南 地的人所做的。你们不可照他们的习俗行。
LEV|18|4|你们要遵行我的典章，谨守我的律例，按此而行。我是耶和华－你们的上帝。
LEV|18|5|你们要谨守我的律例典章；遵行的人就必因此得生。我是耶和华。
LEV|18|6|“任何人都不可亲近骨肉之亲，露其下体。我是耶和华。
LEV|18|7|你父亲的下体，就是你母亲的下体，你不可露；她是你的母亲，不可露她的下体。
LEV|18|8|不可露你继母的下体，就是你父亲的下体。
LEV|18|9|你姊妹的下体，或是同父异母的，或是同母异父的，无论生在家或生在外的，都不可露她们的下体。
LEV|18|10|不可露你孙女或外孙女的下体，因为她们的下体就是你自己的下体。
LEV|18|11|你继母为你父亲所生的女儿是你的姊妹，不可露她的下体。
LEV|18|12|不可露你姑母的下体；她是你父亲的骨肉之亲。
LEV|18|13|不可露你姨母的下体；她是你母亲的骨肉之亲。
LEV|18|14|不可露你叔伯的下体，不可亲近他的妻子；她是你的叔母、伯母。
LEV|18|15|不可露你媳妇的下体，她是你儿子的妻，不可露她的下体。
LEV|18|16|不可露你兄弟妻子的下体，这是你兄弟的下体。
LEV|18|17|不可露妇人的下体，又露她女儿的下体，也不可娶她的孙女或外孙女，露她们的下体；她们是骨肉之亲 。这是邪恶的事。
LEV|18|18|你妻子还活着的时候，不可另娶她的姊妹与她作对，露她姊妹的下体。
LEV|18|19|“不可亲近经期中不洁净的女人，露她的下体。
LEV|18|20|不可跟邻舍的妻交合，因她玷污自己。
LEV|18|21|不可使你儿女经火献给 摩洛 ，也不可亵渎你上帝的名。我是耶和华。
LEV|18|22|不可跟男人同寝，像跟女人同寝；这是可憎恶的事。
LEV|18|23|不可跟兽交合，因它玷污自己。女人也不可站在兽前，与它交合；这是逆性的事。
LEV|18|24|“在这一切的事上，你们都不可玷污自己，因为我在你们面前所逐出的列国，在这一切的事上玷污了自己。
LEV|18|25|连地也玷污了，我惩罚那地的罪孽，地就吐出它的居民来。
LEV|18|26|但你们要遵守我的律例典章。这一切可憎恶的事，无论是本地人或寄居在你们中间的外人，都不可以做。
LEV|18|27|在你们之前居住那地的人做了这一切可憎恶的事，地就玷污了。
LEV|18|28|不要让地因你们玷污了它而把你们吐出来，像吐出在你们之前的国一样。
LEV|18|29|无论是谁，若做了这其中一件可憎恶的事，必从百姓中剪除。
LEV|18|30|你们要遵守我的吩咐，免得你们随从那些可憎的习俗，就是在你们之前的人所做的，玷污了自己。我是耶和华－你们的上帝。”
LEV|19|1|耶和华吩咐 摩西 说：
LEV|19|2|“你要吩咐 以色列 全会众，对他们说：你们要成为圣，因为我耶和华－你们的上帝是神圣的。
LEV|19|3|你们各人都当孝敬父母，也要守我的安息日。我是耶和华－你们的上帝。
LEV|19|4|你们不可转向虚无的神明，也不可为自己铸造神像。我是耶和华－你们的上帝。
LEV|19|5|“你们宰杀祭牲献平安祭给耶和华的时候，要献得使你们可蒙悦纳。
LEV|19|6|这祭物要在献的当天或第二天吃；若有剩到第三天的，就要用火焚烧。
LEV|19|7|第三天若再吃，这祭物是不洁净的，必不蒙悦纳。
LEV|19|8|吃的人必担当自己的罪孽，因为他亵渎了耶和华的圣物，这人必从百姓中剪除。
LEV|19|9|“你们在自己的地收割庄稼时，不可割尽田的角落，也不可拾取庄稼所掉落的。
LEV|19|10|不可摘尽葡萄园的葡萄，也不可拾取葡萄园中掉落的葡萄，要把它们留给穷人和寄居的。我是耶和华－你们的上帝。
LEV|19|11|“你们不可偷盗，不可欺骗，也不可彼此说谎。
LEV|19|12|不可指着我的名起假誓，亵渎你上帝的名。我是耶和华。
LEV|19|13|“不可欺压你的邻舍，也不可偷盗。雇工的工钱不可在你那里过夜，留到早晨。
LEV|19|14|不可咒骂聋子，也不可将绊脚石放在盲人面前。你要敬畏你的上帝。我是耶和华。
LEV|19|15|“你们审判的时候，不可不公正；不可偏护贫穷人，也不可看重有权势人的脸，总要公平审判你的邻舍。
LEV|19|16|不可在百姓中到处搬弄是非，不可陷害邻舍的性命 。我是耶和华。
LEV|19|17|“不可心里恨你的弟兄；要指摘你的邻舍，免得因他承担罪过。
LEV|19|18|不可报仇，也不可埋怨你本国的子民。你要爱邻如己。我是耶和华。
LEV|19|19|“你们要遵守我的律例。不可使你的牲畜与异类交配；不可在你的田地播下两样的种子；也不可穿两种原料做成的衣服。
LEV|19|20|“若有人与女子同寝交合，而她是婢女，许配了丈夫，尚未被赎或得自由，就要受到惩罚，却不可把他们处死，因为婢女还没有得自由。
LEV|19|21|男的要把赎愆祭，就是一只公绵羊牵到耶和华面前，会幕的门口。
LEV|19|22|祭司要用赎愆祭的羊在耶和华面前为他所犯的罪赎罪，他所犯的罪就必蒙赦免。
LEV|19|23|“你们到了 迦南 地，栽种各样的果树，就要把所结的果子当作不洁净的 ；三年之内，你们要把它视为不洁净，是不可吃的。
LEV|19|24|但第四年所结的果子全是圣的，用以赞美耶和华 。
LEV|19|25|第五年，你们就可以吃树上的果子，使树给你们结出更多的果子。我是耶和华－你们的上帝。
LEV|19|26|“你们不可吃带血的食物。不可占卜，也不可观星象。
LEV|19|27|头的周围 不可剃，胡须的周围不可损坏。
LEV|19|28|不可为死人割划自己的身体，也不可在身上刺花纹。我是耶和华。
LEV|19|29|“不可侮辱你的女儿，使她沦为娼妓，免得这地行淫乱，地就充满了邪恶。
LEV|19|30|你们要谨守我的安息日，敬畏我的圣所。我是耶和华。
LEV|19|31|“不可转向招魂的，也不可求问行巫术的，免得被他们玷污。我是耶和华－你们的上帝。
LEV|19|32|“在白发的人面前，你要站起来，要尊敬老人；要敬畏你的上帝，我是耶和华。
LEV|19|33|“若有外人寄居在你们的地上和你同住，不可欺负他。
LEV|19|34|寄居在你们那里的外人，你们要看他如本地人，并要爱他如己，因为你们在 埃及 地也作过寄居的。我是耶和华－你们的上帝。
LEV|19|35|“你们审判的时候，不可用不公正的度量衡。
LEV|19|36|你们要用公正的天平、公正的法码、公正的伊法和公正的欣。我是耶和华－你们的上帝，曾把你们从 埃及 地领出来。
LEV|19|37|你们要谨守我一切的律例典章，遵行它们。我是耶和华。”
LEV|20|1|耶和华吩咐 摩西 说：
LEV|20|2|“你要对 以色列 人说：凡 以色列 人，或是寄居在 以色列 的外人，把自己儿女献给 摩洛 的，必被处死；本地的百姓要用石头打死他。
LEV|20|3|我也要向那人变脸，把他从百姓中剪除，因为他把儿女献给 摩洛 ，玷污了我的圣所，亵渎了我的圣名。
LEV|20|4|那人把儿女献给 摩洛 ，本地的百姓若假装没看见，不把他处死，
LEV|20|5|我就要向这人和他的家人变脸，把他和所有跟随他与 摩洛 行淫的人都从百姓中剪除。
LEV|20|6|“人若转向招魂的和行巫术的，随从他们行淫，我就要向这人变脸，把他从百姓中剪除。
LEV|20|7|你们要使自己分别为圣，要成为圣，因为我是耶和华－你们的上帝。
LEV|20|8|你们要谨守我的律例，遵行它们；我是使你们分别为圣的耶和华。
LEV|20|9|凡咒骂父母的，必被处死；他咒骂了父母，他的血要归在他身上。
LEV|20|10|“凡与有夫之妇行奸淫，就是与邻舍的妻子行奸淫的，奸夫淫妇必被处死。
LEV|20|11|人若与继母同寝，就是露了父亲的下体，二人必被处死，血要归在他们身上。
LEV|20|12|人若与媳妇同寝，二人必被处死；他们行了乱伦的事，血要归在他们身上。
LEV|20|13|男人若跟男人同寝，像跟女人同寝，他们二人行了可憎恶的事，必被处死，血要归在他们身上。
LEV|20|14|人若娶妻，又娶妻子的母亲，这是邪恶的事；要把这三人用火焚烧，在你们中间除去这邪恶。
LEV|20|15|人若与兽交合，必被处死；你们也要杀死那兽。
LEV|20|16|女人若与兽亲近，与它交合，你要把那女人和兽杀死；他们必被处死，血要归在他们身上。
LEV|20|17|“人若娶自己的姊妹，或是同父异母的，或是同母异父的，彼此见了下体，这是可耻的事；他们必在自己百姓眼前被剪除。他露了姊妹的下体，必担当自己的罪孽。
LEV|20|18|若有人跟经期中的妇人同寝，露了她的下体，暴露妇人的血源，妇人也露了自己的血源，二人必从百姓中剪除。
LEV|20|19|不可露姨母或姑母的下体，因为这是露了骨肉之亲的下体，他们必担当自己的罪孽。
LEV|20|20|人若与叔伯之妻同寝，就露了他叔伯的下体，他们必担当自己的罪，必没有子女而死。
LEV|20|21|人若娶了自己兄弟的妻子，就露了他兄弟的下体，这是不洁净的事，他们必没有子女。
LEV|20|22|“你们要谨守我一切的律例典章，遵行它们，免得我领你们去住的那地把你们吐出来。
LEV|20|23|我在你们面前所逐出的国民，你们不可随从他们的风俗。因为他们行了这一切的事，所以我厌恶他们。
LEV|20|24|但我对你们说过，你们要承受他们的土地；我要把这流奶与蜜之地赐给你们，作为你们的产业。我是耶和华－你们的上帝，是把你们从万民中分别出来的。
LEV|20|25|你们要分辨洁净和不洁净的飞禽走兽；不可因我定为不洁净的飞禽走兽，或爬行在土地上的任何生物，使自己成为可憎恶的。
LEV|20|26|你们要归我为圣，因为－我耶和华是神圣的；我把你们从万民中分别出来，作我的子民。
LEV|20|27|“无论男女，是招魂的或行巫术的，他们必被处死。人要用石头打死他们，血要归在他们身上。”
LEV|21|1|耶和华对 摩西 说：“你要告诉 亚伦 子孙作祭司的，对他们说：祭司不可为自己百姓中的死人玷污自己，
LEV|21|2|除非是他的骨肉之亲，他的父母、儿女、兄弟、
LEV|21|3|或未出嫁还是处女的姊妹，因她是至亲，才可以玷污自己。
LEV|21|4|祭司既然在自己百姓中为首，就不可从俗玷污自己 。
LEV|21|5|“不可使头光秃，不可剃除胡须的边缘，也不可割划自己的身体。
LEV|21|6|他们要归上帝为圣，不可亵渎他们上帝的名，因为耶和华的火祭，就是上帝的食物，是他们献的，所以他们要成为圣。
LEV|21|7|“祭司不可娶妓女，或被玷污的女人为妻，也不可娶被休的妇人为妻，因为他是归上帝为圣的。
LEV|21|8|你要使祭司分别为圣，因为他献你上帝的食物。你要以他为圣，因为我是使你们分别为圣 的耶和华，是神圣的。
LEV|21|9|“祭司的女儿若行淫玷污自己，就侮辱了父亲，要用火将她焚烧。
LEV|21|10|“在弟兄中作大祭司的，头上倒了膏油，承接圣职，穿了圣衣，不可蓬头散发，也不可撕裂衣服；
LEV|21|11|不可挨近任何死尸，即使为了父母也不可玷污自己。
LEV|21|12|他不可出圣所，免得亵渎了上帝的圣所，因为在他身上有上帝的膏油为圣冕。我是耶和华。
LEV|21|13|他要娶处女为妻。
LEV|21|14|大祭司不可娶寡妇，被休的妇人，或被玷污的妓女为妻；他只可以娶自己百姓中的处女为妻。
LEV|21|15|他不可在自己百姓中侮辱他的儿女，因为我是使他分别为圣的耶和华。”
LEV|21|16|耶和华吩咐 摩西 说：
LEV|21|17|“你吩咐 亚伦 说：你世世代代的后裔，凡有残疾的都不可近前来献上帝的食物。
LEV|21|18|因为凡有残疾的，无论是失明的、瘸腿的、五官不正的、肢体之一过长的、
LEV|21|19|断脚的、断手的、
LEV|21|20|驼背的、侏儒的、有眼疾的、长癣的、长疥的，或是睾丸压伤的，都不可近前来。
LEV|21|21|亚伦 祭司的后裔，凡有残疾的都不可近前来献耶和华的火祭。他有残疾，不可近前来献上帝的食物。
LEV|21|22|上帝的食物，无论是圣的，或是至圣的，他都可以吃。
LEV|21|23|但他不可进到幔子前，也不可挨近祭坛前，因为他有残疾，免得他亵渎我的圣所。我是使他们分别为圣的耶和华。”
LEV|21|24|于是， 摩西 吩咐了 亚伦 和他的儿子，以及 以色列 众人。
LEV|22|1|耶和华吩咐 摩西 说：
LEV|22|2|“你要吩咐 亚伦 和他子孙说：你们要谨慎处理 以色列 人所分别为圣，归给我的圣物，免得亵渎我的圣名。我是耶和华。
LEV|22|3|你要对他们说：你们世世代代的后裔，凡不洁净，却挨近 以色列 人所分别为圣，归给耶和华的圣物，那人必从我面前剪除。我是耶和华。
LEV|22|4|亚伦 的后裔中，凡有痲疯病的，或患漏症的，都不可吃圣物，直等他洁净了。无论谁摸了那因尸体而不洁净的东西，或遗精的人，
LEV|22|5|或摸到任何使他不洁净的群聚动物或使他不洁净的人，无论那人有什么不洁净，
LEV|22|6|摸了这些的人必不洁净到晚上；若不用水洗身，就不可吃圣物。
LEV|22|7|日落的时候，他就洁净了，然后可以吃圣物，因为这是他的食物。
LEV|22|8|自然死去的或被野兽撕裂的，他不可吃，免得玷污自己。我是耶和华。
LEV|22|9|他们要遵守我的吩咐，免得因亵渎圣物 ，担当自己的罪而死。我是使他们分别为圣的耶和华。
LEV|22|10|“任何外人都不可吃圣物；寄居在祭司家的，或雇工，都不可吃圣物。
LEV|22|11|若是祭司用自己的银钱买来的人，就可以吃圣物；在他家出生的人也可以吃他的食物。
LEV|22|12|祭司的女儿若嫁给外人，就不可吃举祭的圣物。
LEV|22|13|但祭司的女儿若成为寡妇或被休，又没有后裔，她回到父家，好像年轻的时候，就可以吃她父亲的食物。只是任何外人都不可吃它。
LEV|22|14|若有人误吃了圣物，要把圣物加上五分之一交给祭司。
LEV|22|15|祭司不可亵渎 以色列 人献给耶和华的圣物，
LEV|22|16|免得他们因吃圣物而自取罪孽。我是使他们分别为圣的耶和华。”
LEV|22|17|耶和华吩咐 摩西 说：
LEV|22|18|“你要吩咐 亚伦 和他子孙，以及 以色列 众人，对他们说： 以色列 家中的人，或在 以色列 中寄居的 ，若要献供物给耶和华作燔祭，无论是为所许的愿或是甘心献的，
LEV|22|19|就要将一头公的，没有残疾的牛，或绵羊，或山羊献上，这样你们才蒙悦纳。
LEV|22|20|凡有残疾的，你们不可献上，因为这样你们必不蒙悦纳。
LEV|22|21|若有人从牛群或羊群中，将平安祭献给耶和华，无论是为还所许特别的愿，或是甘心献的，所献的必须是健康、无任何残疾的，才蒙悦纳。
LEV|22|22|凡瞎眼的、受伤的、断腿的、溃烂的、长癣的、长疥的，都不可献给耶和华，不可在坛上作为火祭献给耶和华。
LEV|22|23|无论是公牛或小绵羊，若一条腿太长或太短，只可作甘心祭献上；若用来还愿，就不蒙悦纳。
LEV|22|24|凡睾丸损伤，或压碎，或破裂，或阉割的，都不可献给耶和华；不可在你们的地上行这事。
LEV|22|25|从外人的手里得到任何这类的动物，也不可献上作你们上帝的食物；因为它们有缺陷，有残疾，它们必不为你们而蒙悦纳。”
LEV|22|26|耶和华吩咐 摩西 说：
LEV|22|27|“刚出生的公牛，或绵羊，或山羊，七天当跟着它的母亲；从第八天起，可以当供物作为耶和华的火祭，这是蒙悦纳的。
LEV|22|28|无论是牛或羊，不可在同一日宰它和它的小牛小羊。
LEV|22|29|你们宰杀祭牲献感谢祭给耶和华，要献得使你们可蒙悦纳；
LEV|22|30|要在当天吃，一点也不可留到早晨。我是耶和华。
LEV|22|31|“你们要谨守我的诫命，遵行它们。我是耶和华。
LEV|22|32|你们不可亵渎我的圣名；我在 以色列 人中要被尊为圣。我是使你们分别为圣的耶和华，
LEV|22|33|曾把你们从 埃及 地领出来，作你们的上帝。我是耶和华。”
LEV|23|1|耶和华吩咐 摩西 说：
LEV|23|2|“你要吩咐 以色列 人，对他们说：以下是我的节期，是你们要宣告为圣会的耶和华的节期。”
LEV|23|3|“六日要做工，第七日是完全安息的安息日，要有圣会；你们任何工都不可做。这是在你们一切的住处向耶和华当守的安息日。”
LEV|23|4|“以下是你们要按时宣告为圣会的耶和华的节期。”
LEV|23|5|“正月十四日黄昏的时候 ，是向耶和华守的逾越节。
LEV|23|6|这月的十五日是向耶和华守的除酵节；你们要吃无酵饼七日。
LEV|23|7|第一日要有圣会，任何劳动的工都不可做；
LEV|23|8|要将火祭献给耶和华七日。第七日要有圣会，任何劳动的工都不可做。”
LEV|23|9|耶和华吩咐 摩西 说：
LEV|23|10|“你要吩咐 以色列 人，对他们说：你们到了我赐给你们的地，收割庄稼的时候，要把初熟庄稼中的一捆拿来给祭司。
LEV|23|11|他要把这捆在耶和华面前摇一摇，使你们蒙悦纳。祭司要在安息日的次日把这捆摇一摇。
LEV|23|12|摇这捆的那一日，你们要献一只一岁没有残疾的小公绵羊，给耶和华作燔祭。
LEV|23|13|同献的素祭是十分之二伊法调了油的细面，作为献给耶和华馨香的火祭；同献的浇酒祭是四分之一欣酒。
LEV|23|14|无论是饼，是烘熟的谷物，是新穗子，你们都不可吃；直等到你们把这供物带来献给你们上帝的那一天，才可以吃。在你们一切的住处，这要成为你们世世代代永远的定例。”
LEV|23|15|“你们要从安息日的次日，就是献那捆庄稼为摇祭的那日起，计算足足的七个安息日。
LEV|23|16|到第七个安息日的次日，共计五十天，你们要将新的素祭献给耶和华。
LEV|23|17|要从你们的住处取十分之二伊法细面，加酵烤成两个摇祭的饼，作为初熟之物献给耶和华。
LEV|23|18|又要将七只一岁没有残疾的羔羊、一头公牛犊、两只公绵羊和饼一同奉上。这些要和素祭和浇酒祭一同作为燔祭献给耶和华，作馨香的火祭献给耶和华。
LEV|23|19|你们要献一只公山羊为赎罪祭，两只一岁的小公绵羊为平安祭。
LEV|23|20|祭司要把这些和初熟庄稼做成的饼，与两只小公绵羊一同在耶和华面前摇一摇，作为摇祭。这些献给耶和华的圣物是归给祭司的。
LEV|23|21|在这一日，你们要宣告圣会；任何劳动的工都不可做。在你们一切的住处，这要成为你们世世代代永远的定例。
LEV|23|22|“你们在自己的地收割庄稼时，不可割尽田的角落，也不可拾取庄稼所掉落的，要把它们留给穷人和寄居的。我是耶和华－你们的上帝。”
LEV|23|23|耶和华吩咐 摩西 说：
LEV|23|24|“你要吩咐 以色列 人说：七月初一，你们要守为完全安息的日子，要吹角作纪念，当有圣会。
LEV|23|25|任何劳动的工都不可做；要将火祭献给耶和华。”
LEV|23|26|耶和华吩咐 摩西 说：
LEV|23|27|“但是，七月初十是赎罪日；你们要守为圣会，刻苦己心，并要将火祭献给耶和华。
LEV|23|28|在这一日，任何工都不可做；因为这是赎罪日，要在耶和华－你们的上帝面前赎罪。
LEV|23|29|在这一日，凡不刻苦己心的，必从百姓中剪除。
LEV|23|30|凡在这一日做任何工的，我必将他从百姓中除灭。
LEV|23|31|任何工你们都不可做。在你们一切的住处，这要成为你们世世代代永远的定例。
LEV|23|32|你们要守这日为完全安息的安息日，刻苦己心；从这月初九晚上到次日晚上，你们要守为安息日。”
LEV|23|33|耶和华吩咐 摩西 说：
LEV|23|34|“你要吩咐 以色列 人说：这七月十五日是住棚节，要向耶和华守这节七日。
LEV|23|35|第一日当有圣会，任何劳动的工都不可做。
LEV|23|36|要将火祭献给耶和华七日。第八日当守圣会，并要献火祭给耶和华。这是严肃会，任何劳动的工都不可做。
LEV|23|37|“这是耶和华的节期，就是你们要宣告为圣会的节期；要将火祭，就是燔祭、素祭、祭物和浇酒祭，按照每日的规定献给耶和华。
LEV|23|38|除此之外，还有耶和华的安息日，你们献给耶和华的供物，一切的还愿祭，和一切的甘心祭。
LEV|23|39|“但是，从七月十五日起，你们收藏了地的出产之后，要守耶和华的节期七日。第一日为要完全安息，第八日也要完全安息。
LEV|23|40|第一日，你们要拿美好树上的果子、棕树枝、树叶茂密的枝条和河边的柳枝，在耶和华－你们的上帝面前欢乐七日。
LEV|23|41|每年你们要向耶和华守这节七日。你们在七月里所守的节，要成为世世代代永远的定例。
LEV|23|42|你们要住在棚里七日；凡 以色列 家出生的人都要住在棚里，
LEV|23|43|好叫你们世世代代知道，我领 以色列 人出 埃及 地的时候，曾使他们住在棚里。我是耶和华－你们的上帝。”
LEV|23|44|于是， 摩西 向 以色列 人颁布了耶和华的节期。
LEV|24|1|耶和华吩咐 摩西 说：
LEV|24|2|“你要吩咐 以色列 人，把那捣成的纯橄榄油拿来给你，用以点灯，使灯经常点着。
LEV|24|3|在会幕中法柜前的幔子外， 亚伦 从晚上到早晨要在耶和华面前照管这灯。这要成为你们世世代代永远的定例。
LEV|24|4|他要在耶和华面前经常照管纯金 灯台上的灯。”
LEV|24|5|“你要取细面，烤成十二个饼，每个用十分之二伊法。
LEV|24|6|要把饼排成两行 ，每行六个，供在耶和华面前的纯金桌子上。
LEV|24|7|再把纯乳香撒在每行饼上，作为纪念，是献给耶和华为食物的火祭。
LEV|24|8|每个安息日， 亚伦 要把饼不间断地供在耶和华面前。这是 以色列 人永远的约。
LEV|24|9|这饼要归给 亚伦 和他的子孙。他们要在圣处吃这饼，因为在献给耶和华的火祭中，这饼是至圣的，归给他作永远当得的份。”
LEV|24|10|有一个 以色列 妇人的儿子，他父亲是 埃及 人。有一日他出去，到 以色列 人中。这 以色列 妇人的儿子和一个 以色列 人在营里争吵。
LEV|24|11|以色列 妇人的儿子诅咒，亵渎了圣名。有人把他送到 摩西 那里。他的母亲名叫 示罗密 ，是 但 支派 底伯利 的女儿。
LEV|24|12|他们把这人收押在监里，等候耶和华指示的话。
LEV|24|13|耶和华吩咐 摩西 说：
LEV|24|14|“把那诅咒的人带到营外。凡听见的人都要把手放在他头上，全会众要用石头打死他。
LEV|24|15|你要吩咐 以色列 人说：凡诅咒上帝的，必要担当自己的罪。
LEV|24|16|亵渎耶和华名的，必被处死；全会众必须用石头打死他。无论是寄居的，是本地人，他亵渎圣名的时候必被处死。
LEV|24|17|“打死人的，必被处死；
LEV|24|18|打死牲畜的，必赔上牲畜，以命偿命。
LEV|24|19|人若伤害邻舍以致残疾，他怎样做，也要照样向他做：
LEV|24|20|以伤还伤，以眼还眼，以牙还牙。他怎样使人有残疾，也要照样向他做。
LEV|24|21|打死牲畜的，必赔上牲畜；打死人的，必被处死。
LEV|24|22|无论是寄居的，是本地人，都依照同一条例。我是耶和华－你们的上帝。”
LEV|24|23|于是， 摩西 吩咐 以色列 人，他们就把那诅咒的人带到营外，用石头打死。 以色列 人就照耶和华所吩咐 摩西 的做了。
LEV|25|1|耶和华在 西奈山 吩咐 摩西 说：
LEV|25|2|“你要吩咐 以色列 人，对他们说：你们到了我所赐你们那地的时候，地要休耕，向耶和华守安息。
LEV|25|3|你们六年要耕种田地，六年要修整葡萄园，收藏地的出产。
LEV|25|4|第七年，地要守完全安息的安息年，就是向耶和华守安息。你们不可耕种田地，也不可修整葡萄园。
LEV|25|5|不可收割自然生长的庄稼，也不可摘取没有修剪的葡萄树上的葡萄。这年，地要完全安息。
LEV|25|6|地在安息年所长出的，要给你和你的奴仆、使女、雇工，以及寄居在你那里的外人作食物。
LEV|25|7|所有的出产也要给你的牲畜和你地上的走兽作食物。”
LEV|25|8|“你要计算七个安息年，就是七个七年。这就成为你的七个安息年，一共四十九年。
LEV|25|9|七月初十，你要大声吹角；这是赎罪日，你要在全地吹角。
LEV|25|10|你们要以第五十年为圣年，在全地向所有的居民宣告自由。这是你们的禧年，各人的产业要归还自己，各人要归回自己的家。
LEV|25|11|第五十年要作为你们的禧年。你们不可耕种，不可收割自然生长的庄稼，也不可摘取没有修剪的葡萄树上的葡萄。
LEV|25|12|因为这是禧年，是你们的圣年；你们要吃地中自然生长的农作物。
LEV|25|13|“这禧年，你们各人的产业要归还自己。
LEV|25|14|无论你卖什么给邻舍，或从邻舍的手中买什么，彼此不可亏负。
LEV|25|15|你要按照禧年后的年数向邻舍买；他要按照可收成的年数卖给你；
LEV|25|16|年数越多，价钱就越高；年数越少，价钱就越低，因为他卖给你的是收成的数量。
LEV|25|17|你们彼此不可亏负，只要敬畏你的上帝，因为我是耶和华－你们的上帝。”
LEV|25|18|“你们要遵行我的律例，谨守我的典章，遵行它们，就可以在那地上安然居住。
LEV|25|19|地必出产果实，你们可以吃饱，在那地上安然居住。
LEV|25|20|你们若说：‘看哪，第七年我们不耕种，也不收藏农作物，我们吃什么呢？’
LEV|25|21|我必在第六年发令赐福给你们，地就长出三年的农作物来。
LEV|25|22|第八年你们要耕种，也要吃陈粮；等到第九年农作物收成的时候，你们还有陈粮吃。”
LEV|25|23|“地不可以卖断，因为地是我的；你们在我面前是客旅，是寄居的。
LEV|25|24|在你们所得为业的全地，要准许人有权将地赎回。
LEV|25|25|“你的弟兄若渐渐贫穷，卖了他的一些产业，他的至亲就要来把弟兄所卖的赎回。
LEV|25|26|若没有人能为他赎回，他的手头渐渐宽裕，能够赎回，
LEV|25|27|就要计算卖后的年数，把剩余年数的价钱归还给那买主，他的地业便归还自己。
LEV|25|28|若他手头的财力不够赎回，所卖的地就要留在买主的手里，直到禧年。到了禧年，地业要归还卖主。
LEV|25|29|“人若卖城墙内的住宅，卖了以后，一整年内他有权赎回；这是他可以赎回的期限。
LEV|25|30|若他在一整年内不赎回，这有墙之城的房屋就确定永归买主，直到世世代代；在禧年也不必归还。
LEV|25|31|但周围无城墙之村庄的房屋，要看为乡下的田地，可以赎回；到了禧年就要归还。
LEV|25|32|至于 利未 人所得为业的城镇， 利未 人可以随时赎回他们城镇中的房屋。
LEV|25|33|在所得为业的城镇， 利未 人若卖了房屋，又不赎回，到了禧年仍要归还原主，因为 利未 人城镇的房屋是他们在 以色列 人中的产业。
LEV|25|34|但是 利未 人各城郊外之地是不可卖的，因为这是他们永远的产业。”
LEV|25|35|“你的弟兄在你那里若渐渐贫穷，手头缺乏，你就要帮补他，使他与你一同生活，像外人和寄居的一样。
LEV|25|36|不可向他取利息，也不可向他索取高利；要敬畏你的上帝，使你的弟兄与你一同生活。
LEV|25|37|你不可为了利息借钱给他，也不可为了高利而借粮。
LEV|25|38|我是耶和华－你们的上帝，曾领你们从 埃及 地出来，为要把 迦南 地赐给你们，要作你们的上帝。
LEV|25|39|“你的弟兄在你那里若渐渐贫穷，将自己卖给你，你不可叫他像奴仆服事你。
LEV|25|40|他在你那里要像雇工和寄居的，服事你直到禧年。
LEV|25|41|他和他儿女要离开你，一同出去，归回自己的家，回到他祖宗的地业去。
LEV|25|42|因为他们是我的仆人，是我从 埃及 地领出来的。他们不可被卖为奴仆。
LEV|25|43|不可苛刻管辖他，只要敬畏你的上帝。
LEV|25|44|至于你所要的奴仆和使女，可以来自你们四围的列国，你们可以从他们中买奴仆和使女。
LEV|25|45|那些寄居在你们中间的外人和他们的家属，就是在你们地上所生的，你们可以从其中买人；他们要作你们的产业。
LEV|25|46|你们可以把他们遗留给你们后代的子孙，作为永远继承的产业；你们可以使他们作奴仆。至于你们的弟兄 以色列 人，你们彼此不可苛刻管辖。
LEV|25|47|“住在你那里的外人或寄居的，若手头渐渐宽裕，你的弟兄却渐渐贫穷，将自己卖给那外人或寄居的，或外人家族的一支，
LEV|25|48|卖了以后，有权把自己赎回。他弟兄中的一位可以把他赎回。
LEV|25|49|他的叔伯或叔伯的儿子可以赎他。他家族中的骨肉之亲也可以赎他。他自己若手头渐渐宽裕，也可以赎回自己。
LEV|25|50|他要跟买主计算，从卖自己的那年起，算到禧年；所卖的价钱要按照年数计算，就是雇工跟买主在一起的日子。
LEV|25|51|若剩余的年数多，就要按着年数从买价中偿还他的赎价。
LEV|25|52|若到禧年只剩下几年，就要按着年数跟买主计算，偿还他的赎价。
LEV|25|53|他和买主同住，要像按年雇用的工人，买主不可苛刻管辖他。
LEV|25|54|他若不这样被赎，到了禧年，仍要和他的儿女一同出去。
LEV|25|55|因为 以色列 人都是我的仆人，他们是我的仆人，是我领他们从 埃及 地出来的。我是耶和华－你们的上帝。”
LEV|26|1|“你们不可为自己造虚无的神明，不可竖立雕刻的偶像或柱像，也不可在你们的地上安放石像，向它跪拜，因为我是耶和华－你们的上帝。
LEV|26|2|你们要谨守我的安息日，敬畏我的圣所。我是耶和华。
LEV|26|3|“你们若遵行我的律例，谨守我的诫命，实行它们，
LEV|26|4|我必按时降雨给你们，使地长出农作物，田野的树结出果实。
LEV|26|5|你们打谷物要打到摘葡萄的时候，摘葡萄要摘到播种的时候。你们要吃粮食得饱足，在你们的地上安然居住。
LEV|26|6|我要赐平安在地上；你们躺卧，无人惊吓。我要使你们地上的恶兽消灭，刀剑必不穿越你们的地。
LEV|26|7|你们要追赶仇敌，他们必倒在你们刀下。
LEV|26|8|你们五个人要追赶一百人，一百人要追赶一万人；仇敌必在你们面前倒在刀下。
LEV|26|9|我要眷顾你们，使你们生养众多，也要与你们坚立我的约。
LEV|26|10|你们要吃储存的陈粮，又要为新粮清理陈粮。
LEV|26|11|我要在你们中间立我的帐幕，我的心也不厌恶你们。
LEV|26|12|我要行走在你们中间，作你们的上帝，你们要作我的子民。
LEV|26|13|我是耶和华－你们的上帝，曾将你们从 埃及 地领出来，使你们不再作 埃及 人的奴仆；我曾折断你们所负的轭，使你们挺身前行。”
LEV|26|14|“你们若不听从我，不遵行我这一切的诫命，
LEV|26|15|厌弃我的律例，心中厌恶我的典章，不遵行我一切的诫命，背弃了我的约，
LEV|26|16|我就要这样对待你们：我必使惊惶临到你们，使你们患痨病，害热病，以致眼睛失明，身体衰弱。你们要白白撒种，因为仇敌要吃尽你们所种的。
LEV|26|17|我要向你们变脸，使你们败在仇敌的面前。恨恶你们的必管辖你们；无人追赶，你们却要逃跑。
LEV|26|18|如果这样，你们还不听从我，我就要因你们的罪，加重七倍惩罚你们。
LEV|26|19|我必粉碎你们因势力而有的骄傲，又要使你们的天坚如铁，地硬如铜。
LEV|26|20|你们劳力却白费，因为你们的地没有出产，地上的树也不结果实。
LEV|26|21|“你们行事若与我作对，不肯听从我，我就要因你们的罪，加重七倍灾祸击打你们。
LEV|26|22|我要打发野地的走兽到你们中间，夺去你们的儿女，吞灭你们的牲畜，使你们人数减少，道路荒凉。
LEV|26|23|“如果这样，你们还不接受管教归向我，行事与我作对，
LEV|26|24|我就要行事与你们作对，因你们的罪，加重七倍击打你们。
LEV|26|25|我要使刀剑临到你们，报复你们的背约。你们若被赶入城中，我要降瘟疫在你们中间，把你们交在仇敌手中。
LEV|26|26|我要断绝你们粮食的供应 ，使十个女人用一个烤炉给你们烤饼，按配给的定量秤给你们。你们要吃，却吃不饱。
LEV|26|27|“如果这样，你们还不听从我，行事与我作对，
LEV|26|28|我就要向你们发烈怒，行事与你们作对，因你们的罪，加重七倍惩罚你们。
LEV|26|29|你们要吃你们儿子的肉，也要吃你们女儿的肉。
LEV|26|30|我要摧毁你们的丘坛，砍掉你们的香坛，把你们的尸首扔在你们偶像的残骸上。我的心也必厌恶你们，
LEV|26|31|使你们的城镇变成废墟，你们的众圣所变荒凉，我也不闻你们芬芳的香气。
LEV|26|32|我要使这地变荒凉，甚至占领这地的敌人都惊讶。
LEV|26|33|我要把你们驱散到列国中，也要拔刀追赶你们。你们的地要成为荒凉，你们的城镇要变成废墟。
LEV|26|34|“当你们在敌人之地的时候，你们的地要在一切荒凉的日子重享安息；在那时候，地要休息，重享安息。
LEV|26|35|地在一切荒凉的日子都要安息，这是你们住在其上的时候所不能得的安息。
LEV|26|36|至于你们幸存的人，我要使他们在敌人之地心中惊慌，甚至风吹落叶的声音也把他们吓跑。他们要逃避，像人逃避刀剑，虽无人追赶，却要跌倒。
LEV|26|37|虽然无人追赶，他们却要彼此绊倒，像逃避刀剑一样。你们在仇敌面前必站立不住。
LEV|26|38|你们要在列国中灭亡，敌人之地要吞灭你们，
LEV|26|39|你们幸存的人必因自己的罪孽在敌人之地衰残，也要因祖先的罪孽衰残。
LEV|26|40|“他们要承认自己的罪孽和祖先的罪孽，就是背叛我，行事与我作对的过犯。
LEV|26|41|我也行事与他们作对，把他们遣送到敌人之地。那时，他们未受割礼的心若肯谦卑，也服了罪孽的惩罚，
LEV|26|42|我就要记念我与 雅各 的约，记念我与 以撒 的约，与 亚伯拉罕 的约；我也要记念这地。
LEV|26|43|地被他们离弃，因他们不在而荒凉的时候，就要重享安息。他们服了罪孽的惩罚，因为他们厌弃我的典章，心中厌恶我的律例。
LEV|26|44|虽然如此，当他们在敌人之地时，我却不厌弃他们，不厌恶他们，将他们全然灭绝，也不背弃我与他们的约，因为我是耶和华－他们的上帝。
LEV|26|45|我要为他们的缘故记念我与他们祖先的约；我在列国眼前曾把他们的祖先从 埃及 地领出来，为要作他们的上帝。我是耶和华。”
LEV|26|46|这些律例、典章和法度是耶和华在 西奈山 上藉着 摩西 与 以色列 人立的。
LEV|27|1|耶和华吩咐 摩西 说：
LEV|27|2|“你要吩咐 以色列 人，对他们说：人向耶和华许特别的愿，要按照你所估一个人的价钱。
LEV|27|3|你所估的是：二十岁到六十岁男的，按照圣所的舍客勒，估价是五十舍客勒银子。
LEV|27|4|若是女的，估价是三十舍客勒。
LEV|27|5|五岁到二十岁男的，估价是二十舍客勒，女的十舍客勒。
LEV|27|6|一个月到五岁男的，估价是五舍客勒，女的三舍客勒。
LEV|27|7|六十岁以上男的，估价是十五舍客勒，女的十舍客勒。
LEV|27|8|他若贫穷，不能按照你的估价，就要把他带到祭司面前，让祭司为他估价；祭司要按许愿者手头财力所及估价。
LEV|27|9|“许愿要献给耶和华的供物若是牲畜，凡这类献给耶和华的都要成为圣。
LEV|27|10|不可更换，也不可用另一只取代，无论是好的换坏的，或是坏的换好的，都不可。若一定要以牲畜取代牲畜，所许的与所取代的都要成为圣。
LEV|27|11|若牲畜不洁净，不可献给耶和华为供物，就要把牲畜带到祭司面前。
LEV|27|12|祭司要估价；牲畜是好是坏，祭司怎样估定，就是你的估价。
LEV|27|13|许愿者若一定要把它赎回，就要在你的估价上加五分之一。
LEV|27|14|“人将房屋分别为圣，归给耶和华为圣，祭司就要估价。房屋是好是坏，祭司怎样估定，就要以他的估价为准。
LEV|27|15|将房屋分别为圣的人，若要赎回房屋，必须付你所估定的价钱，再加上五分之一，房屋才可以归还给他。
LEV|27|16|“人若将所继承的一块田地分别为圣，归给耶和华，就要按照这地撒种多少来估价；能撒一贺梅珥大麦种子的，是五十舍客勒银子。
LEV|27|17|他若从禧年起将地分别为圣，就要以你的估价为准。
LEV|27|18|倘若他在禧年以后将地分别为圣，祭司就要按照从那时到下一个禧年所剩的年数推算，从你的估价中减掉。
LEV|27|19|将地分别为圣的人若要把地赎回，必须付你所估定的价钱，再加上五分之一，地才可以归还给他。
LEV|27|20|他若不赎回那地，或是将地卖给别人，就不能再赎了。
LEV|27|21|到了禧年，那田地要从买主手中退还，归耶和华为圣，和永献的地一样，要归祭司为业。
LEV|27|22|若分别为圣归耶和华的田地不是继承的，而是买来的，
LEV|27|23|祭司就要依照你的估价，推算到禧年。当天，这人要将你所估的归给耶和华为圣。
LEV|27|24|到了禧年，那田地要退还给卖主，就是继承那地的原主。
LEV|27|25|凡你所估的价钱都要按照圣所的舍客勒：二十季拉是一舍客勒。
LEV|27|26|“头生的，就是牲畜中头生属耶和华的，人不可再将它分别为圣，无论是牛是羊都是耶和华的。
LEV|27|27|头生的牲畜若是不洁净的，就要按照所估定的价钱，再加上五分之一，把它赎回。若不赎回，就要按照你的估价把它卖了。
LEV|27|28|“但一切永献作当灭的，就是人从他所有永献给耶和华作当灭的，无论是人，是牲畜，是他继承的田地，都不可卖，也不可赎。凡永献作当灭的都归耶和华为至圣。
LEV|27|29|凡从人中永献作当灭的都不可赎，必被处死。
LEV|27|30|“地上所有的，无论是地上的种子，是树上的果子，十分之一是耶和华的，是归耶和华为圣的。
LEV|27|31|人若要赎回这十分之一，就要另加五分之一。
LEV|27|32|凡牛群羊群中的十分之一，就是一切从牧人杖下经过的，每第十只要归耶和华为圣。
LEV|27|33|不可追究是好是坏，也不可取代；若一定要取代，所取代的和本来当献的牲畜都要成为圣，不可赎回。”
LEV|27|34|这些是耶和华在 西奈山 为 以色列 人所吩咐 摩西 的命令。
NUM|1|1|以色列 人出 埃及 地后第二年二月初一，耶和华在 西奈 旷野，在会幕中吩咐 摩西 说：
NUM|1|2|“你要按宗族、父家、人名的数目计算 以色列 全会众，数点所有的男丁。
NUM|1|3|以色列 中凡二十岁以上能出去打仗的，你和 亚伦 要按照他们的队伍数点。
NUM|1|4|每支派要有一个人，就是父家的家长跟你们一起。
NUM|1|5|这是帮助你们的人的名字： 属 吕便 的， 示丢珥 的儿子 以利蓿 ；
NUM|1|6|属 西缅 的， 苏利沙代 的儿子 示路蔑 ；
NUM|1|7|属 犹大 的， 亚米拿达 的儿子 拿顺 ；
NUM|1|8|属 以萨迦 的， 苏押 的儿子 拿坦业 ；
NUM|1|9|属 西布伦 的， 希伦 的儿子 以利押 ；
NUM|1|10|约瑟 子孙、属 以法莲 的， 亚米忽 的儿子 以利沙玛 ；属 玛拿西 的， 比大蓿 的儿子 迦玛列 ；
NUM|1|11|属 便雅悯 的， 基多尼 的儿子 亚比但 ；
NUM|1|12|属 但 的， 亚米沙代 的儿子 亚希以谢 ；
NUM|1|13|属 亚设 的， 俄兰 的儿子 帕结 ；
NUM|1|14|属 迦得 的， 丢珥 的儿子 以利雅萨 ；
NUM|1|15|属 拿弗他利 的， 以南 的儿子 亚希拉 。”
NUM|1|16|这些是从会众中选出来的父系支派的领袖，是 以色列 部队的官长。
NUM|1|17|于是， 摩西 和 亚伦 带着这些按名指定的人，
NUM|1|18|在二月初一召集全会众。会众就照他们的宗族、父家、人名的数目，登记二十岁以上的人口。
NUM|1|19|耶和华怎样吩咐 摩西 ，他就照样在 西奈 的旷野数点他们。
NUM|1|20|以色列 的长子， 吕便 子孙的后代，照着宗族、父家、人名的数目，他们的人口凡二十岁以上能出去打仗的男丁，
NUM|1|21|吕便 支派被数的共有四万六千五百名。
NUM|1|22|西缅 子孙的后代，照着宗族、父家、被数 人名的数目，他们的人口凡二十岁以上能出去打仗的男丁，
NUM|1|23|西缅 支派被数的共有五万九千三百名。
NUM|1|24|迦得 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|25|迦得 支派被数的共有四万五千六百五十名。
NUM|1|26|犹大 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|27|犹大 支派被数的共有七万四千六百名。
NUM|1|28|以萨迦 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|29|以萨迦 支派被数的共有五万四千四百名。
NUM|1|30|西布伦 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|31|西布伦 支派被数的共有五万七千四百名。
NUM|1|32|约瑟 子孙属 以法莲 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|33|以法莲 支派被数的共有四万零五百名。
NUM|1|34|玛拿西 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|35|玛拿西 支派被数的共有三万二千二百名。
NUM|1|36|便雅悯 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|37|便雅悯 支派被数的共有三万五千四百名。
NUM|1|38|但 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|39|但 支派被数的共有六万二千七百名。
NUM|1|40|亚设 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|41|亚设 支派被数的共有四万一千五百名。
NUM|1|42|拿弗他利 子孙的后代，照着宗族、父家、人名的数目，凡二十岁以上能出去打仗的，
NUM|1|43|拿弗他利 支派被数的共有五万三千四百名。
NUM|1|44|这些就是被数点的，是 摩西 、 亚伦 和 以色列 十二个领袖所数点的；每一个领袖代表他们的父家。
NUM|1|45|以色列 人被数点的总数， 以色列 中照着父家，凡二十岁以上能出去打仗的，
NUM|1|46|他们被数点的总数是六十万三千五百五十名。
NUM|1|47|利未 人却没有按照父系支派数在其中。
NUM|1|48|耶和华吩咐 摩西 说：
NUM|1|49|“惟独 利未 支派你不可数点，也不可在 以色列 人中计算他们的人口。
NUM|1|50|你要派 利未 人管理法柜的帐幕和其中一切的器具，以及属帐幕的一切。他们要抬帐幕和其中一切的器具，并要办理帐幕的事务，在帐幕的四围安营。
NUM|1|51|帐幕将往前行的时候， 利未 人要拆卸；将驻扎的时候， 利未 人要支搭帐幕。近前来的外人必被处死。
NUM|1|52|以色列 人要按照各自的队伍安营，各归本营，各归本旗。
NUM|1|53|但 利未 人要在法柜帐幕的四围安营，免得愤怒临到 以色列 会众； 利未 人要负责看守法柜的帐幕。”
NUM|1|54|以色列 人就这样做了。凡耶和华所吩咐 摩西 的，他们都照样做了。
NUM|2|1|耶和华吩咐 摩西 和 亚伦 说：
NUM|2|2|“ 以色列 人各人要在自己的旗帜下，按照自己父家的旗号安营，对着会幕的四围安营。
NUM|2|3|“在东边，向日出的方向， 犹大 营按照他们的队伍，在它的旗帜下安营。 犹大 人的领袖是 亚米拿达 的儿子 拿顺 ，
NUM|2|4|他的军队被数的有七万四千六百名。
NUM|2|5|在他旁边安营的是 以萨迦 支派。 以萨迦 人的领袖是 苏押 的儿子 拿坦业 ，
NUM|2|6|他的军队被数的有五万四千四百名。
NUM|2|7|还有 西布伦 支派， 西布伦 人的领袖是 希伦 的儿子 以利押 ，
NUM|2|8|他的军队被数的有五万七千四百名。
NUM|2|9|凡属 犹大 营，照他们队伍被数的共有十八万六千四百名；他们要作第一队往前行。
NUM|2|10|“在南边，按照他们的队伍是 吕便 营的旗帜。 吕便 人的领袖是 示丢珥 的儿子 以利蓿 ，
NUM|2|11|他的军队被数的有四万六千五百名。
NUM|2|12|在他旁边安营的是 西缅 支派。 西缅 人的领袖是 苏利沙代 的儿子 示路蔑 ，
NUM|2|13|他的军队被数的有五万九千三百名。
NUM|2|14|还有 迦得 支派， 迦得 人的领袖是 丢珥 的儿子 以利雅萨 ，
NUM|2|15|他的军队被数的有四万五千六百五十名。
NUM|2|16|凡属 吕便 营，照他们队伍被数的共有十五万一千四百五十名；他们要作第二队往前行。
NUM|2|17|“会幕与 利未 营在诸营中间往前行。他们怎样安营就怎样往前行，各按本位，各归本旗。
NUM|2|18|“在西边，按照他们的队伍是 以法莲 营的旗帜。 以法莲 人的领袖是 亚米忽 的儿子 以利沙玛 ，
NUM|2|19|他的军队被数的有四万零五百名。
NUM|2|20|在他旁边的是 玛拿西 支派。 玛拿西 人的领袖是 比大蓿 的儿子 迦玛列 ，
NUM|2|21|他的军队被数的有三万二千二百名。
NUM|2|22|还有 便雅悯 支派， 便雅悯 人的领袖是 基多尼 的儿子 亚比但 ，
NUM|2|23|他的军队被数的有三万五千四百名。
NUM|2|24|凡属 以法莲 营，照他们队伍被数的共有十万八千一百名；他们要作第三队往前行。
NUM|2|25|“在北边，按照他们的队伍是 但 营的旗帜。 但 人的领袖是 亚米沙代 的儿子 亚希以谢 ，
NUM|2|26|他的军队被数的有六万二千七百名。
NUM|2|27|在他旁边安营的是 亚设 支派。 亚设 人的领袖是 俄兰 的儿子 帕结 ，
NUM|2|28|他的军队被数的有四万一千五百名。
NUM|2|29|还有 拿弗他利 支派， 拿弗他利 人的领袖是 以南 的儿子 亚希拉 ，
NUM|2|30|他的军队被数的有五万三千四百名。
NUM|2|31|凡属 但 营被数的共有十五万七千六百名；他们随着自己的旗帜行在最后。”
NUM|2|32|以上是 以色列 人按照各自的父家被数的，在诸营中按照各自的队伍被数的，共有六十万三千五百五十名。
NUM|2|33|但 利未 人没有数在 以色列 人中，正如耶和华所吩咐 摩西 的。
NUM|2|34|以色列 人就照着耶和华所吩咐 摩西 的做了，在各自的旗帜下安营，随着各自的宗族、父家起行。
NUM|3|1|耶和华在 西奈山 与 摩西 说话的日子， 亚伦 和 摩西 的后代如下：
NUM|3|2|这些是 亚伦 儿子的名字，长子 拿答 ，及 亚比户 、 以利亚撒 、 以他玛 。
NUM|3|3|这些是 亚伦 儿子的名字，都是受膏的祭司，是 摩西 授圣职使他们担任祭司职分的。
NUM|3|4|拿答 、 亚比户 在 西奈 的旷野向耶和华献上凡火的时候，死在耶和华面前。他们没有儿子。 以利亚撒 和 以他玛 在他们的父亲 亚伦 面前担任祭司的职分。
NUM|3|5|耶和华吩咐 摩西 说：
NUM|3|6|“你要带 利未 支派近前来，站在 亚伦 祭司面前伺候他。
NUM|3|7|他们要替他，又替全会众，在会幕前执行任务，办理帐幕的事。
NUM|3|8|他们要看守会幕一切的器具，为 以色列 人执行任务，办理帐幕的事。
NUM|3|9|你要把 利未 人给 亚伦 和他的儿子；他们是从 以色列 人中选出来完全给他的。
NUM|3|10|你要指派 亚伦 和他的儿子谨守祭司的职分；近前来的外人必被处死。”
NUM|3|11|耶和华吩咐 摩西 说：
NUM|3|12|“看哪，我从 以色列 人中选了 利未 人，代替 以色列 人中所有头胎的长子； 利未 人要归我。
NUM|3|13|因为凡头生的是我的；我在 埃及 地击杀所有头生的那日，就把 以色列 中所有头生的，无论是人或牲畜，都分别为圣归我；他们定要属我。我是耶和华。”
NUM|3|14|耶和华在 西奈 的旷野吩咐 摩西 说：
NUM|3|15|“你要照父家、宗族计算 利未 人。凡一个月以上的男子都要数点。”
NUM|3|16|于是 摩西 遵照耶和华的吩咐，按所指示的数点他们。
NUM|3|17|利未 儿子的名字是 革顺 、 哥辖 、 米拉利 。
NUM|3|18|按照宗族， 革顺 儿子的名字是 立尼 、 示每 。
NUM|3|19|按照宗族， 哥辖 的儿子是 暗兰 、 以斯哈 、 希伯伦 、 乌薛 。
NUM|3|20|按照宗族， 米拉利 的儿子是 抹利 、 母示 。按照父家，这些都是 利未 人的宗族。
NUM|3|21|属 革顺 的有 立尼 族、 示每 族，他们是 革顺 人的宗族。
NUM|3|22|他们被数的，一个月以上所有男子的数目共有七千五百名。
NUM|3|23|这 革顺 人的宗族要在西边，在帐幕后面安营。
NUM|3|24|革顺 人父家的领袖是 拉伊勒 的儿子 以利雅萨 。
NUM|3|25|革顺 的子孙在会幕中要看守的是帐幕、罩棚、罩棚的盖、会幕的门帘、
NUM|3|26|帐幕和祭坛周围院子的帷幔和门帘，以及所有需用的绳子。
NUM|3|27|属 哥辖 的有 暗兰 族、 以斯哈 族、 希伯伦 族、 乌薛 族，他们是 哥辖 人的宗族。
NUM|3|28|一个月以上所有男子的数目共有八千六百 名；他们负责看守圣所。
NUM|3|29|哥辖 子孙的宗族要在帐幕的南边安营。
NUM|3|30|哥辖 人父家宗族的领袖是 乌薛 的儿子 以利撒反 。
NUM|3|31|他们要看守的是约柜、供桌、灯台、祭坛、香坛、祭司在圣所内用的器皿、帘子，与一切相关事奉的物件。
NUM|3|32|亚伦 祭司的儿子 以利亚撒 是 利未 人众领袖的主管，他要监督那些负责看守圣所的人。
NUM|3|33|属 米拉利 的有 抹利 族、 母示 族，他们是 米拉利 的宗族。
NUM|3|34|他们被数的，一个月以上所有男子的数目共有六千二百名。
NUM|3|35|米拉利 宗族的领袖是 亚比亥 的儿子 苏列 ，他们要在帐幕的北边安营。
NUM|3|36|米拉利 子孙的职分是看守帐幕的竖板、横木、柱子、带卯眼的座和一切的器具，就是一切相关事奉的物件，
NUM|3|37|以及院子四围的柱子、其上带卯眼的座、橛子和绳子。
NUM|3|38|在帐幕前东边，向日出的方向，安营的是 摩西 、 亚伦 和 亚伦 的儿子。他们负责看守圣所，是为 以色列 人看守的。近前来的外人必被处死。
NUM|3|39|凡被数的 利未 人，就是 摩西 、 亚伦 照耶和华所指示、按宗族所数的，一个月以上所有的男子共有二万二千名。
NUM|3|40|耶和华对 摩西 说：“你要数点 以色列 人中凡一个月以上头生的男子，登记他们的名字。
NUM|3|41|我是耶和华。你要拣选 利未 人归我，代替所有头生的 以色列 人，也取 利未 人的牲畜代替 以色列 人所有头生的牲畜。”
NUM|3|42|摩西 就遵照耶和华所吩咐的，把所有 以色列 人头生的都数点了。
NUM|3|43|按人名的数目，凡一个月以上头生的男子共有二万二千二百七十三名。
NUM|3|44|耶和华吩咐 摩西 说：
NUM|3|45|“你要拣选 利未 人代替所有头生的 以色列 人，也要取 利未 人的牲畜代替 以色列 人的牲畜。 利未 人要归我，我是耶和华。
NUM|3|46|以色列 人头生的男子比 利未 人多了二百七十三名，必须把他们赎出来；
NUM|3|47|按照人丁，照圣所的舍客勒，每人当付五舍客勒，一舍客勒是二十季拉。
NUM|3|48|你要把这些多出来的人的赎银交给 亚伦 和他的儿子。”
NUM|3|49|于是 摩西 从那被 利未 人所赎以外多出来的人取了赎银。
NUM|3|50|从头生的 以色列 人所取的银子，按照圣所的舍客勒，共计一千三百六十五舍客勒。
NUM|3|51|摩西 遵照耶和华指示的话，把赎银交给 亚伦 和他的儿子，正如耶和华所吩咐的。
NUM|4|1|耶和华吩咐 摩西 和 亚伦 说：
NUM|4|2|“你要照宗族、父家计算 利未 人中 哥辖 子孙的人口，
NUM|4|3|就是从三十岁到五十岁，凡前来任职，在会幕里事奉的人。
NUM|4|4|这是 哥辖 子孙在会幕里有关至圣之物的职责。
NUM|4|5|“拔营的时候， 亚伦 和他儿子要进去，把遮掩的幔子取下，用它来遮盖法柜，
NUM|4|6|又用精美皮料盖在上面，铺上纯蓝色的布，再把杠穿上。
NUM|4|7|他们要用蓝色的布铺在供饼的桌上，将盘、碟，以及浇酒祭的杯和壶摆在上面；经常供的饼也要留在桌上。
NUM|4|8|他们要在这些东西的上面铺上朱红色的布，把精美皮料盖在上面，再把杠穿上。
NUM|4|9|他们要用蓝色的布遮盖供职用的灯台、灯台上的灯盏、灯剪、灯盘，以及所有盛油的器皿；
NUM|4|10|又要用精美皮料把灯台和灯台的一切器具包好，放在抬架上。
NUM|4|11|他们要用蓝色的布铺在金坛上，用精美皮料盖在上面，再把杠穿上。
NUM|4|12|要用蓝色的布把圣所供职用的一切器具包好，再用精美皮料盖在上面，放在抬架上。
NUM|4|13|他们要清理祭坛上的灰，用紫色的布铺在坛上；
NUM|4|14|又要把供职用的一切器具，就是祭坛一切的器具，火盆、肉叉、铲子和盘子，都摆在坛上，铺上精美皮料，再把杠穿上。
NUM|4|15|“拔营的时候， 亚伦 和他儿子把圣所和圣所一切的器具盖好之后， 哥辖 的子孙才好来抬，免得他们摸圣物而死；这是 哥辖 子孙在会幕里所当抬的。
NUM|4|16|“祭司 亚伦 的儿子 以利亚撒 所要照管的是点灯的油和香料，以及常献的素祭和膏油。他要照管整个帐幕和其中所有的，以及圣所和圣所的器具。”
NUM|4|17|耶和华吩咐 摩西 和 亚伦 说：
NUM|4|18|“你们不可使 哥辖 人宗族的这一支从 利未 人中剪除。
NUM|4|19|他们挨近至圣之物的时候，要向他们这样做，使他们存活，不致死亡； 亚伦 和他的儿子要进去，分派各人当做的，当抬的。
NUM|4|20|但是他们不可进去观看圣所的拆卸 ，免得死亡。”
NUM|4|21|耶和华吩咐 摩西 说：
NUM|4|22|“你要照父家、宗族计算 革顺 子孙的人口；
NUM|4|23|从三十岁到五十岁，凡前来任职，在会幕里事奉的，都要数点。
NUM|4|24|这是 革顺 人宗族的职责，要做的事，要抬的东西如下：
NUM|4|25|他们要抬帐幕的幔子、会幕和会幕的盖、外层精美皮料的盖、会幕的门帘、
NUM|4|26|帐幕和祭坛周围院子的帷幔和门帘、绳子，以及所有需用的器具；一切与这些东西相关的事务，他们要尽职。
NUM|4|27|革顺 人的子孙一切的事奉，就是所当抬的，所当做的，都要遵照 亚伦 和他儿子的指示；他们所当抬的，你们要派他们负责。
NUM|4|28|这是 革顺 人子孙的宗族在会幕里的事奉；他们要在 亚伦 祭司的儿子 以他玛 的手下尽职。”
NUM|4|29|“至于 米拉利 的子孙，你要照宗族、父家数点他们；
NUM|4|30|从三十岁到五十岁，凡前来任职，在会幕里事奉的，你都要数点。
NUM|4|31|这是他们在会幕里的事奉，他们负责要抬的是帐幕的竖板、横木、柱子和带卯眼的座，
NUM|4|32|院子四围的柱子和其上带卯眼的座、橛子、绳子和一切的器具，与一切相关事奉的物件。你们要按名指定他们要抬的器具。
NUM|4|33|这是 米拉利 子孙的宗族在会幕里的事奉，都在 亚伦 祭司的儿子 以他玛 的手下。”
NUM|4|34|摩西 、 亚伦 和会众的领袖按照宗族、父家数点 哥辖 人的子孙；
NUM|4|35|从三十岁到五十岁，凡前来任职，在会幕里事奉的，
NUM|4|36|按照宗族被数的共有二千七百五十名。
NUM|4|37|这是所有在会幕里事奉的 哥辖 人宗族中被数的，是 摩西 和 亚伦 遵照耶和华藉 摩西 所指示数点的。
NUM|4|38|革顺 子孙被数的，按照宗族、父家，
NUM|4|39|从三十岁到五十岁，凡前来任职，在会幕里事奉的，
NUM|4|40|按照宗族、父家被数的共有二千六百三十名。
NUM|4|41|这是所有在会幕里事奉的 革顺 子孙宗族中被数的，是 摩西 和 亚伦 遵照耶和华的指示所数点的。
NUM|4|42|米拉利 子孙宗族被数的，按照宗族、父家，
NUM|4|43|从三十岁到五十岁，凡前来任职，在会幕里事奉的，
NUM|4|44|按照宗族被数的共有三千二百名。
NUM|4|45|这是 米拉利 子孙宗族中被数的，是 摩西 和 亚伦 遵照耶和华藉 摩西 所指示数点的。
NUM|4|46|摩西 、 亚伦 和 以色列 领袖按照宗族、父家数点 利未 人，
NUM|4|47|从三十岁到五十岁，凡前来任职，在会幕里事奉，做抬物之工的，
NUM|4|48|他们被数的共有八千五百八十名。
NUM|4|49|按照耶和华藉 摩西 所指示的来分派，各人都有自己所做的事、所抬的物；他们就这样被数点，正如耶和华所吩咐 摩西 的。
NUM|5|1|耶和华吩咐 摩西 说：
NUM|5|2|“你要吩咐 以色列 人，把一切患痲疯 的、患漏症的和因尸体而不洁净的，都送到营外去。
NUM|5|3|无论男女你都要送，把他们送到营外，免得他们玷污了他们的营，这是我住在他们中间的地方。”
NUM|5|4|以色列 人就照样做，把他们送到营外去。耶和华怎样吩咐 摩西 ， 以色列 人就照样做了。
NUM|5|5|耶和华吩咐 摩西 说：
NUM|5|6|“你要吩咐 以色列 人：无论男女，若犯了人所常犯的任何罪 ，以致干犯耶和华，那人就有了罪。
NUM|5|7|他要承认所犯的罪，将所亏负人的如数赔偿，另外再加五分之一，交给所亏负的人。
NUM|5|8|那人若没有至亲可接受所赔偿的，所赔偿的就要归耶和华，交给祭司；另外还要献一只赎罪的公羊为他赎罪。
NUM|5|9|以色列 人一切的圣物中，所奉给祭司的一切礼物都要归给祭司。
NUM|5|10|各人自己的圣物归自己，给祭司的要归给祭司。”
NUM|5|11|耶和华吩咐 摩西 说：
NUM|5|12|“你要吩咐 以色列 人，对他们说：若任何人的妻子背离妇道，对丈夫不贞，
NUM|5|13|有人与她同寝交合，这事瞒过她的丈夫，没有被发现；她玷污自己，没有证人指控她，也没有被捉住；
NUM|5|14|丈夫若生了疑忌的心，对妻子起了疑忌，认为她玷污自己；或是丈夫生了疑忌的心，对妻子起了疑忌，虽然她没有玷污自己，
NUM|5|15|这人要带妻子到祭司那里，同时为她带十分之一伊法大麦面粉作供物。不可浇上油，也不可加乳香，因为这是疑忌的素祭，是纪念的素祭，使人记得罪孽。
NUM|5|16|“祭司要使那妇人近前来，站在耶和华面前。
NUM|5|17|祭司要把圣水盛在瓦器里，从帐幕的地上取些尘土，放在水中。
NUM|5|18|祭司要带那妇人站在耶和华面前，使她蓬头散发，再把纪念的素祭，就是疑忌的素祭，放在她的手掌，祭司手里捧着致诅咒的苦水。
NUM|5|19|祭司要叫妇人起誓，对她说：‘若没有人与你同寝，若你未曾背着丈夫做污秽的事，你就能免去这致诅咒的苦水。
NUM|5|20|但你背着丈夫，玷污自己，跟丈夫以外的人同寝。’
NUM|5|21|祭司叫妇人赌咒起誓，祭司对她说：‘当耶和华使你大腿萎缩，肚腹肿胀时，愿耶和华使你在你百姓中成为诅咒和咒骂；
NUM|5|22|愿这致诅咒的水进入你体内，使你肚腹肿胀，大腿萎缩。’妇人要说：‘阿们，阿们。’
NUM|5|23|“祭司要把这诅咒写在册上，然后用苦水涂去，
NUM|5|24|又叫妇人喝这致诅咒的苦水，这诅咒的水要进入她里面，令她痛苦。
NUM|5|25|祭司要从妇人手中取那疑忌的素祭，把素祭在耶和华面前摇一摇，拿到祭坛前；
NUM|5|26|又要从素祭中取出一把，作为纪念，烧在坛上，然后叫妇人喝这水。
NUM|5|27|祭司叫她喝了以后，她若玷污自己，确实对丈夫不贞，这致诅咒的水必进入她里面，令她痛苦，她的肚腹就要肿胀起来，大腿萎缩；这妇人就在她百姓中成为诅咒。
NUM|5|28|这妇人若没有玷污自己，是贞洁的，就要免受这灾，并且能够生育。
NUM|5|29|“这是疑忌的条例。妻子背离丈夫玷污自己，
NUM|5|30|或是丈夫生了疑忌的心，对妻子起了疑忌，祭司要使那妇人站在耶和华面前，在她身上照这条例而行。
NUM|5|31|男人可免罪责；女人必须担当自己的罪孽。”
NUM|6|1|耶和华吩咐 摩西 说：
NUM|6|2|“你要吩咐 以色列 人，对他们说：无论男女，若许了特别的愿，就是拿细耳人的愿，愿意离俗归耶和华，
NUM|6|3|他就要远离清酒烈酒，也不可喝任何清酒烈酒做的醋；不可喝任何葡萄汁，也不可吃鲜葡萄和干葡萄。
NUM|6|4|在一切离俗的日子，任何葡萄树上所结的，甚至果核和果皮，都不可吃。
NUM|6|5|“在他一切许愿离俗的日子，不可用剃刀剃头。在离俗归耶和华的日子未满之前，他要成为圣，要任由头上的发绺生长。
NUM|6|6|在他一切离俗归耶和华的日子，不可挨近死尸。
NUM|6|7|即使他的父母或兄弟姊妹死了，他也不可因他们使自己不洁净，因为他头上有离俗归上帝的记号 。
NUM|6|8|在他一切离俗的日子，他是归耶和华为圣的。
NUM|6|9|“若在他旁边忽然有人死了，因而玷污了他离俗的头，他要在第七日，得洁净的日子剃头。
NUM|6|10|第八日，他要把两只斑鸠或两只雏鸽带到会幕门口，交给祭司。
NUM|6|11|祭司要献一只作赎罪祭，一只作燔祭，为他赎因尸体而有的罪，并要在当日使他的头分别为圣。
NUM|6|12|他要另选离俗归耶和华的日子，牵一只一岁的小公羊来作赎愆祭。先前的那段日子算为无效，因为他在离俗期间被玷污了。
NUM|6|13|“拿细耳人的条例是这样的：离俗的日子满了，祭司要领他到会幕门口，
NUM|6|14|他要将供物献给耶和华，就是一只没有残疾的一岁小公羊作燔祭，一只没有残疾的一岁小母羊作赎罪祭，和一只没有残疾的公绵羊作平安祭，
NUM|6|15|一篮用油调和的无酵细面饼和抹了油的无酵薄饼，以及同献的素祭和浇酒祭。
NUM|6|16|祭司要来到耶和华面前，献上那人的赎罪祭和燔祭。
NUM|6|17|祭司要把公绵羊和那篮无酵饼献给耶和华作平安祭，又要献上同献的素祭和浇酒祭。
NUM|6|18|拿细耳人要在会幕门口剃离俗的头，把离俗头上的发放在平安祭下的火上。
NUM|6|19|他剃了离俗的头以后，祭司要取那煮好的公绵羊的一条前腿，连同篮子里的一块无酵饼和一块无酵薄饼，放在他手掌上。
NUM|6|20|祭司要拿这些在耶和华面前摇一摇，作为摇祭；这和所摇的胸、所举的腿一样是圣物，是归给祭司的。然后拿细耳人才可以喝酒。
NUM|6|21|“这是拿细耳人许愿的条例，除了他手头财力所及之外，他要为离俗献供物给耶和华。他怎样许愿，就当照离俗的条例做。”
NUM|6|22|耶和华吩咐 摩西 说：
NUM|6|23|“你要吩咐 亚伦 和他儿子说：你们要这样为 以色列 人祝福，对他们说：
NUM|6|24|‘愿耶和华赐福给你，保护你。
NUM|6|25|愿耶和华使他的脸光照你，赐恩给你。
NUM|6|26|愿耶和华向你仰脸，赐你平安。’
NUM|6|27|“他们要如此奉我的名为 以色列 人祝福；我也要赐福给他们。”
NUM|7|1|摩西 竖立帐幕后，就用膏抹了帐幕，使它分别为圣，又用膏抹其中的一切器具，以及祭坛和坛上的一切器具，使它们分别为圣。
NUM|7|2|以色列 的领袖，各父家的家长，都前来奉献。他们是各支派的领袖，管理那些被数的人。
NUM|7|3|他们把自己的供物送到耶和华面前，就是六辆篷车和十二头公牛。每两个领袖奉献一辆车，每个领袖奉献一头牛。他们把这些都带到帐幕前。
NUM|7|4|耶和华对 摩西 说：
NUM|7|5|“你要从他们收下这些，作为会幕事奉的用途，照着 利未 人所事奉的交给他们各人。”
NUM|7|6|于是 摩西 收了车和牛，交给 利未 人。
NUM|7|7|他把两辆车和四头牛，照着 革顺 子孙所事奉的交给他们，
NUM|7|8|又把四辆车和八头牛，照着 米拉利 子孙所事奉的交给他们。他们都在 亚伦 祭司的儿子 以他玛 的手下。
NUM|7|9|但没有交给 哥辖 子孙任何东西，因为他们所事奉的是圣物，必须抬在肩头上。
NUM|7|10|用膏抹祭坛的那一天，众领袖前来为献坛奉献；众领袖都在祭坛前献供物。
NUM|7|11|耶和华对 摩西 说：“众领袖为献坛奉献供物，每天要有一个领袖前来奉献。”
NUM|7|12|第一天献供物的是 犹大 支派的 亚米拿达 的儿子 拿顺 。
NUM|7|13|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|14|一个重十舍客勒的金碟子，盛满了香；
NUM|7|15|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|16|一只公山羊作赎罪祭；
NUM|7|17|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 亚米拿达 的儿子 拿顺 的供物。
NUM|7|18|第二天来献的是 以萨迦 的领袖， 苏押 的儿子 拿坦业 。
NUM|7|19|他献为供物的是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|20|一个重十舍客勒的金碟子，盛满了香；
NUM|7|21|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|22|一只公山羊作赎罪祭；
NUM|7|23|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 苏押 的儿子 拿坦业 的供物。
NUM|7|24|第三天是 西布伦 子孙的领袖， 希伦 的儿子 以利押 。
NUM|7|25|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|26|一个重十舍客勒的金碟子，盛满了香；
NUM|7|27|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|28|一只公山羊作赎罪祭；
NUM|7|29|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 希伦 的儿子 以利押 的供物。
NUM|7|30|第四天是 吕便 子孙的领袖， 示丢珥 的儿子 以利蓿 。
NUM|7|31|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|32|一个重十舍客勒的金碟子，盛满了香；
NUM|7|33|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|34|一只公山羊作赎罪祭；
NUM|7|35|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 示丢珥 的儿子 以利蓿 的供物。
NUM|7|36|第五天是 西缅 子孙的领袖， 苏利沙代 的儿子 示路蔑 。
NUM|7|37|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|38|一个重十舍客勒的金碟子，盛满了香；
NUM|7|39|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|40|一只公山羊作赎罪祭；
NUM|7|41|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 苏利沙代 的儿子 示路蔑 的供物。
NUM|7|42|第六天是 迦得 子孙的领袖， 丢珥 的儿子 以利雅萨 。
NUM|7|43|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|44|一个重十舍客勒的金碟子，盛满了香；
NUM|7|45|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|46|一只公山羊作赎罪祭；
NUM|7|47|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 丢珥 的儿子 以利雅萨 的供物。
NUM|7|48|第七天是 以法莲 子孙的领袖， 亚米忽 的儿子 以利沙玛 。
NUM|7|49|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|50|一个重十舍客勒的金碟子，盛满了香；
NUM|7|51|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|52|一只公山羊作赎罪祭；
NUM|7|53|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 亚米忽 的儿子 以利沙玛 的供物。
NUM|7|54|第八天是 玛拿西 子孙的领袖， 比大蓿 的儿子 迦玛列 。
NUM|7|55|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|56|一个重十舍客勒的金碟子，盛满了香；
NUM|7|57|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|58|一只公山羊作赎罪祭；
NUM|7|59|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 比大蓿 的儿子 迦玛列 的供物。
NUM|7|60|第九天是 便雅悯 子孙的领袖， 基多尼 的儿子 亚比但 。
NUM|7|61|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|62|一个重十舍客勒的金碟子，盛满了香；
NUM|7|63|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|64|一只公山羊作赎罪祭；
NUM|7|65|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 基多尼 的儿子 亚比但 的供物。
NUM|7|66|第十天是 但 子孙的领袖， 亚米沙代 的儿子 亚希以谢 。
NUM|7|67|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|68|一个重十舍客勒的金碟子，盛满了香；
NUM|7|69|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|70|一只公山羊作赎罪祭；
NUM|7|71|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 亚米沙代 的儿子 亚希以谢 的供物。
NUM|7|72|第十一天是 亚设 子孙的领袖， 俄兰 的儿子 帕结 。
NUM|7|73|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|74|一个重十舍客勒的金碟子，盛满了香；
NUM|7|75|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|76|一只公山羊作赎罪祭；
NUM|7|77|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 俄兰 的儿子 帕结 的供物。
NUM|7|78|第十二天是 拿弗他利 子孙的领袖， 以南 儿子 亚希拉 。
NUM|7|79|他的供物是：一个重一百三十舍客勒的银盘，一个重七十舍客勒的银碗，都是按照圣所的舍客勒，里面盛满了调油的细面作素祭；
NUM|7|80|一个重十舍客勒的金碟子，盛满了香；
NUM|7|81|一头公牛犊、一只公绵羊、一只一岁的小公羊作燔祭；
NUM|7|82|一只公山羊作赎罪祭；
NUM|7|83|两头公牛、五只公绵羊、五只公山羊、五只一岁的小公羊作平安祭。这是 以南 的儿子 亚希拉 的供物。
NUM|7|84|用膏抹祭坛的那一天， 以色列 的众领袖为献坛所献的是：银盘十二个、银碗十二个、金碟子十二个；
NUM|7|85|一个银盘重一百三十，一个碗七十。一切器皿的银子，按照圣所的舍客勒共二千四百舍客勒。
NUM|7|86|十二个金碟子盛满了香，按照圣所的舍客勒，一个碟子重十舍客勒，所有碟子的金子共一百二十舍客勒。
NUM|7|87|作燔祭的共有公牛十二头、公羊十二只、一岁的小公羊十二只，和同献的素祭，以及作赎罪祭的公山羊十二只；
NUM|7|88|作平安祭的共有公牛二十四头、公绵羊六十只、公山羊六十只、一岁的小公羊六十只。这就是用膏抹坛之后，为献坛的奉献。
NUM|7|89|摩西 进会幕要与耶和华说话的时候，听见法柜的柜盖以上二基路伯中间有对他说话的声音。耶和华向他说话。
NUM|8|1|耶和华吩咐 摩西 说：
NUM|8|2|“你要吩咐 亚伦 ，对他说：点灯的时候，七盏灯都要照亮灯台前面。”
NUM|8|3|亚伦 就照样做了；他点灯，照亮了灯台前面，正如耶和华所吩咐 摩西 的。
NUM|8|4|灯台是这样造的：灯台是用金子锤出来的，连座带花都是锤出来的。 摩西 照着耶和华所指示的样式造了灯台。
NUM|8|5|耶和华吩咐 摩西 说：
NUM|8|6|“你要从 以色列 人中选出 利未 人来，洁净他们。
NUM|8|7|你要这样做来洁净他们：要用洁净的水弹在他们身上，又叫他们用剃刀剃刮全身，洗净衣服，洁净自己。
NUM|8|8|然后他们要取一头公牛犊，以及同献的素祭，就是调油的细面。你要另取一头公牛犊作赎罪祭。
NUM|8|9|你要带 利未 人到会幕前，并且要召集 以色列 全会众。
NUM|8|10|你要把 利未 人带到耶和华面前， 以色列 人要为 利未 人按手。
NUM|8|11|亚伦 要从 以色列 人中将 利未 人奉献 在耶和华面前，作为摇祭，使他们事奉耶和华。
NUM|8|12|利未 人要按手在那两头牛的头上；你要将一头作赎罪祭，一头作燔祭，献给耶和华，为 利未 人赎罪。
NUM|8|13|你也要使 利未 人站在 亚伦 和他儿子面前，将他们奉献给耶和华，作为摇祭。
NUM|8|14|“你从 以色列 人中将 利未 人分别出来， 利未 人就归我了。
NUM|8|15|你洁净了 利未 人，奉献他们作为摇祭之后，他们就可以进会幕事奉。
NUM|8|16|因为他们是从 以色列 人中全然献给我的；我选他们归我，代替 以色列 人中所有头胎的长子。
NUM|8|17|因为 以色列 人中凡头生的，无论是人或牲畜，都是我的。我在 埃及 地击杀所有头生的那日，已将他们分别为圣归我。
NUM|8|18|我选 利未 人代替 以色列 人中所有头生的。
NUM|8|19|我从 以色列 人中将 利未 人给 亚伦 和他的儿子作为赏赐，在会幕中为 以色列 人事奉，又为 以色列 人赎罪，免得 以色列 人因挨近圣所而遭受灾祸。”
NUM|8|20|摩西 、 亚伦 和 以色列 全会众就向 利未 人这样做。关于 利未 人，凡耶和华怎样吩咐 摩西 ， 以色列 人就向他们照样做了。
NUM|8|21|于是 利未 人从罪中洁净自己，洗净衣服。 亚伦 将他们奉献在耶和华面前，作为摇祭，又为他们赎罪，洁净他们。
NUM|8|22|然后 利未 人进去，在 亚伦 和他儿子面前，在会幕中事奉。关于 利未 人，耶和华怎样吩咐 摩西 ，他们就向 利未 人照样做了。
NUM|8|23|耶和华吩咐 摩西 说：
NUM|8|24|“这是有关 利未 人的：二十五岁以上的人都要前来任职，在会幕里事奉。
NUM|8|25|到了五十岁，他们就要从事奉的工作中退休，不再事奉，
NUM|8|26|只可在会幕里辅助他们的弟兄尽责，他们自己不再事奉了。关于 利未 人的职责，你要向他们这样做。”
NUM|9|1|以色列 人出 埃及 地以后，第二年正月，耶和华在 西奈 的旷野吩咐 摩西 说：
NUM|9|2|“ 以色列 人应当在所定的日期守逾越节。
NUM|9|3|你们要在本月十四日黄昏的时候 ，在所定的日期守这节，按照一切的律例典章守节。”
NUM|9|4|于是 摩西 吩咐 以色列 人守逾越节。
NUM|9|5|正月十四日黄昏的时候，他们就在 西奈 的旷野守逾越节。凡耶和华所吩咐 摩西 的， 以色列 人都照样做了。
NUM|9|6|有几个人因尸体成了不洁净，不能在那日守逾越节。当天他们到 摩西 、 亚伦 面前。
NUM|9|7|那些人对他说：“我们因尸体而不洁净，为何禁止我们，不能和 以色列 人在所定的日期献供物给耶和华呢？”
NUM|9|8|摩西 对他们说：“你们稍等，让我去听耶和华对你们有什么吩咐。”
NUM|9|9|耶和华吩咐 摩西 说：
NUM|9|10|“你要吩咐 以色列 人说：你们和你们后代中，若有人因尸体成了不洁净，或出外远行，仍然要向耶和华守逾越节，
NUM|9|11|他们就要在二月十四日黄昏的时候守节，要吃羔羊，以及无酵饼和苦菜。
NUM|9|12|他们不可留一点食物到早晨；羔羊的骨头一根也不可折断。他们要照逾越节的一切律例守这节。
NUM|9|13|但洁净又不出外远行的人若不守逾越节，那人要从百姓中剪除，因为他没有在所定的日期献供物给耶和华，必须担当自己的罪。
NUM|9|14|若有寄居在你们那里的外人要向耶和华守逾越节，他要照逾越节的律例和典章做。无论是寄居的或是本地人，都用同样的律例。”
NUM|9|15|立起帐幕的那日，有云彩遮盖帐幕，就是法柜的帐幕；从晚上到早晨，云彩在帐幕上，形状如火。
NUM|9|16|经常都是这样：云彩遮盖帐幕，夜间云彩形状如火。
NUM|9|17|云彩几时从帐幕上升， 以色列 人就几时起行；云彩在哪里停住， 以色列 人就在哪里安营。
NUM|9|18|以色列 人遵照耶和华的指示起行，也遵照耶和华的指示安营。云彩在帐幕上停留多久，他们就留在营里多久。
NUM|9|19|云彩在帐幕上停留许多日子， 以色列 人就遵照耶和华的吩咐不起行。
NUM|9|20|有时云彩在帐幕上只停了几天，他们就遵照耶和华的指示留在营里，也遵照耶和华的指示起行。
NUM|9|21|有时云彩从晚上留到早晨；早晨云彩上升，他们就起行。无论是白天是黑夜，当云彩上升的时候，他们就要起行。
NUM|9|22|云彩停留在帐幕上，无论是两天，一个月，或更长的日子， 以色列 人就留在营里不起行；但云彩一上升，他们就起行。
NUM|9|23|他们遵照耶和华的指示安营，也遵照耶和华的指示起行。他们遵守耶和华的吩咐，是耶和华藉 摩西 所指示的话。
NUM|10|1|耶和华吩咐 摩西 说：
NUM|10|2|“你要用银子做两枝号筒，把它们锤出来，给你用来召集会众，拔营起行。
NUM|10|3|吹号的时候，全会众要到你那里，聚集在会幕的门口。
NUM|10|4|若只吹一枝，众领袖，就是 以色列 部队的官长，要到你那里聚集。
NUM|10|5|你们大声吹号的时候，东边安营的要起行。
NUM|10|6|第二次大声吹号的时候，南边安营的要起行。起行的时候，要大声吹号；
NUM|10|7|但召集会众的时候，你们要吹号，却不要吹出大声。
NUM|10|8|亚伦 子孙作祭司的要吹这号筒，作为你们世世代代永远的定例。
NUM|10|9|当你们在自己的土地上，与欺压你们的敌人打仗时，要用号筒吹出大声。你们就在耶和华－你们的上帝面前得蒙记念，也必蒙拯救脱离仇敌。
NUM|10|10|在快乐的日子，节期和初一，献燔祭与平安祭的时候，你们要吹号筒，在你们的上帝面前作为纪念。我是耶和华－你们的上帝。”
NUM|10|11|第二年二月二十日，云彩从法柜的帐幕上升。
NUM|10|12|以色列 人离开 西奈 的旷野，一段一段地往前行，云彩停在 巴兰 的旷野。
NUM|10|13|他们遵照耶和华藉 摩西 所指示的，初次往前行。
NUM|10|14|按照队伍首先起行的是 犹大 营旗帜下的人，带队的是 亚米拿达 的儿子 拿顺 。
NUM|10|15|以萨迦 支派带队的是 苏押 的儿子 拿坦业 。
NUM|10|16|西布伦 支派带队的是 希伦 的儿子 以利押 。
NUM|10|17|帐幕拆卸了， 革顺 的子孙和 米拉利 的子孙就抬着帐幕往前行。
NUM|10|18|按照队伍往前行的是 吕便 营旗帜下的人，带队的是 示丢珥 的儿子 以利蓿 。
NUM|10|19|西缅 支派带队的是 苏利沙代 的儿子 示路蔑 。
NUM|10|20|迦得 支派带队的是 丢珥 的儿子 以利雅萨 。
NUM|10|21|哥辖 人抬着圣物往前行。他们未到以前，帐幕已经立好了。
NUM|10|22|按照队伍往前行的是 以法莲 营旗帜下的人，带队的是 亚米忽 的儿子 以利沙玛 。
NUM|10|23|玛拿西 支派带队的是 比大蓿 的儿子 迦玛列 。
NUM|10|24|便雅悯 支派带队的是 基多尼 的儿子 亚比但 。
NUM|10|25|作全营后卫，按队伍往前行的是 但 营旗帜下的人，带队的是 亚米沙代 的儿子 亚希以谢 。
NUM|10|26|亚设 支派带队的是 俄兰 的儿子 帕结 。
NUM|10|27|拿弗他利 支派带队的是 以南 的儿子 亚希拉 。
NUM|10|28|以色列 人就这样按着队伍往前行。
NUM|10|29|摩西 对他岳父 ， 米甸 人 流珥 的儿子 何巴 说：“我们要往前行，到耶和华所说的地方；他曾说：‘我要将这地赐给你们。’现在请你和我们同去，我们必善待你，因为耶和华已经应许赐福气给 以色列 人。”
NUM|10|30|何巴 对他说：“我不去，我要回本地本族去。”
NUM|10|31|摩西 说：“请你不要离开我们，因为你知道我们要在旷野安营，你可以当我们的眼目。
NUM|10|32|你若和我们同去，将来耶和华以什么福气恩待我们，我们也必这样善待你。”
NUM|10|33|以色列 人离开耶和华的山，往前行了三天的路程。耶和华的约柜在前面行了三天的路程，为他们寻找安歇的地方。
NUM|10|34|他们拔营往前行，日间有耶和华的云彩在他们上面。
NUM|10|35|约柜往前行的时候， 摩西 说： “耶和华啊，求你兴起！ 愿你的仇敌溃散！ 愿恨你的人从你面前逃跑！”
NUM|10|36|约柜停住的时候，他说： “ 以色列 千万人的耶和华啊，求你回来 ！”
NUM|11|1|百姓发怨言，恶言传达到耶和华的耳中。耶和华听见了就怒气发作，耶和华的火在他们中间焚烧，烧毁营的外围。
NUM|11|2|百姓向 摩西 哀求， 摩西 祈求耶和华，火就熄了。
NUM|11|3|那地方就叫做 他备拉 ，因为耶和华的火曾在他们中间焚烧。
NUM|11|4|他们中间的闲杂人动了贪欲的心； 以色列 人又再哭着说：“谁给我们肉吃呢？
NUM|11|5|我们记得在 埃及 的时候，不花钱就可以吃鱼，还有黄瓜、西瓜、韭菜、葱、蒜。
NUM|11|6|现在我们的精力枯干了。除了这吗哪以外，在我们眼前什么都没有。”
NUM|11|7|吗哪好像芫荽子，看上去如同树脂的样子。
NUM|11|8|百姓四处走动捡取吗哪，把它用磨磨碎或用臼捣成粉，在锅中煮了做成饼，滋味好像油烤饼的滋味。
NUM|11|9|夜间露水降在营中，吗哪也随着降下。
NUM|11|10|摩西 听见百姓家家户户在帐棚门口哀哭。因此， 耶和华的怒气大大发作， 摩西 看了也不高兴。
NUM|11|11|摩西 对耶和华说：“你为何苦待仆人？我为何不在你眼前蒙恩，竟把这众百姓的担子加在我身上呢？
NUM|11|12|这众百姓岂是我怀的胎，岂是我生下来的呢？你竟对我说：‘把他们抱在怀里，如养育之父抱着吃奶的婴孩，一直抱到你起誓应许给他们祖宗的土地去。’
NUM|11|13|我从哪里拿肉给这众百姓吃呢？他们都向我哭着说：‘给我们肉吃！’
NUM|11|14|我不能独自带领这众百姓，这对我太沉重了。
NUM|11|15|如果你这样待我，倒不如立刻把我杀了吧！我若在你眼前蒙恩，求你不要让我再受这样的苦。”
NUM|11|16|耶和华对 摩西 说：“你要从 以色列 的长老中为我召集七十个人，就是你所认识，作百姓的长老和官长的，领他们到会幕，使他们和你一同站在那里。
NUM|11|17|我要在那里降临，与你说话，把降给你的灵分给他们。他们就和你分担带领百姓的担子，免得你独自承担。
NUM|11|18|你要对百姓说：‘你们要为了明天使自己分别为圣，你们将有肉吃。因你们哭着说：谁给我们肉吃呢？我们在 埃及 多么好！这声音传到了耶和华的耳中，所以他必给你们肉吃。
NUM|11|19|你们不只吃一天、两天、五天、十天、二十天，
NUM|11|20|而是整整一个月，直到肉从你们的鼻孔喷出来，使你们厌恶。因为你们厌弃那住在你们中间的耶和华，在他面前哭着说：我们为何出 埃及 呢？’”
NUM|11|21|摩西 说：“跟我在一起的百姓，步行的男人就有六十万，你还说：‘我要把肉赐给他们，使他们可以整整吃一个月。’
NUM|11|22|难道宰了羊群牛群，就够给他们吗？或者把海中所有的鱼都捕来，就够给他们吗？”
NUM|11|23|耶和华对 摩西 说：“耶和华的膀臂 岂是缩短了吗？现在你要看我的话向你应验不应验。”
NUM|11|24|摩西 出去，把耶和华的话告诉百姓，并从百姓的长老中召集七十个人来，叫他们站在会幕的四围。
NUM|11|25|耶和华在云中降临，对 摩西 说话，把降给他的灵分给那七十个长老。灵停在他们身上的时候，他们就说预言，以后却没有再说了。
NUM|11|26|但有两个人仍在营里，一个名叫 伊利达 ，一个名叫 米达 。他们本是在那些登记的人中，却没有到会幕那里去。灵停在他们身上，他们就在营里说预言。
NUM|11|27|有一个年轻人跑来告诉 摩西 说：“ 伊利达 和 米达 在营里说预言。”
NUM|11|28|嫩 的儿子 约书亚 ，年轻时就作 摩西 的助手 ，说：“请我主 摩西 禁止他们。”
NUM|11|29|摩西 对他说：“你为我的缘故嫉妒吗？惟愿耶和华的百姓都是先知，愿耶和华把他的灵降在他们身上！”
NUM|11|30|于是， 摩西 回到营里去， 以色列 的长老也回去了。
NUM|11|31|有一阵风从耶和华那里刮起，把鹌鹑从海上刮来，散落在营地和周围；一边约有一天的路程，另一边也约有一天的路程，离地面约有二肘。
NUM|11|32|百姓起来，整天整夜，甚至次日一整天，都在捕捉鹌鹑。每人至少捉到十贺梅珥，各自摆在营的四围。
NUM|11|33|但肉在他们牙间还未咀嚼时，耶和华的怒气向百姓发作，用极重的灾祸击杀百姓。
NUM|11|34|那地方就叫 基博罗．哈他瓦 ，因为他们在那里埋葬了贪欲的百姓。
NUM|11|35|百姓从 基博罗．哈他瓦 起程，到 哈洗录 ，就住在 哈洗录 。
NUM|12|1|摩西 娶了 古实 女子为妻。 米利暗 和 亚伦 因他娶了 古实 女子就批评他，
NUM|12|2|他们说：“难道耶和华只与 摩西 说话吗？他不也与我们说话吗？”耶和华听见了。
NUM|12|3|摩西 为人极其谦和，胜过地面上的任何人。
NUM|12|4|忽然，耶和华对 摩西 、 亚伦 和 米利暗 说：“你们三个人都出来，到会幕这里。”他们三个人就出来了。
NUM|12|5|耶和华在云柱中降临，停在会幕门口，叫 亚伦 和 米利暗 。二人就出来，
NUM|12|6|耶和华说：“你们要听我的话：你们中间若有先知，我－耶和华必在异象中向他显现，在梦中与他说话；
NUM|12|7|但我的仆人 摩西 不是这样，他在我全家是尽忠的。
NUM|12|8|我与他面对面说话，清清楚楚，不用谜语，他甚至看见我的形像。你们为何批评我的仆人 摩西 而不惧怕呢？”
NUM|12|9|耶和华向他们怒气发作，就离开了。
NUM|12|10|当云彩从帐幕上离开时，看哪， 米利暗 长了痲疯，像雪那么白。 亚伦 转向 米利暗 ，看哪，她长了痲疯。
NUM|12|11|亚伦 对 摩西 说：“我主啊，求你不要因我们愚昧，因我们犯罪，就将这罪加在我们身上。
NUM|12|12|求你不要使她像那一出母腹、肉已侵蚀了一半的死胎。”
NUM|12|13|于是 摩西 哀求耶和华说：“上帝啊，求你医治她！”
NUM|12|14|耶和华对 摩西 说：“她父亲若吐唾沫在她脸上，她岂不蒙羞七天吗？现在要把她隔离在营外七天，然后才领她回来。”
NUM|12|15|于是 米利暗 被隔离在营外七天；百姓没有起程，直等到 米利暗 回来。
NUM|12|16|以后百姓从 哈洗录 起行，来到 巴兰 的旷野安营。
NUM|13|1|耶和华吩咐 摩西 说：
NUM|13|2|“你要派人去窥探我所赐给 以色列 人的 迦南 地；每个父系支派要派一个人，是他们中间的族长。”
NUM|13|3|摩西 就遵照耶和华的指示，从 巴兰 旷野差派他们去；他们都是 以色列 人中的领袖。
NUM|13|4|这是他们的名字： 属 吕便 支派的， 撒刻 的儿子 沙母亚 。
NUM|13|5|属 西缅 支派的， 何利 的儿子 沙法 。
NUM|13|6|属 犹大 支派的， 耶孚尼 的儿子 迦勒 。
NUM|13|7|属 以萨迦 支派的， 约色 的儿子 以迦 。
NUM|13|8|属 以法莲 支派的， 嫩 的儿子 何西阿 。
NUM|13|9|属 便雅悯 支派的， 拉孚 的儿子 帕提 。
NUM|13|10|属 西布伦 支派的， 梭底 的儿子 迦叠 。
NUM|13|11|属 约瑟 支派，就是 玛拿西 支派的， 稣西 的儿子 迦底 。
NUM|13|12|属 但 支派的， 基玛利 的儿子 亚米利 。
NUM|13|13|属 亚设 支派的， 米迦勒 的儿子 西帖 。
NUM|13|14|属 拿弗他利 支派的， 缚西 的儿子 拿比 。
NUM|13|15|属 迦得 支派的， 玛基 的儿子 臼利 。
NUM|13|16|这些是 摩西 差派去窥探那地之人的名字。 摩西 叫 嫩 的儿子 何西阿 为 约书亚 。
NUM|13|17|摩西 差派他们去窥探 迦南 地，对他们说：“你们上到 尼革夫 那里，上到山区去，
NUM|13|18|看看那地如何：住那里的百姓是强是弱，是多是少，
NUM|13|19|他们所住的地是好是坏，所住的城镇是营地还是堡垒，
NUM|13|20|那地是肥沃还是贫瘠，当中有树木没有。你们要放胆，把那地的果子带些回来。”那时正是葡萄初熟的季节。
NUM|13|21|他们上去窥探那地，从 寻 的旷野到 利合 ，直到 哈马口 。
NUM|13|22|他们从 尼革夫 上去，到了 希伯仑 。在那里有 亚衲 族的 亚希幔 人、 示筛 人和 挞买 人。 希伯仑 的建造比 埃及 的 琐安 早七年。
NUM|13|23|他们到了 以实各谷 ，从那里砍下葡萄树枝，上面有一挂葡萄，两个人用杠抬着，又带了一些石榴和无花果。
NUM|13|24|以色列 人从那里砍下一挂葡萄，所以那地方就叫 以实各谷 。
NUM|13|25|他们窥探那地四十天之后，就回来了。
NUM|13|26|他们来到 巴兰 旷野的 加低斯 ， 摩西 、 亚伦 ，以及 以色列 全会众那里，向他们和全会众报告，又把那地的果子给他们看。
NUM|13|27|他们告诉 摩西 说：“我们到了你派我们去的那地，果然是流奶与蜜之地；这就是那地的果子。
NUM|13|28|但是住那地的百姓很强悍，城镇又大又坚固，我们也在那里看见了 亚衲 族人。
NUM|13|29|亚玛力 人住在 尼革夫 ； 赫 人、 耶布斯 人和 亚摩利 人住在山区； 迦南 人住在沿海一带和 约旦河 旁。”
NUM|13|30|迦勒 在 摩西 面前安抚百姓，说：“我们立刻上去得那地吧！我们必能征服它。”
NUM|13|31|但那些和他同去的人却说：“我们不能上去攻打那些百姓，因为他们比我们强大。”
NUM|13|32|于是探子中有人向 以色列 人散布有关所窥探之地的谣言，说：“我们所走过、所窥探之地是吞没居民之地，并且我们在那里所看见的百姓都身材高大。
NUM|13|33|我们在那里看见巨人，就是巨人中的 亚衲 族人。我们在自己眼中像蚱蜢一样，而在他们眼中，我们也确是这样。”
NUM|14|1|全会众大声喧嚷，那夜百姓哭号。
NUM|14|2|以色列 众人向 摩西 和 亚伦 发怨言，全会众对他们说：“我们宁愿死在 埃及 地，宁愿死在这旷野！
NUM|14|3|耶和华为什么要把我们领到那地，让我们倒在刀下呢？我们的妻子和孩子必成为掳物。我们回 埃及 去岂不更好吗？”
NUM|14|4|他们彼此说：“我们不如选一个领袖，回 埃及 去吧！”
NUM|14|5|摩西 和 亚伦 在 以色列 全会众面前脸伏于地。
NUM|14|6|窥探那地的人中， 嫩 的儿子 约书亚 和 耶孚尼 的儿子 迦勒 撕裂衣服，
NUM|14|7|对 以色列 全会众说：“我们所走过、所窥探之地是极美之地。
NUM|14|8|耶和华若喜爱我们，就必领我们进入那地，把这流奶与蜜之地赐给我们。
NUM|14|9|但你们不可背叛耶和华，也不要怕那地的百姓，因为他们是我们的食物。保护他们的已经离开他们，耶和华却与我们同在。不要怕他们！”
NUM|14|10|当全会众正说着要拿石头打死他们的时候，耶和华的荣光在会幕中向 以色列 众人显现。
NUM|14|11|耶和华对 摩西 说：“这百姓藐视我要到几时呢？我在他们中间行了这一切神迹，他们还不信我要到几时呢？
NUM|14|12|我要用瘟疫击杀他们，使他们不得承受那地。我要使你成为大国，比他们强大。”
NUM|14|13|摩西 对耶和华说：“ 埃及 人必听见，因你曾施展大能，领这百姓从他们中间出来。
NUM|14|14|埃及 人要告诉这地的居民，他们已经听见你─耶和华是在这百姓中间，因为你─耶和华面对面 显示自己，你的云彩停在他们以上。你日间在云柱中，夜间在火柱中，在他们的前面行。
NUM|14|15|你若把这百姓杀了，好像杀一个人那样，那听见你名声的列国必说：
NUM|14|16|‘耶和华因为不能把这百姓领进他向他们起誓应许之地，所以在旷野把他们杀了。’
NUM|14|17|现在求主显出大能，照你说过的话说：
NUM|14|18|‘耶和华不轻易发怒， 且有丰盛的慈爱。 他赦免罪孽和过犯， 万不以有罪的为无罪， 必惩罚人的罪， 从父到子，直到三、四代。’
NUM|14|19|求你照你的大慈爱赦免这百姓的罪孽，好像你从 埃及 到如今饶恕这百姓一样。”
NUM|14|20|耶和华说：“我照着你的话赦免他们。
NUM|14|21|然而，我指着我的永生与遍地充满了耶和华的荣耀起誓：
NUM|14|22|这些人虽然都看过我的荣耀和我在 埃及 与旷野所行的神迹，仍然这十次试探我，不听从我的话，
NUM|14|23|他们绝不能看见我向他们祖宗所起誓应许之地；凡藐视我的，一个也不得看见。
NUM|14|24|惟独我的仆人 迦勒 ，因他另有一个心志，专心跟从我，我要领他进入他所去过的那地；他的后裔必得那地为业。
NUM|14|25|亚玛力 人和 迦南 人住在谷中，明天你们要转回去，沿着 红海 的路往旷野去。”
NUM|14|26|耶和华对 摩西 和 亚伦 说：
NUM|14|27|“这邪恶的会众向我发怨言要到几时呢？ 以色列 人向我发的怨言，我都听见了。
NUM|14|28|你要告诉他们，耶和华说：‘我指着我的永生起誓，我必照你们在我耳中所说的待你们。
NUM|14|29|你们的尸体必倒在这旷野中。你们中间被数点，凡二十岁以上向我发怨言的，
NUM|14|30|必不得进我所起誓应许给你们居住的那地。惟有 耶孚尼 的儿子 迦勒 和 嫩 的儿子 约书亚 才能进去。
NUM|14|31|你们的孩子，就是你们说要成为掳物的，我必领他们进去，他们就得知你们所厌弃的那地。
NUM|14|32|至于你们，你们的尸体必倒在这旷野中；
NUM|14|33|你们的儿女必在旷野游牧四十年，担当你们不信的罪 ，直到你们的尸体在旷野消灭为止。
NUM|14|34|按你们窥探那地的四十日，一年抵一日，你们要担当你们的罪孽四十年，你们就知道我疏远你们了。’
NUM|14|35|我－耶和华说过，我必这样对待这一切聚集对抗我的邪恶会众。他们必在这旷野中消灭，死在这里。”
NUM|14|36|摩西 所差派去窥探那地的人回来，散布有关那地的谣言，使全会众向 摩西 发怨言，
NUM|14|37|这些散布谣言的人都遭受瘟疫，死在耶和华面前。
NUM|14|38|窥探那地的人中，惟有 嫩 的儿子 约书亚 和 耶孚尼 的儿子 迦勒 得以存活。
NUM|14|39|摩西 把这些话告诉 以色列 众人，他们都极其悲哀。
NUM|14|40|他们清晨起来，上到山顶，说：“看哪，我们要上到耶和华所说的地方；因为我们犯了罪。”
NUM|14|41|摩西 说：“你们为何要这样违背耶和华的指示呢？这事必不能顺利。
NUM|14|42|不要上去，因为耶和华不在你们中间，恐怕你们在仇敌面前被击败。
NUM|14|43|亚玛力 人和 迦南 人都在你们面前，你们必倒在刀下。因为你们背离不跟从耶和华，耶和华必不与你们同在。”
NUM|14|44|他们却擅自上到山顶。但耶和华的约柜和 摩西 都没有离开营地。
NUM|14|45|于是 亚玛力 人和住在那山区的 迦南 人下来，击败他们，追击他们直到 何珥玛 。
NUM|15|1|耶和华吩咐 摩西 说：
NUM|15|2|“你要吩咐 以色列 人，对他们说：你们到了我所赐给你们居住的地，
NUM|15|3|你们要从牛群羊群中取牲畜献给耶和华为火祭，无论是燔祭或祭物，为要还所许特别的愿或甘心祭，或节期的祭，作为献给耶和华的馨香之祭，
NUM|15|4|那献供物的要将十分之一伊法细面和四分之一欣油调和作素祭，献给耶和华。
NUM|15|5|无论是燔祭或祭物，要为每只小绵羊预备四分之一欣酒作浇酒祭。
NUM|15|6|要为每只公绵羊预备十分之二伊法细面，和三分之一欣油调和作素祭，
NUM|15|7|又用三分之一欣酒作浇酒祭，献给耶和华为馨香之祭。
NUM|15|8|你预备公牛献给耶和华作燔祭或祭物，为要还所许特别的愿，或平安祭，
NUM|15|9|就要把十分之三伊法细面和半欣油调和作素祭，和公牛一同献上，
NUM|15|10|又用半欣酒作浇酒祭，献给耶和华为馨香的火祭。
NUM|15|11|“献公牛、或公绵羊、或小绵羊、或小山羊，每只都要这样处理；
NUM|15|12|无论你们所献的数目多少，照着数目每只都要这样处理。
NUM|15|13|凡本地人将馨香的火祭献给耶和华，都要照样处理。
NUM|15|14|若有外人寄居在你们那里，或有人世世代代住在你们中间，愿意将馨香的火祭献给耶和华，你们怎样处理，他也要照样处理。
NUM|15|15|至于会众，无论是你们或寄居的外人都要遵守同一条例；这是你们世世代代永远的定例。在耶和华面前，你们怎样，寄居的也要怎样。
NUM|15|16|你们和寄居在你们那里的外人要遵守同一律法，同一典章。”
NUM|15|17|耶和华吩咐 摩西 说：
NUM|15|18|“你要吩咐 以色列 人，对他们说：你们到了我领你们进去的那地，
NUM|15|19|吃那地的粮食时，要把举祭献给耶和华。
NUM|15|20|你们要用初熟的麦子磨面，做成饼当举祭献上。你们要举上，如同举禾场的举祭。
NUM|15|21|你们世世代代要用初熟的麦子磨面，当举祭献给耶和华。
NUM|15|22|“你们若犯了错，不遵守耶和华所吩咐 摩西 的这一切命令，
NUM|15|23|就是耶和华藉 摩西 一切所命令你们的，从耶和华命令的那日直到你们的世世代代，
NUM|15|24|会众因没有察觉而犯了无心之过，全会众就要将一头公牛犊作燔祭，遵照典章把素祭和浇酒祭一同献给耶和华为馨香的祭，又要献一只公山羊作赎罪祭。
NUM|15|25|祭司要为 以色列 全会众赎罪，他们就必蒙赦免，因为这是无心之过。他们要因自己的无心之过，把供物，就是向耶和华当献的火祭和赎罪祭，带到耶和华面前。
NUM|15|26|以色列 全会众和寄居在他们中间的外人就必蒙赦免，因为这是众百姓的无心之过。
NUM|15|27|“若有一个人无意中犯了罪，他就要献一只一岁的母山羊作赎罪祭。
NUM|15|28|这误犯罪的人因无意中犯了罪，祭司要在耶和华面前为他赎罪，他就必蒙赦免。
NUM|15|29|以色列 中的本地人和寄居在他们中间的外人，若无意中犯了罪，都要遵守同一律法。
NUM|15|30|但那故意犯罪的人，无论是本地人是寄居的，亵渎了耶和华，这人必从百姓中剪除。
NUM|15|31|因为他藐视耶和华的话，违背耶和华的命令，这人一定要剪除；他的罪孽要归到自己身上。”
NUM|15|32|以色列 人还在旷野的时候，发现有一个人在安息日捡柴。
NUM|15|33|发现他捡柴的人把他带到 摩西 、 亚伦 以及全会众那里。
NUM|15|34|他们把他收押在监里，因为还不知道要怎样惩罚他。
NUM|15|35|耶和华吩咐 摩西 说：“这人应当处死；全会众要在营外用石头打死他。”
NUM|15|36|于是全会众把他带到营外，用石头打死他，是照耶和华所吩咐 摩西 的。
NUM|15|37|耶和华对 摩西 说：
NUM|15|38|“你吩咐 以色列 人，对他们说，他们世世代代要在衣服边上缝繸子，并在边上的繸子钉一条蓝色带子。
NUM|15|39|你们要佩带这繸子，好叫你们看见它就记起耶和华一切的命令，并且遵行，不随从自己内心和眼目的情欲而跟着行淫。
NUM|15|40|这样，你们就必记得并遵行我一切的命令，成为圣，归你们的上帝。
NUM|15|41|“我是耶和华－你们的上帝，曾把你们从 埃及 地领出来，要作你们的上帝。我是耶和华－你们的上帝。”
NUM|16|1|利未 的曾孙， 哥辖 的孙子， 以斯哈 的儿子 可拉 ，连同 吕便 子孙中 以利押 的儿子 大坍 和 亚比兰 ，与 比勒 的儿子 安 ，带了
NUM|16|2|以色列 人中的二百五十个领袖，就是有名望、从会众中选出来的人，在 摩西 面前一同起来，
NUM|16|3|聚集攻击 摩西 、 亚伦 ，说：“你们太过分了！全会众人人都成为圣，耶和华也在他们中间。你们为什么抬高自己，在耶和华的会众之上呢？”
NUM|16|4|摩西 听见就脸伏于地，
NUM|16|5|对 可拉 和他所有同伙的人说：“到了早晨，耶和华必指示谁是属他的，谁是成为圣的，就准许谁亲近他。他要叫自己所拣选的人亲近他。
NUM|16|6|可拉 和你所有同伙的人哪，你们要这样做：要拿着香炉，
NUM|16|7|明天在耶和华面前把火盛在炉中，把香放在上面。耶和华拣选谁，谁就成为圣。 利未 的子孙哪，你们太过分了！”
NUM|16|8|摩西 又对 可拉 说：“ 利未 的子孙，听吧！
NUM|16|9|以色列 的上帝将你们从 以色列 会众中分别出来，使你们亲近他，在耶和华的帐幕中事奉，并且站在会众面前替他们供职。这对你们岂是小事吗？
NUM|16|10|耶和华已经准许你和你所有的弟兄，就是 利未 的子孙，一同亲近他，你们还要求祭司的职分吗？
NUM|16|11|所以，你和你所有同伙的人聚集是在攻击耶和华。 亚伦 算什么，你们竟向他发怨言？”
NUM|16|12|摩西 派人去叫 以利押 的儿子 大坍 和 亚比兰 。他们却说：“我们不上去！
NUM|16|13|你把我们从流奶与蜜之地领出来，让我们死在旷野，这岂是小事？你还要自立为王管辖我们吗？
NUM|16|14|你根本没有领我们到流奶与蜜之地，也没有给我们田地和葡萄园作为产业。难道你想要挖这些人的眼睛吗？我们不上去！”
NUM|16|15|摩西 非常生气，就对耶和华说：“求你不要接受他们的供物。我并没有夺过他们一匹驴，也没有害过他们中任何一个人。”
NUM|16|16|摩西 对 可拉 说：“明天，你和你所有同伙的人，以及 亚伦 ，都要站在耶和华面前。
NUM|16|17|你们各人要拿一个香炉，把香放在上面，各人带香炉到耶和华面前，共二百五十个；你和 亚伦 也各拿自己的香炉。”
NUM|16|18|于是他们各人拿一个香炉，盛着火，加上香，和 摩西 、 亚伦 一同站在会幕的门口。
NUM|16|19|可拉 召集全会众到会幕门口攻击 摩西 和 亚伦 。这时，耶和华的荣光向全会众显现。
NUM|16|20|耶和华吩咐 摩西 和 亚伦 说：
NUM|16|21|“你们离开这会众，我好立刻把他们灭绝。”
NUM|16|22|摩西 、 亚伦 脸伏于地，说：“上帝，赐万人气息的上帝啊，一人犯罪，你就要向全会众发怒吗？”
NUM|16|23|耶和华吩咐 摩西 说：
NUM|16|24|“你吩咐会众说：‘你们远离 可拉 、 大坍 和 亚比兰 帐棚的周围。’”
NUM|16|25|摩西 起来，到 大坍 、 亚比兰 那里去； 以色列 的长老也都跟着他去。
NUM|16|26|他吩咐会众说：“你们离开这些恶人的帐棚吧！不可碰他们的任何东西，免得你们因他们一切的罪而消灭。”
NUM|16|27|于是会众远离了 可拉 、 大坍 和 亚比兰 的帐棚。 大坍 和 亚比兰 带着妻子、儿女和小孩子出来，站在自己的帐棚门口。
NUM|16|28|摩西 说：“因这件事，你们就必知道这一切事是耶和华差派我做的，并非出于我的心意。
NUM|16|29|这些人的死若和世人无异，或者他们所遭遇的和其他人相同，那么耶和华就不曾差派我了。
NUM|16|30|但是，倘若耶和华创作一件新事，使地开了裂口，把他们和一切属他们的都吞下去，叫他们活活坠落阴间，你们就知道是这些人藐视了耶和华。”
NUM|16|31|摩西 刚说完这些话，他们脚下的地就裂开，
NUM|16|32|地开了裂口，把他们和他们的家眷，以及一切属 可拉 的人和财物，都吞了下去。
NUM|16|33|他们和一切属他们的，都活活坠落阴间；地在他们上面又合拢起来，他们就从会众中灭亡了。
NUM|16|34|在他们四围的 以色列 众人听见他们的叫声，就都逃跑，说：“恐怕地也要把我们吞下去了！”
NUM|16|35|有火从耶和华那里出来，吞灭了那上香的二百五十人。
NUM|16|36|耶和华吩咐 摩西 说：
NUM|16|37|“你要对 亚伦 祭司的儿子 以利亚撒 说，把香炉从火中移开，再把炭火撒在别处，因为这些香炉是分别为圣的。
NUM|16|38|要把那些犯罪自丧己命之人的香炉锤成薄片，用以包祭坛；因为这些本是他们在耶和华面前献过，分别为圣的，可以给 以色列 人作记号。”
NUM|16|39|于是 以利亚撒 祭司把被烧死的人所献的铜香炉拿来；它们被锤出来，用以包坛，
NUM|16|40|给 以色列 人作纪念，为要叫 亚伦 子孙之外的人不得近前来，在耶和华面前烧香，免得他和 可拉 与同他一伙的人一样，正如耶和华藉 摩西 所吩咐的。
NUM|16|41|第二天， 以色列 全会众都向 摩西 、 亚伦 发怨言说：“你们杀了耶和华的百姓了。”
NUM|16|42|会众聚集攻击 摩西 、 亚伦 的时候， 摩西 和 亚伦 转向会幕，看哪，云彩遮盖会幕，耶和华的荣光显现。
NUM|16|43|摩西 、 亚伦 就来到会幕前。
NUM|16|44|耶和华吩咐 摩西 说：
NUM|16|45|“你们离开这会众，我好立刻把他们灭绝。”他们二人就脸伏于地。
NUM|16|46|摩西 对 亚伦 说：“拿你的香炉，把祭坛的火盛在里面，加上香，赶快带到会众那里，为他们赎罪。因为有愤怒从耶和华面前发出，瘟疫已经开始了。”
NUM|16|47|亚伦 照 摩西 所说的拿了香炉，跑到会众中。看哪，瘟疫已经在百姓中开始了。他就加上香，为百姓赎罪。
NUM|16|48|他站在活人和死人之间，瘟疫就止住了。
NUM|16|49|除了因 可拉 事件死的以外，遭瘟疫死的共有一万四千七百人。
NUM|16|50|亚伦 回到会幕门口 ，到 摩西 那里，瘟疫已经止住了。
NUM|17|1|耶和华吩咐 摩西 说：
NUM|17|2|“你要吩咐 以色列 人，从他们当中取杖，每父家一根；从他们所有的领袖，按着父家，共取十二根。你要把各人的名字写在他的杖上，
NUM|17|3|并要把 亚伦 的名字写在 利未 的杖上，因为各父家的家长都有一根杖。
NUM|17|4|你要把这些杖放在会幕里法柜前，我与你们 相会的地方。
NUM|17|5|我所拣选的人，他的杖必发芽。我就平息了 以色列 人向你们所发的怨言，不再达到我这里。”
NUM|17|6|于是， 摩西 吩咐 以色列 人，他们的众领袖就把杖给他，一个领袖一根杖，按照父家一个领袖一根杖，共有十二根； 亚伦 的杖也在其中。
NUM|17|7|摩西 把这些杖放在耶和华面前，在法柜的帐幕里。
NUM|17|8|第二天， 摩西 进到法柜的帐幕去，看哪， 利未 族 亚伦 的杖已经发芽，长了花苞，开了花，也结出熟的杏子！
NUM|17|9|摩西 把所有的杖从耶和华面前拿出来，给 以色列 众人看。他们都看见了，各领袖就把自己的杖拿去。
NUM|17|10|耶和华吩咐 摩西 说：“把 亚伦 的杖放回法柜前，给这些背叛之子留作记号。你就可以平息他们向我所发的怨言，他们也不会死亡。”
NUM|17|11|摩西 就照样做了；耶和华怎样吩咐他，他就照样做。
NUM|17|12|以色列 人对 摩西 说：“看哪，我们死啦！我们灭亡啦！我们全都灭亡啦！
NUM|17|13|凡挨近耶和华帐幕的，就必死亡。我们都要消灭而死吗？”
NUM|18|1|耶和华对 亚伦 说：“你和你的儿子，以及你父家的人，要一同担当干犯圣所的罪孽；你和你的儿子也要担当干犯祭司职分的罪孽。
NUM|18|2|你也要带你弟兄 利未 人，就是你父系支派的人前来，与你联合，服事你。你和你的儿子要一起在法柜的帐幕前；
NUM|18|3|他们要遵守你的吩咐，负责看守整个帐幕，只是不可挨近圣所的器具和祭坛，免得他们和你们都死亡。
NUM|18|4|他们要与你联合，负责看守会幕和帐幕一切的事；只是外人不可挨近你们。
NUM|18|5|你们要负责看守圣所和祭坛，免得愤怒再临到 以色列 人。
NUM|18|6|看哪，我已从 以色列 人中选了你们的弟兄 利未 人，交给你们为赏赐，归给耶和华，为要在会幕里事奉。
NUM|18|7|你和你的儿子要谨守祭司的职分，负责一切关于祭坛和幔子内的事。我把祭司的职分赐给你们，作为赏赐好事奉我；凡挨近的外人必被处死。”
NUM|18|8|耶和华吩咐 亚伦 说：“看哪，我已将归我的举祭，就是 以色列 人一切分别为圣之物，交给你照管；我把受膏的份赐给你和你的子孙，作为永远当得的份。
NUM|18|9|这是至圣供物中所给你的，一切献给我为至圣的素祭、赎罪祭、赎愆祭，其中所有不被火烧的供物，都要归你和你的子孙。
NUM|18|10|你要把它当作至圣之物吃 ；凡男丁都可以吃。你要以这祭物为圣。
NUM|18|11|这也是你的， 以色列 人所献的举祭和摇祭，我已赐给你和你的儿女，作为永远当得的份；你家中任何洁净的人都可以吃。
NUM|18|12|凡最好的新油、最好的新酒和五谷，就是 以色列 人献给耶和华的初熟之物，我都赐给你。
NUM|18|13|凡他们从地上所带来给耶和华的初熟之物也都要归给你。你家中任何洁净的人都可以吃。
NUM|18|14|以色列 中一切永献的都必归给你。
NUM|18|15|他们所有奉给耶和华的，无论是人是牲畜，凡头胎的，都要归给你；但是人的长子，一定要赎出来。不洁净牲畜中头生的，也要赎出来。
NUM|18|16|其中一个月以上所当赎的，要照你的估价，按圣所的舍客勒，付五舍客勒银子将他赎回，一舍客勒是二十季拉。
NUM|18|17|但是头生的牛，或头生的绵羊，或头生的山羊，却不可赎，因为它们都是圣的。要把它们的血洒在祭坛上，把它们的脂肪焚烧，当作馨香的火祭献给耶和华。
NUM|18|18|它们的肉必归你，像被摇的胸、被举的右腿归你一样。
NUM|18|19|凡 以色列 人所献给耶和华圣物中的举祭，我都赐给你和你的儿女，作为永远当得的份。这要成为你和你的后裔在耶和华面前永远的盐 约。
NUM|18|20|耶和华对 亚伦 说：“你在 以色列 人的境内不可有产业，在他们中间也不可有份。在 以色列 人中，我是你的份，你的产业。
NUM|18|21|“至于 利未 的子孙，看哪，我已赐给他们 以色列 所有出产的十分之一为业，作为他们在会幕中事奉的酬劳。
NUM|18|22|以色列 人不可再挨近会幕，免得他们担当罪而死。
NUM|18|23|惟独 利未 人要在会幕中事奉，他们要担当罪孽，作为你们世世代代永远的定例。他们在 以色列 人中不可有产业；
NUM|18|24|因为 以色列 人出产的十分之一，就是献给耶和华为举祭的，我已赐给 利未 人为业。所以我对他们说，他们不可在 以色列 人中有产业。”
NUM|18|25|耶和华吩咐 摩西 说：
NUM|18|26|“你要吩咐 利未 人，对他们说：你们从 以色列 人中所取的十分之一，就是我给你们为业的，要从这十分之一中取十分之一，作为献给耶和华的举祭。
NUM|18|27|这可算为你们的举祭，如同禾场上的谷，酒池中盛满的酒。
NUM|18|28|这样，从 以色列 人中所收取所有的十分之一，你们要从其中取举祭献给耶和华；你们要把献给耶和华的举祭归给 亚伦 祭司。
NUM|18|29|你们要将给你们一切礼物中最好的，就是分别为圣的，献给耶和华为举祭。
NUM|18|30|你要对 利未 人说：当你们把其中最好的献上为举祭之后，这剩下的就算是你们禾场上的农作物，酒池中的酒。
NUM|18|31|你们和你们的家人可以在任何地方吃；这本是你们的赏赐，是你们在会幕里事奉的酬劳。
NUM|18|32|当你们把其中最好的献上为举祭，就不致于因它担当罪。你们不可玷污 以色列 人的圣物，免得死亡。”
NUM|19|1|耶和华吩咐 摩西 和 亚伦 说：
NUM|19|2|“耶和华所吩咐的律法中，其中一条律例这样说：要吩咐 以色列 人，把一头健康、没有残疾、未曾负轭的红母牛牵到你这里来，
NUM|19|3|交给 以利亚撒 祭司。他要把牛牵到营外，人就在他面前把牛宰了。
NUM|19|4|以利亚撒 祭司要用指头蘸这牛的血，向会幕前面弹七次。
NUM|19|5|人要在他眼前焚烧这母牛，牛的皮、肉、血和粪都要焚烧。
NUM|19|6|祭司要把香柏木、牛膝草和朱红色纱都丢在焚烧牛的火中。
NUM|19|7|祭司要洗衣服，用水洗身，然后才可以进营；祭司必不洁净到晚上。
NUM|19|8|焚烧牛的人也要用水洗衣服，用水洗身，必不洁净到晚上。
NUM|19|9|一个洁净的人要收母牛的灰，存放在营外洁净的地方，为 以色列 会众留作除污秽的水之用。这是为除罪用的。
NUM|19|10|收取母牛灰的人要洗衣服，必不洁净到晚上。这要成为 以色列 人和寄居在他们中间的外人永远的定例。
NUM|19|11|“摸了任何人死尸的，必不洁净七天。
NUM|19|12|那人要在第三天和第七天洁净自己，他就洁净了。若他不在第三天和第七天洁净自己，他就不洁净了。
NUM|19|13|凡摸了死尸，就是死了的人的尸体，又不洁净自己的，就玷污了耶和华的帐幕，这人必从 以色列 中剪除；因为那除污秽的水没有洒在他身上，他就不洁净，污秽还在他身上。
NUM|19|14|“若有人死在帐棚里，条例是这样：凡进那帐棚的，和所有在帐棚里的人，都必不洁净七天。
NUM|19|15|凡敞开的，没有用绳子扎好盖子的器皿，也不洁净。
NUM|19|16|任何人在田野里摸了被刀杀的，或自然死的，或人的骨头，或坟墓，就必不洁净七天。
NUM|19|17|要为这不洁净的人拿一些烧好的除罪灰放在器皿里，倒上清水。
NUM|19|18|一个洁净的人要拿牛膝草蘸在这水中，把水弹在帐棚上，和一切器皿以及帐棚内的人身上，又要弹在那摸了骨头，或摸了被杀的或自然死的，或摸了坟墓的人身上。
NUM|19|19|那洁净的人要在第三天和第七天把水弹在不洁净的人身上，在第七天洁净那人。那人要洗衣服，用水洗澡，到晚上就洁净了。
NUM|19|20|但任何不洁净的人，他若不洁净自己，那人要从会中剪除，因为他玷污了耶和华的圣所，除污秽的水没有洒在他身上，他是不洁净的。
NUM|19|21|这要成为你们永远的定例。此外，那弹除污秽水的人也要洗衣服。凡碰除污秽水的，必不洁净到晚上。
NUM|19|22|不洁净的人所摸的任何东西都不洁净；摸了这东西的人必不洁净到晚上。”
NUM|20|1|正月间， 以色列 全会众到了 寻 的旷野；百姓住在 加低斯 。 米利暗 死在那里，也葬在那里。
NUM|20|2|会众没有水，就聚集反对 摩西 和 亚伦 。
NUM|20|3|百姓与 摩西 争闹，说：“我们恨不得与我们的弟兄一同死在耶和华面前。
NUM|20|4|你们为什么领耶和华的会众到这旷野，使我们和我们的牲畜都死在这里呢？
NUM|20|5|你们为什么领我们从 埃及 上来，把我们带到这坏的地方呢？这地方不能撒种，没有无花果树、葡萄树、石榴树，也没有水喝。”
NUM|20|6|摩西 、 亚伦 离开会众面前，到会幕的门口，脸伏于地；耶和华的荣光向他们显现。
NUM|20|7|耶和华吩咐 摩西 说：
NUM|20|8|“你拿着杖去，和你的哥哥 亚伦 召集会众，在他们眼前吩咐磐石涌出水来，水就会从磐石流出，给会众和他们的牲畜喝。”
NUM|20|9|于是 摩西 遵照耶和华所吩咐他的，从耶和华面前拿了杖去。
NUM|20|10|摩西 和 亚伦 召集会众到磐石前。 摩西 对他们说：“听着，你们这些悖逆的人！我们要叫这磐石流出水来给你们吗？”
NUM|20|11|摩西 举起手来，用杖击打磐石两下，就有许多水流出来，会众和他们的牲畜都喝了。
NUM|20|12|但是耶和华对 摩西 、 亚伦 说：“因为你们不信我，没有在 以色列 人眼前尊我为圣，所以你们必不能领这会众进入我所要赐给他们的地去。”
NUM|20|13|这就是 米利巴 水，因 以色列 人与耶和华争闹，耶和华在他们面前显为圣。
NUM|20|14|摩西 从 加低斯 差遣使者到 以东 王那里，说：“你的弟兄 以色列 这样说：‘你知道我们所遭遇的一切困难。
NUM|20|15|我们的祖先曾下到 埃及 ，我们也在 埃及 住了很多年。然而， 埃及 人却恶待我们和我们的祖先。
NUM|20|16|我们哀求耶和华，他垂听了我们的声音，差遣使者把我们从 埃及 领出来。看哪，我们到了你边界的 加低斯城 。
NUM|20|17|求你让我们穿越你的地。我们不走田间和葡萄园，也不喝井里的水。我们只走王的大路，不偏左右，直到过了你的边界。’”
NUM|20|18|但是， 以东 对他说：“你不可从我这里穿越！否则，我要带刀出去攻击你。”
NUM|20|19|以色列 人对他说：“我们只上大道。如果我和我的牲畜喝了你的水，我必付钱给你。我不求别的事，只求让我步行过去。”
NUM|20|20|以东 说：“你不可经过！”他就率领一大群军队，以强硬的手出来攻击 以色列 。
NUM|20|21|这样， 以东 不肯让 以色列 穿越他的境内， 以色列 就转去，离开他了。
NUM|20|22|以色列 全会众从 加低斯 起行，到了 何珥山 。
NUM|20|23|耶和华在 以东 地边界的 何珥山 对 摩西 、 亚伦 说：
NUM|20|24|“ 亚伦 要归到他祖先 那里。他必不得进入我所赐给 以色列 人的地，因为你们在 米利巴 水的事上违背了我的指示。
NUM|20|25|你要带 亚伦 和他的儿子 以利亚撒 上 何珥山 ，
NUM|20|26|把 亚伦 的圣衣脱下，给他的儿子 以利亚撒 穿上。 亚伦 必归去，死在那里。”
NUM|20|27|摩西 就遵照耶和华的吩咐去做，他们在全会众的眼前上了 何珥山 。
NUM|20|28|摩西 把 亚伦 的圣衣脱下，给他的儿子 以利亚撒 穿上， 亚伦 就死在山顶那里。于是， 摩西 和 以利亚撒 下了山。
NUM|20|29|全会众见 亚伦 死了， 以色列 全家就为 亚伦 举哀三十天。
NUM|21|1|住 尼革夫 的 迦南 人的 亚拉得 王，听说 以色列 从 亚他林 路来，就和 以色列 交战，掳去他们一些人。
NUM|21|2|以色列 向耶和华许愿说：“你若把这百姓真的交在我手中，我就把他们的城镇彻底毁灭。”
NUM|21|3|耶和华垂听了 以色列 的声音，把 迦南 人交出来。 以色列 就把 迦南 人和他们的城镇彻底毁灭。因此，那地方名叫 何珥玛 。
NUM|21|4|他们从 何珥山 起行，绕过 以东 地往 红海 那条路走。在路上，百姓心中烦躁。
NUM|21|5|百姓向上帝和 摩西 发怨言，说：“你们为什么把我们从 埃及 领上来 ，使我们死在旷野呢？这里没有粮食，没有水，我们厌恶这淡而无味的食物。”
NUM|21|6|耶和华派火蛇进入百姓当中去咬他们，于是 以色列 中死了许多百姓。
NUM|21|7|百姓到 摩西 那里，说：“我们有罪了，因为我们向耶和华和你发怨言。求你向耶和华祷告，叫蛇离开我们。”于是 摩西 为百姓祷告。
NUM|21|8|耶和华对 摩西 说：“你要造一条火蛇，挂在杆子上。凡被咬的，一望这蛇就必存活。”
NUM|21|9|摩西 就造了一条铜蛇，挂在杆子上。凡被蛇咬的，一望这铜蛇就活了。
NUM|21|10|以色列 人起行，安营在 阿伯 。
NUM|21|11|又从 阿伯 起行，安营在 以耶．亚巴琳 ，在 摩押 对面的旷野，向日出的方向。
NUM|21|12|又从那里起行，安营在 撒烈谷 。
NUM|21|13|从那里再起行，安营在 亚嫩河 的另一边。这 亚嫩河 在旷野，从 亚摩利 人的境内流出来； 亚嫩河 是 摩押 的边界，在 摩押 和 亚摩利 人之间。
NUM|21|14|所以《耶和华的战记》中提到： “ 苏法 的 哇哈伯 ， 亚嫩河 谷，
NUM|21|15|以及 亚珥 地区众河床的斜坡， 都靠近 摩押 的边境。”
NUM|21|16|以色列 人从那里起行，到了 比珥 。从前耶和华对 摩西 说：“召集百姓，我要给他们水”，说的就是这井。
NUM|21|17|当时， 以色列 人唱这首歌： “井啊，涌出水来！ 你们要向它歌唱！
NUM|21|18|这井是领袖用权杖所挖， 是百姓中的贵族用手杖所掘。” 以色列 人从旷野往 玛他拿 去，
NUM|21|19|从 玛他拿 到 拿哈列 ，从 拿哈列 到 巴末 ，
NUM|21|20|从 巴末 到 摩押 地的谷，又到那可以了望旷野的 毗斯迦山 顶。
NUM|21|21|以色列 差遣使者到 亚摩利 人的王 西宏 那里，说：
NUM|21|22|“求你让我们穿越你的地；我们不岔进田间和葡萄园，也不喝井里的水，只走王的大道，直到过了你的边界。”
NUM|21|23|但 西宏 不让 以色列 人穿越他的境内，就召集他的众百姓出到旷野，要攻击 以色列 ，到了 雅杂 与 以色列 交战。
NUM|21|24|以色列 人用刀杀了他，占领了他的地，从 亚嫩河 到 雅博河 ，直到 亚扪 人的边界，因为 亚扪 人的边防坚固。
NUM|21|25|以色列 人夺取这里所有的城镇，就住在 亚摩利 人的城镇中，包括 希实本 和所属的一切乡镇 。
NUM|21|26|希实本 是 亚摩利 王 西宏 的首都； 西宏 曾与先前的 摩押 王交战，从他手中夺取了他所有的地，直到 亚嫩河 。
NUM|21|27|所以那些作诗歌的说： 你们到 希实本 来吧； 愿 西宏 的城被修造建立。
NUM|21|28|因为有火从 希实本 发出， 有火焰从 西宏 的城冒出， 烧毁了 摩押 的 亚珥 ， 亚嫩河 丘坛的主 。
NUM|21|29|摩押 啊，你有祸了！ 基抹 的百姓啊，你们灭亡了！ 基抹 的男子逃亡， 女子被掳， 交给了 亚摩利 王 西宏 。
NUM|21|30|我们射了他们； 希实本 直到 底本 尽都毁灭 。 我们劫掠，直到 挪法 ； 这 挪法 直延到 米底巴 。
NUM|21|31|这样， 以色列 人就住在 亚摩利 人的地。
NUM|21|32|摩西 差派人去窥探 雅谢 ； 以色列 人占领了 雅谢 附近的乡村，赶出那里的 亚摩利 人。
NUM|21|33|后来， 以色列 人转回，往上 巴珊 的路去。 巴珊 王 噩 率领他的众百姓出来，在 以得来 与他们交战。
NUM|21|34|耶和华对 摩西 说：“不要怕他！因为我已将他和他的众百姓，以及他的地都交在你手中。你要待他如同待住在 希实本 的 亚摩利 王 西宏 一样。”
NUM|21|35|于是他们杀了 巴珊 王和他的众子，以及他的众百姓，没有留下一个幸存者，并且占领了他的地。
NUM|22|1|以色列 人起行，在 摩押 平原， 约旦河 东，对着 耶利哥 安营。
NUM|22|2|西拨 的儿子 巴勒 看见 以色列 向 亚摩利 人所做的一切。
NUM|22|3|摩押 因 以色列 百姓这么多，非常惧怕。 摩押 因 以色列 人的缘故就忧惧。
NUM|22|4|摩押 对 米甸 的长老说：“现在这群人要舔尽我们四围的一切，好像牛舔尽田间的草一样。” 那时， 西拨 的儿子 巴勒 作 摩押 王。
NUM|22|5|他派使者往 大河 附近的 毗夺 去，到 比珥 的儿子 巴兰 的家乡 ，召 巴兰 来，说：“看哪，有一群百姓从 埃及 出来；看哪，他们遮满地面，住在我的对面。
NUM|22|6|现在请你来，为我诅咒这百姓，因为他们比我强大，或许我能打败他们，把他们赶出此地。因为我知道，你为谁祝福，谁就得福；你诅咒谁，谁就受诅咒。”
NUM|22|7|摩押 的长老和 米甸 的长老手里拿着占卜的礼金到 巴兰 那里，将 巴勒 的话告诉他。
NUM|22|8|巴兰 对他们说：“今晚你们在这里过夜，我必照着耶和华向我说的话给你们答覆。” 摩押 的官员就在 巴兰 那里住下。
NUM|22|9|上帝临到 巴兰 那里，说：“你这里的这些人是谁？”
NUM|22|10|巴兰 对上帝说：“ 摩押 王 西拨 的儿子 巴勒 送信给我：
NUM|22|11|‘看哪，从 埃及 出来的百姓遮满了地面，现在请你来，为我诅咒他们，或许我能打败他们，把他们赶走。’”
NUM|22|12|上帝对 巴兰 说：“你不可跟他们去，也不可诅咒这百姓，因为他们是蒙福的。”
NUM|22|13|巴兰 早晨起来，对 巴勒 的官员说：“你们回本地去吧，因为耶和华不允许我和你们一起去。”
NUM|22|14|摩押 的官员就起来，到 巴勒 那里，说：“ 巴兰 不肯和我们一起来。”
NUM|22|15|巴勒 又差遣比这些更多，更尊贵的官员。
NUM|22|16|他们来到 巴兰 那里，对他说：“ 西拨 的儿子 巴勒 这样说：‘请你不要再推辞到我这里来！
NUM|22|17|我必使你得极大的尊荣，无论你向我要什么，我都给你。只求你来为我诅咒这百姓。’”
NUM|22|18|巴兰 回答 巴勒 的臣仆说：“ 巴勒 就是将他满屋的金银给我，我也不能做任何大小的事，违背耶和华－我上帝的指示。
NUM|22|19|现在请你们今晚也在这里住下，我好知道耶和华还要对我说什么。”
NUM|22|20|上帝在夜里临到 巴兰 那里，说：“这些人若来求你，你就起来跟他们去吧，只是你必须照着我对你说的话去做。”
NUM|22|21|巴兰 早晨起来，备了驴，就和 摩押 的官员一同去了。
NUM|22|22|上帝因他去就怒气发作；耶和华的使者站在路中间敌对他。他骑着驴，有两个仆人跟随他。
NUM|22|23|驴看见耶和华的使者站在路中间，手里有拔出来的刀，就离开了路，岔入田间。 巴兰 就打驴，要它回到路上。
NUM|22|24|耶和华的使者站在葡萄园的窄路上，这边有墙，那边也有墙。
NUM|22|25|驴看见耶和华的使者，就往墙挤去，把 巴兰 的脚挤到墙上； 巴兰 再打驴。
NUM|22|26|耶和华的使者又往前去，站在狭窄的地方，那里左右都无路可转。
NUM|22|27|驴看见耶和华的使者，就伏在 巴兰 底下。 巴兰 怒气发作，用杖打驴。
NUM|22|28|耶和华使驴开口，对 巴兰 说：“我向你做了什么，你竟打我这三次呢？”
NUM|22|29|巴兰 对驴说：“因为你戏弄我，我恨不得手中有刀，现在就把你杀了。”
NUM|22|30|驴对 巴兰 说：“我不是你从小直到今天所骑的驴吗？我平时有这样待过你吗？” 巴兰 说：“没有。”
NUM|22|31|耶和华使 巴兰 的眼目明亮，他看见耶和华的使者站在路中间，手里有拔出来的刀； 巴兰 就低头俯伏下拜。
NUM|22|32|耶和华的使者对他说：“你为什么这三次打你的驴呢？看哪，我出来敌对你，因为这路在我面前已经偏离了。
NUM|22|33|驴看见我就从我面前回避了这三次；驴若没有回避我，我早把你杀了，留它存活。”
NUM|22|34|巴兰 对耶和华的使者说：“我有罪了。我不知道你站在路中间阻挡我；现在你若看为不好，我就回去。”
NUM|22|35|耶和华的使者对 巴兰 说：“你和这些人去吧！你只要说我对你说的话。”于是 巴兰 和 巴勒 的官员一同去了。
NUM|22|36|巴勒 听见 巴兰 来了，就到 摩押 的城 去迎接他；这城是在边界的 亚嫩河 旁。
NUM|22|37|巴勒 对 巴兰 说：“我不是急切地派人到你那里去召你吗？你为何不到我这里来呢？我岂不能使你得尊荣吗？”
NUM|22|38|巴兰 对 巴勒 说：“看哪，我已经到你这里来了！现在我岂能擅自说什么呢？上帝将什么话放在我口中，我就说什么。”
NUM|22|39|巴兰 和 巴勒 同去，来到 基列．胡琐 。
NUM|22|40|巴勒 宰了牛羊为祭物，送给 巴兰 和陪伴他的官员。
NUM|22|41|到了早晨， 巴勒 领 巴兰 到 巴末．巴力 ，从那里可以看到一部分 以色列 的百姓。
NUM|23|1|巴兰 对 巴勒 说：“你要在这里为我筑七座坛，又要在这里为我预备七头公牛，七只公羊。”
NUM|23|2|巴勒 照 巴兰 的话做了。 巴勒 和 巴兰 在每座坛上献一头公牛，一只公羊。
NUM|23|3|巴兰 对 巴勒 说：“你站在你的燔祭旁边，我要往前去，或许耶和华会向我显现。他指示我什么事，我必告诉你。”于是 巴兰 上到一个光秃的高地。
NUM|23|4|上帝向 巴兰 显现。 巴兰 对他说：“我预备了七座坛，在每座坛上献了一头公牛，一只公羊。”
NUM|23|5|耶和华把话放在 巴兰 口中，说：“你回到 巴勒 那里，要这样说。”
NUM|23|6|他就回到 巴勒 那里，看哪， 巴勒 和 摩押 的众官员站在燔祭旁边。
NUM|23|7|巴兰 唱起诗歌说： “ 巴勒 领我出 亚兰 ， 摩押 王领我出东方的山脉： ‘来啊，为我诅咒 雅各 ； 来啊，怒骂 以色列 。’
NUM|23|8|上帝没有诅咒的， 我焉能诅咒？ 耶和华没有怒骂的， 我岂能怒骂？
NUM|23|9|我从磐石的巅峰看到他， 我从山丘望见他。 看哪，这是独居的民， 不算在列国中。
NUM|23|10|谁能数点 雅各 的尘土？ 谁能计算 以色列 的尘沙 ？ 我愿如正直人之死而死； 我愿如正直人之终而终。”
NUM|23|11|巴勒 对 巴兰 说：“你向我做的是什么呢？我带你来诅咒我的仇敌，看哪，你竟为他们祝福。”
NUM|23|12|他回答说：“耶和华放在我口中的话，我岂能不谨慎地说呢？”
NUM|23|13|巴勒 对他说：“请你跟我到别的地方，在那里可以看见他们。你只能看见他们的一部分，却不能看见全部。请你在那里为我诅咒他们。”
NUM|23|14|于是 巴勒 领 巴兰 到了 琐腓 的田野，上了 毗斯迦山 顶 ，筑了七座坛，在每座坛上献一头公牛，一只公羊。
NUM|23|15|巴兰 对 巴勒 说：“你站在你的燔祭旁边，我要到那边去看看。”
NUM|23|16|耶和华向 巴兰 显现，把话放在他口中，说：“你回到 巴勒 那里，要这样说。”
NUM|23|17|他回到 巴勒 那里，看哪， 巴勒 站在燔祭旁边， 摩押 的官员也和他在一起。 巴勒 对他说：“耶和华说了什么呢？”
NUM|23|18|巴兰 唱起诗歌说： “ 巴勒 啊，起来，听； 西拨 的儿子啊，侧耳听我。
NUM|23|19|上帝非人，必不致说谎， 也非人子，必不致后悔。 他说了岂不照着做呢？ 他发了言岂不实现呢？
NUM|23|20|看哪，我奉命祝福； 上帝赐福，我不能扭转。
NUM|23|21|他未见 雅各 中有灾难 ， 也未见 以色列 中有祸患 。 耶和华－他的上帝和他同在； 在他中间有欢呼王的声音。
NUM|23|22|上帝领他们出 埃及 ， 为 以色列 有如野牛的角。
NUM|23|23|绝没有法术可以伤 雅各 ， 没有占卜可以害 以色列 。 现在，人论及 雅各 ，论及 以色列 必说： ‘上帝成就了何等的事啊！’
NUM|23|24|看哪，这百姓兴起如母狮， 挺身像公狮， 未曾吃猎物， 未曾喝被杀者的血， 绝不躺卧。”
NUM|23|25|巴勒 对 巴兰 说：“你一点也不要诅咒他们，一点也不要为他们祝福！”
NUM|23|26|巴兰 回答 巴勒 说：“我不是告诉过你：‘凡耶和华所说的，我必须遵行’吗？”
NUM|23|27|巴勒 对 巴兰 说：“来，我领你到别的地方，或许上帝喜欢你在那里为我诅咒他们。”
NUM|23|28|巴勒 就领 巴兰 到那可了望旷野的 毗珥山 顶。
NUM|23|29|巴兰 对 巴勒 说：“你要在这里为我筑七座坛，又要在这里为我预备七头公牛，七只公羊。”
NUM|23|30|巴勒 就照 巴兰 的话做，在每座坛上献一头公牛，一只公羊。
NUM|24|1|巴兰 见耶和华喜欢赐福给 以色列 ，就不像前两次去求法术，却面向旷野。
NUM|24|2|巴兰 举目，看见 以色列 人照着支派扎营。上帝的灵就临到他身上，
NUM|24|3|他唱起诗歌说： “ 比珥 的儿子 巴兰 说， 眼目关闭 的人说，
NUM|24|4|听见上帝的言语， 得见全能者的异象， 俯伏着，眼睛却睁开的人说：
NUM|24|5|雅各 啊，你的帐棚何等华美！ 以色列 啊，你的帐幕何其华丽！
NUM|24|6|如连绵的山谷， 如河畔的园子， 如耶和华栽种的沉香树， 又如水边的香柏木。
NUM|24|7|水要从他的桶里流出， 种子要撒在多水之处。 他的王必超越 亚甲 ， 他的国必要振兴。
NUM|24|8|上帝领他出 埃及 ， 为他有如野牛的角。 他要吞灭那敌对他的国， 压碎他们的骨头， 用箭射透他们。
NUM|24|9|他蹲如公狮， 卧如母狮， 谁敢惹他？ 凡为你祝福的，愿他蒙福； 凡诅咒你的，愿他受诅咒。”
NUM|24|10|巴勒 向 巴兰 怒气发作，就紧握拳头 。 巴勒 对 巴兰 说：“我召你来诅咒我的仇敌，看哪，你竟然这三次为他们祝福。
NUM|24|11|如今你赶快回本地去吧！我想使你大得尊荣，看哪，耶和华却阻止你得尊荣。”
NUM|24|12|巴兰 对 巴勒 说：“我不是对你所差遣到我那里的使者说：
NUM|24|13|‘ 巴勒 就是把他满屋的金银给我，我也不能违背耶和华的指示，随自己的心意做好做歹。耶和华说什么，我就说什么。’
NUM|24|14|现在，看哪，我要回到我的百姓那里。来，让我告诉你这百姓日后要怎样对待你的百姓。”
NUM|24|15|他就唱起诗歌说： “ 比珥 的儿子 巴兰 说， 眼目关闭的人说，
NUM|24|16|听见上帝的言语， 明白至高者的知识， 看见全能者的异象， 俯伏着，眼睛却睁开的人说：
NUM|24|17|我看见他，却不在现时； 我望见他，却不在近处。 有星出于 雅各 ， 有杖从 以色列 兴起， 必打破 摩押 的额头， 必毁坏所有的 塞特 人 。
NUM|24|18|以东 将成为产业， 西珥 将成为它敌人的产业 ； 但 以色列 却要得胜。
NUM|24|19|有一位出于 雅各 的，必掌大权， 他要除灭城中的幸存者。”
NUM|24|20|巴兰 看见 亚玛力 人，就唱起诗歌说： “ 亚玛力 是诸国之首， 但它终必永远沉沦 。”
NUM|24|21|巴兰 看见 基尼 人，就唱起诗歌说： “你的住处坚固； 你的巢窝造在岩石中。
NUM|24|22|然而 基尼 族 必被吞灭， 直到何时 亚述 把你掳去？ ”
NUM|24|23|巴兰 又唱起诗歌说： “哀哉！若上帝做这事， 谁能存活呢？
NUM|24|24|有船只 从 基提 边界来到， 要压制 亚述 ， 要压制 希伯 ； 他也必永远沉沦 。”
NUM|24|25|于是 巴兰 起来，回本地去； 巴勒 也回他的路去了。
NUM|25|1|以色列 人住在 什亭 ，百姓开始与 摩押 女子行淫。
NUM|25|2|这些女子请百姓一同为她们的神明献祭，百姓吃了祭物，跪拜她们的神明。
NUM|25|3|以色列 与 巴力．毗珥 联合，耶和华的怒气就向 以色列 发作。
NUM|25|4|耶和华对 摩西 说：“拿下百姓中所有的领袖，对着太阳把他们悬挂在我面前，使我向 以色列 所发的怒气可以平息。”
NUM|25|5|于是 摩西 对 以色列 的审判官说：“你们的人若有与 巴力．毗珥 联合的，你们各人就要把他们杀了。”
NUM|25|6|摩西 和 以色列 全会众在会幕门口哭泣的时候，看哪，有一个 以色列 人，在他们眼前带着一个 米甸 女子，到他弟兄那里。
NUM|25|7|亚伦 祭司的孙子， 以利亚撒 的儿子 非尼哈 看见了，就从会众中起来，手里拿着枪，
NUM|25|8|跟这 以色列 人进入帐棚，刺穿了二人，就是 以色列 人和那女子的肚腹。这样， 以色列 人遭受的瘟疫就停止了。
NUM|25|9|遭瘟疫死的，有二万四千人。
NUM|25|10|耶和华吩咐 摩西 说：
NUM|25|11|“ 亚伦 祭司的孙子， 以利亚撒 的儿子 非尼哈 ，使我的愤怒转离 以色列 人，因为在他们中间，他以我的妒忌为他的妒忌，使我不在妒忌中毁灭 以色列 人。
NUM|25|12|因此，你要说：‘看哪，我将我平安的约赐给他。
NUM|25|13|这是他和他的后裔永远当祭司职任的约，因他为了上帝而妒忌，他为 以色列 人赎罪。’”
NUM|25|14|那与 米甸 女子一起被杀的 以色列 人，名叫 心利 ，是 撒路 的儿子，是 西缅 一个父家的领袖。
NUM|25|15|那被杀的 米甸 女子，名叫 哥斯比 ，是 苏珥 的女儿； 苏珥 是 米甸 一个父家的领袖。
NUM|25|16|耶和华吩咐 摩西 说：
NUM|25|17|“你要苦害 米甸 人，击杀他们；
NUM|25|18|因为他们用诡计苦害你们，在 毗珥 的事上和他们的姊妹， 米甸 领袖的女儿 哥斯比 的事上，欺骗了你们；在瘟疫的日子，这女子因 毗珥 的事件被杀了。”
NUM|26|1|瘟疫过了之后，耶和华对 摩西 和 亚伦 祭司的儿子 以利亚撒 说：
NUM|26|2|“你们要将 以色列 全会众，按他们的父家，凡二十岁以上能出去为 以色列 打仗的，计算总数。”
NUM|26|3|摩西 和 以利亚撒 祭司在 摩押 平原与 耶利哥 相对的 约旦河 边吩咐他们说：
NUM|26|4|“计算你们中间从二十岁以上的人数。”正如耶和华所吩咐 摩西 的。 从 埃及 地出来的 以色列 人如下：
NUM|26|5|以色列 的长子是 吕便 。 吕便 的众子：属 哈诺 的，有 哈诺 族；属 法路 的，有 法路 族；
NUM|26|6|属 希斯伦 的，有 希斯伦 族；属 迦米 的，有 迦米 族。
NUM|26|7|这就是 吕便 的各族；被数的共有四万三千七百三十名。
NUM|26|8|法路 的儿子是 以利押 。
NUM|26|9|以利押 的儿子是 尼母利 、 大坍 、 亚比兰 。这 大坍 、 亚比兰 ，就是从会中选出来，当 可拉 一伙的人向耶和华争闹的时候，一起向 摩西 、 亚伦 争闹的；
NUM|26|10|地开了裂口，吞了他们和 可拉 ， 可拉 一伙的人也一同死亡。当时火吞灭了二百五十个人；他们就成为鉴戒。
NUM|26|11|然而 可拉 的众子没有死亡。
NUM|26|12|按着宗族， 西缅 的众子：属 尼母利 的，有 尼母利 族；属 雅悯 的，有 雅悯 族；属 雅斤 的，有 雅斤 族；
NUM|26|13|属 谢拉 的，有 谢拉 族；属 扫罗 的，有 扫罗 族。
NUM|26|14|这就是 西缅 的各族，共有二万二千二百名。
NUM|26|15|按着宗族， 迦得 的众子：属 洗分 的，有 洗分 族；属 哈基 的，有 哈基 族；属 书尼 的，有 书尼 族；
NUM|26|16|属 阿斯尼 的，有 阿斯尼 族；属 以利 的，有 以利 族；
NUM|26|17|属 亚律 的，有 亚律 族；属 亚列利 的，有 亚列利 族。
NUM|26|18|这就是 迦得 子孙的各族；他们被数的共有四万零五百名。
NUM|26|19|犹大 的儿子是 珥 和 俄南 。 珥 和 俄南 死在 迦南 地。
NUM|26|20|按着宗族， 犹大 的众子：属 示拉 的，有 示拉 族；属 法勒斯 的，有 法勒斯 族；属 谢拉 的，有 谢拉 族。
NUM|26|21|法勒斯 的众子：属 希斯仑 的，有 希斯仑 族；属 哈母勒 的，有 哈母勒 族。
NUM|26|22|这就是 犹大 的各族；他们被数的共有七万六千五百名。
NUM|26|23|按着宗族， 以萨迦 的众子：属 陀拉 的，有 陀拉 族；属 普瓦 的，有 普瓦 族；
NUM|26|24|属 雅述 的，有 雅述 族；属 伸仑 的，有 伸仑 族。
NUM|26|25|这就是 以萨迦 的各族；他们被数的共有六万四千三百名。
NUM|26|26|按着宗族， 西布伦 的众子：属 西烈 的，有 西烈 族；属 以伦 的，有 以伦 族；属 雅利 的，有 雅利 族。
NUM|26|27|这就是 西布伦 的各族；他们被数的共有六万零五百名。
NUM|26|28|按着宗族， 约瑟 的儿子有 玛拿西 、 以法莲 。
NUM|26|29|玛拿西 的众子：属 玛吉 的，有 玛吉 族； 玛吉 生 基列 ；属 基列 的，有 基列 族。
NUM|26|30|这就是 基列 的众子：属 伊以谢 的，有 伊以谢 族；属 希勒 的，有 希勒 族；
NUM|26|31|属 亚斯烈 的，有 亚斯烈 族；属 示剑 的，有 示剑 族；
NUM|26|32|属 示米大 的，有 示米大 族；属 希弗 的，有 希弗 族。
NUM|26|33|希弗 的儿子 西罗非哈 没有儿子，只有女儿。 西罗非哈 的女儿的名字是 玛拉 、 挪阿 、 曷拉 、 密迦 、 得撒 。
NUM|26|34|这就是 玛拿西 的各族；他们被数的共有五万二千七百名。
NUM|26|35|这就是按着宗族， 以法莲 的众子：属 书提拉 的，有 书提拉 族；属 比结 的，有 比结 族；属 他罕 的，有 他罕 族。
NUM|26|36|这就是 书提拉 的众子：属 以兰 的，有 以兰 族。
NUM|26|37|这就是 以法莲 子孙的各族；他们被数的共有三万二千五百名。按着宗族，以上这些都是 约瑟 的子孙。
NUM|26|38|按着宗族， 便雅悯 的众子：属 比拉 的，有 比拉 族；属 亚实别 的，有 亚实别 族；属 亚希兰 的，有 亚希兰 族；
NUM|26|39|属 书反 的，有 书反 族；属 户反 的，有 户反 族。
NUM|26|40|比拉 的儿子是 亚勒 、 乃幔 ；属 亚勒 的 ，有 亚勒 族；属 乃幔 的，有 乃幔 族。
NUM|26|41|按着宗族，这就是 便雅悯 的子孙；他们被数的共有四万五千六百名。
NUM|26|42|这就是按着宗族， 但 的众子：属 书含 的，有 书含 族。按着宗族，这就是 但 的各族。
NUM|26|43|按照他们被数的， 书含 全宗族共有六万四千四百名。
NUM|26|44|按着宗族， 亚设 的众子：属 音拿 的，有 音拿 族；属 亦施韦 的，有 亦施韦 族；属 比利亚 的，有 比利亚 族。
NUM|26|45|比利亚 的众子：属 希别 的，有 希别 族；属 玛结 的，有 玛结 族。
NUM|26|46|亚设 的女儿名叫 西拉 。
NUM|26|47|这就是 亚设 子孙的各族；他们被数的共有五万三千四百名。
NUM|26|48|按着宗族， 拿弗他利 的众子：属 雅薛 的，有 雅薛 族；属 沽尼 的，有 沽尼 族；
NUM|26|49|属 耶色 的，有 耶色 族；属 示冷 的，有 示冷 族。
NUM|26|50|按着宗族，这就是 拿弗他利 的各族；他们被数的共有四万五千四百名。
NUM|26|51|这就是 以色列 人中被数的，共有六十万零一千七百三十名。
NUM|26|52|耶和华吩咐 摩西 说：
NUM|26|53|“你要按着人名的数目，将地分给这些人为产业。
NUM|26|54|人多的要多给他们产业，人少的要少给他们产业；各照被数的人数分配产业。
NUM|26|55|此外，要以抽签来分地，按着父系各支派的名字承受产业。
NUM|26|56|要根据抽签，看人数的多寡，给他们分配产业。”
NUM|26|57|这就是按着宗族，被数的 利未 人：属 革顺 的，有 革顺 族；属 哥辖 的，有 哥辖 族；属 米拉利 的，有 米拉利 族。
NUM|26|58|这就是 利未 的宗族： 立尼 族、 希伯伦 族、 玛利 族、 母示 族、 可拉 族。 哥辖 生 暗兰 。
NUM|26|59|暗兰 的妻子名叫 约基别 ，是 利未 的女儿，是 利未 在 埃及 所生的。她给 暗兰 生了 亚伦 、 摩西 ，和他们的姊姊 米利暗 。
NUM|26|60|亚伦 生 拿答 、 亚比户 、 以利亚撒 、 以他玛 。
NUM|26|61|拿答 、 亚比户 在耶和华面前献凡火的时候死了。
NUM|26|62|利未 人中，凡一个月以上所有被数的男子，共有二万三千名。他们没有数在 以色列 人中；因为在 以色列 人中，没有分给他们产业。
NUM|26|63|这些是 摩西 和 以利亚撒 祭司所数的；他们在 摩押 平原与 耶利哥 相对的 约旦河 边数点 以色列 人。
NUM|26|64|这些被数的人中，没有一个是 摩西 和 亚伦 祭司先前在 西奈 旷野所数的 以色列 人，
NUM|26|65|因为耶和华论到他们说：“他们必死在旷野。”所以，除了 耶孚尼 的儿子 迦勒 和 嫩 的儿子 约书亚 以外，他们一个也没有存留。
NUM|27|1|约瑟 的儿子 玛拿西 的宗族中，有 玛拿西 的玄孙， 玛吉 的曾孙， 基列 的孙子， 希弗 的儿子 西罗非哈 的女儿，名叫 玛拉 、 挪阿 、 曷拉 、 密迦 、 得撒 。她们前来，
NUM|27|2|站在会幕门口，在 摩西 和 以利亚撒 祭司，以及众领袖与全会众面前，说：
NUM|27|3|“我们的父亲死在旷野。他没有与 可拉 同伙聚集攻击耶和华，是在自己的罪中死的；他没有儿子。
NUM|27|4|为什么因我们的父亲没有儿子就把他的名从他族中除掉呢？求你们在我们父亲的兄弟中分给我们产业。”
NUM|27|5|于是， 摩西 将她们的案件呈到耶和华面前。
NUM|27|6|耶和华对 摩西 说：
NUM|27|7|“ 西罗非哈 的女儿说得有理。你定要在她们父亲的兄弟中，把地分给她们为业，把她们父亲的产业传给她们。
NUM|27|8|你也要吩咐 以色列 人说：‘人死了，若没有儿子，就要把他的产业传给他的女儿。
NUM|27|9|他若没有女儿，就要把他的产业给他的兄弟。
NUM|27|10|他若没有兄弟，就要把他的产业给他父亲的兄弟。
NUM|27|11|他父亲若没有兄弟，就要把他的产业给他族中最近的亲属继承为业。’”这要作 以色列 人的律例典章，是照耶和华所吩咐 摩西 的。
NUM|27|12|耶和华对 摩西 说：“你上这 亚巴琳山脉 ，看我所赐给 以色列 人的地。
NUM|27|13|看了以后，你也必归到你祖先 那里，像你哥哥 亚伦 归去一样。
NUM|27|14|因为你们在 寻 的旷野，当会众争闹的时候，违背了我的命令，在取水之事上没有在会众眼前尊我为圣。”这水就是 寻 的旷野中， 加低斯 的 米利巴 水。
NUM|27|15|摩西 对耶和华说：
NUM|27|16|“愿耶和华，赐万人气息的上帝，立一个人治理会众，
NUM|27|17|可以在他们面前出入，引导他们进出，免得耶和华的会众如同没有牧人的羊群一般。”
NUM|27|18|耶和华对 摩西 说：“ 嫩 的儿子 约书亚 是一个有圣灵的人；你要领他来，为他按手，
NUM|27|19|使他站在 以利亚撒 祭司和全会众面前，在他们眼前委派他，
NUM|27|20|又将你的尊荣给他一些，好使 以色列 全会众都听从他。
NUM|27|21|他要站在 以利亚撒 祭司面前； 以利亚撒 要凭乌陵的判断，在耶和华面前为他求问。他和 以色列 全会众都要照 以利亚撒 的指示出入。”
NUM|27|22|于是 摩西 照耶和华所吩咐他的，将 约书亚 领来，使他站在 以利亚撒 祭司和全会众面前，
NUM|27|23|为他按手，委派他，是照耶和华藉 摩西 所说的。
NUM|28|1|耶和华吩咐 摩西 说：
NUM|28|2|“你要吩咐 以色列 人说：‘你们要按时把我的供物，就是献给我作馨香火祭的食物，献给我。’
NUM|28|3|要对他们说：‘这是当献给耶和华的火祭：每天两只没有残疾一岁的小公羊，作为经常献的燔祭。
NUM|28|4|早晨献第一只小公羊，黄昏献第二只小公羊；
NUM|28|5|又用十分之一伊法细面和四分之一欣捣成的油，调和作为素祭。
NUM|28|6|这是在 西奈山 上规定为经常献的燔祭，是献给耶和华为馨香的火祭。
NUM|28|7|为每只小公羊，要有四分之一欣的浇酒祭；在圣所中，你要将醇酒献给耶和华作浇酒祭。
NUM|28|8|黄昏你献第二只小公羊，要照早晨的素祭和同献的浇酒祭献上，作为馨香的火祭，献给耶和华。’”
NUM|28|9|“在安息日，要献两只没有残疾，一岁的小公羊、十分之二伊法调了油的细面为素祭，和同献的浇酒祭。
NUM|28|10|除了经常献的燔祭和同献的浇酒祭之外，这是每一个安息日当献的燔祭。”
NUM|28|11|“每月初一，要将两头公牛犊、一只公绵羊、七只没有残疾一岁的小公羊，献给耶和华为燔祭。
NUM|28|12|为每头公牛，要用十分之三伊法调了油的细面作为素祭；为那只公绵羊，要用十分之二伊法调了油的细面作为素祭；
NUM|28|13|为每只小公羊，要用十分之一伊法调了油的细面作为素祭。这是馨香的燔祭，是献给耶和华的火祭。
NUM|28|14|每头公牛要有半欣的浇酒祭，每只公绵羊三分之一欣的浇酒祭，每只小公羊四分之一欣的浇酒祭。这是一年之中每月初一当献的燔祭。
NUM|28|15|除了经常献的燔祭和同献的浇酒祭之外，又要将一只公山羊，献给耶和华为赎罪祭。”
NUM|28|16|“正月十四日是向耶和华守的逾越节。
NUM|28|17|这月十五日是节期，要吃无酵饼七日。
NUM|28|18|第一日要有圣会，任何劳动的工都不可做。
NUM|28|19|要把火祭，就是两头公牛犊，一只公绵羊、七只一岁的小公羊，都要没有残疾的，献给耶和华为燔祭。
NUM|28|20|要同时献调了油的细面为素祭：每头公牛要献十分之三伊法；每只公绵羊要献十分之二伊法；
NUM|28|21|为那七只小公羊，每只要献十分之一伊法。
NUM|28|22|此外，要献一只公山羊作赎罪祭，为你们赎罪。
NUM|28|23|除了早晨经常献的燔祭之外，你们也要献这些祭。
NUM|28|24|一连七天，在经常献的燔祭和同献的浇酒祭之外，每天要这样把馨香火祭的食物献给耶和华。
NUM|28|25|第七日要有圣会，任何劳动的工都不可做。”
NUM|28|26|“七七初熟节，就是你们献初熟谷物给耶和华为素祭的那一天，要宣告圣会；任何劳动的工都不可做。
NUM|28|27|要将两头公牛犊，一只公绵羊，七只一岁的小公羊，作为馨香的燔祭献给耶和华。
NUM|28|28|要同时献调了油的细面为素祭：每头公牛要献十分之三伊法；每只公绵羊要献十分之二伊法；
NUM|28|29|为那七只小公羊，每只要献十分之一伊法。
NUM|28|30|此外，要献一只公山羊为你们赎罪。
NUM|28|31|除了经常献的燔祭和同献的素祭，你们也要献上这些没有残疾的，和同献的浇酒祭。”
NUM|29|1|“七月初一，你们当有圣会；任何劳动的工都不可做，是你们当守为吹角的日子。
NUM|29|2|你们要将一头公牛犊、一只公绵羊、七只一岁的小公羊，都是没有残疾的，献给耶和华为馨香的燔祭。
NUM|29|3|要同时献调了油的细面为素祭：每头公牛要献十分之三伊法；每只公绵羊要献十分之二伊法；
NUM|29|4|为那七只小公羊，每只要献十分之一伊法。
NUM|29|5|此外，要献一只公山羊作赎罪祭，为你们赎罪。
NUM|29|6|除了初一的燔祭和同献的素祭、经常献的燔祭与同献的素祭，以及同献的浇酒祭以外，这些都照例作为馨香的火祭献给耶和华。”
NUM|29|7|“七月初十，你们当有圣会；要刻苦己心，任何工都不可做。
NUM|29|8|要将一头公牛犊、一只公绵羊、七只一岁的小公羊，都是没有残疾的，献给耶和华为馨香的燔祭。
NUM|29|9|要同时献调了油的细面为素祭：每头公牛要献十分之三伊法；每只公绵羊要献十分之二伊法；
NUM|29|10|为那七只小公羊，每只要献十分之一伊法。
NUM|29|11|又要献一只公山羊为赎罪祭。这是在赎罪祭和经常献的燔祭，以及同献的素祭和浇酒祭以外所献的。”
NUM|29|12|“七月十五日，你们当有圣会；任何劳动的工都不可做，要向耶和华守节七天。
NUM|29|13|要将十三头公牛犊、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，献上作火祭，是献给耶和华馨香的燔祭。
NUM|29|14|要同时献调了油的细面为素祭：为那十三头公牛犊，每头要献十分之三伊法；为那两只公绵羊，每只要献十分之二伊法；
NUM|29|15|为那十四只小公羊，每只要献十分之一伊法。
NUM|29|16|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|17|“第二日要献十二头公牛犊、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，
NUM|29|18|并为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|19|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|20|“第三日要献十一头公牛、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，
NUM|29|21|并为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|22|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|23|“第四日要献十头公牛、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，
NUM|29|24|并为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|25|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|26|“第五日要献九头公牛、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，
NUM|29|27|并为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|28|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|29|“第六日要献八头公牛、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，
NUM|29|30|并为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|31|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|32|“第七日要献七头公牛、两只公绵羊、十四只一岁的小公羊，都是没有残疾的，
NUM|29|33|并为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|34|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|35|“第八日你们当有严肃会；任何劳动的工都不可做；
NUM|29|36|要将一头公牛、一只公绵羊、七只一岁的小公羊，都是没有残疾的，献上作火祭，是献给耶和华馨香的燔祭。
NUM|29|37|要为公牛、公绵羊和小公羊，按数照例奉献同献的素祭和浇酒祭。
NUM|29|38|又要献一只公山羊为赎罪祭。这是在经常献的燔祭、同献的素祭和浇酒祭以外所献的。
NUM|29|39|“这些祭要在你们的节期献给耶和华，都是在所许的愿和甘心献的以外所献的，作为你们的燔祭、素祭、浇酒祭和平安祭。”
NUM|29|40|于是， 摩西 照耶和华所吩咐他的一切话告诉 以色列 人。
NUM|30|1|摩西 对 以色列 各支派的领袖说：“这是耶和华所吩咐的话：
NUM|30|2|人若向耶和华许愿或起誓，要约束自己，就不可食言，必须照口中所出的一切话去做。
NUM|30|3|女子年轻，还在父家的时候，若向耶和华许愿，要约束自己，
NUM|30|4|她父亲听见她所许的愿和约束自己的话，却向她默默不言，她所许的愿和约束自己的话就都有效。
NUM|30|5|但是，若她父亲在听见的日子不允许她一切所许的愿和约束自己的话，这就不算为有效；耶和华也必赦免她，因为她的父亲不允许。
NUM|30|6|她若已出嫁，有愿在身，或口中出了约束自己的冒失话，
NUM|30|7|她丈夫听见了，却在听见的日子向她默默不言，她所许的愿和约束自己的话就都有效。
NUM|30|8|但是，若她丈夫在听见的日子不允许，丈夫就废了她所许的愿和口中所出约束自己的冒失话；耶和华也必赦免她。
NUM|30|9|寡妇或被休的妇人所许的愿，她所有约束自己的话，都是有效的。
NUM|30|10|她若在丈夫家里许了愿或起了誓，要约束自己，
NUM|30|11|丈夫听见了，却向她默默不言，没有不允许，她所许的愿和约束自己的话就都有效。
NUM|30|12|她丈夫听见的日子，若把这些全废了，她口中一切所许的愿或约束自己的话就不算为有效。她丈夫已把这些都废了，耶和华也必赦免她。
NUM|30|13|凡她所许的愿和刻苦约束自己所起的誓，丈夫可以坚立，也可以废去。
NUM|30|14|倘若她丈夫天天向她默默不言，这就算是坚立她一切所许的愿或约束自己的话；因为丈夫在听见的日子向她默默不言，就算是坚立了这些话。
NUM|30|15|但她丈夫听见了，以后若再废了这些话，就要担当妇人的罪孽。”
NUM|30|16|这是关于丈夫待妻子，父亲待女儿，女儿年轻还在父家，耶和华所吩咐 摩西 的条例。
NUM|31|1|耶和华吩咐 摩西 说：
NUM|31|2|“你要为 以色列 人向 米甸 人报仇，然后归到你祖先 那里。”
NUM|31|3|摩西 吩咐百姓说：“要在你们中间叫人带兵器去攻击 米甸 ，为耶和华向 米甸 报仇。
NUM|31|4|从 以色列 众支派中，每支派要派一千人去打仗。”
NUM|31|5|于是从 以色列 千万人中，每支派征召一千人，一共一万二千名，带着兵器预备打仗。
NUM|31|6|摩西 派他们去打仗，每支派一千人；又派 以利亚撒 祭司的儿子 非尼哈 同去； 非尼哈 手里拿着圣所的器皿和吹号的号筒。
NUM|31|7|他们遵照耶和华所吩咐 摩西 的，与 米甸 打仗，杀了所有的男丁。
NUM|31|8|在所杀的人中，他们杀了 米甸 的王，就是 以未 、 利金 、 苏珥 、 户珥 、 利巴 五个 米甸 的王，又用刀杀了 比珥 的儿子 巴兰 。
NUM|31|9|以色列 人掳了 米甸 的妇女和孩童，抢夺他们一切的牲畜、牛羊和所有的财物，
NUM|31|10|又用火焚烧了他们所住的一切城镇和所有的营寨。
NUM|31|11|以色列 人把一切掳物和掠物，连人和牲畜都带走，
NUM|31|12|将俘虏、掠物、掳物带到 摩押 平原，在 约旦河 边与 耶利哥 相对的营地，交给 摩西 和 以利亚撒 祭司，以及 以色列 的会众。
NUM|31|13|摩西 和 以利亚撒 祭司，以及会众中所有的领袖，都出营迎接他们。
NUM|31|14|摩西 向打仗回来的军官，就是千夫长和百夫长发怒。
NUM|31|15|摩西 对他们说：“你们要让这所有的妇女活着吗？
NUM|31|16|看哪，正是这些妇女，因 巴兰 的话，在 毗珥 的事上导致 以色列 人背叛耶和华，以致耶和华的会众遭遇瘟疫。
NUM|31|17|现在，你们要杀所有的男孩，也要把所有曾与男人同房共寝的女子都杀了。
NUM|31|18|但那些未曾与男人同房共寝的女孩，你们可以让她们存活。
NUM|31|19|你们和你们所掳来的人，要住在营外七天；凡杀了人的，和一切摸了尸体的，要在第三日和第七日洁净自己。
NUM|31|20|你们也要洁净一切的衣服，以及用皮革、山羊毛和木头做的任何东西。”
NUM|31|21|以利亚撒 祭司对打仗回来的士兵说：“耶和华所吩咐 摩西 律法中的条例是这样：
NUM|31|22|金、银、铜、铁、锡、铅，
NUM|31|23|凡能耐火的，你们要使它经过火，它就洁净，然而还要用除污秽的水来洁净它；凡不能耐火的，你们要使它经过水。
NUM|31|24|第七日，你们要洗衣服，才为洁净，然后可以进营。”
NUM|31|25|耶和华对 摩西 说：
NUM|31|26|“你和 以利亚撒 祭司，以及会众的各父系家长，要计算所掳掠的人和牲畜的总数。
NUM|31|27|要把所掳掠的分成两半：一半给那出去打仗的精兵，一半给全会众。
NUM|31|28|再从那出去打仗的战士所得的人、牛、驴、羊中，每五百取一，献给耶和华为贡物。
NUM|31|29|要从他们那一半中取出这些，交给 以利亚撒 祭司，作为耶和华的举祭。
NUM|31|30|又要从 以色列 人的那一半中，就是从人、牛、驴、羊，各样牲畜中，每五十取一，交给照管耶和华帐幕的 利未 人。”
NUM|31|31|于是 摩西 和 以利亚撒 祭司遵照耶和华所吩咐 摩西 的做了。
NUM|31|32|除了士兵所夺的财物以外，所掳来的有羊六十七万五千只，
NUM|31|33|牛七万二千头，
NUM|31|34|驴六万一千匹；
NUM|31|35|至于人，就是未曾与男人同房共寝的女子，总共三万二千名。
NUM|31|36|出去打仗之人的那分，就是他们所得的一半，共计羊三十三万七千五百只，
NUM|31|37|其中归耶和华为贡物的羊，六百七十五只；
NUM|31|38|牛三万六千头，其中归耶和华为贡物的七十二头；
NUM|31|39|驴三万零五百匹，其中归耶和华为贡物的六十一匹；
NUM|31|40|人一万六千名，其中归耶和华的三十二名。
NUM|31|41|摩西 把贡物，就是归给耶和华的举祭，交给 以利亚撒 祭司，是照耶和华所吩咐 摩西 的。
NUM|31|42|以色列 人所得的另一半，是 摩西 从打仗的人取来分给他们的。
NUM|31|43|会众的这一半有羊三十三万七千五百只，
NUM|31|44|牛三万六千头，
NUM|31|45|驴三万零五百匹，
NUM|31|46|人一万六千名。
NUM|31|47|无论是人或牲畜， 摩西 都每五十取一，交给照管耶和华帐幕的 利未 人，是照耶和华所吩咐 摩西 的。
NUM|31|48|带领众军队的军官，就是千夫长、百夫长，进到 摩西 那里，
NUM|31|49|对他说：“你的仆人已经计算属下战士的总数，一个也没有少。
NUM|31|50|如今我们把各人所得的金器，就是脚链子、手镯、打印的戒指、耳环、项链，都送给耶和华为供物，好在耶和华面前为我们赎罪。”
NUM|31|51|摩西 和 以利亚撒 祭司就收了他们的金子，就是各样的首饰。
NUM|31|52|千夫长、百夫长所献给耶和华为举祭的金子共有一万六千七百五十舍客勒。
NUM|31|53|打仗的人都把自己所掠夺的各自留下。
NUM|31|54|摩西 和 以利亚撒 祭司收了千夫长、百夫长的金子，就带进会幕，好使 以色列 人在耶和华面前蒙记念。
NUM|32|1|吕便 子孙和 迦得 子孙的牲畜极其众多。他们看到 雅谢 地和 基列 地；看哪，这是可牧放牲畜的地方。
NUM|32|2|吕便 子孙和 迦得 子孙就到 摩西 和 以利亚撒 祭司，以及会众的领袖那里，说：
NUM|32|3|“ 亚他录 、 底本 、 雅谢 、 宁拉 、 希实本 、 以利亚利 、 示班 、 尼波 、 比稳 ，
NUM|32|4|就是耶和华在 以色列 会众面前所攻取之地，是可牧放牲畜之地，而你的仆人也有牲畜。”
NUM|32|5|又说：“我们若在你眼前蒙恩，求你把这地给我们为业；不要领我们过 约旦河 。”
NUM|32|6|摩西 对 迦得 子孙和 吕便 子孙说：“难道你们的弟兄去打仗，你们却留在这里吗？
NUM|32|7|你们为什么使 以色列 人灰心，不渡过去，进入耶和华所赐给他们的那地呢？
NUM|32|8|我从 加低斯．巴尼亚 派你们的父执之辈去窥探那地时，他们就曾这样做过。
NUM|32|9|他们上到 以实各谷 ，窥探了那地之后，竟然使 以色列 人灰心，不愿进入耶和华所赐给他们的地。
NUM|32|10|当日，耶和华的怒气发作，起誓说：
NUM|32|11|‘凡从 埃及 上来二十岁以上的人，断不得看见我对 亚伯拉罕 、 以撒 、 雅各 起誓应许之地，因为他们没有专心跟从我；
NUM|32|12|惟有 基尼洗 族 耶孚尼 的儿子 迦勒 ，还有 嫩 的儿子 约书亚 可以看见，因为他们专心跟从耶和华。’
NUM|32|13|耶和华的怒气向 以色列 发作，使他们在旷野飘流四十年，直到在耶和华眼前作恶的那一代都消灭了。
NUM|32|14|看哪，你们这一伙罪人，竟然接续你们父执之辈，再增加耶和华对 以色列 所发的怒气。
NUM|32|15|你们若转离不跟从他，他要再把 以色列 人撇在旷野；这样，你们就使这众百姓灭亡了。”
NUM|32|16|他们挨近 摩西 ，说：“我们要在这里为牲畜筑圈，为孩童建城。
NUM|32|17|我们自己却要带兵器，急速行在 以色列 人的前面，领他们直到他们的地方。我们的孩童可以留在坚固的城内，躲避当地的居民。
NUM|32|18|我们必不回自己的家，直等到 以色列 人各自承受了自己的产业。
NUM|32|19|我们不和他们在 约旦河 那边分产业，因为我们的产业是在 约旦河 的东边。”
NUM|32|20|摩西 对他们说：“你们若要这么做，若要在耶和华面前带着兵器出去打仗，
NUM|32|21|你们中间所有带兵器的人都要在耶和华面前过 约旦河 ，直到耶和华把仇敌从他面前赶出去。
NUM|32|22|那地在耶和华面前被征服以后，你们方可回来。这样，你们向耶和华和 以色列 才算为无罪，这地也必在耶和华面前归你们为业。
NUM|32|23|倘若你们不这样做，看哪，你们就得罪了耶和华，当知道你们的罪必找上你们。
NUM|32|24|如今你们可以为孩童建城，为羊群筑圈，但你们口所讲出来的话，必须实践。”
NUM|32|25|迦得 子孙和 吕便 子孙对 摩西 说：“你的仆人们必照我主所吩咐的去做。
NUM|32|26|我们的孩子、妻子、牛羊和所有的牲畜都要留在 基列 的各城。
NUM|32|27|但你的仆人，凡能带兵器上战场的，都要照我主所说的话，在耶和华面前渡过去打仗。”
NUM|32|28|于是， 摩西 为他们吩咐 以利亚撒 祭司和 嫩 的儿子 约书亚 ，以及 以色列 人各支派父系的领袖。
NUM|32|29|摩西 对他们说：“ 迦得 子孙和 吕便 子孙，凡带兵器在耶和华面前去打仗的，若与你们一同渡过 约旦河 ，那地被你们征服以后，你们就要把 基列 地给他们为业。
NUM|32|30|倘若他们不带兵器与你们一同渡过去，他们就要在 迦南 地你们中间得产业。”
NUM|32|31|迦得 子孙和 吕便 子孙回答说：“耶和华怎样吩咐仆人，我们就必照样做。
NUM|32|32|我们自己必带着兵器，在耶和华面前渡过去，进入 迦南 地，好使我们在 约旦河 这边得到我们的产业。”
NUM|32|33|摩西 把 亚摩利 王 西宏 的国和 巴珊 王 噩 的国，就是他们的国土和周围的城镇，都给了 迦得 子孙和 吕便 子孙，以及 约瑟 的儿子 玛拿西 半个支派。
NUM|32|34|迦得 子孙建造了 底本 、 亚他录 、 亚罗珥 、
NUM|32|35|亚他录．朔反 、 雅谢 、 约比哈 、
NUM|32|36|伯．宁拉 、 伯．哈兰 ，都是坚固城，并筑有羊圈。
NUM|32|37|吕便 子孙建造了 希实本 、 以利亚利 、 基列亭 、
NUM|32|38|尼波 、 巴力．免 （名字是改了的）、 西比玛 ；他们给建造的城另起别名。
NUM|32|39|玛拿西 的儿子 玛吉 的子孙往 基列 去，占了那地，赶出那里的 亚摩利 人。
NUM|32|40|摩西 把 基列 赐给 玛拿西 的儿子 玛吉 ，他就住在那里。
NUM|32|41|玛拿西 的子孙 睚珥 占了 基列 的城镇，就称这些城镇为 哈倭特．睚珥 。
NUM|32|42|挪巴 占了 基纳 和 基纳 的乡镇，就照自己的名字称 基纳 为 挪巴 。
NUM|33|1|这是 以色列 人按着队伍，在 摩西 、 亚伦 的手下，出 埃及 地的行程。
NUM|33|2|摩西 遵照耶和华的指示记录他们每段行程的起点，这些行程的起点如下：
NUM|33|3|第一个月，就是正月十五日，逾越的第二天，他们从 兰塞 起行，在所有 埃及 人的眼前抬起头 来出去了。
NUM|33|4|那时， 埃及 人正埋葬他们的长子，就是耶和华在他们中间所击杀的；耶和华也惩治了他们的众神明。
NUM|33|5|以色列 人从 兰塞 起行，安营在 疏割 。
NUM|33|6|从 疏割 起行，安营在旷野边上的 以倘 。
NUM|33|7|从 以倘 起行，转向 巴力．洗分 对面的 比．哈希录 ，安营在 密夺 。
NUM|33|8|从 比．哈希录 起行，经过海，进入旷野，在 以倘 的旷野走了三天的路程，就安营在 玛拉 。
NUM|33|9|从 玛拉 起行，来到 以琳 ， 以琳 有十二股水泉，七十棵棕树，就安营在那里。
NUM|33|10|从 以琳 起行，安营在 红海 边。
NUM|33|11|从 红海 边起行，安营在 汛 的旷野。
NUM|33|12|从 汛 的旷野起行，安营在 脱加 。
NUM|33|13|从 脱加 起行，安营在 亚录 。
NUM|33|14|从 亚录 起行，安营在 利非订 ；在那里，百姓没有水喝。
NUM|33|15|从 利非订 起行，安营在 西奈 的旷野。
NUM|33|16|从 西奈 的旷野起行，安营在 基博罗．哈他瓦 。
NUM|33|17|从 基博罗．哈他瓦 起行，安营在 哈洗录 。
NUM|33|18|从 哈洗录 起行，安营在 利提玛 。
NUM|33|19|从 利提玛 起行，安营在 临门．帕烈 。
NUM|33|20|从 临门．帕烈 起行，安营在 立拿 。
NUM|33|21|从 立拿 起行，安营在 勒撒 。
NUM|33|22|从 勒撒 起行，安营在 基希拉他 。
NUM|33|23|从 基希拉他 起行，安营在 沙斐山 。
NUM|33|24|从 沙斐山 起行，安营在 哈拉大 。
NUM|33|25|从 哈拉大 起行，安营在 玛吉希录 。
NUM|33|26|从 玛吉希录 起行，安营在 他哈 。
NUM|33|27|从 他哈 起行，安营在 他拉 。
NUM|33|28|从 他拉 起行，安营在 密加 。
NUM|33|29|从 密加 起行，安营在 哈摩拿 。
NUM|33|30|从 哈摩拿 起行，安营在 摩西录 。
NUM|33|31|从 摩西录 起行，安营在 比尼．亚干 。
NUM|33|32|从 比尼．亚干 起行，安营在 曷．哈及甲 。
NUM|33|33|从 曷．哈及甲 起行，安营在 约巴他 。
NUM|33|34|从 约巴他 起行，安营在 阿博拿 。
NUM|33|35|从 阿博拿 起行，安营在 以旬．迦别 。
NUM|33|36|从 以旬．迦别 起行，安营在 寻 的旷野，就是 加低斯 。
NUM|33|37|从 加低斯 起行，安营在 以东 地边界的 何珥山 。
NUM|33|38|以色列 人出 埃及 地后四十年，五月初一， 亚伦 祭司遵照耶和华的指示，上 何珥山 ，死在那里。
NUM|33|39|亚伦 死在 何珥山 的时候一百二十三岁。
NUM|33|40|住在 迦南 地 尼革夫 的 迦南 人 亚拉得 王听说 以色列 人来了。
NUM|33|41|以色列 人从 何珥山 起行，安营在 撒摩拿 。
NUM|33|42|从 撒摩拿 起行，安营在 普嫩 。
NUM|33|43|从 普嫩 起行，安营在 阿伯 。
NUM|33|44|从 阿伯 起行，安营在 摩押 境内的 以耶．亚巴琳 。
NUM|33|45|从 以耶．亚巴琳 起行，安营在 底本．迦得 。
NUM|33|46|从 底本．迦得 起行，安营在 亚门．低比拉太音 。
NUM|33|47|从 亚门．低比拉太音 起行，安营在 尼波 前面的 亚巴琳山脉 。
NUM|33|48|从 亚巴琳山脉 起行，安营在 约旦河 边， 耶利哥 对面的 摩押 平原。
NUM|33|49|他们在 摩押 平原，沿着 约旦河 安营，从 伯．耶施末 直到 亚伯．什亭 。
NUM|33|50|耶和华在 约旦河 边， 耶利哥 对面的 摩押 平原吩咐 摩西 说：
NUM|33|51|“你要吩咐 以色列 人说：你们过 约旦河 进 迦南 地的时候，
NUM|33|52|要从你们面前赶出那地所有的居民，摧毁他们一切的石像和铸成的偶像，也要拆毁他们一切的丘坛。
NUM|33|53|你们要占领那地，住在那里，因我已把那地赐给你们为业。
NUM|33|54|你们要按照宗族抽签，承受土地：人多的要多给他们产业；人少的要少给他们产业。抽到何地给何人，那地就属于他。你们要按照父系的支派承受产业。
NUM|33|55|倘若你们不把那地的居民从你们面前赶出去，那留下的居民就必成为你们眼中的刺，肋下的荆棘，也必在你们所住的地上扰乱你们；
NUM|33|56|我想要怎样待他们，也必照样待你们。”
NUM|34|1|耶和华吩咐 摩西 说：
NUM|34|2|“你要吩咐 以色列 人，对他们说：你们到了 迦南 地，这就是归你们为业的地， 迦南 地和它四周的边界：
NUM|34|3|你们的南边是从 寻 的旷野起，沿着 以东 的边界；南边的地界从 盐海 东边开始，
NUM|34|4|绕过 亚克拉滨 斜坡的南边，经过 寻 ，直通到 加低斯．巴尼亚 的南边，又通到 哈萨．亚达 ，经过 押们 ，
NUM|34|5|从 押们 转向 埃及 溪谷，直通到海。
NUM|34|6|“你们西边的地界要以 大海 为边界；这就是你们西边的地界。
NUM|34|7|“你们北边的地界要从 大海 开始划界，直到 何珥山 ，
NUM|34|8|从 何珥山 划到 哈马口 ，直通到 西达达 ，
NUM|34|9|又通到 西斐仑 ，直达 哈萨．以难 。这就是你们北边的地界。
NUM|34|10|“东边的地界，你们要从 哈萨．以难 开始划界，直到 示番 ，
NUM|34|11|这地界要从 示番 下到 亚延 东边的 利比拉 ，这地界要下延到 基尼烈海 的东边，
NUM|34|12|这地界又下到 约旦河 ，直通到 盐海 。这就是你们的地和它四围的边界。”
NUM|34|13|摩西 吩咐 以色列 人说：“这就是耶和华吩咐抽签给九个半支派承受为业的地。
NUM|34|14|因为 吕便 子孙的支派按着父家、 迦得 子孙的支派按着父家，和 玛拿西 半个支派已经得到了他们的产业：
NUM|34|15|这两个半支派已经在 耶利哥 对面， 约旦河 东边，向日出的方向承受了产业。”
NUM|34|16|耶和华吩咐 摩西 说：
NUM|34|17|“这是为你们分地为业的人的名字： 以利亚撒 祭司和 嫩 的儿子 约书亚 。
NUM|34|18|你要从每个支派中选一个领袖来分配产业。
NUM|34|19|这些人的名字如下： 犹大 支派， 耶孚尼 的儿子 迦勒 。
NUM|34|20|西缅 子孙的支派， 亚米忽 的儿子 示母利 。
NUM|34|21|便雅悯 支派， 基斯伦 的儿子 以利达 。
NUM|34|22|但 子孙支派的领袖， 约利 的儿子 布基 。
NUM|34|23|约瑟 的子孙， 玛拿西 子孙支派的领袖： 以弗 的儿子 汉尼业 。
NUM|34|24|以法莲 子孙支派的领袖： 拾弗但 的儿子 基摩利 。
NUM|34|25|西布伦 子孙支派的领袖： 帕纳 的儿子 以利撒番 。
NUM|34|26|以萨迦 子孙支派的领袖： 阿散 的儿子 帕铁 。
NUM|34|27|亚设 子孙支派的领袖： 示罗米 的儿子 亚希忽 。
NUM|34|28|拿弗他利 子孙支派的领袖： 亚米忽 的儿子 比大黑 。”
NUM|34|29|这些就是耶和华所吩咐，在 迦南 地为 以色列 人分产业的人。
NUM|35|1|耶和华在 约旦河 边， 耶利哥 对面的 摩押 平原吩咐 摩西 说：
NUM|35|2|“你吩咐 以色列 人，要从所得为业的地中把一些城给 利未 人居住，也要把这些城四围的郊野给 利未 人。
NUM|35|3|这些城镇要归他们居住，郊外可以给他们牧放牛羊、牲畜和所有的动物。
NUM|35|4|你们给 利未 人城的郊外，要从城墙量起，四围往外量一千肘。
NUM|35|5|你们要往东量二千肘，往南量二千肘，往西量二千肘，往北量二千肘为边界，以城为中心；这城镇的郊外要归给他们。”
NUM|35|6|“你们给 利未 人的城镇中，要设立六座逃城，让误杀人的可以逃到那里。此外还要给他们四十二座城。
NUM|35|7|所以，给 利未 人的城一共有四十八座，连同城的郊外都给他们。
NUM|35|8|从 以色列 人所得的产业中给 利未 人的这些城镇，多的要多给，少的要少给；各支派要按照所承受为业之地的多少把城镇给 利未 人。”
NUM|35|9|耶和华吩咐 摩西 说：
NUM|35|10|“你要吩咐 以色列 人，对他们说：你们过了 约旦河 ，进入 迦南 地，
NUM|35|11|要指定几座城，作为你们的逃城，使误杀人的可以逃到那里。
NUM|35|12|这些城要作为逃避报仇者的城，使误杀人的不至于死，等他站在会众面前受审判。
NUM|35|13|“你们指定的城，是要作你们的六座逃城。
NUM|35|14|约旦河 东指定三座， 迦南 地也指定三座，作为逃城。
NUM|35|15|这六座城要给 以色列 人和他们中间的外人，以及寄居者，作为逃城，让误杀人的可以逃到那里。
NUM|35|16|“倘若人用铁器打死人，他是故意杀人的；故意杀人的必被处死。
NUM|35|17|若用手中可以致命的石头打死人，他是故意杀人的；故意杀人的必被处死。
NUM|35|18|若用手中可以致命的木器打死人，他是故意杀人的；故意杀人的必被处死。
NUM|35|19|报血仇者可以亲自杀死那故意杀人的；他一找到凶手，就可以杀死他。
NUM|35|20|人若因怨恨把人推倒，或埋伏等着丢东西砸人，以至于死，
NUM|35|21|或因仇恨用手打死人，打人的必被处死，他是故意杀人的；报血仇者一遇见凶手就可以杀死他。
NUM|35|22|“人若不是出于仇恨，把人推倒，或不是埋伏等着丢东西砸人，
NUM|35|23|或是在不注意的时候，用可以致命的石头扔在人身上，以至于死，彼此没有仇恨，也无意害对方，
NUM|35|24|会众就要照着这些典章，在杀人者和报血仇者中间审判。
NUM|35|25|会众要救这误杀人的脱离报血仇者的手，送他回到他曾逃入的逃城那里。他要住在城中，直到受圣膏的大祭司去世。
NUM|35|26|但误杀人的，无论什么时候，若离开了他所逃入的逃城边界，
NUM|35|27|报血仇者在逃城边界外遇见他，把凶手杀了，报血仇者就没有流人血之罪。
NUM|35|28|因为误杀人的应该住在逃城里，直到大祭司去世。大祭司去世以后，误杀人的才可以回到他所得为业之地。
NUM|35|29|在你们一切的住处，这些都要作为你们世世代代的律例典章。
NUM|35|30|“无论谁杀了人，必须凭几个证人的口，才可把那故意杀人的处死；只凭一个证人，不足以判人死。
NUM|35|31|那犯死罪的杀人犯，你们不可收赎价来代替他的命；他必须被处死。
NUM|35|32|那逃到逃城的人，你们不可向他收赎价，使他在大祭司未死以先回本地居住。
NUM|35|33|这样，你们就不会污秽所住之地，因为血能使地污秽；若有血流在地上，除非流那杀人者的血，否则那地就不得洁净。
NUM|35|34|你们不可玷污所住之地，就是我住在当中的地，因为我－耶和华住在 以色列 人中间。”
NUM|36|1|约瑟 子孙的宗族， 玛拿西 的孙子， 玛吉 的儿子 基列 ，他父系宗族的领袖来到 摩西 和作领袖的 以色列 众父系家长面前，说：
NUM|36|2|“耶和华曾吩咐我主抽签分地给 以色列 人为业，我主也遵照耶和华的吩咐，把我们兄弟 西罗非哈 的产业给他的女儿。
NUM|36|3|她们若嫁给 以色列 别个支派的人，必拿走我们祖宗所遗留的产业，加在她们丈夫支派的产业上。这样，我们抽签所得的产业就要减少了。
NUM|36|4|到了 以色列 人的禧年，她们的产业就必加在她们丈夫支派的产业上。这样，我们祖宗支派的产业就要减少了。”
NUM|36|5|摩西 照耶和华的指示吩咐 以色列 人说：“ 约瑟 子孙支派的人说得有理。
NUM|36|6|关于 西罗非哈 的女儿们，这是耶和华吩咐的话说：‘她们可以随意嫁人，只是必须嫁给同宗，她们父亲支派的人。
NUM|36|7|这样， 以色列 人的产业就不会从这支派转到另一个支派，因为 以色列 人要各自守住祖宗支派的产业。
NUM|36|8|凡在 以色列 支派中得了产业的女儿，必须嫁给同宗，她们父亲支派的人，好使 以色列 人各自承受他们祖宗的产业。
NUM|36|9|产业不可从一个支派转到另一个支派，因为 以色列 支派的人要各自守住自己的产业。’”
NUM|36|10|耶和华怎样吩咐 摩西 ， 西罗非哈 的女儿就照样做。
NUM|36|11|西罗非哈 的女儿 玛拉 、 得撒 、 曷拉 、 密迦 、 挪阿 都嫁给她们叔伯的儿子。
NUM|36|12|她们嫁给了 约瑟 儿子 玛拿西 子孙宗族的人；她们的产业保留在同宗，她们父亲的支派中。
NUM|36|13|这是耶和华在 约旦河 边， 耶利哥 对面的 摩押 平原，藉着 摩西 吩咐 以色列 人的命令和典章。
DEUT|1|1|以下是 摩西 在 约旦河 东的旷野， 疏弗 对面的 亚拉巴 ，就是在 巴兰 、 陀弗 、 拉班 、 哈洗录 、 底撒哈 之间，向 以色列 众人所说的话。
DEUT|1|2|从 何烈山 经过 西珥山 到 加低斯．巴尼亚 要十一天的路程。
DEUT|1|3|第四十年十一月初一， 摩西 照耶和华所吩咐他一切有关 以色列 人的话，都告诉他们。
DEUT|1|4|那时，他已经击败了住 希实本 的 亚摩利 王 西宏 和住 亚斯她录 、 以得来 的 巴珊 王 噩 。
DEUT|1|5|摩西 在 约旦河 东的 摩押 地讲解这律法，说：
DEUT|1|6|“耶和华－我们的上帝在 何烈山 吩咐我们说：你们住在这山上已经够久了。
DEUT|1|7|要起行，转到 亚摩利 人的山区和附近的地区，就是 亚拉巴 、山区、 谢非拉 、 尼革夫 、沿海一带， 迦南 人的地和 黎巴嫩 ，直到 大河 ，就是 幼发拉底河 。
DEUT|1|8|看，我将这地摆在你们面前。你们要进去得这地，就是耶和华向你们列祖 亚伯拉罕 、 以撒 、 雅各 起誓要赐给他们和他们后裔为业之地。”
DEUT|1|9|“那时，我对你们说：‘我独自一人无法承担你们的事。
DEUT|1|10|耶和华－你们的上帝使你们增多。看哪，你们今日好像天上的星那样多。
DEUT|1|11|惟愿耶和华－你们列祖的上帝使你们更增加千倍，照他所应许你们的赐福给你们。
DEUT|1|12|但你们的担子，你们的重任，以及你们的争讼，我独自一人怎能承担呢？
DEUT|1|13|你们要按着各支派选出有智慧、明辨是非、为人所知的人来，我就立他们为你们的领袖。’
DEUT|1|14|你们回答我说：‘你说要做的事很好！’
DEUT|1|15|我就将你们各支派的领袖，就是有智慧、为人所知的人，立他们为领袖，作你们各支派的千夫长、百夫长、五十夫长、十夫长等官长，来管理你们。
DEUT|1|16|“当时，我吩咐你们的审判官说：‘你们听讼，无论是弟兄之间的诉讼，或与寄居者之间的诉讼，都要秉公判断。
DEUT|1|17|审判的时候不可看人的情面；无论大小，你们都要听讼。不可因人而惧怕，因为审判是上帝的事。你们当中若有难断的案件，可以呈到我这里，让我来听讼。’
DEUT|1|18|那时，我已经把你们所当做的事都吩咐你们了。”
DEUT|1|19|“我们照着耶和华－我们上帝所吩咐的，从 何烈山 起行，经过你们所看见那一切大而可怕的旷野，往 亚摩利 人的山区去，到了 加低斯．巴尼亚 。
DEUT|1|20|我对你们说：‘你们已经到了耶和华－我们上帝所赐给我们的 亚摩利 人之山区。
DEUT|1|21|看，耶和华－你的上帝已将那地摆在你面前，你要照耶和华－你列祖的上帝所说的，上去得那地为业。不要惧怕，也不要惊惶。’
DEUT|1|22|你们都来到我这里，说：‘让我们先派人去，为我们窥探那地，把我们上去该走的路线和该进的城镇回报我们。’
DEUT|1|23|这话我看为美，就从你们中间选取十二个人，每支派一人。
DEUT|1|24|于是他们起身上山区去，到 以实各谷 ，窥探那地。
DEUT|1|25|他们的手带着那地的一些果子，下到我们这里，回报我们说：‘耶和华－我们的上帝所赐给我们的是美地。’
DEUT|1|26|“你们却不肯上去，竟违背了耶和华─你们上帝的指示，
DEUT|1|27|在帐棚内发怨言说：‘耶和华因为恨我们，所以将我们从 埃及 地领出来，要把我们交在 亚摩利 人的手中，除灭我们。
DEUT|1|28|我们上哪里去呢？我们的弟兄使我们胆战心惊 ，说那里的百姓比我们又大又高 ，那里的城镇又大，城墙又坚固，如天一样高，并且我们在那里看见 亚衲 族人。’
DEUT|1|29|我就对你们说：‘不要惊惶，也不要怕他们。
DEUT|1|30|在你们前面行的耶和华－你们的上帝必为你们争战，正如他在 埃及 ，在你们眼前为你们所做的一样；
DEUT|1|31|并且你们在旷野所行的一切路上，也看见了耶和华─你们的上帝背着你们，如同人背自己的儿子一样，直到你们来到这地方。’
DEUT|1|32|你们在这事上却不信耶和华─你们的上帝。
DEUT|1|33|他一路行在你们前面，为你们寻找安营的地方；他夜间在火中，日间在云中，指示你们当走的路。”
DEUT|1|34|“耶和华听见你们的怨言，就发怒，起誓说：
DEUT|1|35|‘这邪恶世代的人，一个也不得看见我起誓要赐给你们列祖的美地；
DEUT|1|36|惟有 耶孚尼 的儿子 迦勒 必得看见，并且我要将他所踏过的地赐给他和他的子孙，因为他专心跟从我。’
DEUT|1|37|耶和华也因你们的缘故向我发怒，说：‘你也不得进入那地。
DEUT|1|38|那侍候你， 嫩 的儿子 约书亚 必得进入那地。你要勉励他，因为他要使 以色列 承受那地为业。
DEUT|1|39|你们的孩子，你们说要成为掳物的，就是今日尚不知善恶的儿女，必进入那地。我要将那地赐给他们，他们必得为业。
DEUT|1|40|至于你们，要转回，从 红海 的路往旷野去。’
DEUT|1|41|“你们回答我说：‘我们得罪了耶和华！现在我们愿遵照耶和华─我们上帝一切所吩咐的上去争战。’于是你们各人带着兵器，以为很容易就能上到山区去。
DEUT|1|42|耶和华对我说：‘你对他们说：不要上去，也不要争战，因我不在你们中间，恐怕你们在仇敌面前被击败。’
DEUT|1|43|我就告诉了你们，你们却不听从，竟违背耶和华的指示，擅自上到山区去。
DEUT|1|44|住在那山区的 亚摩利 人像蜂群一样出来迎击你们，追赶你们，在 西珥 击败你们，直到 何珥玛 。
DEUT|1|45|你们就回来，在耶和华面前哭泣；耶和华却不听你们的声音，也不向你们侧耳。
DEUT|1|46|你们照着所停留的日子，在 加低斯 停留了许多日子。”
DEUT|2|1|“我们转回，从 红海 的路往旷野去，正如耶和华所吩咐我的。我们在 西珥山 绕行了许多日子。
DEUT|2|2|耶和华对我说：
DEUT|2|3|‘你们绕行这山已经够久了，要转向北方。
DEUT|2|4|你要吩咐百姓说：你们弟兄 以扫 的子孙住在 西珥 ，你们要经过他们的边界。他们必惧怕你们，但你们要分外谨慎。
DEUT|2|5|不可向他们挑战；他们的地，连脚掌可踏之处，我都不给你们，因我已将 西珥山 赐给 以扫 为业。
DEUT|2|6|你们要用钱向他们买粮吃，也要用钱向他们买水喝。
DEUT|2|7|因为耶和华─你的上帝在你手里所做的一切事上已赐福给你。你走这大旷野，他都知道。这四十年，耶和华─你的上帝与你同在，因此你一无所缺。’
DEUT|2|8|“于是，我们经过我们弟兄 以扫 子孙所住的 西珥 ，从 亚拉巴 的路，经过 以拉他 、 以旬．迦别 ，转向 摩押 旷野的路去。
DEUT|2|9|耶和华对我说：‘不可侵犯 摩押 ，也不可向他们挑战。他们的地，我不赐给你为业，因我已将 亚珥 赐给 罗得 的子孙为业。’
DEUT|2|10|先前， 以米 人住在那里，百姓又大又多，像 亚衲 人一样高大。
DEUT|2|11|他们跟 亚衲 人一样，也算是 利乏音 人，但 摩押 人却称他们为 以米 人。
DEUT|2|12|从前， 何利 人也住在 西珥 ，但 以扫 的子孙把他们除灭，占领了他们的地，接续他们在那里居住，如同 以色列 在耶和华赐给他们为业之地所做的一样。
DEUT|2|13|‘现在，起来，过 撒烈溪 ！’于是我们过了 撒烈溪 。
DEUT|2|14|从离开 加低斯．巴尼亚 到渡过 撒烈溪 ，这段时期共三十八年，直到这一代的战士都从营中灭尽，正如耶和华向他们所起的誓。
DEUT|2|15|耶和华的手也攻击他们，将他们从营中除灭，直到灭尽。
DEUT|2|16|“百姓中所有的战士灭尽死亡以后，
DEUT|2|17|耶和华吩咐我说：
DEUT|2|18|‘你今日要经过 摩押 的边界 亚珥 ，
DEUT|2|19|走到 亚扪 人之地。不可侵犯他们，也不可向他们挑战。 亚扪 人的地，我不赐给你们为业，因我已将那地赐给 罗得 的子孙为业。’
DEUT|2|20|那地也算是 利乏音 人之地，因为先前 利乏音 人住在那里， 亚扪 人称他们为 散送冥 人。
DEUT|2|21|那里的百姓又大又多，像 亚衲 人一样高大，但耶和华从 亚扪 人面前除灭他们， 亚扪 人就占领他们的地，接续他们在那里居住。
DEUT|2|22|这正如耶和华从前为住在 西珥 的 以扫 子孙，将 何利 人从他们面前除灭，使他们得了 何利 人的地，接续他们在那里居住，直到今日一样。
DEUT|2|23|亚卫 人先前住在乡村直到 迦萨 ；从 迦斐托 出来的 迦斐托 人将 亚卫 人除灭，接续他们在那里居住。
DEUT|2|24|你们起来往前去，过 亚嫩谷 。看哪，我已将 亚摩利 人 希实本 王 西宏 和他的地交在你手中，你要开始去得他的地为业，向他挑战。
DEUT|2|25|从今日起，我要让天下万民因你惊慌惧怕，听见你的名声，就因你发颤伤恸。”
DEUT|2|26|“我从 基底莫 的旷野派遣使者到 希实本 王 西宏 那里，用和平的话说：
DEUT|2|27|‘求你让我穿越你的地，我走路的时候，只走大路，不偏左右。
DEUT|2|28|你可以卖粮给我吃，卖水给我喝；只要让我步行过去，
DEUT|2|29|就如住在 西珥 的 以扫 子孙和住在 亚珥 的 摩押 人待我一样，等我过了 约旦河 ，进入耶和华－我们上帝所赐给我们的地。’
DEUT|2|30|但 希实本 王 西宏 不肯让我们从他那里经过，因为耶和华－你的上帝使他性情顽梗，内心刚硬，为要把他交在你手中，像今日一样。
DEUT|2|31|耶和华对我说：‘看，我已开始把 西宏 和他的地交给你了，你要开始得他的地为业。’
DEUT|2|32|“ 西宏 和他的众百姓出来迎击我们，在 雅杂 与我们交战。
DEUT|2|33|耶和华－我们的上帝把他交给我们，我们就杀了他和他的众儿子，以及他所有的百姓。
DEUT|2|34|那时，我们夺了他一切的城镇，毁灭各城的男人、女人、孩子，没有留下一个幸存者。
DEUT|2|35|只有牲畜和所夺各城的财物，我们都取为自己的掠物。
DEUT|2|36|从 亚嫩谷 旁的 亚罗珥 和谷中的城，直到 基列 ，没有一座城是高得我们不能攻取的；耶和华－我们的上帝把它们全都交给我们了。
DEUT|2|37|只有 亚扪 人之地， 雅博河 沿岸，以及山区的城镇，你没有挨近，这全是耶和华－我们上帝所吩咐的。”
DEUT|3|1|“我们又转回，朝 巴珊 的路上去。 巴珊 王 噩 和他的众百姓出来迎击我们，在 以得来 与我们交战。
DEUT|3|2|耶和华对我说：‘不要怕他！因我已把他和他的众百姓，以及他的地，都交在你手中；你要待他像从前待住在 希实本 的 亚摩利 王 西宏 一样。’
DEUT|3|3|于是耶和华－我们的上帝也把 巴珊 王 噩 和他的众百姓都交在我们手中；我们杀了他，没有给他留下一个幸存者。
DEUT|3|4|那时，我们夺了他一切的城镇，共六十座，没有一座城不被我们所夺，这是 亚珥歌伯 的全境， 巴珊 王 噩 的国度。
DEUT|3|5|这些坚固的城都有高的城墙，有门有闩，此外，还有许多无城墙的乡村。
DEUT|3|6|我们把这些都毁灭了，像从前待 希实本 王 西宏 一样，毁灭各城的男人、女人、孩子；
DEUT|3|7|只有一切牲畜和城中的财物，我们取为自己的掠物。
DEUT|3|8|那时，我们从两个 亚摩利 王的手里把 约旦河 东边的地夺过来，从 亚嫩谷 直到 黑门山 ，
DEUT|3|9|这 黑门山 ， 西顿 人称为 西连 ， 亚摩利 人称为 示尼珥 。
DEUT|3|10|我们夺了平原的各城、 基列 全地、 巴珊 全地，直到 撒迦 和 以得来 ，都是 巴珊 王 噩 国内的城镇。
DEUT|3|11|利乏音 人所剩下的只有 巴珊 王 噩 。看哪，他的床是铁床，按照人肘的度量，长九肘，宽四肘，现今不是在 亚扪 人的 拉巴 吗？”
DEUT|3|12|“那时，我们得了这地。从 亚嫩谷 旁的 亚罗珥 起，连同 基列 山区的一半和境内的城镇，我都给了 吕便 人和 迦得 人。
DEUT|3|13|基列 其余的地和 巴珊 全地，就是 噩 的国度，我给了 玛拿西 半支派。 亚珥歌伯 全境就是 巴珊 全地，也称为 利乏音 人之地。
DEUT|3|14|玛拿西 的子孙 睚珥 占领了 亚珥歌伯 全境，直到 基述 人和 玛迦 人的边界，就按自己的名字称这些地，就是 巴珊 ，为 哈倭特．睚珥 ，直到今日。
DEUT|3|15|我又将 基列 给了 玛吉 。
DEUT|3|16|我给了 吕便 人和 迦得 人从 基列 到 亚嫩谷 ，以谷的中央为界，直到 亚扪 人边界的 雅博河 ；
DEUT|3|17|还有 亚拉巴 和靠近 约旦河 之地，从 基尼烈 直到 亚拉巴海 ，就是 盐海 ，以及 毗斯迦山 斜坡的山脚东边之地。
DEUT|3|18|“那时，我吩咐你们说：‘耶和华－你们的上帝已将这地赐给你们为业；你们所有的勇士都要带着兵器，在你们的弟兄 以色列 人前面过去。
DEUT|3|19|但你们的妻子、孩子、牲畜，可以住在我所赐给你们的各城里，我知道你们有许多牲畜。
DEUT|3|20|等到耶和华让你们的弟兄像你们一样，得享太平，他们在 约旦河 另一边，也得了耶和华－你们的上帝所赐给他们的地，你们各人才可以回到我所赐给你们为业之地。’
DEUT|3|21|那时，我吩咐 约书亚 说：‘你亲眼看见了耶和华－你们的上帝向这两个王一切所做的事，耶和华也必向你所要去的各国照样做。
DEUT|3|22|不要怕他们，因为那为你们争战的是耶和华－你们的上帝。’”
DEUT|3|23|“那时，我恳求耶和华说：
DEUT|3|24|‘主耶和华啊，你已开始将你的伟大和你大能的手显给你仆人看。在天上，在地下，有什么神明能像你行事，像你有大能的作为呢？
DEUT|3|25|求你让我过去，看 约旦河 另一边的美地，就是那佳美的山区和 黎巴嫩 。’
DEUT|3|26|但耶和华因你们的缘故向我发怒，不应允我。耶和华对我说：‘你够了吧！不要再向我提这事。
DEUT|3|27|你上 毗斯迦山 顶去，向东、西、南、北举目，用你的眼睛观看，因为你必不能过这 约旦河 。
DEUT|3|28|你却要吩咐 约书亚 ，勉励他，使他壮胆，因为他必在这百姓前面过去，使他们承受你所要观看之地。’
DEUT|3|29|于是我们停留在 伯．毗珥 对面的谷中。”
DEUT|4|1|“现在， 以色列 啊，听我所教导你们的律例典章，要遵行，好使你们存活，得以进入耶和华－你们列祖之上帝所赐给你们的地，承受为业。
DEUT|4|2|我吩咐你们的话，你们不可加添，也不可删减，好叫你们遵守耶和华－你们上帝的命令，就是我所吩咐你们的。
DEUT|4|3|你们已亲眼看见耶和华因 巴力．毗珥 所做的。凡随从 巴力．毗珥 的人，耶和华－你的上帝都从你中间除灭了。
DEUT|4|4|只有你们这紧紧跟随耶和华－你们上帝的人，今日全都存活。
DEUT|4|5|看，我照着耶和华－我的上帝所吩咐我的，将律例和典章教导你们，使你们在所要进去得为业的地上遵行。
DEUT|4|6|你们要谨守遵行；这就是你们在万民眼前的智慧和聪明。他们听见这一切律例，必说：‘这大国的人真是有智慧，有聪明！’
DEUT|4|7|哪一大国有神明与他们相近，像耶和华－我们的上帝在我们求告他的时候与我们相近呢？
DEUT|4|8|哪一大国有这样公义的律例典章，像我今日在你们面前所颁布的这一切律法呢？
DEUT|4|9|“但你要谨慎，殷勤保守你的心灵，免得忘记你亲眼所看见的事，又免得在你一生的年日这些事离开你的心，总要把它们传给你的子子孙孙。
DEUT|4|10|你在 何烈山 站在耶和华－你上帝面前的那日，耶和华对我说：‘你为我召集百姓，我要叫他们听见我的话，使他们活在世上的日子，可以学习敬畏我，又可以教导他们的儿女。’
DEUT|4|11|那时，你们近前来，站在山下；山上有火燃烧，直冲天顶，并有黑暗、密云、幽暗。
DEUT|4|12|耶和华从火焰中对你们说话，你们听见说话的声音，只有声音，却没有看见形像。
DEUT|4|13|他将所吩咐你们当守的约指示你们，就是十条诫命 ，并将诫命写在两块石版上。
DEUT|4|14|那时，耶和华吩咐我将律例典章教导你们，使你们在所要过去得为业的地上遵行。”
DEUT|4|15|“所以，你们为自己的缘故要分外谨慎；因为耶和华在 何烈山 ，从火中对你们说话的那日，你们没有看见任何形像。
DEUT|4|16|惟恐你们的行为败坏，为自己雕刻任何形状的偶像，无论是男像或女像，
DEUT|4|17|或地上任何走兽的像，或任何飞在空中有翅膀的鸟的像，
DEUT|4|18|或地上任何爬行动物的像，或地底下任何水中鱼的像。
DEUT|4|19|又恐怕你向天举目，看见耶和华－你的上帝为天下万民所摆列的日月星辰，就是天上的万象，就被诱惑去敬拜它们，事奉它们。
DEUT|4|20|耶和华将你们从 埃及 带领出来，脱离铁炉，是要你们成为他产业的子民，像今日一样。
DEUT|4|21|“耶和华又因你们的缘故向我发怒，起誓不容我过 约旦河 ，不让我进入耶和华－你上帝所赐你为业的那美地。
DEUT|4|22|我只好死在这地，不能过 约旦河 ；但你们必过去得那美地。
DEUT|4|23|你们要谨慎，免得忘记耶和华－你们的上帝与你们所立的约，为自己雕刻任何形状的偶像，就是耶和华－你上帝所禁止的，
DEUT|4|24|因为耶和华－你的上帝是吞灭的火，是忌邪 的上帝。
DEUT|4|25|“你们在那地住久了，生子生孙，若行为败坏，为自己雕刻任何形状的偶像，行耶和华－你上帝眼中看为恶的事，惹他发怒，
DEUT|4|26|我今日呼天唤地向你们作见证，你们在过 约旦河 得为业的地上必迅速灭亡！你们在那地的日子必不长久，必全然灭绝。
DEUT|4|27|耶和华必将你们分散在万民中；在耶和华领你们到的列国中，你们剩下的人丁稀少。
DEUT|4|28|在那里，你们必事奉人手所造的神明，它们是木头，是石头，不能看，不能听，不能吃，不能闻。
DEUT|4|29|你们在那里必寻求耶和华－你的上帝。你若尽心尽性寻求他，就必寻见。
DEUT|4|30|日后你在患难中，当这一切的事临到你，你必归回耶和华－你的上帝，听从他的话。
DEUT|4|31|耶和华－你的上帝是有怜悯的上帝，他不撇下你，不灭绝你，也不忘记他起誓与你列祖所立的约。
DEUT|4|32|“你去问，在你先前的时代，自从上帝造人在地上以来，从天这边到天那边，曾有过或听过这样的大事吗？
DEUT|4|33|有哪些百姓听见上帝在火中说话的声音，像你听见了还能存活呢？
DEUT|4|34|上帝何曾为自己尝试从别的国中领出一国的子民来，用考验、神迹、奇事、战争、大能的手、伸出来的膀臂和大可畏的事，像耶和华－你们的上帝在 埃及 ，在你们眼前为你们所做的一切事呢？
DEUT|4|35|这是要显给你看，使你知道，惟有耶和华他是上帝，除他以外，再没有别的了。
DEUT|4|36|他从天上使你听见他的声音，为要教导你，又在地上使你看见他的烈火，并且听见他从火中所说的话。
DEUT|4|37|因为他爱你的列祖，拣选他们的后裔 ，亲自用大能领你出了 埃及 ，
DEUT|4|38|要将比你强大的列国从你面前赶出，领你进去，把他们的地赐你为业，像今日一样。
DEUT|4|39|所以，今日你要知道，也要记在心里，天上地下惟有耶和华他是上帝，再没有别的了。
DEUT|4|40|我今日吩咐你的律例诫命，你要遵守，使你和你的后裔可以得福，并使你的日子一直在耶和华－你上帝赐你的地上得以长久。”
DEUT|4|41|“那时， 摩西 在 约旦河 东边，向日出的方向，指定三座城，
DEUT|4|42|使那素无仇恨、无意中杀了邻舍的凶手，可以逃到这三座城中的一座，就得存活：
DEUT|4|43|属 吕便 人的是旷野平坦之地的 比悉 ，属 迦得 人的是 基列 的 拉末 ，属 玛拿西 人的是 巴珊 的 哥兰 。”
DEUT|4|44|这是 摩西 在 以色列 人面前颁布的律法。
DEUT|4|45|这些法度、律例、典章是 摩西 在 以色列 人出 埃及 后对他们说的，
DEUT|4|46|在 约旦河 东 伯毗珥 对面的谷中，在住 希实本 的 亚摩利 王 西宏 之地；这 西宏 是 摩西 和 以色列 人出 埃及 后所击杀的。
DEUT|4|47|他们得了他的地，又得了 巴珊 王 噩 的地，就是两个 亚摩利 王，在 约旦河 东，向日出方向的地：
DEUT|4|48|从 亚嫩谷 旁的 亚罗珥 ，直到 西云山 ，就是 黑门山 ，
DEUT|4|49|还有 约旦河 东的整个 亚拉巴 ，向日出方向，直到 亚拉巴海 ，靠近 毗斯迦山 斜坡的山脚。
DEUT|5|1|摩西 召集 以色列 众人，对他们说：“ 以色列 啊，要听我今日在你们耳中所吩咐的律例典章，要学习，谨守遵行。
DEUT|5|2|耶和华－我们的上帝在 何烈山 与我们立约。
DEUT|5|3|这约耶和华不是与我们列祖立的，而是与我们，就是今日在这里还活着的人立的。
DEUT|5|4|耶和华在山上，从火中，面对面与你们说话。
DEUT|5|5|那时我站在耶和华和你们之间，要将耶和华的话传给你们，因为你们惧怕那火，没有上山。他说：
DEUT|5|6|“‘我是耶和华－你的上帝，曾将你从 埃及 地为奴之家领出来。
DEUT|5|7|“‘除了我以外，你不可有别的神。
DEUT|5|8|“‘不可为自己雕刻偶像，也不可做什么形像，仿佛上天、下地和地底下水中的百物。
DEUT|5|9|不可跪拜那些像，也不可事奉它们，因为我耶和华－你的上帝是忌邪 的上帝。恨我的，我必惩罚他们的罪，自父及子，直到三、四代；
DEUT|5|10|爱我、守我诫命的，我必向他们施慈爱，直到千代。
DEUT|5|11|“‘不可妄称耶和华－你上帝的名，因为妄称耶和华名的，耶和华必不以他为无罪。
DEUT|5|12|“‘当守安息日为圣日，正如耶和华－你上帝所吩咐的。
DEUT|5|13|六日要劳碌做你一切的工，
DEUT|5|14|但第七日是向耶和华－你的上帝当守的安息日。这一日，你和你的儿女、仆婢、牛、驴、牲畜，以及你城里寄居的客旅，都不可做任何的工，使你的仆婢可以和你一样休息。
DEUT|5|15|你要记念你在 埃及 地作过奴仆，耶和华－你的上帝用大能的手和伸出来的膀臂领你从那里出来。因此，耶和华－你的上帝吩咐你守安息日。
DEUT|5|16|“‘当孝敬父母，正如耶和华－你上帝所吩咐的，使你得福，并使你的日子在耶和华－你上帝所赐给你的地上得以长久。
DEUT|5|17|“‘不可杀人。
DEUT|5|18|“‘不可奸淫。
DEUT|5|19|“‘不可偷盗。
DEUT|5|20|“‘不可做假见证陷害你的邻舍。
DEUT|5|21|“‘不可贪恋你邻舍的妻子；也不可贪图你邻舍的房屋、田地、仆婢、牛驴，以及他一切所有的。’
DEUT|5|22|“这些话是耶和华在山上，从火焰、密云、幽暗中，大声吩咐你们全会众的，再没有加添别的话了。他把这些话写在两块石版上，交给我。
DEUT|5|23|山被火焰烧着，你们听见从黑暗中发出的声音，那时，你们各支派的领袖和长老都挨近我。
DEUT|5|24|你们说：‘看哪，耶和华－我们的上帝将他的荣耀和他的伟大显给我们看，我们也听见他从火中发出的声音。今日我们看到上帝与人说话，人还活着。
DEUT|5|25|现在这大火将要吞灭我们，我们何必死呢？若再听见耶和华我们上帝的声音，我们就必死。
DEUT|5|26|凡血肉之躯，有谁像我们一样，听见了永生上帝从火中讲话的声音还能活着呢？
DEUT|5|27|求你近前去，听耶和华－我们上帝所要说的一切话，将耶和华－我们上帝对你说的话都传给我们，我们就听从遵行。’
DEUT|5|28|“你们对我说的话，耶和华都听见了。耶和华对我说：‘这百姓对你说的话，我听见了；他们所说的都对。
DEUT|5|29|惟愿他们存这样的心敬畏我，常遵守我一切的诫命，使他们和他们的子孙永远得福。
DEUT|5|30|你去对他们说：你们回帐棚去吧！
DEUT|5|31|至于你，可以站在我这里，我要将一切诫命、律例、典章传给你。你要教导他们，使他们在我赐他们为业的地上遵行。’
DEUT|5|32|所以，你们要照耶和华－你们上帝所吩咐的谨守遵行，不可偏离左右。
DEUT|5|33|你们要走耶和华－你们的上帝所吩咐的一切道路，使你们可以存活得福，并使你们的日子在所要承受的地上得以长久。”
DEUT|6|1|“这是耶和华－你们的上帝所吩咐要教导你们的诫命、律例、典章，叫你们在所要过去得为业的地上遵行，
DEUT|6|2|好叫你和你的子孙在一生的日子都敬畏耶和华－你的上帝，谨守他的一切律例、诫命，就是我所吩咐你的，使你的日子得以长久。
DEUT|6|3|以色列 啊，你要听，要谨守遵行，使你可以在那流奶与蜜之地得福，人数极其增多，正如耶和华－你列祖的上帝所应许你的。
DEUT|6|4|“ 以色列 啊，你要听！耶和华－我们的上帝是独一的主 。
DEUT|6|5|你要尽心、尽性、尽力爱耶和华－你的上帝。
DEUT|6|6|我今日吩咐你的这些话都要记在心上，
DEUT|6|7|也要殷勤教导你的儿女。无论你坐在家里，走在路上，躺下，起来，都要吟诵。
DEUT|6|8|要系在手上作记号，戴在额上 作经匣 ；
DEUT|6|9|又要写在你房屋的门框上和你的城门上。
DEUT|6|10|“耶和华－你的上帝必领你进他向你列祖 亚伯拉罕 、 以撒 、 雅各 起誓要给你的地。那里有又大又美的城镇，不是你建造的；
DEUT|6|11|有装满各样美物的房屋，不是你装满的；有挖成的水井，不是你挖的；有葡萄园、橄榄园，不是你栽植的；你吃了而且饱足。
DEUT|6|12|你要谨慎，免得你忘记领你从 埃及 地为奴之家出来的耶和华。
DEUT|6|13|你要敬畏耶和华－你的上帝，事奉他，奉他的名起誓。
DEUT|6|14|不可随从别神，就是你们四围民族的众神明，
DEUT|6|15|因为在你中间的耶和华－你的上帝是忌邪 的上帝，恐怕耶和华－你上帝的怒气向你发作，把你从地上除灭。
DEUT|6|16|“你们不可试探耶和华－你们的上帝，像你们在 玛撒 那样试探他。
DEUT|6|17|要谨慎遵守耶和华－你们上帝的诫命，和他所吩咐的法度、律例。
DEUT|6|18|耶和华眼中看为正直和美善的事，你都要遵行，使你得福，可以进去得耶和华向你列祖起誓应许的美地，
DEUT|6|19|可以从你面前赶出你所有的仇敌，正如耶和华所说的。
DEUT|6|20|“日后，你的儿子问你说：‘耶和华－我们上帝吩咐你们的法度、律例、典章是什么意思呢？’
DEUT|6|21|你要告诉你的儿子说：‘我们在 埃及 作过法老的奴仆，耶和华用大能的手将我们从 埃及 领出来。
DEUT|6|22|在我们眼前，他施行重大可怕的神迹奇事对付 埃及 、法老和他的全家。
DEUT|6|23|他将我们从那里领出来，为要领我们进入他向我们列祖起誓应许之地，把这地赐给我们。
DEUT|6|24|耶和华又吩咐我们遵行这一切的律例，敬畏耶和华－我们的上帝，使我们一生得福，得以存活，像今日一样。
DEUT|6|25|我们若照耶和华－我们上帝所吩咐的，在他面前谨守遵行这一切诫命，这就是我们的义了。’”
DEUT|7|1|“耶和华－你的上帝领你进入你要得为业之地，从你面前赶出许多国家，就是比你更强大的七个国家： 赫 人、 革迦撒 人、 亚摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人。
DEUT|7|2|当耶和华－你的上帝把他们交给你，你击杀他们的时候，你要完全消灭他们，不可与他们立约，也不可怜惜他们。
DEUT|7|3|不可与他们结亲；不可将你的女儿嫁给他的儿子，也不可叫你的儿子娶他的女儿。
DEUT|7|4|因为他必使你的儿女离弃我，去事奉别神，以致耶和华的怒气向你们发作，迅速将你除灭。
DEUT|7|5|你们却要这样处置他们：拆毁他们的祭坛，打碎他们的柱像，砍断他们的 亚舍拉 ，用火焚烧他们雕刻的偶像。
DEUT|7|6|“因为你是属于耶和华－你上帝神圣的子民；耶和华－你的上帝从地面上的万民中拣选你，作自己宝贵的子民。
DEUT|7|7|耶和华专爱你们，拣选你们，并非因你们人数比任何民族多，其实你们的人数在各民族中是最少的。
DEUT|7|8|因为耶和华爱你们，又因要遵守他向你们列祖所起的誓，耶和华就用大能的手领你们出来，救赎你脱离为奴之家，脱离 埃及 王法老的手。
DEUT|7|9|所以，你知道耶和华－你的上帝，他是上帝，是信实的上帝。他向爱他、守他诫命的人守约施慈爱，直到千代；
DEUT|7|10|向恨他的人，他必当面报应，消灭他们。凡恨他的，他必当面报应，绝不迟延。
DEUT|7|11|所以，你要谨守我今日所吩咐你的诫命、律例、典章，遵行它们。”
DEUT|7|12|“你们若听从这些典章，谨守遵行，耶和华－你的上帝必照他向你列祖所起的誓，对你守约，施慈爱。
DEUT|7|13|他必爱你，赐福给你，使你人数增多，也必在他向你列祖起誓要给你的地上赐福给你身所生的，你地所产的，你的五谷、新酒和新的油，以及你的牛犊、羔羊。
DEUT|7|14|你必蒙福胜过万民；你没有不育的男人和不孕的女人，牲畜也没有不生育的。
DEUT|7|15|耶和华必使一切的疾病远离你；你所知道 埃及 各样的恶疾，他不加在你身上，反要加在所有恨你的人身上。
DEUT|7|16|你要吞灭耶和华－你的上帝交给你的各民族，你的眼目不可顾惜他们。你也不可事奉他们的神明，因为这必成为你的圈套。
DEUT|7|17|“你若心里说，这些国的人数比我多，我怎能赶出他们呢？
DEUT|7|18|你不必怕他们，要牢牢记住耶和华－你上帝向法老和 埃及 全地所行的事，
DEUT|7|19|你亲眼见过的大考验、神迹、奇事、大能的手和伸出来的膀臂，都是耶和华－你上帝领你出来所施行的。耶和华－你的上帝也必照样处置你所惧怕的各民族，
DEUT|7|20|并且耶和华－你的上帝必派瘟疫 攻击他们，直到那剩下而躲起来的人都从你面前灭亡。
DEUT|7|21|不要因他们惊恐，因为耶和华－你的上帝在你中间是大而可畏的上帝。
DEUT|7|22|耶和华－你的上帝必将这些国从你面前渐渐赶出；你不可迅速把他们消灭，免得野地的走兽多起来危害你。
DEUT|7|23|耶和华－你的上帝必将他们交给你，大大扰乱他们，直到他们被除灭。
DEUT|7|24|他又要将他们的君王交在你手中，你必从天下除去他们的名；必无一人能在你面前站立得住，直到你把他们除灭了。
DEUT|7|25|你们要用火焚烧他们神明的雕刻偶像；不可贪爱偶像上的金银，也不可私自收起来，免得你因此陷入圈套，因为这是耶和华－你上帝所憎恶的。
DEUT|7|26|你不可把可憎之物带进你的家，否则，你就像它一样成为当毁灭的。你要彻底憎恨它，极其厌恶它，因为这是当毁灭的。”
DEUT|8|1|“我今日所吩咐你的一切诫命，你们要谨守遵行，好使你们存活，人数增多，可以进去得耶和华向你们列祖起誓应许的那地。
DEUT|8|2|你要记得，这四十年耶和华─你的上帝在旷野一路引导你，是要磨炼你，考验你，为要知道你的心如何，是否愿意遵守他的诫命。
DEUT|8|3|他磨炼你，任你饥饿，将你和你列祖所不认识的吗哪赐给你吃，使你知道，人活着，不是单靠食物，乃是靠耶和华口里所出的一切话。
DEUT|8|4|这四十年，你身上的衣服没有穿破，你的脚也没有肿。
DEUT|8|5|你心里要知道，耶和华─你的上帝管教你，像人管教儿女一样。
DEUT|8|6|你要谨守耶和华─你上帝的诫命，遵行他的道，敬畏他。
DEUT|8|7|“耶和华─你的上帝必领你进入美地，那地有河流，有泉源和深渊的水从谷中和山上流出。
DEUT|8|8|那地有小麦、大麦、葡萄树、无花果树、石榴树，那地也有橄榄油和蜂蜜。
DEUT|8|9|那地没有缺乏，你在那里有食物吃，一无所缺；那地的石头是铁，山中可以挖铜。
DEUT|8|10|你吃得饱足，要称颂耶和华─你的上帝，因为他将那美地赐给你。”
DEUT|8|11|“你要谨慎，免得忘记耶和华─你的上帝，不守他的诫命、典章、律例，就是我今日吩咐你的。
DEUT|8|12|免得你吃得饱足，建造上好的房屋，住在其中，
DEUT|8|13|你的牛羊增多，你的金银增多，你拥有的一切全都增多，
DEUT|8|14|于是你的心高傲，忘记耶和华─你的上帝。他曾将你从 埃及 地为奴之家领出来，
DEUT|8|15|曾引领你经过那大而可怕的旷野，有火蛇、蝎子、干旱无水之地。他也曾为你使水从坚硬的磐石中流出来，
DEUT|8|16|又在旷野将你列祖所不认识的吗哪赐给你吃，为要磨炼你，考验你，终久使你享福。
DEUT|8|17|你心里说：‘这财富是我的力量、我手的能力得来的。’
DEUT|8|18|你要记得耶和华─你的上帝，因为得财富的能力是他给你的，为要坚守他向你列祖起誓所立的约，像今日一样。
DEUT|8|19|你若忘记耶和华─你的上帝，随从别神，事奉它们，敬拜它们，我今日警告你们，你们必定灭亡。
DEUT|8|20|耶和华在你们面前怎样使列国灭亡，你们也必照样灭亡，因为你们不听从耶和华─你们上帝的话。”
DEUT|9|1|“ 以色列 啊，你要听！你今日要过 约旦河 ，进去占领比你更强大的列国，那里的城镇又大，城墙又坚固，如天一样高。
DEUT|9|2|那里的百姓是 亚衲 族人，又高又壮，是你所知道的；你也听说过：‘谁能在 亚衲 族人面前站立得住呢？’
DEUT|9|3|你今日应当知道，耶和华─你的上帝在你前面渡过去，如同吞噬的火，要除灭他们，并要在你面前将他们制伏，使你可以赶出他们，速速消灭他们，正如耶和华向你所说的。
DEUT|9|4|“耶和华─你的上帝将他们从你面前赶出以后，你心里不可说：‘耶和华领我得这地是因我的义。’其实，耶和华将这些国家从你面前赶出去是因他们的恶。
DEUT|9|5|你能进去得他们的地，并不是因你的义，也不是因你心里正直，而是因这些国家的恶，耶和华─你的上帝才把他们从你面前赶出去，为了应验耶和华向你列祖 亚伯拉罕 、 以撒 、 雅各 起誓应许的话。
DEUT|9|6|“你当知道，耶和华─你的上帝将这美地赐你为业，并不是因你的义；你本是硬着颈项的百姓。
DEUT|9|7|你要记得，不要忘记，你在旷野怎样惹耶和华－你的上帝发怒。自从你出了 埃及 地的那日，直到你们来到这地方，你们常常悖逆耶和华。
DEUT|9|8|你们在 何烈山 惹耶和华发怒，耶和华对你们动怒，甚至要除灭你们。
DEUT|9|9|我上了山，要领受两块石版，就是耶和华与你们立约的版。那时我在山上住了四十昼夜，没有吃饭，也没有喝水。
DEUT|9|10|耶和华把那两块石版交给我，是上帝用指头写成的；版上是耶和华在大会的那一天，在山上从火中对你们所说的一切话。
DEUT|9|11|过了四十昼夜，耶和华把那两块石版，就是约版，交给我。
DEUT|9|12|耶和华对我说：‘起来，赶快从这里下去！因为你从 埃及 领出来的百姓已经败坏了；他们这么快偏离了我所吩咐的道，为自己铸造偶像。’
DEUT|9|13|“耶和华对我说：‘我看这百姓，看哪，他们是硬着颈项的百姓。
DEUT|9|14|你且由着我，我要除灭他们，从天下涂去他们的名，我要使你成为比他们更大更强的国。’
DEUT|9|15|于是我转身下山，山上有火燃烧，两块约版在我双手中。
DEUT|9|16|我观看，看哪，你们得罪了耶和华－你们的上帝，为自己铸成了一头牛犊，迅速偏离了耶和华所吩咐你们的道，
DEUT|9|17|我拿着那两块石版，从我双手中扔出去，在你们眼前把它们摔碎了。
DEUT|9|18|因为你们所犯的一切罪，做了耶和华眼中看为恶的事，惹他发怒，我就像从前一样俯伏在耶和华面前四十昼夜，没有吃饭，没有喝水。
DEUT|9|19|我很害怕，因为耶和华向你们大发烈怒，要除灭你们。但那一次耶和华又应允了我。
DEUT|9|20|耶和华也向 亚伦 非常生气，甚至要除灭他；那时我也为 亚伦 祈祷。
DEUT|9|21|我把那使你们犯罪所铸的牛犊拿来，用火焚烧，捣碎后再磨成粉末，好像灰尘。我把这灰尘撒在从山上流下来的溪水中。
DEUT|9|22|“你们在 他备拉 、 玛撒 、 基博罗．哈他瓦 又惹耶和华发怒。
DEUT|9|23|耶和华叫你们离开 加低斯．巴尼亚 ，说：‘你们上去得我所赐给你们的地。’那时，你们违背了耶和华－你们上帝的指示，不信服他，不听从他的话。
DEUT|9|24|自从我认识你们的日子以来，你们常常悖逆耶和华。
DEUT|9|25|“我因耶和华说要除灭你们，就在耶和华面前俯伏四十昼夜，像我以前俯伏一样。
DEUT|9|26|我向耶和华祈祷，说：‘主耶和华啊，求你不要灭绝你的百姓，你的产业。他们是你用大能救赎，用你强有力的手从 埃及 领出来的。
DEUT|9|27|求你记念你的仆人 亚伯拉罕 、 以撒 、 雅各 ，不看这百姓的顽梗、邪恶、罪愆，
DEUT|9|28|免得你领我们出来的那地之人说：耶和华因为不能将这百姓领进他所应许之地，又因恨他们，所以领他们出去，要在旷野杀他们。
DEUT|9|29|其实他们是你的百姓，你的产业，是你用大能和伸出的膀臂领出来的。’”
DEUT|10|1|“那时，耶和华对我说：‘你要凿出两块石版，和先前的一样，上山到我这里来。你也要造一个木柜。
DEUT|10|2|我要把你先前摔碎的版上所写的字，写在这版上；你要把这版放在柜里。’
DEUT|10|3|于是我用金合欢木造了一个柜子，又凿出两块石版，和先前的一样。我手里拿着这两块版上山。
DEUT|10|4|耶和华将那大会之日、在山上从火中所吩咐你们的十条诫命，照先前所写的写在这版上。耶和华把它们交给我。
DEUT|10|5|我转身下山，将这版放在我所造的柜里，现今这版还在那里，正如耶和华所吩咐我的。
DEUT|10|6|（ 以色列 人从 比罗比尼．亚干 起行，来到 摩西拉 ， 亚伦 死在那里，就葬在那里。他的儿子 以利亚撒 接续他担任祭司的职分。
DEUT|10|7|他们从那里起行，来到 谷歌大 ，又从 谷歌大 来到 约巴他 ，有溪水之地。
DEUT|10|8|那时，耶和华将 利未 支派分别出来，抬耶和华的约柜，又侍立在耶和华面前事奉他，奉他的名祝福，直到今日。
DEUT|10|9|因此， 利未 没有像他的弟兄有产业，耶和华是他的产业，正如耶和华－你上帝所应许他的。）
DEUT|10|10|“我又像先前一样在山上停留了四十昼夜。这一次耶和华也应允我，不将你灭绝。
DEUT|10|11|耶和华对我说：‘起来，走在百姓前面，领他们进去得我向他们列祖起誓要给他们的地。’”
DEUT|10|12|“ 以色列 啊，现在耶和华－你的上帝向你要的是什么呢？只要你敬畏耶和华－你的上帝，遵行他一切的道，爱他，尽心尽性事奉耶和华－你的上帝，
DEUT|10|13|遵守耶和华的诫命律例，就是我今日所吩咐你的，为要使你得福。
DEUT|10|14|看哪，天和天上的天，地和地上所有的，都属耶和华－你的上帝。
DEUT|10|15|然而，耶和华专爱你的列祖，爱他们，从万民中拣选你们，就是他们的后裔，像今日一样。
DEUT|10|16|所以你们的心要受割礼，不可再硬着颈项。
DEUT|10|17|因为耶和华－你们的上帝是万神之神，万主之主，是伟大、强有力、可畏的上帝，不看人的情面，也不受贿赂。
DEUT|10|18|他为孤儿寡妇伸冤，爱护寄居的，赐给他衣食。
DEUT|10|19|所以你们要爱护寄居的，因为你们在 埃及 地也作过寄居的。
DEUT|10|20|你要敬畏耶和华－你的上帝，事奉他，紧紧跟随他，奉他的名起誓。
DEUT|10|21|他是你当赞美的，是你的上帝，为你做了大而可畏的事，这些是你亲眼见过的。
DEUT|10|22|你的列祖七十人下 埃及 ，现在耶和华－你的上帝却使你如同天上的星那样多。”
DEUT|11|1|“你要爱耶和华－你的上帝，天天遵守他的吩咐、律例、典章、诫命。
DEUT|11|2|今日你们应当知道，而不是你们的儿女，因为他们不知道，也没有见过耶和华─你们上帝的管教、他的伟大、他大能的手和伸出来的膀臂，
DEUT|11|3|以及他在 埃及 向 埃及 王法老和其全地所行的神迹奇事；
DEUT|11|4|他怎样对待 埃及 的军队、马和战车，他们追赶你们的时候，耶和华怎样用 红海 的水淹没他们，消灭了他们，直到今日；
DEUT|11|5|他在旷野怎样待你们，直到你们来到这地方，
DEUT|11|6|以及他怎样待 吕便 子孙， 以利押 的儿子 大坍 、 亚比兰 ，地怎样在 以色列 人中开了裂口，吞了他们和他们的家眷，帐棚，以及跟他们在一起所有活着的。
DEUT|11|7|惟有你们亲眼见过耶和华所做的一切大事。”
DEUT|11|8|“所以，你们要遵守我今日所吩咐的一切诫命，使你们刚强，可以进去得你们所要得的那地，就是你们将过河到那里要得的，
DEUT|11|9|也使你们的日子，在耶和华向你们列祖起誓要给他们和他们后裔的地上得以长久，那是流奶与蜜之地。
DEUT|11|10|你要进去得为业的那地，不像你出来的 埃及 地。在 埃及 ，你撒种后，要用脚浇灌，像浇灌菜园一样。
DEUT|11|11|你们要过去得为业的那地乃是有山有谷、天上的雨水滋润之地，
DEUT|11|12|是耶和华－你上帝所眷顾的地；从岁首到年终，耶和华－你上帝的眼目时常看顾那地。
DEUT|11|13|“你们若留心听从我今日所吩咐你们的诫命，爱耶和华－你们的上帝，尽心尽性事奉他，
DEUT|11|14|我 必按时降下雨水在你们的地上，就是秋雨和春雨，使你们可以收藏五谷、新酒和新的油，
DEUT|11|15|也必使田野为你的牲畜长出草来；这样，你必吃得饱足。
DEUT|11|16|你们要谨慎，免得心受诱惑，转去事奉别神，敬拜它们，
DEUT|11|17|以致耶和华的怒气向你们发作，使天封闭不下雨，使地不出产，使你们在耶和华所赐给你们的美地上速速灭亡。
DEUT|11|18|“你们要将我这些话存在心里，留在意念中，系在手上作记号，戴在额上 作经匣。
DEUT|11|19|你们也要将这些话教导你们的儿女，无论坐在家里，行在路上，躺下，起来，都要讲论，
DEUT|11|20|又要写在房屋的门框上和你的城门上。
DEUT|11|21|这样，你们和你们子孙的日子必在耶和华向你们列祖起誓要给他们的地上得以增多，如天地之长久。
DEUT|11|22|你们若留心谨守遵行我所吩咐这一切的诫命，爱耶和华－你们的上帝，遵行他一切的道，紧紧跟随他，
DEUT|11|23|他必从你们面前赶出这一切国家，你们也要占领比你们更大更强的国家。
DEUT|11|24|凡你们脚掌所踏之地都必归于你们；从旷野到 黎巴嫩 ，从 幼发拉底 大河，直到西边的海，都要成为你们的疆土。
DEUT|11|25|必无一人能在你们面前站立得住；耶和华－你们的上帝必照他所说的，使惧怕惊恐临到你们所踏的全地。
DEUT|11|26|“看，我今日将祝福与诅咒都陈明在你们面前。
DEUT|11|27|你们若听从耶和华─你们上帝的诫命，就是我今日所吩咐你们的，就必蒙福。
DEUT|11|28|你们若不听从耶和华─你们上帝的诫命，偏离我今日所吩咐你们的道，去随从你们所不认识的别神，就必受诅咒。
DEUT|11|29|当耶和华－你的上帝领你进入要得为业的那地，你就要在 基利心山 上宣布祝福，在 以巴路山 上宣布诅咒。
DEUT|11|30|这二座山岂不是在 约旦河 的那边，日落的方向，在住 亚拉巴 的 迦南 人之地， 吉甲 的前面，靠近 摩利 橡树吗？
DEUT|11|31|你们过 约旦河 ，进去得耶和华－你们的上帝所赐你们为业之地；当你们占领它，在那地居住的时候，
DEUT|11|32|你们要谨守遵行我今日在你们面前颁布的一切律例典章。”
DEUT|12|1|“你们活在世上的日子，在耶和华─你列祖的上帝所赐你为业的地上，你们要谨守遵行这些律例典章：
DEUT|12|2|你们占领的国家所事奉他们众神明的地方，无论是在高山，在小山，在一切的青翠树下，你们要彻底毁坏；
DEUT|12|3|要拆毁他们的祭坛，打碎他们的柱像，用火焚烧他们的 亚舍拉 ，砍断他们神明的雕刻偶像，并要从那地方除去他们的名。
DEUT|12|4|你们不可那样敬拜耶和华－你们的上帝。
DEUT|12|5|但耶和华－你们的上帝在你们各支派中选择何处作为立他名的居所，你们就要到那里求问，
DEUT|12|6|将你们的燔祭、祭物、十一奉献、手中的举祭、还愿祭、甘心祭，以及牛群羊群中头生的，都带到那里。
DEUT|12|7|在那里，你们和你们的全家都可以在耶和华─你们上帝的面前吃，并且因你们手所做的一切蒙耶和华－你的上帝赐福而欢乐。
DEUT|12|8|你们不可做像我们今日在这里所做的，各人行自己眼中看为正的一切事；
DEUT|12|9|因为你们现在还没有进入耶和华－你上帝所赐你的安息，所给你的产业。
DEUT|12|10|你们过了 约旦河 ，住在耶和华─你们上帝给你们承受为业的地；他又使你们得享太平，不受四围一切仇敌扰乱，使你们安然居住。
DEUT|12|11|那时你们要将我所吩咐你们的燔祭、祭物、十一奉献、手中的举祭，和向耶和华许愿的一切上好的祭，都带到耶和华─你们上帝所选择立他名的居所。
DEUT|12|12|你们和儿女、仆婢，以及住在你们城里，没有与你们一起分得产业的 利未 人，都要在耶和华－你们的上帝面前欢乐。
DEUT|12|13|你要谨慎，不可在自己所看中的各处献燔祭。
DEUT|12|14|惟独耶和华从你的一个支派中所选择的地方，你要在那里献燔祭，在那里遵行我一切所吩咐你的。
DEUT|12|15|“然而，你在各城里都可以照着耶和华－你上帝所赐给你的福分，随心所欲宰牲吃肉；无论洁净的人不洁净的人都可以吃，就如吃羚羊和鹿的肉一样。
DEUT|12|16|只是血，你不可吃，要把它倒在地上，如同倒水一样。
DEUT|12|17|你的五谷、新酒和新油的十分之一，或是牛群羊群中头生的，或是你的许愿祭、甘心祭和手中的举祭，都不可在你的城里吃，
DEUT|12|18|必须在耶和华－你的上帝面前吃，在耶和华－你上帝所选择的地方，你和儿女、仆婢，以及住在你城里的 利未 人都可以吃，并要因你手所做的一切，在耶和华－你上帝面前欢乐。
DEUT|12|19|你要谨慎，在你所住的地上，你永不可离弃 利未 人。
DEUT|12|20|“耶和华－你的上帝照他的应许扩张你疆土的时候，你心里想要吃肉，说：‘我要吃肉’，就可以随心所欲吃肉。
DEUT|12|21|耶和华－你上帝选择立他名的地方若离你太远，你可以照我所吩咐的，将耶和华赐给你的牛羊取些宰了，随心所欲在你的城里吃。
DEUT|12|22|其实，就如吃羚羊和鹿的肉一样，你要这样吃它，无论洁净的人不洁净的人都可以一起吃。
DEUT|12|23|但是你要坚定，不可吃血，因为血是生命；不可将生命与肉一起吃。
DEUT|12|24|你不可吃血，要把它倒在地上，如同倒水一样。
DEUT|12|25|不可吃血，好让你和你的子孙可以得福，因为你行了耶和华眼中看为正的事。
DEUT|12|26|只是你分别为圣的物和你所还的愿，都要带到耶和华所选择的地方去。
DEUT|12|27|你的燔祭，连肉带血，都要献在耶和华－你上帝的坛上。祭物的血要倒在耶和华－你上帝的坛上；肉你可以吃。
DEUT|12|28|你要谨守听从我所吩咐的一切话，好让你和你的子孙可以永远得福，因为你行耶和华－你上帝眼中看为善、看为正的事。”
DEUT|12|29|“耶和华－你上帝把你要进去赶出的列国从你面前剪除，并且你得了他们的地为业居住，
DEUT|12|30|那时你要谨慎，在他们从你面前被除灭之后，你不可受引诱随从他们，也不可求问他们的神明，说：‘这些国家怎样事奉他们的神明，我也要照样做。’
DEUT|12|31|你不可向耶和华－你的上帝这样做，因为他们向他们的神明做了耶和华所憎恨、所厌恶的一切事，甚至将自己的儿女用火焚烧，献给他们的神明。
DEUT|12|32|凡我所吩咐你们的事，你们都要谨守遵行，不可加添，也不可删减。”
DEUT|13|1|“你中间若有先知或是做梦的人起来，向你显神迹奇事，
DEUT|13|2|他对你说的神迹奇事应验了，说：‘我们去随从别神，事奉它们吧。’那是你不认识的。
DEUT|13|3|你不可听那先知或是那做梦之人的话，因为这是耶和华－你们的上帝考验你们，要知道你们是否尽心尽性爱耶和华－你们的上帝。
DEUT|13|4|你们要顺从耶和华－你们的上帝，敬畏他，谨守他的诫命，听从他的话，事奉他，紧紧跟随他。
DEUT|13|5|那先知或那做梦的人要被处死，因为他出言悖逆那领你们出 埃及 地、救赎你脱离为奴之家的耶和华－你们的上帝，要引诱你离开耶和华－你上帝吩咐你要行的道。这样，你就把恶从你中间除掉。
DEUT|13|6|“你的同胞兄弟，或是你的儿女，或是你怀中的妻，或是如同自己性命的朋友，若暗中引诱你，说：‘我们去事奉别神吧。’那是你和你列祖所不认识的，
DEUT|13|7|你四围列国的神明，无论是离你近或离你远，从地这边到地那边，
DEUT|13|8|你都不可附和他，也不要听从他。你的眼不可顾惜他，不可怜悯他，也不可袒护他。
DEUT|13|9|你务必杀他；你先下手，然后众百姓才下手，把他处死。
DEUT|13|10|要用石头打死他，因为他想引诱你离开那领你出 埃及 地为奴之家的耶和华－你的上帝。
DEUT|13|11|全 以色列 都要听见而害怕，不敢在你中间再行这样的恶事了。
DEUT|13|12|“若你听见人说，在耶和华－你上帝所赐给你居住的城镇中的一座，
DEUT|13|13|有些无赖之徒从你中间出来，引诱本城的居民，说：‘我们去事奉别神吧。’那是你们不认识的，
DEUT|13|14|你就要调查，探听，细心询问。看哪，是真的，确实有这可憎的事在你中间发生，
DEUT|13|15|你务必用刀杀那城里的居民，把城里所有的，连牲畜都用刀灭尽。
DEUT|13|16|你要把从城里所夺取的一切财物堆在广场中，用火将那城和其中夺取的一切财物全烧给耶和华－你的上帝。那城要永远成为废墟，不得重建。
DEUT|13|17|那当毁灭的物一点都不可粘你的手，好让耶和华转回，不向你发烈怒，却恩待你，怜悯你，照他向你列祖所起的誓使你人数增多；
DEUT|13|18|因为你听从耶和华－你上帝的话，遵守我今日所吩咐你的一切诫命，行耶和华－你上帝眼中看为正的事。”
DEUT|14|1|“你们是耶和华─你们上帝的儿女。不可为了死人割划自己，也不可使额上 光秃；
DEUT|14|2|因为你是属于耶和华－你上帝神圣的子民，耶和华从地面上的万民中拣选了你，作自己宝贵的子民。”
DEUT|14|3|“凡可憎的物， 你都不可吃。
DEUT|14|4|可吃的牲畜是：牛、绵羊、山羊、
DEUT|14|5|鹿、羚、麃子、野山羊、瞪羚、羚羊、山绵羊。
DEUT|14|6|凡蹄分两瓣，分趾蹄而又反刍食物的牲畜，你们都可以吃。
DEUT|14|7|但那反刍或分蹄之中不可吃的是：骆驼、兔子、石獾，虽然反刍却不分蹄，对你们是不洁净的；
DEUT|14|8|猪，虽然分蹄却不反刍，对你们也是不洁净的。它们的肉，你们一点都不可吃；它们的尸体，你们也不可摸。
DEUT|14|9|“水中可吃的是这些：凡有鳍有鳞的都可以吃；
DEUT|14|10|凡无鳍无鳞的都不可吃，对你们是不洁净的。
DEUT|14|11|“凡洁净的鸟，你们都可以吃。
DEUT|14|12|不可吃的是：雕、狗头雕、红头雕、
DEUT|14|13|鹯、小鹰、鹞鹰的类群，
DEUT|14|14|各种乌鸦的类群、
DEUT|14|15|鸵鸟、夜鹰、鱼鹰、鹰的类群、
DEUT|14|16|鸮鸟、猫头鹰、角鸱、
DEUT|14|17|鹈鹕、秃雕、鸬鹚、
DEUT|14|18|鹳、鹭鸶的类群、戴鵀与蝙蝠。
DEUT|14|19|凡有翅膀却爬行的群聚动物对你们是不洁净的，都不可吃。
DEUT|14|20|凡洁净的鸟，你们都可以吃。
DEUT|14|21|“凡自然死去的动物，你们都不可吃，可以给城里寄居的人吃，或卖给外人，因为你是属于耶和华－你上帝神圣的子民。 “不可用母山羊的奶来煮它的小山羊。”
DEUT|14|22|“每年，你务必从你播种的一切收成，田地所出产的，取十分之一献上。
DEUT|14|23|要在耶和华－你上帝面前，就是他选择那里作为他名居所的地方，吃你所献十分之一的五谷、新酒和新的油，以及牛群羊群中头生的，好让你天天学习敬畏耶和华－你的上帝。
DEUT|14|24|当耶和华－你的上帝赐福给你的时候，耶和华－你上帝选择立他名的地方若离你太远，路途太长，使你不能把这东西带到那里去，
DEUT|14|25|你可以把它换成银子，把银子包起来，拿在手中，往耶和华－你上帝所选择的地方去。
DEUT|14|26|在那里，你可以随心所欲用银子或买牛羊，或买清酒烈酒，或买任何你心所想的。你和你的全家要在耶和华－你上帝面前吃喝欢乐。
DEUT|14|27|“住在你城里的 利未 人，你不可离弃他，因为他在你那里没有分得产业。
DEUT|14|28|每三年的最后一年，你要把那一年收成的十分之一取出来，积存在你的城中；
DEUT|14|29|那没有与你一起分得产业的 利未 人，和城里的寄居者，以及孤儿寡妇，都可以前来，吃得饱足，好让耶和华－你的上帝在你手里所做的一切事上赐福给你。”
DEUT|15|1|“每七年的最后一年，你要施行豁免。
DEUT|15|2|豁免的方式是这样：凡债主要把手里所借给邻舍的全豁免，不可向邻舍和弟兄追讨，因为耶和华的豁免已经宣告了。
DEUT|15|3|你可以向外邦人追讨；但你弟兄欠你的，无论是什么，你都要放手豁免。
DEUT|15|4|其实，在你中间不会有贫穷人；因为在耶和华－你上帝所赐你为业的地上，耶和华必大大赐福给你。
DEUT|15|5|只要你留心听从耶和华－你上帝的话，谨守遵行我今日所吩咐你这一切的命令，
DEUT|15|6|因为耶和华－你的上帝会照他所应许你的赐福给你，你必借给许多国家，却不需要去借贷；你要管辖许多国家，它们却不能管辖你。
DEUT|15|7|“在耶和华－你上帝所赐给你的地上，任何一座城里，你弟兄中若有一个贫穷人，你不可硬着心，袖手不帮助你贫穷的弟兄。
DEUT|15|8|你总要伸手帮助他，照他所缺乏的借给他，补他的不足。
DEUT|15|9|你要谨慎，不可心起恶念，说：‘第七年的豁免年快到了’，你就冷眼看你贫穷的弟兄，什么都不给他。他若为你的缘故求告耶和华，你就有罪了。
DEUT|15|10|你要慷慨解囊，给他的时候不要心疼，因为耶和华－你的上帝必为这事，在你一切的工作上和你手所做的一切赐福给你。
DEUT|15|11|因为地上的贫穷人永远不会断绝，所以我吩咐你说：‘总要伸手帮助你地上困苦贫穷的弟兄。’”
DEUT|15|12|“你弟兄中，若有一个 希伯来 男人或 希伯来 女人卖给你，已服事你六年，到了第七年就要让他自由离开你。
DEUT|15|13|你让他自由离开的时候，不可让他空手而去，
DEUT|15|14|要从你的羊群、禾场、压酒池中取一些，慷慨地送给他；耶和华－你的上帝怎样赐福给你，你也要照样给他。
DEUT|15|15|要记得你在 埃及 地作过奴仆，耶和华－你的上帝救赎了你。为此，我今日将这事吩咐你。
DEUT|15|16|他若对你说：‘我不愿意离开你’，因为他爱你和你的家，并且他在你那里很好，
DEUT|15|17|你要拿锥子在门上穿透他的耳朵，他就永远成为你的奴仆了。你待婢女也要这样。
DEUT|15|18|你让他从你那里自由离开的时候，不要看作困难，因为他已服事你六年，相当于雇工双倍的工钱。这样，耶和华－你的上帝必在你所做的一切事上赐福给你。”
DEUT|15|19|“你牛群羊群中头生的，凡是公的，都要分别为圣，归给耶和华－你的上帝。头生的牛，不可用它来耕作；头生的羊，不可剪它的毛。
DEUT|15|20|这头生的，你和你全家每年要到耶和华所选择的地方，在耶和华－你上帝面前吃。
DEUT|15|21|这头生的若有残疾，瘸腿的或瞎眼的，若有任何严重缺陷，都不可献给耶和华－你的上帝。
DEUT|15|22|你们可以在城里吃，洁净的人和不洁净的人都可以吃，就如吃羚羊和鹿一样。
DEUT|15|23|只是它的血，你不可吃，要倒在地上，如同倒水一样。”
DEUT|16|1|“你要守亚笔月，向耶和华－你的上帝守逾越节，因为在亚笔月，耶和华－你的上帝在夜间领你出 埃及 。
DEUT|16|2|你当在那里，耶和华选择作为他名居所的地方，从羊群牛群中，将逾越节的祭牲献给耶和华－你的上帝。
DEUT|16|3|这祭牲不可和有酵的东西一起吃。因为你曾匆忙离开 埃及 地，你要吃无酵饼，就是困苦饼七日，好让你一生的年日记得你从 埃及 地出来的那一日。
DEUT|16|4|在你全境内，七日不可见到酵母。第一日晚上所献的肉，一点也不可留到早晨。
DEUT|16|5|你不可在耶和华－你上帝所赐的各城中，任何一座城里，献逾越节的祭，
DEUT|16|6|只可在那里，耶和华－你上帝选择作为他名居所的地方，在晚上日落的时候，就是你出 埃及 的时候，献逾越节的祭。
DEUT|16|7|你要在耶和华－你上帝所选择的地方把肉烤来吃，次日早晨就回到你的帐棚去。
DEUT|16|8|你要吃无酵饼六日，第七日要向耶和华－你的上帝守严肃会，不可做工。”
DEUT|16|9|“你要计算七个七日：从你用镰刀开始收割庄稼时算起，一共七个七日。
DEUT|16|10|你要向耶和华－你的上帝守七七节，按照耶和华－你上帝所赐你的福，献上你手里的甘心祭。
DEUT|16|11|你和你的儿女、仆婢，以及住在你城里的 利未 人、在你中间寄居的和孤儿寡妇，都要在那里，耶和华－你上帝选择作为他名居所的地方，在耶和华－你上帝面前欢乐。
DEUT|16|12|你要记得你在 埃及 作过奴仆，也要谨守遵行这些律例。”
DEUT|16|13|“你收藏了禾场和压酒池的出产以后，就要守住棚节七日。
DEUT|16|14|在节期中，你和你的儿女、仆婢，以及住在你城里的 利未 人、寄居的和孤儿寡妇，都要欢乐。
DEUT|16|15|在耶和华所选择的地方，你要向耶和华－你的上帝守节七日，因为耶和华－你的上帝要在你一切的收成上和你手里所做的一切赐福给你，你就非常欢乐。
DEUT|16|16|“你所有的男丁要在除酵节、七七节、住棚节，一年三次，在耶和华－你上帝所选择的地方朝见他，不可空手朝见耶和华。
DEUT|16|17|各人要按自己手中的能力，照耶和华－你上帝所赐你的福，奉献礼物。”
DEUT|16|18|“你要在耶和华－你上帝所赐的各城中，为各支派设立审判官和官长。他们要按公义的判断审判百姓，
DEUT|16|19|不可屈枉正直，不可看人的情面，也不可接受贿赂，因为贿赂能使智慧人的眼睛变瞎，又能曲解义人的证词。
DEUT|16|20|公正！你要追求公正，好使你存活，承受耶和华－你上帝所赐你的地。”
DEUT|16|21|“你为耶和华－你的上帝筑坛，不可在坛旁栽种任何树木作 亚舍拉 ，
DEUT|16|22|也不可为自己设立柱像，这是耶和华－你的上帝所憎恨的。”
DEUT|17|1|“凡有残疾，有任何恶疾的牛羊，你都不可献给耶和华－你的上帝，因为这是耶和华－你上帝所憎恶的。
DEUT|17|2|“在你中间，在耶和华－你上帝所赐你的各城中，任何一座城里，若有男人或女人做了耶和华－你上帝眼中看为恶的事，违背了他的约，
DEUT|17|3|去事奉别神，敬拜它们，或拜太阳，或拜月亮，或拜天上的万象，是我 不曾吩咐的。
DEUT|17|4|有人告诉你，你也听见了，就要细心探听。看哪，是真的，确实有这可憎的事在 以色列 中发生，
DEUT|17|5|你就要将行这恶事的男人或女人拉到城门外，用石头把这男人或女人处死。
DEUT|17|6|要凭两个证人或三个证人的口，才可以把他处死，不可只凭一个证人的口处死他。
DEUT|17|7|证人要先动手，然后众百姓也动手把他处死。这样，你就把恶从你中间除掉。
DEUT|17|8|“你城中若有难以判断的案件，涉及流血，诉讼，或殴打等争讼的事，你就要起来，上到那里，耶和华－你上帝所选择的地方，
DEUT|17|9|去见 利未 家的祭司和当时的审判官，求问他们，他们必将判决指示你。
DEUT|17|10|他们在耶和华所选择的地方指示你的判决，你要执行，谨守遵行他们一切所教导你的。
DEUT|17|11|要按照所教导你的律法、所告诉你的典章去执行；他们指示你的判决，你不可偏离左右。
DEUT|17|12|若有人擅自行事，不听从那侍立在耶和华－你上帝那里事奉的祭司，或不听从审判官，那人就要处死。这样，你就把恶从 以色列 中除掉。
DEUT|17|13|众百姓听见了都要害怕，不再擅自行事了。”
DEUT|17|14|“你到了耶和华－你上帝所赐你的地，得了那地居住在其中的时候，若说：‘我要立王治理我，像我四围所有的国家一样’，
DEUT|17|15|你一定要立耶和华－你上帝所拣选的人为你的王。要从你弟兄中立一人为你的王，不可立你弟兄之外的外邦人治理你。
DEUT|17|16|只是王不可为自己加添马匹，也不可为加添马匹使百姓回 埃及 去，因耶和华曾对你们说：‘不可再回那条路去。’
DEUT|17|17|王不可为自己多立妃嫔，免得他的心偏离；也不可为自己多积金银。
DEUT|17|18|他登了国度的王位之后，要在 利未 家的祭司面前，将这律法书为自己抄写一份在书卷上。
DEUT|17|19|这书要存在他那里，他一生的年日要诵读，好使他学习敬畏耶和华－他的上帝，谨守遵行这律法书上的一切话和这些律例，
DEUT|17|20|免得他的心向弟兄高傲，偏离了这诫命，或向右或向左。这样，他和他的子孙就可以长久作王治理 以色列 。”
DEUT|18|1|“ 利未 家的祭司和 利未 全支派在 以色列 中没有分得产业；他们可以吃耶和华的火祭，那是他的产业。
DEUT|18|2|他在弟兄中没有产业；耶和华是他的产业，正如耶和华所应许他的。
DEUT|18|3|祭司从百姓当得的权益是这样：凡献牛或羊为祭物的，要把前腿、两腮和胃给祭司。
DEUT|18|4|初收的五谷、新酒和新的油，以及初剪的羊毛，也要给他。
DEUT|18|5|因为耶和华－你的上帝从你众支派中拣选他，使他和他子孙永远奉耶和华的名侍立，事奉。
DEUT|18|6|“ 利未 人若离开他在 以色列 中所居住的任何一座城，一心愿意到耶和华所选择的地方，
DEUT|18|7|就要在那里奉耶和华－他上帝的名事奉，正如他的众弟兄 利未 人在耶和华面前侍立一样。
DEUT|18|8|除了卖祖产所得的以外，他们 要吃同等分量的祭物。”
DEUT|18|9|“你到了耶和华－你上帝所赐你之地，不可学那些国家行可憎恶的事。
DEUT|18|10|你中间不可有人使儿女经火，也不可有占卜的、观星象的、行法术的 、行邪术的、
DEUT|18|11|施符咒的、招魂的、行巫术的和求问死人的。
DEUT|18|12|凡做这些事的都是耶和华所憎恶的；因这可憎恶的事，耶和华－你的上帝把他们从你面前赶出去。
DEUT|18|13|你要向耶和华－你的上帝作完全人。
DEUT|18|14|你所要赶出的那些国家都听从观星象的和占卜的，但是耶和华－你的上帝从来不准你这样做。”
DEUT|18|15|“耶和华－你的上帝要从你弟兄中给你兴起一位先知像我，你们要听他。
DEUT|18|16|这正如你在 何烈山 大会的那日向耶和华－你的上帝所求的一切，说：‘求你不要再叫我听见耶和华－我上帝的声音，也不要再叫我看见这大火，免得我死亡。’
DEUT|18|17|耶和华对我说：‘他们说得对。
DEUT|18|18|我必在他们弟兄中给他们兴起一位先知像你。我要将当说的话放在他口里；他要将我一切所吩咐的都告诉他们。
DEUT|18|19|谁不听从他奉我名所说的话，我必亲自向他追究。
DEUT|18|20|若有先知擅自奉我的名说了我未曾吩咐他说的话，或是奉别神的名说话，那先知就必处死。’
DEUT|18|21|你心里若说：‘我们怎能知道那话是耶和华未曾吩咐的呢？’
DEUT|18|22|先知奉耶和华的名说话，所说的若没有实现，或不应验，这话就是耶和华未曾吩咐的，而是那先知擅自说的，你不必怕他。”
DEUT|19|1|“耶和华－你的上帝将列国剪除，他们的地耶和华－你上帝已赐给你，你又赶出他们，并且住在他们的城镇和房屋，
DEUT|19|2|那时，你要在耶和华－你上帝所赐你为业的地上，为自己指定三座城。
DEUT|19|3|你要预备道路，将耶和华－你上帝使你承受为业的地分为三区，使任何一个杀人的可以逃到那里去。
DEUT|19|4|“杀人的逃到那里得以存活的案例是这样：凡素无仇恨，无意中杀了邻舍的，
DEUT|19|5|就如人与邻舍同入林中伐木，手拿斧子一砍，本想砍下树木，斧头却脱了把，飞落在邻舍身上，以致那人死去，这人就可以逃到那些城中的一座，得以存活，
DEUT|19|6|免得报血仇的心中发火，去追赶那杀了人的，因为路途遥远就能追上他，把他杀死。其实他是不该死的，因为他与被杀者素无仇恨。
DEUT|19|7|所以我吩咐你说，要为自己指定三座城。
DEUT|19|8|耶和华－你的上帝若照他向你列祖所起的誓扩张你的疆土，将所应许赐你列祖的全地给你，
DEUT|19|9|你若谨守遵行我今日所吩咐的这一切诫命，爱耶和华－你的上帝，天天遵行他的道，就要在这三座城之外，再添三座城，
DEUT|19|10|免得无辜人的血流在耶和华－你上帝所赐你为业的地中间，血就归到你身上了。
DEUT|19|11|“若有人恨他的邻舍，埋伏等着，起来击杀他，把他杀死，然后逃到这些城中的一座，
DEUT|19|12|他本城的长老就要派人去，从那里把他带出来，交在报血仇者的手中，把他处死。
DEUT|19|13|你的眼不可顾惜他，要从 以色列 中除掉流无辜血的罪，使你得福。”
DEUT|19|14|“在耶和华－你上帝所赐你承受为业，所分得的地上，不可挪移你邻舍的地界，因为这是前人所定的。”
DEUT|19|15|“人无论犯什么罪，作什么恶，不可单凭一个人的见证，总要凭两个证人的口或三个证人的口才可定案。
DEUT|19|16|若有人怀恶意，起来作证，控告他人犯法，
DEUT|19|17|这两个争讼的人就要站在耶和华面前，和当时的祭司与审判官面前，
DEUT|19|18|审判官要细心调查。看哪，证人作的是伪证，要用伪证陷害弟兄，
DEUT|19|19|你们就要对付他如同他想要对付的弟兄一样。这样，你就把恶从你中间除掉。
DEUT|19|20|其他的人听见就害怕，不敢在你中间再行这样的恶事了。
DEUT|19|21|你的眼不可顾惜，要以命偿命，以眼还眼，以牙还牙，以手还手，以脚还脚。”
DEUT|20|1|“你出去与仇敌作战，若看见马匹、战车，以及比你更多的士兵，不要怕他们，因为领你出 埃及 地的耶和华－你的上帝与你同在。
DEUT|20|2|你们将要上阵的时候，祭司要来，向士兵宣告，
DEUT|20|3|对他们说：‘ 以色列 啊，要听！你们今日将要与仇敌作战，不要心惊胆战，不要惧怕战兢，也不要因他们惊慌，
DEUT|20|4|因为与你们同去的是耶和华－你们的上帝，他要为你们与仇敌作战，拯救你们。’
DEUT|20|5|官长也要向士兵宣告说：‘谁建了新的房屋尚未奉献，他可以回家去，免得他阵亡，别人去奉献。
DEUT|20|6|谁栽植了葡萄园尚未享用所结的果子，他可以回家去，免得他阵亡，别人去享用。
DEUT|20|7|谁与女子订了婚尚未迎娶，他可以回家去，免得他阵亡，别人去娶。’
DEUT|20|8|官长要继续对士兵说：‘谁惧怕，心惊胆战，可以回家去，免得他弟兄的心像他的心一样消沉。’
DEUT|20|9|官长向士兵宣告完毕，军官就率领士兵去了。
DEUT|20|10|“你来到一座城，要攻城之前，先向它宣告和平。
DEUT|20|11|那城若愿意以和平回应，给你开城，城里所有的人就要为你做苦工，服事你。
DEUT|20|12|若那城拒绝和平，却要与你打仗，你就要围困那城。
DEUT|20|13|耶和华－你的上帝把那城交在你手里时，你就要用刀杀尽城里的男丁。
DEUT|20|14|至于妇女、孩童、牲畜和城里所有的，你都可以取为自己的掠物。从仇敌所掠夺的，就是耶和华－你上帝所赐给你的，你都可以享用。
DEUT|20|15|离你很远的各城，就是不属于这些国家的城镇，你都要这样对待他们。
DEUT|20|16|但是这些民族的城镇，就是耶和华－你上帝所赐给你的产业，其中凡有气息的，一个都不可存留。
DEUT|20|17|你要照耶和华－你上帝所吩咐的，将这些 赫 人、 亚摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人全都灭绝，
DEUT|20|18|免得他们教导你们去行一切可憎恶的事，就是他们向自己神明所行的，使你们得罪耶和华－你们的上帝。
DEUT|20|19|“你若围困一座城，需要攻打许多日子才能夺取，就不可用斧头砍坏树木。你可以吃树上的果子，却不可把树砍下来。田间的树木岂是人，让你去围攻的吗？
DEUT|20|20|只有那些你知道不能生产食物的树才可以毁坏；你可以把它们砍下来造攻城的工具，攻打那与你打仗的城，直到把城攻下。”
DEUT|21|1|“在耶和华－你上帝所赐你为业的地上，若发现有人被杀，暴尸野地，不知道是谁杀的，
DEUT|21|2|长老和审判官 就要出去，从尸体那里量起，量到四围的城镇，
DEUT|21|3|看哪一座城最靠近这尸体，那城的几位长老就要取一头未曾耕地、未曾负轭的母牛犊；
DEUT|21|4|那城的长老要把这母牛犊牵到流着溪水、未曾耕耘、未曾撒种的山谷去，在谷中打断它的颈项。
DEUT|21|5|利未 人祭司要近前来，因为耶和华－你的上帝拣选他们来事奉他，奉耶和华的名祝福，并且有任何的争讼和殴打，都由他们的口判决。
DEUT|21|6|离尸体最近的那座城的每位长老要在山谷中，在颈项被打断的母牛犊上面洗手，
DEUT|21|7|声明说：‘我们的手未曾流这人的血；我们的眼也未曾看见这事。
DEUT|21|8|耶和华啊，求你赦免你所救赎的百姓 以色列 ，不要让无辜的血归在你的百姓 以色列 中间。’这样，他们流血的罪就必得赦免。
DEUT|21|9|你行了耶和华眼中看为正的事，就可以从你中间除掉无辜的血。”
DEUT|21|10|“你出去与仇敌作战的时候，耶和华－你的上帝将他交在你手中，你就掳了他为俘虏。
DEUT|21|11|若你在被掳的人中看见美丽的女子，喜欢她，要娶她为妻，
DEUT|21|12|就可以带她到你家去。她要剪头发，修指甲，
DEUT|21|13|脱去被掳时所穿的衣服，住在你家里为自己父母哀哭一个月。然后，你就可以与她同房；你作她的丈夫，她作你的妻子。
DEUT|21|14|以后你若不喜欢她，就要让她自由离开，绝不可为钱把她卖了，也不可把她当奴隶看待，因为你已经占有过她。”
DEUT|21|15|“人若有两个妻子，一个是他宠爱的，另一个是失宠的 ，她们都给他生了儿子，但长子是他失宠妻子生的；
DEUT|21|16|到了分产业给儿子的时候，不可将自己宠爱的妻子所生的儿子立为长子，在他失宠妻子所生的长子之上。
DEUT|21|17|他必须认失宠妻子所生的儿子为长子，在所有的产业中给他双分，因为这儿子是他壮年时生的，长子的名分应当是他的。”
DEUT|21|18|“人若有顽梗忤逆的儿子，不听从父母的话，他们虽然惩戒他，他还是不听从他们，
DEUT|21|19|父母就要抓住他，带他出去到当地的城门，本城的长老那里，
DEUT|21|20|对本城的长老说：‘我们这个儿子顽梗忤逆，不听从我们的话，是贪食好酒的人。’
DEUT|21|21|然后，城里的众人就要用石头将他打死。这样，你就把恶从你中间除掉，全 以色列 听见了都要害怕。”
DEUT|21|22|“人若犯了死罪被处死，你把他挂在木头上，
DEUT|21|23|不可让尸体留在木头上过夜，一定要当日把他埋葬，因为被挂的人是上帝所诅咒的。你不可玷污耶和华－你上帝所赐你为业的地。”
DEUT|22|1|“你若看见弟兄的牛或羊迷了路，不可避开它们，总要把它们牵回来交给你的弟兄。
DEUT|22|2|你弟兄若离你远，或是你不认识他，你就要牵到你家，留在你那里，等你的弟兄来寻找就还给他。
DEUT|22|3|你弟兄所失落的，无论是驴，衣服，或任何东西，你若发现，都要这样做，不能避开。
DEUT|22|4|你若看见你弟兄的牛或驴在路上跌倒了，不可避开它们，总要帮助他把牛或驴拉起来。
DEUT|22|5|“妇女不可穿戴男子所穿戴的，男人也不可穿妇女的衣服，因为这样做是耶和华－你上帝所憎恶的。
DEUT|22|6|“你若路上看见鸟窝，无论在树上或地上，里头有小鸟或有蛋，母鸟伏在小鸟或蛋上，你不可连母鸟带小鸟一起拿去。
DEUT|22|7|总要放母鸟走，只可以取小鸟。这样你就可以享福，日子得以长久。
DEUT|22|8|“你若建造新房屋，要在屋顶安栏杆，免得有人从屋顶掉下来，血就归于你家。
DEUT|22|9|“不可在你的葡萄园里栽种别的种子，免得你栽种所结的和葡萄园的果子都成了圣物。
DEUT|22|10|不可并用牛和驴来耕地。
DEUT|22|11|不可穿羊毛和细麻混合做成的衣服。
DEUT|22|12|“你要在所披外衣的四个边上缝繸子。”
DEUT|22|13|“人若娶妻，与她同房后恨恶她，
DEUT|22|14|捏造她行可耻的事，把丑名加在她身上，说：‘我娶了这女人，亲近她，却发现她没有贞洁的凭据’。
DEUT|22|15|女方的父母就要把这女子贞洁的凭据拿出去，到城门的本城长老那里。
DEUT|22|16|女方的父亲要对长老说：‘我把女儿嫁给这人，他却恨恶她，
DEUT|22|17|看哪，他捏造可耻的事，说：我发现你女儿没有贞洁的凭据。但是，这就是我女儿贞洁的凭据。’父母要把那布铺在本城长老的面前。
DEUT|22|18|那城的长老要拿住那人，惩罚他，
DEUT|22|19|罚他一百银子，给女方的父亲，因为他把丑名加在 以色列 一个少女身上。这女子仍是他的妻子，那人终身不可休她。
DEUT|22|20|但若这事是真的，找不到女子贞洁的凭据，
DEUT|22|21|他们就要把这女子带到她父家的门口，城里的人要用石头打死她，因为她在父家犯了淫乱，在 以色列 中做了可耻的事。这样，你就把恶从你中间除掉。
DEUT|22|22|“若发现有人与有夫之妇同寝，就要将奸夫淫妇一起处死。这样，你就把恶从 以色列 中除掉。
DEUT|22|23|“若一女子是处女，已经许配了人，有男子在城里遇见她，与她同寝，
DEUT|22|24|你们就要把这二人带到那城的城门口，用石头打死他们。处死女子是因为她虽然在城里， 却没有喊叫；处死男子是因为他玷污了邻舍的妻子。这样，你就把恶从你中间除掉。
DEUT|22|25|“若有男子在野地遇见已经许配人的女子，抓住她与她同寝，只要处死那与女子同寝的男子。
DEUT|22|26|不可对女子处刑，这女子没有该死的罪。这案件就好比人起来攻击邻舍，把他杀了一样。
DEUT|22|27|因为男子是在野地遇见她，这已经许配了人的女子虽然喊叫，却没有人救她。
DEUT|22|28|“若有男子遇见没有许配人的少女，抓住她与她同寝，被人发现，
DEUT|22|29|这男子就要拿五十银子给女子的父亲，并要娶她为妻，终身不可休她，因为他玷污了这女子。
DEUT|22|30|“人不可娶继母为妻，不可掀开父亲衣服的下边 。”
DEUT|23|1|“凡外肾损伤的，或被阉割的，不可入耶和华的会。
DEUT|23|2|“私生子不可入耶和华的会；甚至到第十代，也不可入耶和华的会。
DEUT|23|3|“ 亚扪 人或 摩押 人不可入耶和华的会；甚至到第十代，也永不可入耶和华的会。
DEUT|23|4|因为你们出 埃及 的时候，他们没有拿食物和水在路上迎接你们，并且雇了 美索不达米亚 的 毗夺 人， 比珥 的儿子 巴兰 来诅咒你。
DEUT|23|5|然而耶和华－你的上帝不愿听 巴兰 ，耶和华－你的上帝为你使诅咒变为祝福，因为耶和华－你的上帝爱你。
DEUT|23|6|你一生一世永不可为他们求平安和福气。
DEUT|23|7|“不可憎恶 以东 人，因为他是你的弟兄。不可憎恶 埃及 人，因为你曾在他的地上作过寄居的。
DEUT|23|8|他们所生的第三代子孙可以入耶和华的会。”
DEUT|23|9|“你出兵攻打敌人，要远离一切恶事。
DEUT|23|10|“你中间若有人因夜间梦遗而不洁净，就要出到营外，不可入营。
DEUT|23|11|到了傍晚，他要用水洗澡，等到日落才可以入营。
DEUT|23|12|“你要在营外划定一个地方，你可以出去在那里方便。
DEUT|23|13|在你器械中当有一把锹；你出营外便溺以后，要用它挖洞，转身掩盖排泄物。
DEUT|23|14|因为耶和华－你的上帝在你营中走动，要拯救你，将仇敌交给你，所以你的营应当圣洁，免得他见你那里有污秽之物就转身离开你。”
DEUT|23|15|“你不可把从主人身边逃到你那里的奴仆，交回给他的主人，
DEUT|23|16|要让他在你那里与你同住，由他在你的城镇中选择一个自己喜欢的地方居住，不可欺负他。
DEUT|23|17|“ 以色列 的女子中不可作神庙娼妓； 以色列 的男子中也不可作神庙娼妓。
DEUT|23|18|妓女和男娼 的赏金，都不可带进耶和华－你上帝的殿中还愿，因为两者都是耶和华－你上帝所憎恶的。
DEUT|23|19|“你借给你弟兄的，无论是钱财是粮食，或任何可生利息的财物，都不可取利。
DEUT|23|20|借给外邦人可以取利，但借给你的弟兄就不可取利；好让耶和华－你的上帝在你去得为业的地上和你手里所做的一切，赐福给你。
DEUT|23|21|“你向耶和华－你的上帝许愿，不可迟延还愿，因为耶和华－你的上帝必定向你追讨，你就有罪了。
DEUT|23|22|你若不许愿，倒没有罪。
DEUT|23|23|你嘴唇所说的，你亲口承诺的，要照你甘心向耶和华－你上帝许的愿谨守遵行。
DEUT|23|24|“你进入邻舍的葡萄园，可以随意吃葡萄，直到饱足，却不可装在器皿中。
DEUT|23|25|你进入邻舍的庄稼中，可以用手摘麦穗，却不可用镰刀割取庄稼。”
DEUT|24|1|“人若娶妻，作了她的丈夫，发现她有不合宜的事不喜欢她，而写休书交在她手中，打发她离开夫家，
DEUT|24|2|妇人若离开夫家以后，去嫁别人，
DEUT|24|3|后夫若恨恶她，写休书交在她手中，打发她离开夫家，又或者娶她为妻的后夫死了，
DEUT|24|4|那休她的前夫就不可在妇人玷污之后再娶她为妻，因为这是耶和华所憎恶的。不可使耶和华－你上帝所赐为业之地蒙受玷污。
DEUT|24|5|“人若娶了新娘，不可从军出征，也不可派他办理任何事情。他可以在家清闲一年，使他所娶的妻快活。
DEUT|24|6|“不可拿人的石磨或上面的磨石作抵押，因为这是拿人的命作抵押。
DEUT|24|7|“若发现有人绑架 以色列 人中的一个弟兄，把他当奴隶对待，或把他卖了，那绑架人的就必处死。这样，你就把恶从你中间除掉。
DEUT|24|8|“关于痲疯 的灾病，你们要谨慎，照 利未 家的祭司一切所指教你们的留心遵行。我怎样吩咐他们，你们要照样遵行。
DEUT|24|9|要记得，在你们出 埃及 后的路途中，耶和华－你的上帝向 米利暗 所做的事。
DEUT|24|10|“你借给邻舍，无论是什么，不可进他家拿抵押品。
DEUT|24|11|要站在外面，等那借贷的人把抵押品拿出来交给你。
DEUT|24|12|他若是困苦的人，你不可用他的抵押品盖着睡觉。
DEUT|24|13|日落的时候，总要把抵押品还给他，让他用那件外衣盖着睡觉，他就为你祝福。这在耶和华－你的上帝面前就是你的义行了。
DEUT|24|14|“困苦贫穷的雇工，无论是你的弟兄，或是住在你境内，在你城里寄居的，你都不可欺负他 。
DEUT|24|15|要当日给他工钱，不可等到日落，因为他困苦，需要靠工钱过活，免得他因你的缘故求告耶和华，罪就归于你了。
DEUT|24|16|“不可因儿子处死父亲，也不可因父亲处死儿子；各人要因自己的罪被处死。
DEUT|24|17|“不可对寄居的和孤儿屈枉正直，也不可拿寡妇的衣服作抵押。
DEUT|24|18|要记得你曾在 埃及 作过奴仆，耶和华－你的上帝从那里救赎了你，所以我吩咐你遵行这事。
DEUT|24|19|“你在田间收割庄稼，若忘了一捆在田间，就不要再回去拿，要留给寄居的、孤儿和寡妇；好让耶和华－你的上帝在你手里所做的一切，赐福给你。
DEUT|24|20|你打了橄榄树，枝上剩下的不可再打，要留给寄居的、孤儿和寡妇。
DEUT|24|21|你摘葡萄园的葡萄，掉落的不可拾取，要留给寄居的、孤儿和寡妇。
DEUT|24|22|你要记得你曾在 埃及 地作过奴仆，所以我吩咐你遵行这事。
DEUT|25|1|“人与人若有争讼，要求审判，当宣判义人为义，恶人有罪的时候，
DEUT|25|2|恶人若该受责打，审判官就要叫他当着面，伏在地上，按他的罪照数责打。
DEUT|25|3|只能打四十下，不可加多；多过这数目就是在你眼中作贱你的弟兄了。
DEUT|25|4|“牛在踹谷的时候，不可笼住它的嘴。”
DEUT|25|5|“兄弟住在一起，若其中一个死了，没有儿子，死者的妻子就不可出去嫁给陌生人。她丈夫的兄弟应当尽兄弟的本分，娶她为妻，与她同房。
DEUT|25|6|妇人生的长子要归在已故兄弟的名下，免得他的名在 以色列 中涂去了。
DEUT|25|7|那人若不情愿娶他兄弟的妻子，他兄弟的妻子就要上到城门长老那里，说：‘我丈夫的兄弟拒绝在 以色列 中为他的兄弟留名，不愿意为我尽兄弟的本分。’
DEUT|25|8|本城的长老就要召那人来，跟他谈话。若他坚持说：‘我不情愿娶她。’
DEUT|25|9|他兄弟的妻子就要在长老眼前来到那人跟前，脱下他脚上的鞋，吐唾沫在他脸上，回应说：‘凡不为兄弟建立家室的都要这样待他。’
DEUT|25|10|在 以色列 中，他要以‘脱鞋之家’闻名。”
DEUT|25|11|“若有人和弟兄争斗，其中一人的妻子近前去，为了救丈夫脱离那打丈夫之人的手，伸手抓住那人的下体，
DEUT|25|12|你就要砍断妇人的手，你的眼不可顾惜。
DEUT|25|13|“你袋中不可有一大一小两样的法码。
DEUT|25|14|你家里不可有一大一小两样的伊法 。
DEUT|25|15|当用准确公正的法码和伊法，好使你的日子在耶和华－你上帝所赐你的地上得以长久。
DEUT|25|16|因为行这一切不义之事的人都是耶和华－你上帝所憎恶的。”
DEUT|25|17|“你要记得你们出 埃及 的时候， 亚玛力 在路上怎样对待你，
DEUT|25|18|在路上迎击你，趁你疲乏困倦时击杀所有在你后面软弱的人；并不敬畏上帝。
DEUT|25|19|所以，当耶和华－你的上帝使你不被四围一切仇敌扰乱，在耶和华－你上帝赐你为业的地上得享平静的时候，你要把 亚玛力 的名从天下涂去；你不可忘记这事。”
DEUT|26|1|“你进去得了耶和华－你上帝所赐你为业的地，并且居住在那里的时候，
DEUT|26|2|就要从耶和华－你上帝所赐你的地上，将收成的各种初熟土产取一些来，盛在筐子里，带到那里，耶和华－你上帝选择作为他名居所的地方，
DEUT|26|3|到当时的祭司那里，对他说：‘我今日向耶和华－你的上帝宣认，我已来到耶和华向我们列祖起誓要赐给我们的地。’
DEUT|26|4|祭司就从你手里把筐子接过来，供在耶和华－你上帝的祭坛前。
DEUT|26|5|你要在耶和华－你上帝面前告白说：‘我的祖先原是一个流亡的 亚兰 人，带着稀少的人丁下到 埃及 寄居。在那里，他却成了又大又强、人数众多的国。
DEUT|26|6|埃及 人恶待我们，迫害我们，将苦工加在我们身上。
DEUT|26|7|于是我们哀求耶和华我们列祖的上帝。耶和华听见我们的声音，看见我们所受的困苦、劳役和欺压，
DEUT|26|8|耶和华就用大能的手和伸出来的膀臂，以及大而可畏的事和神迹奇事，领我们出了 埃及 ，
DEUT|26|9|将我们领进这地方，把这流奶与蜜之地赐给我们。
DEUT|26|10|耶和华啊，看哪，现在我把你所赐我地上初熟的土产供上。’随后你要把筐子供在耶和华－你上帝面前，向耶和华－你的上帝下拜。
DEUT|26|11|你和 利未 人，以及在你中间寄居的，要因耶和华－你上帝所赐你和你家的一切福分欢乐。
DEUT|26|12|“每逢第三年，就是捐十分之一的那年，你从你一切土产中取了十分之一，要分给 利未 人、寄居的、孤儿和寡妇，使他们在你的城镇中可以吃得饱足。
DEUT|26|13|你又要在耶和华－你上帝面前说：‘我已将圣物从家里拿出来，给了 利未 人、寄居的、孤儿和寡妇，是遵照你吩咐我的一切命令。你的命令，我没有违背，也没有忘记。
DEUT|26|14|我守丧的时候，没有吃这圣物，不洁净的时候，也没有拿出来，又没有把它献给死人。我听从了耶和华－我上帝的话，都照你一切所吩咐的做了。
DEUT|26|15|求你从天上，从你的圣所垂看，赐福给你的百姓 以色列 和你向我们列祖起誓所赐给我们的这片土地，就是流奶与蜜之地。’”
DEUT|26|16|“耶和华－你的上帝今日吩咐你遵行这些律例典章，所以你要尽心尽性谨守遵行。
DEUT|26|17|你今日宣认耶和华为你的上帝，承诺遵行他的道，谨守他的律例、诫命、典章，听从他的话。
DEUT|26|18|耶和华今日照他所应许你的，也认你为他宝贵的子民，叫你谨守他的一切诫命，
DEUT|26|19|要使你得称赞、美名、尊荣，超乎他所造的万国之上，并且照他所应许的，使你归耶和华－你的上帝为神圣的子民。”
DEUT|27|1|摩西 和 以色列 的众长老吩咐百姓说：“你们要遵守我今日所吩咐的一切诫命。
DEUT|27|2|你们过了 约旦河 ，到耶和华－你上帝所赐给你的地，当日要竖立几块大石头，涂上石灰。
DEUT|27|3|当你过了河，进入耶和华－你上帝所赐给你流奶与蜜之地，正如耶和华－你列祖的上帝所应许你的，你要把这律法的一切话写在石头上。
DEUT|27|4|你们过了 约旦河 ，就要在 基利心山 上照我今日所吩咐的，把这些石头竖立起来，涂上石灰。
DEUT|27|5|你在那里要为耶和华－你的上帝筑一座石坛，却不可动用铁器在石头上。
DEUT|27|6|要用没有凿过的石头筑耶和华－你上帝的坛，在坛上将燔祭献给耶和华－你的上帝，
DEUT|27|7|又要献平安祭，在那里吃，在耶和华－你的上帝面前欢乐。
DEUT|27|8|你要将这律法的一切话清楚地写在石头上。”
DEUT|27|9|摩西 和 利未 家的祭司吩咐 以色列 众人说：“ 以色列 啊，你要静默倾听！你今日已成为耶和华－你上帝的子民了。
DEUT|27|10|你要听从耶和华－你上帝的话，遵行他的诫命律例，就是我今日所吩咐你的。”
DEUT|27|11|当日， 摩西 吩咐百姓说：
DEUT|27|12|“你们过了 约旦河 ， 西缅 、 利未 、 犹大 、 以萨迦 、 约瑟 和 便雅悯 等支派的人要站在 基利心山 上为百姓祝福。
DEUT|27|13|吕便 、 迦得 、 亚设 、 西布伦 、 但 和 拿弗他利 等支派的人要站在 以巴路山 上宣布诅咒。
DEUT|27|14|利未 人要大声对 以色列 众人说：
DEUT|27|15|“‘凡制造耶和华所憎恶的偶像，无论是雕刻的，是铸造的，就是工匠用手造的，或暗中设置的，这人必受诅咒！’众百姓要回应说：‘阿们！’
DEUT|27|16|“‘轻慢父母的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|17|“‘挪移邻舍地界的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|18|“‘引领瞎子走错路的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|19|“‘对寄居的、孤儿和寡妇屈枉正直的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|20|“‘与继母同寝的，必受诅咒！因为他掀开父亲衣服的下边。’众百姓要说：‘阿们！’
DEUT|27|21|“‘与兽交合的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|22|“‘与同父异母，或同母异父的姊妹同寝的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|23|“‘与岳母同寝的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|24|“‘暗中击杀邻舍的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|25|“‘受贿赂击杀人而流无辜之血的，必受诅咒！’众百姓要说：‘阿们！’
DEUT|27|26|“‘不坚守遵行这律法之话的，必受诅咒！’众百姓要说：‘阿们！’”
DEUT|28|1|“你若留心听从耶和华－你上帝的话，谨守遵行他的一切诫命，就是我今日所吩咐你的，他必使你超乎地上的万国之上。
DEUT|28|2|你若听从耶和华－你上帝的话，这一切的福气必临到你身上，追随你：
DEUT|28|3|你在城里必蒙福，在田间也必蒙福。
DEUT|28|4|你身所生的，你地所产的，你牲畜所生的，牛犊、羔羊，都必蒙福。
DEUT|28|5|你的筐子和你的揉面盆都必蒙福。
DEUT|28|6|你出也蒙福，入也蒙福。
DEUT|28|7|“耶和华必使那起来攻击你的仇敌在你面前溃败。他们从一条路来攻击你，必在你面前从七条路逃跑。
DEUT|28|8|在你仓房里，以及你手所做的一切，耶和华必发令赐福给你。耶和华－你上帝也必在所赐你的地上赐福给你。
DEUT|28|9|你若谨守耶和华－你上帝的诫命，遵行他的道，他必照他向你所起的誓立你为自己神圣的子民。
DEUT|28|10|地上的万民见你归在耶和华的名下，就必惧怕你。
DEUT|28|11|在耶和华向你列祖起誓应许赐你的土地上，他必使你身所生的，牲畜所生的，地所产的，都丰富有余。
DEUT|28|12|耶和华必为你敞开天上的宝库，按时降雨在你的地上。他必赐福你手里所做的一切。你必借给许多国家，却不必去借贷。
DEUT|28|13|你若听从耶和华－你上帝的诫命，就是我今日所吩咐你的，谨守遵行，耶和华就必使你作首不作尾，居上不居下，
DEUT|28|14|只要你不偏左右，不背离我今日所吩咐你的一切话，也不随从别神，事奉它们。”
DEUT|28|15|“你若不听从耶和华－你上帝的话，不谨守遵行他的一切诫命律例，就是我今日所吩咐你的，这一切的诅咒必临到你身上，追随你：
DEUT|28|16|你在城里必受诅咒，在田间也必受诅咒。
DEUT|28|17|你的筐子和你的揉面盆都必受诅咒。
DEUT|28|18|你身所生的，你地所产的，以及牛犊、羔羊，都必受诅咒。
DEUT|28|19|你出也受诅咒，入也受诅咒。
DEUT|28|20|耶和华因你作恶离弃他，必在你手里所做的一切，使诅咒、困扰、责罚临到你，直到你被除灭，直到你迅速灭亡。
DEUT|28|21|耶和华必使瘟疫紧贴着你，直到他把你从所进去得为业的地上灭绝。
DEUT|28|22|耶和华要用痨病、热病、发炎、高烧、刀剑 、焚风 和霉烂攻击你；这些要追赶你，直到你灭亡。
DEUT|28|23|你头上的天要变成铜，下面的地要化为铁。
DEUT|28|24|耶和华要使那降在你地上的雨变为灰尘，尘土从天落在你身上，直到你被除灭。
DEUT|28|25|“耶和华必使你在仇敌面前溃败。你从一条路去攻击他们，必从七条路逃跑。地上万国必因你而惊骇。
DEUT|28|26|你的尸首必给空中的飞鸟和地上的走兽作食物，却无人哄赶。
DEUT|28|27|耶和华必用 埃及 人的疮、溃疡、癣和疥攻击你，使你不得医治。
DEUT|28|28|耶和华必用癫狂、眼瞎、心惊攻击你。
DEUT|28|29|你必在午间摸索，好像盲人在黑暗中摸索。你的道路必不亨通，天天受人欺压、抢夺，无人搭救。
DEUT|28|30|你聘了妻子，别人必与她同寝；你建了房屋，却不得住在其内；你栽植了葡萄园，却不得享用所结的果子。
DEUT|28|31|你的牛在你眼前宰了，你吃不到它的肉；你的驴在你眼前被人抢夺，却讨不回来；你的羊被敌人拿走，无人帮助你。
DEUT|28|32|你的儿女被交给别国的民；你的眼目终日切望，甚至失明，你的手却无能为力。
DEUT|28|33|你地所产的和你劳力所得的，必被你所不认识的百姓吃尽。你天天只被欺负，受压制，
DEUT|28|34|甚至你因眼中所见的景象而疯狂。
DEUT|28|35|耶和华必攻击你，使你膝上腿上，从脚掌到头顶，都长满了毒疮，无法医治。
DEUT|28|36|“耶和华必将你和你所立统治你的王，领到你和你列祖不认识的国去；在那里你必事奉别神，就是木头和石头。
DEUT|28|37|你在耶和华赶你到的万民中，要令人惊骇，成为笑柄，被人讥诮。
DEUT|28|38|你撒在田里的种子虽多，收的却少，因为蝗虫把它吃光了。
DEUT|28|39|你栽植修整葡萄园，却没有酒喝，也不得储存，因为虫子把它吃了。
DEUT|28|40|你全境有橄榄树，却得不到油抹身，因为你的橄榄都掉光了。
DEUT|28|41|你生儿育女，却不属于你，因为他们必被掳去。
DEUT|28|42|你所有的树木和你地里的出产必被蝗虫吃尽了。
DEUT|28|43|在你中间寄居的必上升高过你，高而又高；你必下降，低而又低。
DEUT|28|44|他必借给你，你却不能借给他；他必作首，你必作尾。
DEUT|28|45|这一切的诅咒必临到你，追赶你，赶上你，直到把你除灭，因为你不听从耶和华－你上帝的话，不遵守他吩咐的诫命律例。
DEUT|28|46|这些诅咒必在你和你后裔身上成为神迹奇事，直到永远！
DEUT|28|47|因为你富裕的时候，不以欢喜快乐的心事奉耶和华－你的上帝，
DEUT|28|48|所以你必在饥饿、干渴、赤身、缺乏中事奉仇敌，那是耶和华派来攻击你的。他必把铁轭加在你的颈项上，直到把你除灭。
DEUT|28|49|耶和华要从远方、地极之处带一国来，如鹰飞来攻击你；这国的语言，你听不懂。
DEUT|28|50|这国的人面貌凶恶，不给长者面子，也不恩待年轻人。
DEUT|28|51|他们必吃你牲畜所生的和你土地所产的，直到你被除灭。你的五谷、新酒和新的油，以及牛犊、羔羊，他都不给你留下，直到使你灭亡。
DEUT|28|52|他们必在你的各城围困你，直到你在全地所倚靠、高大坚固的城墙都倒塌。他们必在耶和华－你上帝所赐给你全地的各城围困你。
DEUT|28|53|你在仇敌围困的窘迫中，必吃你本身所生的，就是耶和华－你上帝所赐给你的儿女之肉。
DEUT|28|54|你中间，连那温和文雅的人都必冷眼恶待自己的兄弟和怀中的妻子，以及他所剩下其余的儿女，
DEUT|28|55|不把所吃儿女的肉分一点给他们任何一个人，因为在被仇敌围困、陷入窘迫的各城中，他已经一无所剩了。
DEUT|28|56|你中间柔顺娇嫩的妇人，甚至因柔顺娇嫩脚不肯踏地的妇人，也必冷眼恶待她怀中的丈夫和自己的儿女。
DEUT|28|57|在被仇敌围困、陷入窘迫的城镇中，她因缺乏一切，就要暗中把从她两腿中间出来的胞衣和所生下的儿女吃了。
DEUT|28|58|“这书上所写律法的一切话，是叫你敬畏耶和华－你上帝尊荣可畏的名，你若不谨守遵行，
DEUT|28|59|耶和华就必将奇异的灾害，就是严重持久的灾害和长期难治的疾病，加在你和你后裔的身上。
DEUT|28|60|他必使你所畏惧、 埃及 一切的疾病临到你，紧贴着你，
DEUT|28|61|没有写在这律法书上的各样疾病、灾害，耶和华也必降在你身上，直到你被除灭。
DEUT|28|62|你们虽然曾像天上的星那样多，却因不听从耶和华－你上帝的话，所剩的人丁就稀少了。
DEUT|28|63|耶和华先前怎样喜爱善待你们，使你们增多，耶和华也要照样喜爱消灭你们，使你们灭绝。你们必从所要进去得为业的地上被拔除。
DEUT|28|64|耶和华必把你们分散在万民中，从地的这边到地的另一边，在那里你必事奉你和你列祖不认识的神明，就是木头和石头。
DEUT|28|65|在那些国中，你必得不到安宁，脚掌也没有安歇之处；耶和华却要使你在那里心中发颤，眼目失明，精神沮丧。
DEUT|28|66|你的一生悬空不安；你昼夜恐惧，生命没有保障。
DEUT|28|67|你因心中的恐惧，眼睛所见的景象，早晨必说：‘但愿现在是晚上！’晚上必说：‘但愿现在是早晨！’
DEUT|28|68|耶和华要用船把你送回 埃及 去，走那我曾告诉你不再看见的路；在那里你们必卖身给你的仇敌作奴婢，却没有人要买。”
DEUT|29|1|耶和华在 何烈山 与 以色列 人立约以外，这是耶和华在 摩押 地吩咐 摩西 与 以色列 人立约的话。
DEUT|29|2|摩西 召全 以色列 来，对他们说：“耶和华在 埃及 地，在你们眼前向法老和他众臣仆，以及他的全地所做的一切事，你们都看见了，
DEUT|29|3|就是你亲眼看见的大考验，那些神迹和大奇事。
DEUT|29|4|但耶和华到今日还没有使你们心能明白，眼能看见，耳能听见。
DEUT|29|5|我领你们在旷野四十年，你们身上的衣服没有穿破，脚上的鞋也没有穿坏；
DEUT|29|6|你们没有吃饼，也没有喝清酒烈酒，好让你们知道‘我─耶和华是你们的上帝’。
DEUT|29|7|你们来到这地方， 希实本 王 西宏 和 巴珊 王 噩 出来迎击我们，与我们交战，我们击败了他们，
DEUT|29|8|取了他们的地，给 吕便 支派、 迦得 支派和 玛拿西 半支派为业。
DEUT|29|9|所以你们要谨守这约的话，遵行它们，好使你们在一切所做的事上亨通。
DEUT|29|10|“今日你们全都要站在耶和华－你们的上帝面前，就是各领袖、族长 、长老、官长、 以色列 所有的男子、
DEUT|29|11|你们的妻子儿女、你营中寄居的，从为你砍柴到为你挑水的人，
DEUT|29|12|为要使你进入耶和华－你上帝的约，就是耶和华－你上帝今日向你起誓所立的；
DEUT|29|13|这样，他今日要立你作他的子民，他作你的上帝，是照他向你所应许的，又照他向你列祖 亚伯拉罕 、 以撒 、 雅各 所起的誓。
DEUT|29|14|我不单单与你们立这约，起这誓，
DEUT|29|15|就是今日与我们一同站在耶和华－我们上帝面前的，而且也包括今日不在我们这里的人。
DEUT|29|16|“你们知道，我们曾住过 埃及 地，也经过列国，从他们中间穿越。
DEUT|29|17|你们也见过他们的可憎之物，他们木、石、金、银的偶像。
DEUT|29|18|惟恐你们中间有人，或男或女，或宗族或支派，今日心里偏离耶和华－我们的上帝，去事奉那些国的神明，又怕你们中间有根长出苦菜和茵蔯来。
DEUT|29|19|这样的人听见这诅咒的话，心里还庆幸，说：‘我虽然随着顽固的心行事，却还是平安无事。’以致有水的和无水的都消灭了。
DEUT|29|20|耶和华必不愿饶恕他；耶和华的怒气与妒忌必向他如烟冒出，将这书上所写的一切诅咒都加在他身上，耶和华也要从天下涂去他的名。
DEUT|29|21|耶和华又必照着写在律法书上，约中的一切诅咒，将他从 以色列 众支派中分别出来，使他遭受祸害。
DEUT|29|22|你们的后代，就是接续你们兴起的子孙，和远方来的外邦人，看见这地的灾祸，以及耶和华所降于这地的疾病，
DEUT|29|23|遍地都被硫磺和盐所侵蚀，不能耕种，没有出产，连草都长不出来，好像耶和华在怒气和愤怒中所倾覆的 所多玛 、 蛾摩拉 、 押玛 、 洗扁 一样，
DEUT|29|24|万国必说：‘耶和华为什么向此地这样做呢？为什么要大发烈怒呢？’
DEUT|29|25|人必说：‘这是因为这地的人离弃了耶和华─他们列祖的上帝领他们出 埃及 地的时候与他们所立的约，
DEUT|29|26|去事奉别神，敬拜他们所不认识的神明，这是耶和华未曾允许的。
DEUT|29|27|所以耶和华的怒气向这地发作，将这书上所写的一切诅咒都降在这地上。
DEUT|29|28|耶和华在怒气、愤怒、大恼恨中将他们从本地拔出来，扔到别的地上，像今日一样。’
DEUT|29|29|“隐秘的事是属耶和华─我们上帝的，但明显的事是永远属我们和我们子孙的，为要叫我们遵行这律法上的一切话。”
DEUT|30|1|“当这一切的事，就是我摆在你面前的祝福和诅咒临到你的时候，你在耶和华－你上帝赶逐你去的万国中，心里回想这些事，
DEUT|30|2|你和你的子孙若尽心尽性归向耶和华－你的上帝，照我今日一切所吩咐你的，听从他的话，
DEUT|30|3|耶和华－你的上帝就必怜悯你，使你这被掳的子民归回。耶和华－你的上帝必转回，从分散你到的万民中把你召集回来。
DEUT|30|4|你就是被赶逐到天涯，耶和华－你的上帝也必从那里召集你，从那里领你回来。
DEUT|30|5|耶和华－你的上帝必领你进入你列祖所得的地，你必得着这地为业。他必善待你，使你增多，胜过你的列祖。
DEUT|30|6|耶和华－你的上帝要使你的心和你后裔的心受割礼，好叫你尽心尽性爱耶和华－你的上帝，使你可以存活。
DEUT|30|7|耶和华－你的上帝必将这一切诅咒加在你仇敌和恨恶你、迫害你的人身上。
DEUT|30|8|你必回转，听从耶和华的话，遵行他的一切诫命，就是我今日所吩咐你的。
DEUT|30|9|耶和华－你的上帝必使你手里所做的一切，以及你身所生的，牲畜所生的，土地所产的都丰富有余，而且顺利；耶和华必再喜爱善待你，正如他喜爱你的列祖一样，
DEUT|30|10|只要你听从耶和华－你上帝的话，谨守这律法书上所写的诫命律例，尽心尽性归向耶和华－你的上帝。”
DEUT|30|11|“我今日所吩咐你的诫命，对你并不困难，也不太远；
DEUT|30|12|不是在天上，使你说：‘谁为我们上天去取来给我们，使我们听了可以遵行呢？’
DEUT|30|13|也不是在海的那边，使你说：‘谁为我们渡海到另一边，去取来给我们，使我们听了可以遵行呢？’
DEUT|30|14|因这话离你很近，就在你口中，在你心里，使你可以遵行。
DEUT|30|15|“看，我今日将生死祸福摆在你面前。
DEUT|30|16|我今日所吩咐你的 ，就是要爱耶和华－你的上帝，遵行他的道，谨守他的诫命、律例、典章，使你可以存活，增多，而且耶和华－你的上帝必在你所要进去得为业的地上赐福给你。
DEUT|30|17|倘若你的心偏离，不肯听从，却被引诱去敬拜别神，事奉它们，
DEUT|30|18|我今日向你们申明，你们必定灭亡；在你过 约旦河 进去得为业的地上，你的日子必不长久。
DEUT|30|19|我今日呼天唤地向你作见证：我已经将生与死，祝福与诅咒，摆在你面前。所以你要拣选生命，好使你和你的后裔都得存活。
DEUT|30|20|要爱耶和华－你的上帝，听从他的话，紧紧跟随他，因为他是你的生命，必使你的日子得以长久，可以在耶和华向你列祖 亚伯拉罕 、 以撒 、 雅各 起誓要给他们的地上居住。”
DEUT|31|1|摩西 去把这些话吩咐 以色列 众人 ，
DEUT|31|2|对他们说：“我已经一百二十岁了，现在不能照常出入。耶和华曾对我说：‘你不得过这 约旦河 。’
DEUT|31|3|耶和华－你的上帝必在你面前过河，把这些国从你面前除灭，你就必得他们的地。 约书亚 要在你面前过河，是照耶和华所吩咐的。
DEUT|31|4|耶和华必对待他们，如同从前待他所除灭的 亚摩利 人的王 西宏 与 噩 ，以及他们的国一样。
DEUT|31|5|耶和华必将他们交在你们面前，你们要照我所吩咐的一切命令待他们。
DEUT|31|6|你们当刚强壮胆，不要害怕，也不要畏惧他们，因为耶和华－你的上帝必与你同去；他必不撇下你，也不丢弃你。”
DEUT|31|7|摩西 召了 约书亚 来，在 以色列 众人眼前对他说：“你当刚强壮胆！因为你要和这百姓一同进入 耶和华向他们列祖起誓要给他们的地，你也要使他们承受那地为业。
DEUT|31|8|耶和华必在你前面行，他必亲自与你同在，必不撇下你，也不丢弃你。你不要惧怕，也不要惊惶。”
DEUT|31|9|摩西 写下这律法，交给抬耶和华约柜的 利未 人祭司和 以色列 的众长老。
DEUT|31|10|摩西 吩咐他们说：“每逢七年的最后一年，就是定期的豁免年，在住棚节的时候，
DEUT|31|11|当 以色列 众人来到耶和华－你上帝所选择的地方朝见他的时候，你要在 以色列 众人面前念这律法给他们听。
DEUT|31|12|要召集百姓，男人、女人、孩子，和在你城里寄居的，叫他们都得以听见，好学习敬畏耶和华－你们的上帝，谨守遵行这律法的一切话。
DEUT|31|13|他们的儿女，就是那未曾认识的，也可以听，学习敬畏耶和华－你们的上帝；你们一生的日子，在你们过 约旦河 得为业的地上，都要这样做。”
DEUT|31|14|耶和华对 摩西 说：“看哪，你的死期已近了。要召 约书亚 来，和你一起站在会幕里，我好吩咐他。”于是 摩西 和 约书亚 去站在会幕里。
DEUT|31|15|耶和华在会幕里，在云柱中显现，云柱停在会幕门口的上面。
DEUT|31|16|耶和华对 摩西 说：“看哪，你必和你的祖先同睡。这百姓要起来，在他们所要去的地上，在那地的人中，随从外邦的神明行淫，离弃我，违背我与他们所立的约。
DEUT|31|17|那时，我的怒气必向他们发作，我必离弃他们，转脸不顾他们，以致他们被吞灭，并有许多的祸患灾难临到他们。在那日，人必说：‘这些祸患临到我，岂不是因为我的上帝不在我中间吗？’
DEUT|31|18|在那日，因人偏向别神所行的一切恶事，我必定转脸不顾。
DEUT|31|19|现在你们要写下这首歌，教导 以色列 人，放在他们口中，使这首歌成为我指责 以色列 人的见证。
DEUT|31|20|因为我将他们领进我向他们列祖起誓应许那流奶与蜜之地，他们在那里吃得饱足，长得肥胖，就偏向别神，事奉它们，藐视我，背弃我的约。
DEUT|31|21|当许多祸患灾难临到他们的时候，这首歌必在他们面前作见证，因为他们后裔的口必吟诵不忘。我未领他们到我所起誓应许之地以先，他们所怀的意念我都知道了。”
DEUT|31|22|当日 摩西 就写了一首歌，教导 以色列 人。
DEUT|31|23|耶和华吩咐 嫩 的儿子 约书亚 说：“你当刚强壮胆，因为你必领 以色列 人进入我所起誓应许他们的地，我必与你同在。”
DEUT|31|24|当 摩西 把这律法的话写完在书上，到完成的时候，
DEUT|31|25|摩西 吩咐抬耶和华约柜的 利未 人说：
DEUT|31|26|“把这律法书拿来，放在耶和华－你们上帝的约柜旁，可以在那里作指责你们的见证。
DEUT|31|27|因为我知道你们是悖逆的，是硬着颈项的。看哪，我今日还活着与你们同在，你们尚且悖逆耶和华，何况我死后呢？
DEUT|31|28|你们要召集你们支派的众长老和官长到我这里来，我好把这些话说给他们听，并且呼唤天地见证他们的不是。
DEUT|31|29|我知道我死后你们必全然败坏，偏离我所吩咐你们的道。日后必有祸患临到你们，因为你们做了耶和华眼中看为恶的事，以你们手中所做的惹他发怒。”
DEUT|31|30|摩西 把这首歌的话，从头到尾吟诵给 以色列 全会众听。
DEUT|32|1|“诸天哪，要侧耳听我说话； 愿地聆听我口中的言语。
DEUT|32|2|我的教导要淋漓如雨， 我的言语要滴落如露， 如细雨降在嫩草上， 如甘霖降在蔬菜中。
DEUT|32|3|因为我要宣扬耶和华的名， 你们要把伟大归给我们的上帝。
DEUT|32|4|“他是磐石，他的作为完全， 他一切所行的都公平； 他是信实无伪的上帝， 又公义，又正直。
DEUT|32|5|这乖僻弯曲的世代 向他行了败坏的事； 因着他们的弊病， 不再是他的儿女。
DEUT|32|6|愚昧无知的百姓啊， 你们这样报答耶和华吗？ 他岂不是你的父，创造了你吗？ 他造了你，坚立你。
DEUT|32|7|你当回想上古之日， 思念历代之年； 问你的父亲，他必告诉你； 问你的长者，他必向你述说。
DEUT|32|8|至高者将地业赐给列国， 将世人分开， 他按照神明 的数目， 为万民划定疆界。
DEUT|32|9|因为耶和华的份是他的百姓， 他的产业就是 雅各 。
DEUT|32|10|“耶和华在旷野之地， 在空旷，野兽吼叫之荒地遇见他， 就环绕他，看顾他， 保护他，如同保护眼中的瞳人。
DEUT|32|11|鹰怎样搅动巢窝， 在雏鹰上面飞翔， 展开双翅接住雏鹰， 背在两翼之上，
DEUT|32|12|耶和华也照样独自引导他， 并无外邦神明与他同在。
DEUT|32|13|耶和华使他驰骋在地的高处， 他吃田间的出产； 耶和华使他从岩石中吃蜜， 从坚石中吸油，
DEUT|32|14|也吃牛的乳酪、羊的奶、 羔羊的脂肪， 巴珊 所出的公绵羊和山羊， 和上好的麦子。 你要喝葡萄汁酿的美酒。
DEUT|32|15|“ 耶书仑 渐渐肥胖，能踼跳。 你长得肥胖，粗壮，丰润。 他离弃造他的上帝， 轻看救他的磐石。
DEUT|32|16|他们用外邦神明惹上帝妒忌， 以可憎之物惹他发怒。
DEUT|32|17|他们祭祀鬼魔，而非上帝， 是他们不认识的神明， 是近来新兴的， 是你们列祖所不畏惧的。
DEUT|32|18|你轻忽生你的磐石， 忘记生产你的上帝。
DEUT|32|19|“耶和华看见了， 因他儿女惹动他就抛弃他们，
DEUT|32|20|说：‘我要转脸离开他们， 看他们的结局如何。 他们是极乖谬的世代， 是不忠实的儿女。
DEUT|32|21|他们以那不是上帝的激起我妒忌， 以虚无的神明 惹我发怒。 我也要以不成国的激起你们嫉妒， 我要以愚顽的国惹起你们发怒。
DEUT|32|22|因为我的怒火焚烧， 直烧到极深的阴间， 吞噬地和地的出产， 连山的根基也烧着了。
DEUT|32|23|“‘我要把祸患堆在他们身上， 我用尽我的箭射向他们：
DEUT|32|24|饿死人的饥荒、 灼人的热症、 痛苦的灾害。 我要叫野兽用牙齿咬他们， 叫土中爬行的用毒液害他们。
DEUT|32|25|外有刀剑使人丧亡， 内有惊恐， 少男少女是如此， 吃奶的、白发的也是如此。
DEUT|32|26|我曾说，我要粉碎他们， 使他们的名 从人间消失。
DEUT|32|27|惟恐仇敌挑衅， 他们的敌人误解， 说，我们的手得胜了， 这一切并非耶和华做的。’
DEUT|32|28|“因为他们是缺乏智谋的国家， 他们里面毫无聪明。
DEUT|32|29|惟愿他们有智慧，能明白这事， 他们就会想到自己的结局。
DEUT|32|30|若非他们的磐石卖了他们， 若非耶和华交出他们， 一人岂能追赶千人， 二人焉能使万人逃跑呢？
DEUT|32|31|甚至我们的仇敌都承认， 他们的磐石不如我们的磐石。
DEUT|32|32|他们的葡萄树是 所多玛 的葡萄树， 是 蛾摩拉 田园所长的； 他们的葡萄是毒葡萄， 整串都是苦的。
DEUT|32|33|他们的酒是大蛇的毒液， 是毒蛇剧烈的毒汁。
DEUT|32|34|“这岂不都存放在我这里， 封存在我库房中吗？
DEUT|32|35|伸冤报应在我 ， 到了时候他们会失脚。 因为他们遭难的日子近了， 他们的厄运快要临到。
DEUT|32|36|耶和华见他的百姓毫无能力， 无论是为奴的、自由的，都没有存留， 就必为他们伸冤， 为自己的仆人发怜悯。
DEUT|32|37|他必说：‘他们的神明， 他们所投靠的磐石，在哪里呢？
DEUT|32|38|吃了他们祭牲脂肪的， 喝了他们浇酒祭之酒的， 叫那些神明站出来帮助你们， 作为你们的保障吧！
DEUT|32|39|“‘如今，看！我，惟有我是上帝 ； 我以外并无别神。 我使人死，我使人活； 我击伤人，也医治人， 没有人能从我手中救出来。
DEUT|32|40|我向天举手， 我凭我的永生起誓说：
DEUT|32|41|我若磨我闪亮的刀， 我的手掌握审判权， 就必报复我的敌人， 报应那些恨我的人。
DEUT|32|42|我要使我的箭饮血而醉， 就是被杀被掳之人的血； 我的刀也要吃肉， 就是仇敌披发头颅 的肉。’
DEUT|32|43|“列国啊，当与耶和华的子民一同欢呼 ； 因为他要为他仆人 所流的血伸冤， 报应他的敌人 ， 救赎他的土地和他的子民 。”
DEUT|32|44|摩西 和 嫩 的儿子 约书亚 前来把这首歌的一切话吟诵给百姓听。
DEUT|32|45|摩西 向 以色列 众人吟诵完了这一切话，
DEUT|32|46|对他们说：“我今日以这一切话警戒你们，你们都要记在心中，要吩咐你们的子孙谨守遵行这律法上一切的话。
DEUT|32|47|因为这不是与你们无关的空话，而是你们的生命；因遵行这话，你们的日子必在你们过 约旦河 得为业的地上得以长久。”
DEUT|32|48|就在那日，耶和华吩咐 摩西 说：
DEUT|32|49|“你上 摩押 地的 亚巴琳山脉 ，到面对 耶利哥 的 尼波山 去，看我所要赐给 以色列 人为业的 迦南 地。
DEUT|32|50|你必死在你所登的山上，归到你祖先 那里，像你哥哥 亚伦 死在 何珥山 上，归到他祖先 那里一样。
DEUT|32|51|因为你们在 以色列 人中得罪了我，在 寻 的旷野， 加低斯 的 米利巴 水那里，在 以色列 人中没有尊我为圣。
DEUT|32|52|我所赐给 以色列 人的地，你只可从对面观看，却不得进到那里去。”
DEUT|33|1|这是神人 摩西 未死以前为 以色列 人的祝福。
DEUT|33|2|他说： “耶和华从 西奈 来， 从 西珥 向他们显现， 从 巴兰山 发出光辉； 从万万圣者中来临 ， 从他右手向他们发出烈火的律法 。
DEUT|33|3|他实在疼爱万民。 他的众圣徒都在你手中， 他们坐在你的脚下， 领受你的言语。”
DEUT|33|4|摩西 将律法传给我们， 作为 雅各 会众的产业。
DEUT|33|5|“耶和华 在 耶书仑 作王； 百姓的众领袖和 以色列 各支派一同欢聚。
DEUT|33|6|愿 吕便 存活，不致死亡， 虽然他的人丁稀少。
DEUT|33|7|关于 犹大 ，他这么说： ‘耶和华啊，求你垂听 犹大 的声音， 引导他归回他的百姓中。 他曾用手为自己争战， 你必帮助他攻击敌人。’
DEUT|33|8|关于 利未 ，他说： ‘愿你的土明和乌陵都在你的虔诚人那里 。 你在 玛撒 曾考验他， 在 米利巴 水与他争论。
DEUT|33|9|关于自己的父母，他说：我未曾关注。 他的弟兄，他不承认， 他的儿女，他也不认识， 因为 利未 人遵行你的话， 谨守你的约。
DEUT|33|10|他们将你的典章教导 雅各 ， 将你的律法教导 以色列 。 他们奉上香让你闻， 把全牲的燔祭献在你坛上。
DEUT|33|11|求耶和华赐福给他的财物 ， 悦纳他手里的工作。 求你刺透起来攻击他的人的腰， 使那些恨恶他的人不再起来。’
DEUT|33|12|关于 便雅悯 ，他说： ‘耶和华所亲爱的必同耶和华安然居住， 耶和华终日庇护他， 他也住在耶和华两肩之中 。’
DEUT|33|13|关于 约瑟 ，他说： ‘愿他的地蒙耶和华赐福， 得天上的甘露， 地下的泉源；
DEUT|33|14|得太阳下的美果， 月光中的佳谷；
DEUT|33|15|得古老山岳的至宝， 永恒山岭的宝物；
DEUT|33|16|得地的宝物和其中所充满的， 得住在荆棘中者的喜悦。 愿这些福都临到 约瑟 的头上， 临到那与兄弟有分别之人的头顶上。
DEUT|33|17|他是牛群中头生的， 大有威严； 他的双角是野牛的角， 用以抵触万民，直到地极。 这对角是 以法莲 的万万， 这对角是 玛拿西 的千千。’
DEUT|33|18|关于 西布伦 ，他说： ‘ 西布伦 哪，你出外可以欢喜。 以萨迦 啊，你在帐棚里可以快乐。
DEUT|33|19|他们要召集万民到山上， 在那里献公义的祭。 因为他们要吸取海里的财富， 沙中隐藏的珍宝。’
DEUT|33|20|关于 迦得 ，他说： ‘那使 迦得 扩张的，当受称颂！ 迦得 卧如母狮， 撕裂膀臂和头皮。
DEUT|33|21|他为自己看中了最好的， 因为那是为掌权者所存留的一份。 他与百姓的领袖同来 ， 执行耶和华的公义 和耶和华为 以色列 所立的典章。’
DEUT|33|22|关于 但 ，他说： ‘ 但 是小狮子， 从 巴珊 跳出来。’
DEUT|33|23|关于 拿弗他利 ，他说： ‘ 拿弗他利 啊，你享足恩宠， 满得耶和华的福， 可以得西方和南方为业。’
DEUT|33|24|关于 亚设 ，他说： ‘愿 亚设 在众子中蒙福 ， 愿他得他弟兄的喜悦， 可以把脚蘸在油中。
DEUT|33|25|你的门闩是铁的，是铜的。 只要你有多少日子，你就有多少力量 。’
DEUT|33|26|“ 耶书仑 哪，没有谁能比上帝！ 他腾云，大显威荣， 从天空来帮助你。
DEUT|33|27|亘古的上帝是避难所， 下面有永久的膀臂。 他从你面前赶走仇敌， 说：‘毁灭吧！’
DEUT|33|28|因此， 以色列 独自安然居住， 雅各 的泉源在五谷新酒之地， 他的天也滴下露水。
DEUT|33|29|以色列 啊，你有福了！ 蒙耶和华拯救的百姓啊，谁能像你？ 他是帮助你的盾牌， 是你威荣的刀剑。 你的仇敌要屈身就你； 你却要践踏他们的背脊 。”
DEUT|34|1|摩西 从 摩押 平原登上 尼波山 ，到了 耶利哥 对面的 毗斯迦山 顶。耶和华把全地指给他看：从 基列 到 但 ，
DEUT|34|2|拿弗他利 全地， 以法莲 、 玛拿西 的地， 犹大 全地直到西边的海，
DEUT|34|3|尼革夫 ，从棕树城 耶利哥 的平原到 琐珥 。
DEUT|34|4|耶和华对他说：“这就是我向 亚伯拉罕 、 以撒 、 雅各 起誓应许之地，说：‘我必将这地赐给你的后裔。’现在我使你亲眼看见了，你却不得过到那里去。”
DEUT|34|5|于是耶和华的仆人 摩西 死在 摩押 地那里，正如耶和华所说的。
DEUT|34|6|耶和华将他葬在 摩押 地， 伯．毗珥 对面的谷中，只是到今日，没有人知道他的坟墓。
DEUT|34|7|摩西 死的时候一百二十岁，眼目没有昏花，力量没有衰退。
DEUT|34|8|以色列 人在 摩押 平原为 摩西 哀哭了三十天，为 摩西 哀哭居丧的日期才结束。
DEUT|34|9|嫩 的儿子 约书亚 ，因为 摩西 曾为他按手，他就被智慧的灵充满。 以色列 人听从他，照着耶和华所吩咐 摩西 的去做。
DEUT|34|10|以后， 以色列 中再没有兴起一位先知像 摩西 的，他是耶和华面对面所认识的。
DEUT|34|11|耶和华差派他在 埃及 地，向法老和他的一切臣仆，以及他的全地，行了各样神迹奇事，
DEUT|34|12|又在 以色列 众人眼前显出大能的手，行了一切大而可畏的事。
JOSH|1|1|耶和华的仆人 摩西 死了以后，耶和华对 摩西 的助手 嫩 的儿子 约书亚 说：
JOSH|1|2|“我的仆人 摩西 死了。现在你要起来，和众百姓过这 约旦河 ，往我所要赐给 以色列 人的地去。
JOSH|1|3|凡你们脚掌所踏之地，我都照我所应许 摩西 的话赐给你们了。
JOSH|1|4|从旷野和这 黎巴嫩 ，直到 大河 ，就是 幼发拉底河 ， 赫 人的全地，又到 大海 日落的方向，都要作你们的疆土。
JOSH|1|5|你一生的日子，必无人能在你面前站立得住。我怎样与 摩西 同在，也必照样与你同在；我必不撇下你，也不丢弃你。
JOSH|1|6|你当刚强壮胆，因为你必使这百姓承受那地为业，就是我向他们列祖起誓要给他们的地。
JOSH|1|7|只要刚强，大大壮胆，谨守遵行我仆人 摩西 所吩咐你的一切律法，不可偏离左右，使你无论往哪里去， 都可以顺利。
JOSH|1|8|这律法书不可离开你的口，总要昼夜思想 ，好使你谨守遵行这书上所写的一切话。如此，你的道路就可以亨通，凡事顺利。
JOSH|1|9|我岂没有吩咐你吗？你当刚强壮胆，不要惧怕，也不要惊惶，因为你无论往哪里去，耶和华你的上帝必与你同在。”
JOSH|1|10|于是， 约书亚 吩咐百姓的官长说：
JOSH|1|11|“你们要走遍营中，吩咐百姓说：‘当预备食物， 因为三日之内你们要过这 约旦河 ，进去得耶和华－你们上帝赐给你们为业之地。’”
JOSH|1|12|约书亚 对 吕便 人、 迦得 人和 玛拿西 半支派的人说：
JOSH|1|13|“你们要记得耶和华的仆人 摩西 所吩咐你们的话说：‘耶和华－你们的上帝使你们得享安宁，必将这地赐给你们。’
JOSH|1|14|你们的妻子、孩子和牲畜可以留在 约旦河 东、 摩西 所给你们的地。但你们中间所有大能的勇士都要带着兵器，在你们的弟兄前面过去，你们要帮助他们。
JOSH|1|15|等到耶和华使你们的弟兄和你们一样得享平静，并且得着耶和华－你们上帝所赐他们为业之地的时候，你们才可以回到你们所得之地，承受为业，就是耶和华的仆人 摩西 在 约旦河 东、向日出的方向所给你们的地。”
JOSH|1|16|他们回答 约书亚 说：“凡你吩咐我们的，我们都必做；凡你差我们去的地方，我们都必去。
JOSH|1|17|我们在一切事上怎样听从 摩西 ，也必照样听从你。惟愿耶和华－你的上帝与你同在，像与 摩西 同在一样。
JOSH|1|18|无论什么人违背你的命令，不听从你所吩咐他的一切话，就必处死。你只要刚强壮胆！”
JOSH|2|1|嫩 的儿子 约书亚 从 什亭 暗中派两个人作探子，说：“你们去窥探那地和 耶利哥 。”于是二人去了，来到一个名叫 喇合 的妓女家里，在那里睡觉。
JOSH|2|2|有人告诉 耶利哥 王说：“看哪，今夜有 以色列 人到这里来窥探此地。”
JOSH|2|3|耶利哥 王派人到 喇合 那里， 说：“你要交出那来到你这里、进了你家的人，因为他们来是要窥探全地。”
JOSH|2|4|但女人已把二人藏起来，却说：“那两个人确实到我这里来过，他们从哪里来，我却不知道。
JOSH|2|5|天黑、要关城门的时候，他们就出去了。他们往哪里去我也不知道。你们赶快去追他们，就必追上。”
JOSH|2|6|其实，这女人已经领二人上了屋顶，把他们藏在她摆列在屋顶的的亚麻梗中。
JOSH|2|7|那些人就往 约旦河 的路上追赶他们，直到渡口。追赶他们的人一出去，城门就关了。
JOSH|2|8|二人还没有睡之前，女人就上屋顶，到他们那里，
JOSH|2|9|对他们说：“我知道耶和华已经把这地赐给你们了，并且我们也都惧怕你们。这地所有的居民在你们面前都融化了。
JOSH|2|10|因为我们听见你们出 埃及 的时候，耶和华怎样在你们前面使 红海 的水干了，并且你们怎样处置 约旦河 东的两个 亚摩利 王， 西宏 和 噩 ，把他们完全消灭。
JOSH|2|11|我们一听见就胆战心惊 ，人人因你们的缘故勇气全失。耶和华－你们的上帝是天上地下的上帝。
JOSH|2|12|现在我既然恩待你们，求你们指着耶和华向我起誓，你们也要恩待我的父家。请你们给我一个确实的凭据，
JOSH|2|13|要救活我的父母、兄弟、姊妹，和所有属他们的，拯救我们的性命脱离死亡。”
JOSH|2|14|那二人对她说：“我们愿意以性命来替你们死。你们若不泄漏我们这件事，当耶和华将这地赐给我们的时候，我们必以慈爱和诚信待你。”
JOSH|2|15|于是女人用绳子把二人从窗户缒下去，因为她的屋子是在城墙边上，她也住在城墙上。
JOSH|2|16|她对他们说：“你们暂且往山上去，免得追赶的人遇见你们。要在那里躲藏三天，等追赶的人回来，你们才可以走自己的路。”
JOSH|2|17|二人对她说：“你叫我们所起的誓与我们无关，
JOSH|2|18|除非，看哪，当我们来到这地的时候，你把这条朱红线绳子系在缒我们下去的窗户上，并要叫你的父母、兄弟和你父的全家都聚集在你家中。
JOSH|2|19|凡离开你家门往街上去的，他的血必归到自己头上，与我们无关；凡在你家里的，若有人下手害他，他的血就归到我们头上。
JOSH|2|20|你若泄漏我们这件事，你叫我们所起的誓 就与我们无关了。”
JOSH|2|21|女人说：“就照你们的话吧！”于是她送他们走了，就把朱红绳子系在窗户上。
JOSH|2|22|二人离开，到山上去，在那里停留三天，直等到追赶的人回去。追赶的人一路寻找，却找不着。
JOSH|2|23|二人回来，下了山，过了河，来到 嫩 的儿子 约书亚 那里，向他报告他们所遭遇的一切事。
JOSH|2|24|他们对 约书亚 说：“耶和华果然将那全地交在我们手中了，并且那地所有的居民在我们面前都融化了。”
JOSH|3|1|约书亚 清早起来，和 以色列 众人起行，离开 什亭 ，来到 约旦河 ，过河以前住在那里。
JOSH|3|2|过了三天，官长走遍营中，
JOSH|3|3|吩咐百姓说：“当你们看见 利未 家的祭司抬着耶和华－你们上帝的约柜的时候，你们就要起行离开所住的地方，跟着约柜走，
JOSH|3|4|使你们知道所当走的路，因为这条路是你们从来没有走过的。只是你们要与约柜相隔约二千肘，不可太靠近约柜。”
JOSH|3|5|约书亚 吩咐百姓说：“你们要使自己分别为圣，因为明天耶和华必在你们中间行奇事。”
JOSH|3|6|约书亚 对祭司说：“你们抬起约柜，在百姓的前面过去。”于是他们抬起约柜，走在百姓前面。
JOSH|3|7|耶和华对 约书亚 说：“从今日起，我必使你在 以色列 众人眼前被尊为大，使他们知道我怎样与 摩西 同在，也必照样与你同在。
JOSH|3|8|你要吩咐抬约柜的祭司说：‘你们到了 约旦河 的水边，要在 约旦河 中站着。’”
JOSH|3|9|约书亚 对 以色列 人说：“你们近前，到这里来，听耶和华－你们上帝的话。”
JOSH|3|10|约书亚 说：“你们因这事会知道永生的上帝在你们中间，他必从你们面前赶出 迦南 人、 赫 人、 希未 人、 比利洗 人、 革迦撒 人、 亚摩利 人、 耶布斯 人。
JOSH|3|11|看哪！全地之主的约柜必在你们的前面过去，到 约旦河 里。
JOSH|3|12|现在， 你们要从 以色列 支派中选出十二个人，每支派一人。
JOSH|3|13|当抬耶和华全地之主约柜的祭司，脚掌踏入 约旦河 水里的时候， 约旦河 的水，就是从上往下流的水，必然中断，竖立成垒。”
JOSH|3|14|百姓起行离开帐棚过 约旦河 的时候，抬约柜的祭司在百姓的前面。
JOSH|3|15|那时正是收割的日子， 约旦河 的水涨满两岸。抬约柜的人到了 约旦河 ，抬约柜的祭司脚一入水边，
JOSH|3|16|那从上往下流的水就在很远的地方，在 撒拉但 旁边的 亚当城 那里停住，竖立成垒；那往 亚拉巴海 ，就是 盐海 下流的水全然中断。于是，百姓在 耶利哥 的对面过了河。
JOSH|3|17|抬耶和华约柜的祭司在 约旦河 中的干地上稳稳站着， 以色列 众人都从干地上过去，直到全国都过了 约旦河 。
JOSH|4|1|当全国都过了 约旦河 ，耶和华对 约书亚 说：
JOSH|4|2|“你要从百姓中选出十二个人，每支派一人，
JOSH|4|3|吩咐他们说：‘你们从这里，从 约旦河 中祭司的脚稳稳站立的地方，取十二块石头 ，一起带过去，放在你们今夜住宿的地方。’”
JOSH|4|4|于是 约书亚 召集了他从 以色列 人中所选的十二个人，每支派一人。
JOSH|4|5|约书亚 对他们说：“你们要过去，到 约旦河 中，耶和华－你们上帝的约柜前面，按 以色列 人支派的数目，每人各取一块石头扛在肩上。
JOSH|4|6|这些石头在你们中间将成为记号。日后，你们的子孙问你们说：‘这些石头对你们有什么意思呢？’
JOSH|4|7|你们就对他们说：‘这是因为 约旦河 的水在耶和华的约柜前中断；约柜过 约旦河 的时候， 约旦河 的水就中断了。这些石头要作 以色列 人永远的纪念。’”
JOSH|4|8|以色列 人就照 约书亚 所吩咐的做了。他们按 以色列 人支派的数目，从 约旦河 中取了十二块石头，正如耶和华所吩咐 约书亚 的。他们把石头带过去，到他们所住宿的地方，就放在那里。
JOSH|4|9|约书亚 另外把十二块石头立在 约旦河 的中间，在抬约柜祭司的脚站立的地方；直到今日，石头还在那里。
JOSH|4|10|抬约柜的祭司站在 约旦河 的中间，直到耶和华命令 约书亚 告诉百姓的一切事办完为止，正如 摩西 所吩咐 约书亚 的一切话。 于是，百姓急速过了河。
JOSH|4|11|全体百姓都过了河之后，耶和华的约柜和祭司才过去，到百姓的前面。
JOSH|4|12|吕便 人、 迦得 人、 玛拿西 半支派的人都照 摩西 所吩咐他们的，带着兵器在 以色列 人的前面过去。
JOSH|4|13|约有四万带兵器的军队在耶和华面前过去，到 耶利哥 的平原，准备上阵。
JOSH|4|14|在那日，耶和华使 约书亚 在 以色列 众人眼前被尊为大。在他一生的年日中，百姓敬服他，像从前敬服 摩西 一样。
JOSH|4|15|耶和华对 约书亚 说：
JOSH|4|16|“你吩咐抬法柜的祭司从 约旦河 上来。”
JOSH|4|17|约书亚 就吩咐祭司说：“你们从 约旦河 上来。”
JOSH|4|18|抬耶和华约柜的祭司从 约旦河 中上来，脚掌一落干地， 约旦河 的水就流回原处，仍旧涨满两岸。
JOSH|4|19|正月初十，百姓从 约旦河 上来，就在 耶利哥 东边的 吉甲 安营。
JOSH|4|20|约书亚 把他们从 约旦河 取来的那十二块石头立在 吉甲 ，
JOSH|4|21|对 以色列 人说：“日后，你们的子孙问他们的父亲说：‘这些石头是什么意思呢？’
JOSH|4|22|你们就让你们的子孙知道，说：‘ 以色列 人曾走干地过这 约旦河 。’
JOSH|4|23|因为耶和华－你们的上帝在你们前面使 约旦河 的水干了，直到你们过来，就如耶和华－你们的上帝从前在我们前面使 红海 干了，直到我们过来一样，
JOSH|4|24|要使地上万民都知道，耶和华的手大有能力，也要使你们天天敬畏耶和华－你们的上帝。”
JOSH|5|1|约旦河 西 亚摩利 人的众王和靠海 迦南 人的众王，听见耶和华在 以色列 人前面使 约旦河 的水干了，直到他们过了河 ，众王因 以色列 人的缘故都胆战心惊，勇气全失。
JOSH|5|2|那时，耶和华对 约书亚 说：“你要造火石刀，第二次为 以色列 人行割礼。”
JOSH|5|3|约书亚 就造了火石刀，在 哈尔拉勒山 为 以色列 人行割礼。
JOSH|5|4|约书亚 行割礼的原因是这样：从 埃及 出来的众百姓，所有能打仗的男丁，出了 埃及 以后，都死在旷野的路上。
JOSH|5|5|这些从 埃及 出来的众百姓都受过割礼；但是那些出 埃及 以后，在旷野的路上所生的众百姓却没有受过割礼。
JOSH|5|6|以色列 人在旷野走了四十年，直到那从 埃及 出来，全国能打仗的人都消灭了，因为他们没有听从耶和华的话。耶和华曾向他们起誓，必不容许他们看见耶和华向他们列祖起誓要给我们的地，就是流奶与蜜之地。
JOSH|5|7|他们的子孙，就是耶和华兴起接续他们的，都没有受过割礼；因为在路上他们没有受割礼， 约书亚 就为他们行割礼。
JOSH|5|8|全国的人都受了割礼，留在营中自己的地方，直到痊愈。
JOSH|5|9|耶和华对 约书亚 说：“我今日将 埃及 的羞辱从你们身上除掉了。”因此，那地方名叫 吉甲 ，直到今日。
JOSH|5|10|以色列 人在 吉甲 安营。正月十四日晚上，他们在 耶利哥 的平原守逾越节。
JOSH|5|11|逾越节的第二日，他们吃了当地的出产，就在那一天，吃了无酵饼和烘过的谷物。
JOSH|5|12|他们吃了当地出产的第二日，吗哪就停止了。 以色列 人不再有吗哪了。那一年，他们就吃 迦南 地的出产。
JOSH|5|13|约书亚 靠近 耶利哥 的时候，举目观看，看哪，有一个人站在他对面，手里拿着拔出来的刀。 约书亚 到他那里，对他说：“你是属我们的，还是属我们敌人的呢？”
JOSH|5|14|他说：“不，我现在来是要作耶和华军队的元帅。” 约书亚 就脸伏于地下拜，说：“我主有什么话，请吩咐仆人吧！”
JOSH|5|15|耶和华军队的元帅对 约书亚 说：“把你脚上的鞋脱下来，因为你所站的地方是圣的。” 约书亚 就照着做了。
JOSH|6|1|耶利哥 的城门因 以色列 人的缘故，关得严紧，无人出入。
JOSH|6|2|耶和华对 约书亚 说：“看，我已经把 耶利哥城 和 耶利哥 王，以及大能的勇士，都交在你手中。
JOSH|6|3|你们要围绕这城，所有的士兵绕城一次，六日你都要这样做。
JOSH|6|4|七个祭司要拿七个羊角走在约柜前。到了第七日，你们要围绕这城七次，祭司也要吹角。
JOSH|6|5|羊角声拖长的时候，你们一听见角声，众百姓要大声呼喊，城墙就必倒塌，各人要往前直上。”
JOSH|6|6|嫩 的儿子 约书亚 召了祭司来，对他们说：“你们抬起约柜来，要有七个祭司拿七个羊角在耶和华的约柜前。”
JOSH|6|7|他又对百姓说：“你们向前去围绕那城，带兵器的要在耶和华的约柜前过去。”
JOSH|6|8|按照 约书亚 对百姓所说的，七个祭司拿了七个羊角在耶和华面前过去，他们吹着角，耶和华的约柜在他们后面跟着。
JOSH|6|9|带兵器的走在吹角的祭司前面，后队跟着约柜走，号角继续在吹。
JOSH|6|10|约书亚 吩咐百姓说：“你们不可呼喊，不可让人听见你们的声音，连一句话也不可出你们的口，直到我对你们说‘呼喊’的那日，你们才呼喊。”
JOSH|6|11|这样， 约书亚 使耶和华的约柜围绕那城，把城绕了一次。然后，众人回到营里，就在营里住宿。
JOSH|6|12|约书亚 清早起来，祭司又抬起耶和华的约柜。
JOSH|6|13|七个祭司拿七个羊角，走在耶和华的约柜前，他们吹着角；带兵器的走在他们前面，后队跟着耶和华的约柜走，号角继续在吹。
JOSH|6|14|第二日，他们再把城围绕一次，就回营里去。六日都是这样做。
JOSH|6|15|第七日清早黎明时，他们起来，以同样的方式围绕城七次；惟独这一日他们围绕城七次。
JOSH|6|16|到了第七次，祭司吹角的时候， 约书亚 对百姓说：“呼喊吧，因为耶和华已经把城交给你们了！
JOSH|6|17|这城和其中所有的都要永献给耶和华作当毁灭的，只有妓女 喇合 与她家中所有的可以存活，因为她隐藏了我们所派的使者。
JOSH|6|18|但你们务必谨慎，不可取那当灭的物，免得你们受诅咒，取了那当灭的物，使 以色列 全营成为诅咒而遭受灾祸。
JOSH|6|19|只有金子、银子和铜铁的器皿都要归耶和华为圣，放入耶和华的库房中。”
JOSH|6|20|于是百姓呼喊，祭司吹角。百姓一听见角声就大声呼喊，城墙随着倒塌。百姓上去进城，各人往前直上，把城夺取。
JOSH|6|21|他们把城中所有的，无论男女老少，牛羊和驴，都用刀杀尽。
JOSH|6|22|约书亚 对窥探这地的两个人说：“你们进那妓女的家，照你们向她所起的誓，将那女人和她所有的都从那里带出来。”
JOSH|6|23|两个作过探子的青年进去，把 喇合 与她的父母、兄弟，和她所有的带出来，他们把她所有的亲属都带出来，安置在 以色列 的营外。
JOSH|6|24|他们用火焚烧了那城和其中所有的，只有金子、银子和铜铁的器皿都放在耶和华殿的库房中。
JOSH|6|25|至于妓女 喇合 和她父家，以及她所有的， 约书亚 保存了他们的性命。她就住在 以色列 中，直到今日，因为她隐藏了 约书亚 派来窥探 耶利哥 的使者。
JOSH|6|26|当时， 约书亚 叫众人起誓说：“凡兴起重修这 耶利哥城 的，当在耶和华面前受诅咒。 他立根基的时候，必丧长子， 安城门的时候，必丧幼子。”
JOSH|6|27|耶和华与 约书亚 同在， 约书亚 的名声传遍全地。
JOSH|7|1|以色列 人在当灭之物上犯了罪。 犹大 支派中， 谢拉 的曾孙， 撒底 的孙子， 迦米 的儿子 亚干 取了当灭之物，耶和华的怒气就向 以色列 人发作。
JOSH|7|2|约书亚 从 耶利哥 派人往 伯特利 东边，靠近 伯．亚文 的 艾城 去，对他们说：“你们上去窥探那地。”那些人就上去窥探 艾城 。
JOSH|7|3|他们回到 约书亚 那里，对他说：“众百姓不必都上去，只要二、三千人上去就能攻取 艾城 ；不必劳动众百姓都上去，因为他们人少。”
JOSH|7|4|于是百姓中约有三千人上那里去，但他们竟在 艾城 的人面前逃跑。
JOSH|7|5|艾城 的人击杀他们约三十六人，从城门前追赶他们，直到 示巴琳 ，在下坡的地方击败他们。他们都胆战心惊，融化如水。
JOSH|7|6|约书亚 和 以色列 的长老就撕裂衣服，在耶和华的约柜前脸伏于地，直到晚上。他们把灰撒在头上。
JOSH|7|7|约书亚 说：“唉！主耶和华啊，你为什么领这百姓过 约旦河 ，把我们交在 亚摩利 人手中，使我们灭亡呢？我们不如住在 约旦河 的那边！
JOSH|7|8|主啊，求求你， 以色列 人既在仇敌面前转身逃跑，我还有什么可说的呢？
JOSH|7|9|迦南 人和这地所有的居民听见了就必围困我们，把我们的名从地上除去。那时，你为你至大的名要怎样做呢？”
JOSH|7|10|耶和华对 约书亚 说：“起来！你的脸为何这样俯伏呢？
JOSH|7|11|以色列 犯了罪，又违背了我所吩咐他们的约，又取了当灭之物。他们又偷窃，又行诡诈，又把那当灭的物与自己的器皿放在一起。
JOSH|7|12|因此， 以色列 人在仇敌面前站立不住。他们在仇敌面前转身逃跑，因为他们成了当灭的物。你们若不把当灭的物从你们中间除掉，我就不再与你们同在了。
JOSH|7|13|你起来，去叫百姓分别为圣，说：‘你们要为了明天使自己分别为圣，因为耶和华－ 以色列 的上帝这样说： 以色列 啊，在你中间有当灭的物；你们若不把你们中间当灭之物除掉，你在仇敌面前必站立不住！’
JOSH|7|14|到了早晨，你们要按着支派近前来。耶和华所选的支派，要按着宗族近前来；耶和华所选的宗族，要按着家族近前来；耶和华所选的家族，要按着男丁，一个一个近前来。
JOSH|7|15|被选的人有当灭之物在他那里，他和他所有的必被火焚烧，因为他违背了耶和华的约，又因他在 以色列 中做了愚妄的事。”
JOSH|7|16|于是， 约书亚 清早起来，召 以色列 按着支派近前来。选出来的是 犹大 支派。
JOSH|7|17|他召 犹大 的宗族近前来，选出来的是 谢拉 宗族。他召 谢拉 宗族，按着男丁 ，一个一个近前来，选出来的是 撒底 。
JOSH|7|18|他召 撒底 的家族，按着男丁，一个一个近前来，就选出 犹大 支派， 谢拉 的曾孙， 撒底 的孙子， 迦米 的儿子 亚干 。
JOSH|7|19|约书亚 对 亚干 说：“我儿，我劝你将荣耀归给耶和华－ 以色列 的上帝，在他面前认罪，把你所做的事告诉我，不可向我隐瞒。”
JOSH|7|20|亚干 回答 约书亚 说：“我实在得罪了耶和华－ 以色列 的上帝。这是我所做的：
JOSH|7|21|我在所夺取的财物中看见一件美好的 示拿 外袍，二百舍客勒银子，一条重五十舍客勒的金子。我贪爱这些物件，就拿去了。看哪，这些东西都埋在我帐棚内的地里，银子在外袍底下。”
JOSH|7|22|约书亚 就派使者跑到 亚干 的帐棚里。看哪，那件外袍藏在他的帐棚里，银子在外袍底下。
JOSH|7|23|他们从帐棚里把这些东西取出来，拿到 约书亚 和 以色列 众人 那里，倒在耶和华面前。
JOSH|7|24|约书亚 和 以色列 众人把 谢拉 的曾孙 亚干 和那银子、那件外袍、那条金子，以及 亚干 的儿女、牛、驴、羊、帐棚，和他所有的，都带着上到 亚割谷 去。
JOSH|7|25|约书亚 说：“你为什么给我们招惹灾祸呢？今日耶和华必使你遭受灾祸。”于是 以色列 众人用石头打死他，用火焚烧他们，把石头扔在其上。
JOSH|7|26|众人在 亚干 身上堆了一大堆石头，直存到今日。于是耶和华转意，不发他的烈怒。因此，那地方名叫 亚割谷 ，直到今日。
JOSH|8|1|耶和华对 约书亚 说：“不要惧怕，也不要惊惶。你起来，率领所有作战的士兵上 艾城 去。看，我已经把 艾城 的王和他的百姓、他的城，以及他的地，都交在你手里。
JOSH|8|2|你怎样处置 耶利哥 和 耶利哥 的王，也当照样处置 艾城 和 艾城 的王。只是城内所夺的财物和牲畜，你们可以取为自己的掠物。你要在城的后面设下伏兵。
JOSH|8|3|于是， 约书亚 和所有作战的士兵都起来，上 艾城 去。 约书亚 选了三万大能的勇士，夜间派遣他们前去，
JOSH|8|4|吩咐他们说：“看，你们要在城的后面埋伏，不可离城太远，各人都要准备。
JOSH|8|5|我与我所带领的众士兵要向城前进。城里的人像上一次那样出来迎击我们的时候，我们就在他们面前逃跑。
JOSH|8|6|他们会出来追赶我们，直到我们引诱他们远离那城。因为他们必说：‘这些人像上次那样在我们面前逃跑。’所以我们要在他们面前逃跑 。
JOSH|8|7|那时，你们就从埋伏的地方起来，夺取那城，因为耶和华－你们的上帝必把城交在你们的手里。
JOSH|8|8|你们夺了城以后，要放火烧城，照耶和华的话去做。看，这是我吩咐你们的。”
JOSH|8|9|于是， 约书亚 派遣他们前去。他们行军到埋伏的地方，伏在 伯特利 和 艾城 的中间，就是 艾城 的西边。这夜， 约书亚 在士兵中间过夜。
JOSH|8|10|约书亚 清早起来，点齐士兵。他和 以色列 的长老在百姓前面上 艾城 去。
JOSH|8|11|所有跟他一起作战的士兵都上去，向前逼近，来到城前，就在 艾城 北边安营。 约书亚 与 艾城 之间隔着一个山谷。
JOSH|8|12|他选了约五千人，安排他们埋伏在 伯特利 和 艾城 的中间，就是 艾城 的西边。
JOSH|8|13|于是，他们布署军队，就是城北的全军和城西的伏兵。当夜 约书亚 进入山谷之中。
JOSH|8|14|艾城 的王看见了，就和城里的人清早起来，急忙出去，他和所有的士兵到了所定的地点，在 亚拉巴 前，迎击 以色列 ，与之交战；王并不知道城的后面有伏兵。
JOSH|8|15|约书亚 和 以色列 众人在他们面前装败，往旷野的路逃跑。
JOSH|8|16|城内所有的百姓都被召来追赶他们。 艾城 的人追赶 约书亚 的时候，就被引诱远离了城。
JOSH|8|17|艾城 和 伯特利 没有一人不出来追赶 以色列 人的。他们撇下敞开的城门，去追赶 以色列 人。
JOSH|8|18|耶和华对 约书亚 说：“你向 艾城 伸出手里的标枪，因为我要把那城交在你手里。” 约书亚 就向那城伸出手里的标枪。
JOSH|8|19|他一伸手，伏兵立刻从埋伏的地方冲出来，直攻入城，夺了它，立刻放火烧城。
JOSH|8|20|艾城 的人回头，往后一看，看哪，城中烟气冲天，他们向这边或那边都无处可逃。往旷野逃跑的百姓就转身攻击那些追赶他们的人。
JOSH|8|21|约书亚 和 以色列 众人见伏兵已经夺了城，城中烟气上腾，就转身击杀 艾城 的人。
JOSH|8|22|伏兵也出城追击他们，他们就被 以色列 人前后夹攻，四面受敌。于是 以色列 人击杀他们，没有留下一个幸存者，也没有一个逃脱。
JOSH|8|23|以色列 人生擒了 艾城 的王，把他解到 约书亚 那里。
JOSH|8|24|以色列 人在田间和旷野杀尽了追赶他们的 艾城 所有的居民。他们全倒在刀下，直到灭尽。 以色列 众人就回到 艾城 ，用刀杀了城中的人。
JOSH|8|25|当日杀死的人，连男带女共有一万二千，这也是 艾城 所有的人。
JOSH|8|26|约书亚 没有收回手里所伸出来的标枪，直到他灭绝 艾城 所有的居民。
JOSH|8|27|只是牲畜和城内所夺的财物， 以色列 人都照耶和华所吩咐 约书亚 的话，取为自己的掠物。
JOSH|8|28|约书亚 焚烧 艾城 ，使城成为永远的废墟，直到今日还是荒凉。
JOSH|8|29|他把 艾城 的王挂在树上，直到晚上。日落的时候， 约书亚 吩咐人把尸首从树上取下来，丢在城门口，并在尸首上堆了一大堆石头，直存到今日。
JOSH|8|30|那时， 约书亚 在 以巴路山 上为耶和华－ 以色列 的上帝筑一座坛。
JOSH|8|31|这坛是照耶和华的仆人 摩西 吩咐 以色列 人，用没有动过铁器的整块石头所筑的，正如 摩西 律法书上所写的。他们在这坛上给耶和华奉献燔祭，又宰牲作为平安祭。
JOSH|8|32|约书亚 在那里，当着 以色列 人面前，将 摩西 所写的律法抄写在石头上。
JOSH|8|33|以色列 众人，无论是本地人或寄居的，都和他们的长老、官长和审判官，站在约柜两旁，在抬耶和华约柜的 利未 家的祭司面前，一半对着 基利心山 ，一半对着 以巴路山 ，照耶和华的仆人 摩西 先前所吩咐的，为 以色列 百姓祝福。
JOSH|8|34|随后， 约书亚 将律法上祝福和诅咒的话，照着律法书上一切所写的，宣读一遍。
JOSH|8|35|摩西 所吩咐的一切话， 约书亚 在 以色列 全会众和妇女、孩童，以及住在他们中间的外人面前，没有一句不宣读的。
JOSH|9|1|约旦河 西，住山区、低地和沿 大海 一带直到 黎巴嫩 的诸王，就是 赫 人、 亚摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人的诸王，听见这事，
JOSH|9|2|就都聚集，同心合意要与 约书亚 和 以色列 人作战。
JOSH|9|3|基遍 的居民听见 约书亚 向 耶利哥 和 艾城 所做的事，
JOSH|9|4|就设诡计，假扮使者 出去。他们拿旧布袋和破裂补过的旧皮酒袋驮在驴上，
JOSH|9|5|将补过的旧鞋穿在脚上，把旧衣服穿在身上，作食物的饼都又干又长了霉 。
JOSH|9|6|他们到 吉甲 营中 约书亚 那里，对他和 以色列 人说：“我们是从远地来的，现在求你与我们立约。”
JOSH|9|7|以色列 人对 希未 人说：“或许你是住在我附近的。若是这样，我怎能和你立约呢？”
JOSH|9|8|他们对 约书亚 说：“我们是你的仆人。” 约书亚 对他们说：“你们是什么人？是从哪里来的？”
JOSH|9|9|他们对他说：“你的仆人是因耶和华－你上帝的名从极远之地来的。我们听见他的名声，他在 埃及 所做的一切，
JOSH|9|10|以及他向 约旦河 东的两个 亚摩利 王， 希实本 王 西宏 和在 亚斯她录 的 巴珊 王 噩 所做的一切。
JOSH|9|11|我们的长老和我们当地所有的居民对我们说：‘你们手里要带着路上用的干粮去迎接 以色列 人，对他们说：我们是你们的仆人。现在求你们与我们立约。’
JOSH|9|12|我们出来要往你们这里来的那日，这从我们家里带出来的饼是热的；看哪，现在这饼又干又长了霉。
JOSH|9|13|这些皮酒袋，我们盛酒的时候还是新的；看哪，现在已经破裂了。我们这些衣服和鞋，因为路途非常遥远，也都穿旧了。”
JOSH|9|14|以色列 人收下他们的一些食物，但是没有求问耶和华的指示。
JOSH|9|15|于是 约书亚 与他们建立和好关系，与他们立约，让他们存活；会众的领袖也向他们起誓。
JOSH|9|16|以色列 人与他们立约之后，过了三天才听说他们是近邻，住在附近。
JOSH|9|17|以色列 人起行，第三天就到了他们的城镇，他们的城镇是 基遍 、 基非拉 、 比录 和 基列．耶琳 。
JOSH|9|18|因为会众的领袖已经指着耶和华－ 以色列 的上帝向他们起誓，所以 以色列 人不击杀他们。全会众就向领袖发怨言。
JOSH|9|19|众领袖对全会众说：“我们已经指着耶和华－ 以色列 的上帝向他们起誓，现在我们不能碰他们。
JOSH|9|20|我们要这样对待他们，让他们存活，免得因我们向他们所起的誓而愤怒临到我们。”
JOSH|9|21|领袖对会众说：“让他们活着吧。”于是他们照领袖所说的，为全会众作劈柴挑水的人。
JOSH|9|22|约书亚 召了他们来，对他们说：“你们为什么欺骗我们说：‘我们离你们很远’呢？其实你们就住在我们附近。
JOSH|9|23|现在你们当受诅咒！你们中间必不断有人作奴仆，为我上帝的殿作劈柴挑水的人。”
JOSH|9|24|他们回答 约书亚 说：“因为确实有人告诉你的仆人，耶和华－你的上帝曾吩咐他的仆人 摩西 ，把这全地赐给你们，并要在你们面前除灭这地所有的居民。我们因你们的缘故很怕自己丧命，就做了这事。
JOSH|9|25|现在，看哪，我们在你手中，你看怎样待我们是好的，是对的，就这样做吧！”
JOSH|9|26|于是 约书亚 就这样对待他们，他救了他们脱离 以色列 人的手， 以色列 人没有杀他们。
JOSH|9|27|那日， 约书亚 分派他们到耶和华选择的地方，为会众和耶和华的坛劈柴挑水，直到今日。
JOSH|10|1|耶路撒冷 王 亚多尼．洗德 听见 约书亚 夺了 艾城 ，彻底毁灭，处置 艾城 和 艾城 的王像处置 耶利哥 和 耶利哥 的王一样，又听见 基遍 的居民与 以色列 人立了和约，住在他们中间，
JOSH|10|2|耶路撒冷 人就很惧怕，因为 基遍 是一座大城，如京城一样，比 艾城 更大，并且城内的人都是勇士。
JOSH|10|3|耶路撒冷 王 亚多尼．洗德 派人去见 希伯仑 王 何咸 、 耶末 王 毗兰 、 拉吉 王 雅非亚 和 伊矶伦 王 底璧 ，说：
JOSH|10|4|“求你们上来帮助我，我们好攻打 基遍 ，因为它与 约书亚 和 以色列 人立了和约。”
JOSH|10|5|于是五个 亚摩利 王，就是 耶路撒冷 王、 希伯仑 王、 耶末 王、 拉吉 王和 伊矶伦 王，联合上去，率领他们所有的军队，对着 基遍 安营，要攻打 基遍 。
JOSH|10|6|基遍 人就派人到 吉甲 的营中 约书亚 那里，说：“不要袖手不顾你的仆人，求你赶快上来拯救我们，帮助我们，因为住山区 亚摩利 人的诸王已经联合来攻击我们。”
JOSH|10|7|于是 约书亚 和所有跟他一起作战的士兵，以及大能的勇士，从 吉甲 上去。
JOSH|10|8|耶和华对 约书亚 说：“不要怕他们， 因为我已将他们交在你手里，他们没有一人能在你面前站立得住。”
JOSH|10|9|约书亚 就连夜从 吉甲 上去，猛然袭击他们。
JOSH|10|10|耶和华使他们在 以色列 人面前溃乱。 约书亚 在 基遍 大大击杀他们，在 伯．和仑 的上坡路上追赶他们，击杀他们，直到 亚西加 和 玛基大 。
JOSH|10|11|他们在 以色列 人面前逃跑。正在 伯．和仑 下坡的时候，耶和华从天上降下大冰雹 在他们身上，直降到 亚西加 ，打死他们。被冰雹打死的，比 以色列 人用刀杀死的还多。
JOSH|10|12|当耶和华将 亚摩利 人交给 以色列 人的那一日， 约书亚 向耶和华说话，在 以色列 人眼前说： “太阳啊，停在 基遍 ； 月亮啊，停在 亚雅仑谷 。”
JOSH|10|13|太阳就停住，月亮就止住， 直到国民向敌人报仇。 这事岂不是写在《雅煞珥书》上吗？太阳停在天空当中，没有急速下落，约有一整天。
JOSH|10|14|在这日以前，这日以后，耶和华听人的声音，没有像这日的，这是因为耶和华为 以色列 作战。
JOSH|10|15|约书亚 和跟他一起的 以色列 众人回到 吉甲 的营中。
JOSH|10|16|那五个王逃跑，躲在 玛基大 洞里。
JOSH|10|17|有人告诉 约书亚 说：“那五个王已经找到了，都躲在 玛基大 洞里。”
JOSH|10|18|约书亚 说：“你们把几块大石头滚到洞口，派人在那里看守他们。
JOSH|10|19|你们却不可停留，要追赶你们的仇敌，从后面攻击他们，不让他们进到自己的城镇，因为耶和华－你们的上帝已经把他们交在你们手里。”
JOSH|10|20|约书亚 和 以色列 人彻底击败他们，直到把他们灭尽，只剩下少许的人逃进坚固的城。
JOSH|10|21|众百姓就安然回到 玛基大 营中 ，到 约书亚 那里。没有人敢向 以色列 人饶舌。
JOSH|10|22|约书亚 说：“打开洞口，把那五个王从洞里带出来，到我这里。”
JOSH|10|23|众人就这样做，把那五个王，就是 耶路撒冷 王、 希伯仑 王、 耶末 王、 拉吉 王和 伊矶伦 王，从洞里带出来，到 约书亚 那里。
JOSH|10|24|他们带出那五个王到 约书亚 那里的时候， 约书亚 就召了 以色列 众人来，对和他同去的军官说：“你们近前来，把脚踏在这些王的颈项上。”他们就近前来，把脚踏在这些王的颈项上。
JOSH|10|25|约书亚 对他们说：“你们不要惧怕，也不要惊惶。当刚强壮胆，因为耶和华必这样处置你们要攻打的所有仇敌。”
JOSH|10|26|随后， 约书亚 把这五个王杀死，挂在五棵树上。他们就被挂在树上，直到晚上。
JOSH|10|27|日落的时候， 约书亚 吩咐人把尸首从树上取下来，丢在他们躲过的洞里，把几块大石头放在洞口，直存到今日。
JOSH|10|28|当日， 约书亚 夺了 玛基大 ，用刀击杀城中的人和王，把城中所有人完全灭尽，没有留下一个幸存者。他处置 玛基大 王，像从前处置 耶利哥 王一样。
JOSH|10|29|约书亚 和跟他一起的 以色列 众人从 玛基大 往 立拿 去，攻打 立拿 。
JOSH|10|30|耶和华将 立拿 和 立拿 的王也交在 以色列 人手里。 约书亚 攻打这城，用刀击杀了城中所有的人，没有留下一个幸存者。他处置 立拿 王，像从前处置 耶利哥 王一样。
JOSH|10|31|约书亚 和跟他一起的 以色列 众人从 立拿 往 拉吉 去，对着 拉吉 安营，攻打这城。
JOSH|10|32|耶和华将 拉吉 交在 以色列 人的手里。第二日 约书亚 就夺了 拉吉 ，用刀击杀了城中所有的人，正如他向 立拿 一切所做的。
JOSH|10|33|那时 基色 王 何兰 上来帮助 拉吉 ， 约书亚 就把他和他的百姓都击杀了，没有留下一个幸存者。
JOSH|10|34|约书亚 和跟他一起的 以色列 众人从 拉吉 往 伊矶伦 去，对着 伊矶伦 安营，攻打这城。
JOSH|10|35|当日 约书亚 就夺了城，用刀击杀了城中的人。那日， 约书亚 把城中所有的人完全灭尽，正如他向 拉吉 一切所做的。
JOSH|10|36|约书亚 和跟他一起的 以色列 众人从 伊矶伦 上 希伯仑 去，攻打这城，
JOSH|10|37|夺了 希伯仑 ，用刀击败 希伯仑 、它的王和属它的一切城镇，以及城中所有的人；他没有留下一个幸存者，正如他向 伊矶伦 所做的，把城中所有的人完全灭尽。
JOSH|10|38|约书亚 和跟他一起的 以色列 众人回到 底璧 ，攻打这城，
JOSH|10|39|夺了 底璧 和属它的一切城镇，又擒获它的王，用刀把城中所有的人完全灭尽，没有留下一个幸存者。他处置 底璧 和它的王，像从前处置 希伯仑 ，处置 立拿 和它的王一样。
JOSH|10|40|这样， 约书亚 击败全地的人，就是山区、 尼革夫 、低地、山坡的人，和那里的众王，没有留下一个幸存者。他把凡有气息的完全灭尽，正如耶和华－ 以色列 的上帝所吩咐的。
JOSH|10|41|约书亚 从 加低斯．巴尼亚 攻到 迦萨 ，又攻打 歌珊 全地，直到 基遍 。
JOSH|10|42|约书亚 一举击败了这些王，夺了他们的地，因为耶和华－ 以色列 的上帝为 以色列 作战。
JOSH|10|43|于是 约书亚 和跟他一起的 以色列 众人回到 吉甲 的营中。
JOSH|11|1|夏琐 王 耶宾 听见了，就派人到 玛顿 王 约巴 、 伸仑 王、 押煞 王，
JOSH|11|2|和北方山区、 基尼烈 南边的 亚拉巴 、低地、西边 多珥 山冈 的诸王，
JOSH|11|3|以及东方和西方的 迦南 人、山区的 亚摩利 人、 赫 人、 比利洗 人、 耶布斯 人，和 黑门山 下 米斯巴 地的 希未 人那里。
JOSH|11|4|他们和他们的众军都出来，一大队人马，多如海边的沙，并有极多的战车战马。
JOSH|11|5|众王组成联军，来到 米伦 水边一同安营，要与 以色列 作战。
JOSH|11|6|耶和华对 约书亚 说：“你不要怕他们。明日这时，我必把他们全部交给 以色列 人杀灭。你要砍断他们马的蹄筋，用火焚烧他们的战车。”
JOSH|11|7|于是 约书亚 和所有跟他一起作战的士兵，来到 米伦 水边，突然攻击他们。
JOSH|11|8|耶和华将他们交在 以色列 人手里， 以色列 人就击杀他们，追赶他们到 西顿 大城，到 米斯利弗．玛音 ，直到东边 米斯巴 的山谷。 以色列 人击杀他们，没有留下一个幸存者。
JOSH|11|9|约书亚 照耶和华所吩咐他的去做，砍断他们马的蹄筋，用火焚烧他们的战车。
JOSH|11|10|那时， 约书亚 转回，夺了 夏琐 ，用刀杀了 夏琐 王。先前 夏琐 在这些王国中是为首的。
JOSH|11|11|以色列 人用刀击杀城中所有的人，把他们完全灭尽；凡有气息的，没有留下一个。 约书亚 又用火焚烧 夏琐 。
JOSH|11|12|约书亚 夺了这些王的一切城镇，擒获了这些王，用刀杀了他们，把他们完全灭尽，正如耶和华的仆人 摩西 所吩咐的。
JOSH|11|13|至于造在山冈上的城镇，除了 夏琐 以外， 以色列 人都没有焚烧。 约书亚 只焚烧了 夏琐 。
JOSH|11|14|从那些城镇所夺的财物和牲畜， 以色列 人都取为自己的掠物。至于所有的人，他们都用刀杀了，直到灭尽；凡有气息的，没有留下一个。
JOSH|11|15|耶和华怎样吩咐他的仆人 摩西 ， 摩西 就这样吩咐 约书亚 ， 约书亚 也照样做了。凡耶和华所吩咐 摩西 的， 约书亚 没有一件偏离不做的。
JOSH|11|16|约书亚 夺了那全地，就是山区、整个 尼革夫 、 歌珊 全地、低地、 亚拉巴 、 以色列 的山区和山下的低地，
JOSH|11|17|从上 西珥 的 哈拉山 ，直到 黑门山 下面 黎巴嫩 平原的 巴力．迦得 。他擒获了那里的众王，把他们杀死。
JOSH|11|18|约书亚 和这些王作战了很长的一段日子。
JOSH|11|19|除了 希未 人 基遍 的居民之外，没有一城与 以色列 人讲和，都是 以色列 人作战夺来的。
JOSH|11|20|因为耶和华的意思是要使他们的心刚硬，来与 以色列 人作战，好使他们全被杀灭，不蒙怜悯，反被除灭，正如耶和华所吩咐 摩西 的。
JOSH|11|21|那时 约书亚 来到，剪除了住山区、 希伯仑 、 底璧 、 亚拿伯 、整个 犹大 山区和 以色列 山区的 亚衲 族人。 约书亚 把他们和他们的城镇尽都毁灭。
JOSH|11|22|以色列 人的地中没有留下一个 亚衲 族人，只有一些还留在 迦萨 、 迦特 和 亚实突 。
JOSH|11|23|这样， 约书亚 照着耶和华所吩咐 摩西 的一切话夺了那全地，就按着 以色列 支派所得的份把地分给他们为业。于是国中太平，没有战争了。
JOSH|12|1|这些是 以色列 人在 约旦河 东，向日出的方向，从 亚嫩谷 直到 黑门山 ，以及东边 亚拉巴 的整个地区所击杀的王和所得的地：
JOSH|12|2|有住 希实本 的 亚摩利 王 西宏 ，他统治的地从 亚嫩谷 边的 亚罗珥 起，包括谷中之城和 基列 的一半，直到 亚扪 人边界的 雅博河 ，
JOSH|12|3|以及从东边的 亚拉巴 ，直到 基尼烈海 ，又向东通过 伯．耶施末 的路，直到 亚拉巴 的海，就是 盐海 ，再往南直到 毗斯迦山 斜坡的山脚。
JOSH|12|4|又有 巴珊 王 噩 ，他是 利乏音 人所剩下的，住在 亚斯她录 和 以得来 。
JOSH|12|5|他统治的地是 黑门山 、 撒迦 、 巴珊 全地，直到 基述 人和 玛迦 人的边界，以及 基列 的一半，直到 希实本 王 西宏 的边界。
JOSH|12|6|这两个王是耶和华的仆人 摩西 和 以色列 人所击杀的。耶和华的仆人 摩西 把他们的地赐给 吕便 人、 迦得 人和 玛拿西 半支派的人为业。
JOSH|12|7|这些是 约书亚 和 以色列 人在 约旦河 西所击杀的诸王，他们的地从 黎巴嫩 平原的 巴力．迦得 ，直上到 西珥 的 哈拉山 。 约书亚 按着 以色列 支派所得的份把这地分给他们为业，
JOSH|12|8|就是 赫 人、 亚摩利 人、 迦南 人、 比利洗 人、 希未 人、 耶布斯 人的地，包括山区、低地、 亚拉巴 、山坡、旷野和 尼革夫 。
JOSH|12|9|这些王是： 耶利哥 王一人， 靠近 伯特利 的 艾城 王一人，
JOSH|12|10|耶路撒冷 王一人， 希伯仑 王一人，
JOSH|12|11|耶末 王一人， 拉吉 王一人，
JOSH|12|12|伊矶伦 王一人， 基色 王一人，
JOSH|12|13|底璧 王一人， 基德 王一人，
JOSH|12|14|何珥玛 王一人， 亚拉得 王一人，
JOSH|12|15|立拿 王一人， 亚杜兰 王一人，
JOSH|12|16|玛基大 王一人， 伯特利 王一人，
JOSH|12|17|他普亚 王一人， 希弗 王一人，
JOSH|12|18|亚弗 王一人， 拉沙仑 王一人，
JOSH|12|19|玛顿 王一人， 夏琐 王一人，
JOSH|12|20|伸仑．米仑 王一人 ， 押煞 王一人，
JOSH|12|21|他纳 王一人， 米吉多 王一人，
JOSH|12|22|基低斯 王一人， 靠近 迦密 的 约念 王一人，
JOSH|12|23|多珥 山冈 的 多珥 王一人， 吉甲 的 戈印 王一人，
JOSH|12|24|得撒 王一人， 共三十一个王。
JOSH|13|1|约书亚 年纪老迈，耶和华对他说：“你年纪老迈了，还有极多剩下的未得之地。
JOSH|13|2|这是剩下的地： 非利士 人的全境和一切属于 基述 人的，
JOSH|13|3|是从 埃及 东边的 西曷河 往北，直到 以革伦 的边界，算是属 迦南 人的地，那里有 非利士 人五个领袖统治 迦萨 人、 亚实突 人、 亚实基伦 人、 迦特 人、 以革伦 人；还有属于 亚卫 人的，
JOSH|13|4|在南边；还有 迦南 人的全地，以及 西顿 人的 米亚拉 到 亚弗 ，直到 亚摩利 人的边界；
JOSH|13|5|还有 迦巴勒 人的地，以及向日出方向的 黎巴嫩 全地，从 黑门山 下的 巴力．迦得 ，直到 哈马口 ；
JOSH|13|6|从 黎巴嫩 直到 米斯利弗．玛音 ，一切山区的居民，就是所有的 西顿 人，我必在 以色列 人面前赶走他们。你只管照我所吩咐的，抽签将这地分给 以色列 人为业。
JOSH|13|7|现在你要把这地分给九个支派和 玛拿西 半个支派为业。
JOSH|13|8|吕便 、 迦得 二支派已经和 玛拿西 另外半个支派得了产业，就是耶和华的仆人 摩西 在 约旦河 东所赐给他们的：
JOSH|13|9|从 亚嫩谷 边的 亚罗珥 和谷中之城， 米底巴 的整个平原，直到 底本 ；
JOSH|13|10|还有在 希实本 作王的 亚摩利 王 西宏 的诸城，直到 亚扪 人的边界；
JOSH|13|11|还有 基列 ， 基述 人和 玛迦 人的边界，整个 黑门山 、整个 巴珊 ，直到 撒迦 ；
JOSH|13|12|还有在 亚斯她录 和 以得来 作王的 巴珊 王 噩 的整个国土， 噩 是 利乏音 人惟一存留的。 摩西 击败了这些人，把他们赶走。
JOSH|13|13|以色列 人却没有赶走 基述 人和 玛迦 人； 基述 人和 玛迦 人仍住在 以色列 中，直到今日。
JOSH|13|14|只是 利未 支派， 摩西 没有分产业给他们。他们的产业是献给耶和华－ 以色列 上帝的火祭，正如耶和华对他们说的。
JOSH|13|15|摩西 按着 吕便 支派的宗族分产业给他们。
JOSH|13|16|他们的地界是 亚嫩谷 边的 亚罗珥 和谷中之城，靠近 米底巴 的整个平原；
JOSH|13|17|还有 希实本 和属 希实本 平原的各城， 底本 、 巴末．巴力 、 伯．巴力．勉 、
JOSH|13|18|雅杂 、 基底莫 、 米法押 、
JOSH|13|19|基列亭 、 西比玛 、谷中山冈上的 细列．沙辖 、
JOSH|13|20|伯．毗珥 、 毗斯迦山 斜坡、 伯．耶施末 ；
JOSH|13|21|还有平原的各城，和 亚摩利 王 西宏 的整个国土。这 西宏 曾在 希实本 作王， 摩西 把他和 米甸 的族长 以未 、 利金 、 苏珥 、 户珥 、 利巴 击杀了；他们都是属 西宏 的领袖，曾住在这地。
JOSH|13|22|以色列 人杀了这些人时，也用刀杀了 比珥 的儿子占卜的 巴兰 。
JOSH|13|23|吕便 人的地界就是 约旦河 和靠近 约旦河 的地。以上是 吕便 人按着宗族所得为业的城镇和所属的村庄。
JOSH|13|24|摩西 按着 迦得 支派的宗族分产业给他们。
JOSH|13|25|他们的地界是 雅谢 和 基列 的各城，以及 亚扪 人之地的一半，直到 拉巴 前面的 亚罗珥 ；
JOSH|13|26|还有从 希实本 到 拉抹．米斯巴 和 比多宁 ，又从 玛哈念 到 底璧 的边界，
JOSH|13|27|和谷中的 伯．亚兰 、 伯．宁拉 、 疏割 、 撒分 ，就是 希实本 王 西宏 国土中其余的地，以及 约旦河 与靠近 约旦河 的地，直到 基尼烈海 的边缘，都在 约旦河 东。
JOSH|13|28|以上是 迦得 人按着宗族所得为业的城镇和所属的村庄。
JOSH|13|29|摩西 分产业给 玛拿西 半支派，这是按着 玛拿西 半支派的宗族分的。
JOSH|13|30|他们的地界是从 玛哈念 起，包括整个 巴珊 全地，就是 巴珊 王 噩 的整个国土，以及在 巴珊 、 睚珥 的一切城镇，共六十个；
JOSH|13|31|还有 基列 的一半，以及 巴珊 国的王 噩 的 亚斯她录 和 以得来 两座城。这些地是按着宗族分给 玛拿西 儿子 玛吉 子孙的，就是给 玛吉 一半子孙的。
JOSH|13|32|以上是 摩西 在 约旦河 东， 耶利哥 对面的 摩押 平原所分配的产业。
JOSH|13|33|只是 利未 支派， 摩西 没有把产业分给他们。耶和华－ 以色列 的上帝是他们的产业，正如耶和华对他们说的。
JOSH|14|1|这是 以色列 人在 迦南 地所得的产业，就是祭司 以利亚撒 和 嫩 的儿子 约书亚 ，以及 以色列 人各支派父系的领袖所分给他们的。
JOSH|14|2|他们照耶和华藉 摩西 所吩咐的，抽签分产业给九个半支派。
JOSH|14|3|摩西 在 约旦河 东已经分了产业给另外两个半支派。但是，他在他们中间没有分产业给 利未 人。
JOSH|14|4|因 约瑟 的子孙成了两个支派，就是 玛拿西 和 以法莲 。虽然他们没有分地给 利未 人，却给 利未 人城镇居住，以及城镇的郊外供他们牧养牲畜，安置财物。
JOSH|14|5|耶和华怎样吩咐 摩西 ， 以色列 人就照样做，把地分了。
JOSH|14|6|犹大 人来到 吉甲 ， 约书亚 那里， 基尼洗 族 耶孚尼 的儿子 迦勒 对 约书亚 说：“耶和华在 加低斯．巴尼亚 指着我和你对神人 摩西 所说的话，你都知道。
JOSH|14|7|耶和华的仆人 摩西 从 加低斯．巴尼亚 差派我窥探这地的时候，我刚四十岁。我把心里的话向他报告。
JOSH|14|8|虽然同我上去的众弟兄使百姓胆战心惊，我仍然专心跟从耶和华－我的上帝。
JOSH|14|9|那日， 摩西 起誓说：‘你脚所踏之地必要归你和你的子孙永远为业，因为你专心跟从耶和华－我的上帝。’
JOSH|14|10|现在，看哪，耶和华照他所说的使我活了这四十五年。当 以色列 人在旷野飘流的时候，耶和华曾对 摩西 说了这话。现在，看哪，我已经八十五岁了。
JOSH|14|11|现今我还很健壮，像 摩西 差派我去的那天一样；无论是战争，是出入，我现在的力量和那时的力量一样。
JOSH|14|12|请你将耶和华那日所说的这山区给我。那日你也曾听说，这里有 亚衲 族人，以及宽大坚固的城，或许耶和华会照他所说的与我同在，我就把他们赶出去。”
JOSH|14|13|于是 约书亚 为 耶孚尼 的儿子 迦勒 祝福，把 希伯仑 给他为业。
JOSH|14|14|所以 希伯仑 成了 基尼洗 族 耶孚尼 的儿子 迦勒 的产业，直到今日，因为他专心跟从耶和华－ 以色列 的上帝。
JOSH|14|15|希伯仑 从前名叫 基列．亚巴 ； 亚巴 是 亚衲 族最尊贵的人。于是国中太平，没有战争了。
JOSH|15|1|犹大 支派按着宗族抽签所得之地是在最南端，到 以东 的边界，往南直到 寻 的旷野。
JOSH|15|2|他们南边的地界是从 盐海 的顶端，就是朝南的海湾开始，
JOSH|15|3|通到 亚克拉滨 斜坡的南边，经过 寻 ，上到 加低斯．巴尼亚 的南边，又经过 希斯仑 ，上到 亚达珥 ，转到 甲加 ，
JOSH|15|4|再经过 押们 ，顺着 埃及 溪谷，这地界直通到海为止。这就是你们 南边的地界。
JOSH|15|5|东边的地界是从 盐海 到 约旦河 口。北边的地界是从 约旦河 口的海湾开始，
JOSH|15|6|这地界上到 伯．曷拉 ，经过 伯．亚拉巴 的北边，这地界上到 吕便 之子 波罕 的磐石。
JOSH|15|7|这地界是从 亚割谷 往北上到 底璧 ，直向 亚都冥 斜坡对面的 吉甲 ，就是河的南边，这地界再经过 隐．示麦 泉，直通到 隐．罗结 。
JOSH|15|8|这地界又上到 欣嫩子谷 ， 耶布斯 斜坡的南方， 耶布斯 就是 耶路撒冷 ，这地界又上到 欣嫩谷 西边对面的山顶，就是在 利乏音谷 的最北端。
JOSH|15|9|这地界又从山顶延伸到 尼弗多亚 水泉，通到 以弗仑山 的城镇，这地界又延伸到 巴拉 ， 巴拉 就是 基列．耶琳 。
JOSH|15|10|这地界又从 巴拉 往西绕到 西珥山 ，经过 耶琳山 斜坡的北边， 耶琳 就是 基撒仑 ，从那里又下到 伯．示麦 ，经过 亭拿 ，
JOSH|15|11|这地界通到 以革伦 斜坡的北边。这地界又延伸到 施基仑 ，经过 巴拉山 到 雅比聂 ，这地界直通到海为止。
JOSH|15|12|西边的地界就是 大海 和沿海一带之地。这是 犹大 人按着宗族所得之地四围的边界。
JOSH|15|13|约书亚 照耶和华所指示的，把 犹大 人中的一份土地，就是 基列．亚巴 ，分给 耶孚尼 的儿子 迦勒 。 亚巴 是 亚衲 族的祖先， 基列．亚巴 就是 希伯仑 。
JOSH|15|14|迦勒 从那里赶出 亚衲 的三族，就是 亚衲 族的 示筛 人、 亚希幔 人和 挞买 人。
JOSH|15|15|他又从那里上去，攻击 底璧 的居民，这 底璧 从前名叫 基列．西弗 。
JOSH|15|16|迦勒 说：“谁能攻打 基列．西弗 ，夺取那城，我就把我女儿 押撒 嫁给他。”
JOSH|15|17|迦勒 兄弟 基纳斯 的儿子 俄陀聂 夺取了那城， 迦勒 就把女儿 押撒 嫁给他。
JOSH|15|18|押撒 来的时候，催促丈夫向她父亲要一块田。 押撒 一下驴， 迦勒 就对她说：“你要什么？”
JOSH|15|19|她说：“求你给我福分；你既然把我安置在 尼革夫 地，求你也给我水泉。”她父亲就把上泉和下泉都赐给她。
JOSH|15|20|这是 犹大 支派按着宗族所得的产业。
JOSH|15|21|犹大 支派最南端，靠近 以东 边界的城镇，是 甲薛 、 以得 、 雅姑珥 、
JOSH|15|22|基拿 、 底摩拿 、 亚大达 、
JOSH|15|23|基低斯 、 夏琐 、 以提楠 、
JOSH|15|24|西弗 、 提鍊 、 比亚绿 、
JOSH|15|25|夏琐．哈大他 、 加略．希斯仑 ， 加略．希斯仑 就是 夏琐 ，
JOSH|15|26|亚曼 、 示玛 、 摩拉大 、
JOSH|15|27|哈萨．迦大 、 黑实门 、 伯．帕列 、
JOSH|15|28|哈萨．书亚 、 别是巴 、 比斯约他 、
JOSH|15|29|巴拉 、 以因 、 以森 、
JOSH|15|30|伊勒多腊 、 基失 、 何珥玛 、
JOSH|15|31|洗革拉 、 麦玛拿 、 三撒拿 、
JOSH|15|32|利巴勿 、 实忻 、 亚因 、 临门 ，共二十九座城，还有所属的村庄。
JOSH|15|33|在低地有 以实陶 、 琐拉 、 亚实拿 、
JOSH|15|34|撒挪亚 、 隐．干宁 、 他普亚 、 以楠 、
JOSH|15|35|耶末 、 亚杜兰 、 梭哥 、 亚西加 、
JOSH|15|36|沙拉音 、 亚底他音 、 基底拉 、 基底罗他音 ，共十四座城，还有所属的村庄。
JOSH|15|37|又有 洗楠 、 哈大沙 、 麦大．迦得 、
JOSH|15|38|底连 、 米斯巴 、 约帖 、
JOSH|15|39|拉吉 、 波斯加 、 伊矶伦 、
JOSH|15|40|迦本 、 拉幔 、 基提利 、
JOSH|15|41|基低罗 、 伯．大衮 、 拿玛 、 玛基大 ，共十六座城，还有所属的村庄。
JOSH|15|42|又有 立拿 、 以帖 、 亚珊 、
JOSH|15|43|益弗他 、 亚实拿 、 尼悉 、
JOSH|15|44|基伊拉 、 亚革悉 、 玛利沙 ，共九座城，还有所属的村庄。
JOSH|15|45|又有 以革伦 和所属的乡镇 与村庄，
JOSH|15|46|从 以革伦 直到海，一切靠近 亚实突 之地，以及所属的村庄、
JOSH|15|47|亚实突 和所属的乡镇与村庄， 迦萨 和所属的乡镇与村庄，到 埃及 溪谷，直到 大海 以及沿海一带之地。
JOSH|15|48|在山区有 沙密 、 雅提珥 、 梭哥 、
JOSH|15|49|大拿 、 基列．萨拿 ， 基列．萨拿 就是 底璧 ，
JOSH|15|50|亚拿伯 、 以实提莫 、 亚念 、
JOSH|15|51|歌珊 、 何仑 、 基罗 ，共十一座城，还有所属的村庄。
JOSH|15|52|又有 亚拉 、 度玛 、 以珊 、
JOSH|15|53|雅农 、 伯．他普亚 、 亚非加 、
JOSH|15|54|宏他 、 基列．亚巴 ， 基列．亚巴 就是 希伯仑 ， 洗珥 ，共九座城，还有所属的村庄。
JOSH|15|55|又有 玛云 、 迦密 、 西弗 、 淤他 、
JOSH|15|56|耶斯列 、 约甸 、 撒挪亚 、
JOSH|15|57|该隐 、 基比亚 、 亭拿 ，共十座城，还有所属的村庄。
JOSH|15|58|又有 哈忽 、 伯．夙 、 基突 、
JOSH|15|59|玛腊 、 伯．亚诺 、 伊勒提君 ，共六座城，还有所属的村庄。
JOSH|15|60|又有 基列．巴力 ， 基列．巴力 就是 基列．耶琳 ， 拉巴 ，共两座城，还有所属的村庄。
JOSH|15|61|在旷野有 伯．亚拉巴 、 密丁 、 西迦迦 、
JOSH|15|62|匿珊 、 盐城 、 隐．基底 ，共六座城，还有所属的村庄。
JOSH|15|63|至于住 耶路撒冷 的 耶布斯 人， 犹大 人不能把他们赶出去。于是， 耶布斯 人与 犹大 人同住在 耶路撒冷 ，直到今日。
JOSH|16|1|约瑟 的子孙抽签所得之地是从靠近 耶利哥 的 约旦河 起，以 耶利哥 东边的河水为边界，经过旷野，从 耶利哥 上去，直到 伯特利 的山区；
JOSH|16|2|从 伯特利 又到 路斯 ，经过 亚基 人的边界，直到 亚大录 ；
JOSH|16|3|又往西，下到 押利提 人的边界，到 下伯．和仑 的边界，到 基色 ，直通到海为止。
JOSH|16|4|约瑟 的儿子 玛拿西 、 以法莲 得了地业。
JOSH|16|5|以法莲 子孙的地界，按着宗族所得的如下：他们地业的东界，是从 亚大录．亚达 到 上伯．和仑 ，
JOSH|16|6|这地界直通到海。在北边，这地界是从 密米他 ，向东绕到 他纳．示罗 ，又经过 雅挪哈 的东边，
JOSH|16|7|从 雅挪哈 下到 亚大录 和 拿拉 ，再到 耶利哥 ，直到 约旦河 为止。
JOSH|16|8|这地界又从 他普亚 ，顺着 加拿河 往西延伸，直通到海为止。这就是 以法莲 支派按着宗族所得的地业。
JOSH|16|9|在 玛拿西 人地业的一切城镇和所属的村庄中，也保留一些城镇给 以法莲 的子孙。
JOSH|16|10|他们却没有赶出住在 基色 的 迦南 人。 迦南 人就住在 以法莲 人中，成为服劳役的仆人，直到今日。
JOSH|17|1|玛拿西 是 约瑟 的长子，这是他的支派抽签所得之地。 玛拿西 的长子， 基列 的父亲 玛吉 ，因为是勇士，就得了 基列 和 巴珊 。
JOSH|17|2|玛拿西 其余的子孙，就是 亚比以谢 的子孙， 希勒 的子孙， 亚斯烈 的子孙， 示剑 的子孙， 希弗 的子孙， 示米大 的子孙，都按着宗族抽签得了地。这都是 约瑟 的儿子 玛拿西 子孙中各宗族的男丁。
JOSH|17|3|玛拿西 的玄孙， 玛吉 的曾孙， 基列 的孙子， 希弗 的儿子 西罗非哈 没有儿子，只有女儿。他的女儿名叫 玛拉 、 挪阿 、 曷拉 、 密迦 、 得撒 。
JOSH|17|4|她们来到 以利亚撒 祭司和 嫩 的儿子 约书亚 以及众领袖面前，说：“耶和华曾吩咐 摩西 在我们兄弟中分产业给我们。”于是 约书亚 照耶和华的指示，在她们叔伯中，把产业分给她们。
JOSH|17|5|除了 约旦河 东的 基列 和 巴珊 地之外，还有十份的地业是属于 玛拿西 的，
JOSH|17|6|因为 玛拿西 支派的女子也在男子中分得产业。 基列 地属于 玛拿西 其余的子孙。
JOSH|17|7|玛拿西 的地界是从 亚设 起，到 示剑 前面的 密米他 ，往右 到 隐．他普亚 居民之地。
JOSH|17|8|他普亚 地归于 玛拿西 ，只是 玛拿西 边界的 他普亚城 却归于 以法莲 子孙。
JOSH|17|9|这地界从那里下到 加拿河 。河南边的城镇虽然在 玛拿西 境内，却是属于 以法莲 的。 玛拿西 的地界是在河的北边直通到海为止。
JOSH|17|10|南边属于 以法莲 ，北边属于 玛拿西 ，以海为界；北边达到 亚设 ，东边达到 以萨迦 。
JOSH|17|11|玛拿西 在 以萨迦 和 亚设 境内，有 伯．善 和所属的乡镇， 以伯莲 和所属的乡镇， 多珥 和所属乡镇的居民；还有 隐．多珥 和所属乡镇的居民， 他纳 和所属乡镇的居民， 米吉多 和所属乡镇的居民，共三个山冈 。
JOSH|17|12|只是 玛拿西 的子孙不能赶出这些城镇的居民， 迦南 人仍坚持住在那地。
JOSH|17|13|以色列 人强盛的时候，就叫 迦南 人做苦工，没有把他们全然赶走。
JOSH|17|14|约瑟 的子孙对 约书亚 说：“耶和华到如今这样赐福给我，我百姓众多，你为什么只给我抽一签，分一份的土地为业呢？”
JOSH|17|15|约书亚 对他们说：“如果你百姓众多，而 以法莲 山区太窄小，那么你可以上 比利洗 人和 利乏音 人之地的树林中，在那里开垦。”
JOSH|17|16|约瑟 的子孙说：“那山区容不下我们，而且住平原的 迦南 人，就是住 伯．善 和所属的乡镇，以及住在 耶斯列 平原的人，都有铁的战车。”
JOSH|17|17|约书亚 对 约瑟 家，就是 以法莲 和 玛拿西 人，说：“你百姓众多，并且强大，不可只有一签而已。
JOSH|17|18|那山区也要归你，虽然是树林，你可以去开垦，边缘之地也必归你。 迦南 人纵然强盛，有铁的战车，你也能把他们赶出去。”
JOSH|18|1|以色列 全会众都聚集在 示罗 ，把会幕设立在那里。那地已经被他们征服了。
JOSH|18|2|以色列 人中剩下七个支派还没有分得他们的地业。
JOSH|18|3|约书亚 对 以色列 人说：“耶和华－你们列祖的上帝所赐给你们的地，你们耽延不去得，要到几时呢？
JOSH|18|4|你们每支派要选三个人，我好派他们去，他们要起身走遍那地，按照各支派应得的地业写明，然后回到我这里来。
JOSH|18|5|他们要把地分成七份。 犹大 在南方，住在他的境内。 约瑟 家在北方，住在他们的境内。
JOSH|18|6|你们把地划成七份之后，就要把所写的带到我这里来。我要在耶和华－我们的上帝面前，为你们抽签。
JOSH|18|7|利未 人在你们中间没有分得地业，因为耶和华祭司的职分就是他们的产业。 迦得 支派、 吕便 支派和 玛拿西 半支派已经在 约旦河 东得了地业，是耶和华的仆人 摩西 给他们的。”
JOSH|18|8|那些去划地的人起来正要去的时候， 约书亚 吩咐他们说：“你们去走遍那地，把地划分以后，就回到我这里来。我要在 示罗 这里，在耶和华面前为你们抽签。”
JOSH|18|9|那些人就去了，走遍那地，按照城镇把地划成七份，写在册上，回到 示罗 营中 约书亚 那里。
JOSH|18|10|约书亚 就在 示罗 ，在耶和华面前为他们抽签。 约书亚 按照 以色列 人的支派，在那里把地分给他们。
JOSH|18|11|便雅悯 支派，按着宗族抽签所得之地，是在 犹大 子孙和 约瑟 子孙之间。
JOSH|18|12|他们北边的地界是从 约旦河 起，上到 耶利哥 斜坡的北边，再往西上到山区，直到 伯．亚文 的旷野。
JOSH|18|13|这地界从那里往南经过 路斯 ，直到 路斯 的斜坡， 路斯 就是 伯特利 ，又下到 亚他录．亚达 ，直到 下伯．和仑 南边的山。
JOSH|18|14|这地界往西延伸，又转向南，从 伯．和仑 南边对面的山，直通到 犹大 人的城 基列．巴力 ， 基列．巴力 就是 基列．耶琳 。这就是西边的地界。
JOSH|18|15|南边是从 基列．耶琳 的顶端为起点，这地界往西 通到 尼弗多亚 水泉，
JOSH|18|16|这地界又下到 欣嫩子谷 对面山的边缘，就是 利乏音谷 的北边；又下到 欣嫩谷 ，沿着 耶布斯 斜坡的南边，下到 隐．罗结 ；
JOSH|18|17|又往北转弯，通到 隐．示麦 ，直到 亚都冥 斜坡对面的 基利绿 ，又下到 吕便 之子 波罕 的磐石，
JOSH|18|18|又往北经过 亚拉巴 对面的斜坡 ，下到 亚拉巴 。
JOSH|18|19|这地界又经过 伯．曷拉 斜坡的北边，直通到 盐海 的北湾，就是 约旦河 的南端为止。这就是南边的地界。
JOSH|18|20|东边的地界是 约旦河 。这是 便雅悯 人按着宗族，照着他们四围的边界所得的地业。
JOSH|18|21|便雅悯 支派按着宗族所得的城镇就是： 耶利哥 、 伯．曷拉 、 伊麦．基悉 、
JOSH|18|22|伯．亚拉巴 、 洗玛脸 、 伯特利 、
JOSH|18|23|亚文 、 巴拉 、 俄弗拉 、
JOSH|18|24|基法．阿摩尼 、 俄弗尼 和 迦巴 ，共十二座城，以及所属的村庄；
JOSH|18|25|又有 基遍 、 拉玛 、 比录 、
JOSH|18|26|米斯巴 、 基非拉 、 摩撒 、
JOSH|18|27|利坚 、 伊利毗勒 、 他拉拉 、
JOSH|18|28|洗拉 、 以利弗 、 耶布斯 ， 耶布斯 就是 耶路撒冷 ， 基比亚 、 基列 ，共十四座城，以及所属的村庄。这是 便雅悯 人按着宗族所得的地业。
JOSH|19|1|第二签是 西缅 ，是 西缅 支派的人按着宗族抽出的，他们所得的地业是在 犹大 人地业的中间。
JOSH|19|2|他们所得为业之地是： 别是巴 ，或名 示巴 ， 摩拉大 、
JOSH|19|3|哈萨．书亚 、 巴拉 、 以森 、
JOSH|19|4|伊勒多腊 、 比土力 、 何珥玛 、
JOSH|19|5|洗革拉 、 伯．玛加博 、 哈萨．苏撒 、
JOSH|19|6|伯．利巴勿 、 沙鲁险 ，共十三座城，还有所属的村庄；
JOSH|19|7|又有 亚因 、 利门 、 以帖 、 亚珊 ，共四座城，还有所属的村庄；
JOSH|19|8|以及这些城镇周围一切的村庄，直到 巴拉．比珥 ，就是 尼革夫 的 拉玛 。这是 西缅 支派的人按着宗族所得的地业。
JOSH|19|9|西缅 人的地业取自 犹大 人的土地，因为 犹大 人所得的份过多，所以 西缅 人从 犹大 人的地业中取了地业。
JOSH|19|10|第三签是 西布伦 人按着宗族抽到的。他们地业的边界延伸到 撒立 。
JOSH|19|11|他们的地界往西，上到 玛拉拉 ，达到 大巴设 ，又达到 约念 前面的河。
JOSH|19|12|又从 撒立 往东转到向日出的方向，经过 吉斯绿．他泊 的边界，到 大比拉 ，又上到 雅非亚 。
JOSH|19|13|又从那里往东，经过 迦特．希弗 ，到 以特．加汛 ，通到 临门 ，延伸到 尼亚 。
JOSH|19|14|这地界在北边绕过 尼亚 ，到 哈拿顿 ，直通到 伊弗他．伊勒谷 ，
JOSH|19|15|包括 加他 、 拿哈拉 、 伸仑 、 以大拉 、 伯利恒 ，共十二座城，还有所属的村庄。
JOSH|19|16|这些城镇和所属的村庄是 西布伦 人按着宗族所得的地业。
JOSH|19|17|第四签是 以萨迦 ，是 以萨迦 人按着宗族抽出的。
JOSH|19|18|他们的地界是到 耶斯列 、 基苏律 、 书念 、
JOSH|19|19|哈弗连 、 示按 、 亚拿哈拉 、
JOSH|19|20|拉璧 、 基善 、 亚别 、
JOSH|19|21|利篾 、 隐．干宁 、 隐．哈大 、 伯．帕薛 。
JOSH|19|22|这地界达到 他泊 、 沙哈洗玛 、 伯．示麦 ，他们的地界直通到 约旦河 为止，共十六座城，还有所属的村庄。
JOSH|19|23|这些城镇和所属的村庄是 以萨迦 支派的人按着宗族所得的地业。
JOSH|19|24|第五签是 亚设 支派的人按着宗族抽出的。
JOSH|19|25|他们的地界是 黑甲 、 哈利 、 比田 、 押煞 、
JOSH|19|26|亚拉米勒 、 亚末 、 米沙勒 ，往西达到 迦密 ，又到 希曷．立纳 ，
JOSH|19|27|又转到向日出方向的 伯．大衮 ，达到 细步纶 ；又往北到 伊弗他．伊勒谷 ，到 伯．以墨 和 尼业 ，也通到 迦步勒 的左边 ，
JOSH|19|28|又到 义伯仑 、 利合 、 哈们 、 加拿 ，直到 西顿 大城。
JOSH|19|29|这地界转到 拉玛 ，直到坚固的 推罗城 。这地界又转到 何萨 ，靠近 亚革悉 一带的地方 ，直通到海为止。
JOSH|19|30|又有 乌玛 、 亚弗 、 利合 ，共二十二座城，还有所属的村庄。
JOSH|19|31|这些城镇和所属的村庄是 亚设 支派的人按着宗族所得的地业。
JOSH|19|32|第六签是 拿弗他利 人，是 拿弗他利 人按着宗族抽出的。
JOSH|19|33|他们的地界是从 希利弗 ，从 撒拿音 的橡树、 亚大米．尼吉 和 雅比聂 ，直到 拉共 ，直通到 约旦河 为止。
JOSH|19|34|这地界往西转到 亚斯纳．他泊 ，从那里通到 户割 ，南边达到 西布伦 ，西边达到 亚设 ，向日出的方向达到 约旦河 的 犹大 。
JOSH|19|35|坚固的城有 西丁 、 侧耳 、 哈末 、 拉甲 、 基尼烈 、
JOSH|19|36|亚大玛 、 拉玛 、 夏琐 、
JOSH|19|37|基低斯 、 以得来 、 隐．夏琐 、
JOSH|19|38|以利稳 、 密大．伊勒 、 和琏 、 伯．亚纳 、 伯．示麦 ，共十九座城，还有所属的村庄。
JOSH|19|39|这些城镇和所属的村庄是 拿弗他利 支派的人按着宗族所得的地业。
JOSH|19|40|但 支派，按着宗族，抽到第七签。
JOSH|19|41|他们地业的边界是 琐拉 、 以实陶 、 伊珥．示麦 、
JOSH|19|42|沙拉宾 、 亚雅仑 、 伊提拉 、
JOSH|19|43|以伦 、 亭拿 、 以革伦 、
JOSH|19|44|伊利提基 、 基比顿 、 巴拉 、
JOSH|19|45|伊胡得 、 比尼．比拉 、 迦特．临门 、
JOSH|19|46|美．耶昆 、 拉昆 ，以及 约帕 对面的地界。
JOSH|19|47|当 但 的子孙失去他们疆土的时候，就上去攻取 利善 ，用刀击杀城中的人，得了那城，住在城中，以他们祖先 但 的名字将 利善 改名为 但 。
JOSH|19|48|这些城镇和所属的村庄是 但 支派的人按着宗族所得的地业。
JOSH|19|49|以色列 人按着疆土完成了地业的分配，就在他们中间把地给 嫩 的儿子 约书亚 为业。
JOSH|19|50|他们照着耶和华的指示，把 约书亚 所要的城，就是 以法莲 山区的 亭拿．西拉 给了他。 约书亚 修建那城，住在城中。
JOSH|19|51|这就是 以利亚撒 祭司和 嫩 的儿子 约书亚 ，以及 以色列 人各支派父系的领袖，在 示罗 会幕的门口，耶和华面前抽签所分的地业。这样， 他们就完成了分地的事。
JOSH|20|1|耶和华吩咐 约书亚 说：
JOSH|20|2|“你吩咐 以色列 人说：‘你们要照我藉 摩西 所吩咐你们的，为自己设立逃城，
JOSH|20|3|使那无意中误杀人的，可以逃到那里。这些要作为你们逃避报血仇者的城。
JOSH|20|4|杀人者要逃到这些城中的一座，站在城门口，把他的事情陈诉给那城的长老听。他们就要接他入城，给他地方，让他住在他们中间。
JOSH|20|5|若是报血仇者追上了他，长老不可把他交在报血仇者的手里，因为他是无意中杀了邻舍的，并非过去彼此之间有仇恨。
JOSH|20|6|他要住在那城里，直到他站在会众面前受审判；等到当时的大祭司死后，杀人者才可以回到本城本家，就是他所逃出来的那城。’”
JOSH|20|7|于是， 以色列 人划分 拿弗他利 山区 加利利 的 基低斯 、 以法莲 山区的 示剑 和 犹大 山区的 基列．亚巴 ， 基列．亚巴 就是 希伯仑 。
JOSH|20|8|他们在 约旦河 的另一边，就是 耶利哥 的东边，从 吕便 支派中，在旷野的平原设立 比悉 ，从 迦得 支派中设立 基列 的 拉末 ，从 玛拿西 支派中设立 巴珊 的 哥兰 。
JOSH|20|9|这都是为 以色列 众人和在他们中间寄居的外人所指定的城镇，使凡误杀人者可以逃到那里，不至于死在报血仇者的手中，直到他站在会众面前受审判 。
JOSH|21|1|利未 人的众族长近前来到 以利亚撒 祭司和 嫩 的儿子 约书亚 ，以及 以色列 人各支派父系的领袖那里，
JOSH|21|2|在 迦南 地的 示罗 对他们说：“从前耶和华曾藉着 摩西 吩咐给我们城镇居住，以及城镇的郊外供我们牧养牲畜。”
JOSH|21|3|于是 以色列 人照耶和华的指示，从自己的地业中，把这些城镇和城镇的郊外给了 利未 人。
JOSH|21|4|哥辖 族抽了签。 利未 人中 亚伦 祭司的子孙，从 犹大 支派、 西缅 支派、 便雅悯 支派的地业中，抽签得了十三座城。
JOSH|21|5|哥辖 其余的子孙，从 以法莲 支派、 但 支派、 玛拿西 半支派宗族的地业中，抽签得了十座城。
JOSH|21|6|革顺 的子孙，从 以萨迦 支派、 亚设 支派、 拿弗他利 支派、住 巴珊 的 玛拿西 半支派宗族的地业中，抽签得了十三座城。
JOSH|21|7|米拉利 的子孙，按着宗族，从 吕便 支派、 迦得 支派、 西布伦 支派的地业中，得了十二座城。
JOSH|21|8|以色列 人照耶和华藉 摩西 所吩咐的，把这些城镇和城镇的郊外，抽签给 利未 人。
JOSH|21|9|他们从 犹大 支派和 西缅 支派的地业中，给了以下所记名字的各城，
JOSH|21|10|就是给 利未 人 哥辖 宗族的 亚伦 子孙，因为他们抽到第一签：
JOSH|21|11|把 犹大 山区的 基列．亚巴 ，就是 希伯仑 ，和四围的郊野给了他们。 亚巴 是 亚衲 族的祖先。
JOSH|21|12|但是，这城的田地和所属的村庄却给了 耶孚尼 的儿子 迦勒 为业。
JOSH|21|13|他们把 希伯仑 ，就是误杀人的逃城和城的郊外，给了 亚伦 祭司的子孙；又给了 立拿 和城的郊外、
JOSH|21|14|雅提珥 和城的郊外、 以实提莫 和城的郊外、
JOSH|21|15|何仑 和城的郊外、 底璧 和城的郊外、
JOSH|21|16|亚因 和城的郊外、 淤他 和城的郊外，以及 伯．示麦 和城的郊外，共九座城，都是从这二支派中分出来的。
JOSH|21|17|又从 便雅悯 支派的地业中给了 基遍 和城的郊外、 迦巴 和城的郊外、
JOSH|21|18|亚拿突 和城的郊外，以及 亚勒们 和城的郊外，共四座城。
JOSH|21|19|亚伦 子孙作祭司的共有十三座城，以及城的郊外。
JOSH|21|20|利未 人 哥辖 的宗族，就是 哥辖 其余的子孙，抽签所得的城是从 以法莲 支派来的。
JOSH|21|21|他们把 以法莲 山区的 示剑 ，就是误杀人的逃城和城的郊外给了 哥辖 其余的子孙；又给了 基色 和城的郊外、
JOSH|21|22|基伯先 和城的郊外，以及 伯．和仑 和城的郊外，共四座城。
JOSH|21|23|又从 但 支派的地业中给了 伊利提基 和城的郊外、 基比顿 和城的郊外、
JOSH|21|24|亚雅仑 和城的郊外，以及 迦特．临门 和城的郊外，共四座城。
JOSH|21|25|又从 玛拿西 半支派的地业中给了 他纳 和城的郊外，以及 迦特．临门 和城的郊外，共两座城。
JOSH|21|26|哥辖 其余的子孙共有十座城，以及城的郊外。
JOSH|21|27|利未 人宗族中 革顺 的子孙，从 玛拿西 半支派的地业中所得的是 巴珊 的 哥兰 ，就是误杀人的逃城和城的郊外，以及 比．施提拉 和城的郊外，共两座城。
JOSH|21|28|从 以萨迦 支派的地业中所得的是 基善 和城的郊外、 大比拉 和城的郊外、
JOSH|21|29|耶末 和城的郊外，以及 隐．干宁 和城的郊外，共四座城。
JOSH|21|30|从 亚设 支派的地业中所得的是 米沙勒 和城的郊外、 押顿 和城的郊外、
JOSH|21|31|黑甲 和城的郊外，以及 利合 和城的郊外，共四座城。
JOSH|21|32|从 拿弗他利 支派的地业中所得的是 加利利 的 基低斯 ，就是误杀人的逃城和城的郊外、 哈末．多珥 和城的郊外，以及 加珥坦 和城的郊外，共三座城。
JOSH|21|33|革顺 人按着宗族共有十三个城，以及城的郊外。
JOSH|21|34|其余的 利未 人，就是 米拉利 的子孙，按着宗族从 西布伦 支派的地业中所得的是 约念 和城的郊外、 加珥他 和城的郊外、
JOSH|21|35|丁拿 和城的郊外，以及 拿哈拉 和城的郊外，共四座城。
JOSH|21|36|从 吕便 支派的地业中所得的是 比悉 和城的郊外、 雅杂 和城的郊外、
JOSH|21|37|基底莫 和城的郊外，以及 米法押 和城的郊外，共四座城。
JOSH|21|38|从 迦得 支派的地业中所得的是 基列 的 拉末 ，就是误杀人的逃城和城的郊外、 玛哈念 和城的郊外、
JOSH|21|39|希实本 和城的郊外，以及 雅谢 和城的郊外，共四座城。
JOSH|21|40|利未 宗族其余的人，就是 米拉利 的子孙，按着宗族抽签所得的，共十二座城。
JOSH|21|41|利未 人在 以色列 人的地业中所得的城，共四十八个，还有城的郊外。
JOSH|21|42|这些城的四围都有郊野，每个城都是如此。
JOSH|21|43|这样，耶和华将从前向他们列祖起誓要给他们的全地赐给 以色列 人，他们就得了为业，住在其中。
JOSH|21|44|耶和华照着向他们列祖起誓所应许的一切，赐给他们全境安宁。他们所有的仇敌，没有一个能在他们面前站立得住。耶和华把所有仇敌都交在他们手中。
JOSH|21|45|耶和华应许赐福给 以色列 家的话，一句都没有落空，全都应验了。
JOSH|22|1|此后， 约书亚 召了 吕便 人、 迦得 人和 玛拿西 半支派的人来，
JOSH|22|2|对他们说：“耶和华的仆人 摩西 所吩咐你们的，你们都遵守了；我吩咐你们的话，你们也都听从了。
JOSH|22|3|你们这许多日子，都没有撇弃你们的弟兄，直到今日，并且遵守了耶和华你们上帝所吩咐的命令。
JOSH|22|4|如今耶和华－你们的上帝已经照着他所应许的，使你们的弟兄得享安宁。你们现在可以返回自己的帐棚，回到耶和华的仆人 摩西 在 约旦河 东所赐给你们为业之地。
JOSH|22|5|只是务要谨守遵行耶和华的仆人 摩西 所吩咐你们的诫命和律法，爱耶和华－你们的上帝，行他一切的道，守他的诫命，紧紧跟随他，尽心尽性事奉他。”
JOSH|22|6|于是 约书亚 为他们祝福，送他们回去，他们就回到自己的帐棚去了。
JOSH|22|7|摩西 在 巴珊 曾把地业分给 玛拿西 的半支派；然后 约书亚 在 约旦河 的西岸，在他们弟兄中，又把地业分给 玛拿西 的另外半支派。 约书亚 送他们回帐棚的时候，为他们祝福，
JOSH|22|8|对他们说：“你们要把许多财物，许多牲畜，和金、银、铜、铁，以及许多衣服，带回你们的帐棚去，要把你们从仇敌夺来的东西分给你们的众弟兄。”
JOSH|22|9|于是 吕便 人、 迦得 人、 玛拿西 半支派的人从 迦南 地的 示罗 起行，离开 以色列 人，回到他们已得为业的 基列 地，就是他们照耶和华藉 摩西 所吩咐而得的。
JOSH|22|10|吕便 人、 迦得 人和 玛拿西 半支派的人到了 迦南 地的 约旦河 一带地方，就在 约旦河 那里筑了一座坛，一座高大壮观的坛。
JOSH|22|11|以色列 人听见了，说：“看哪， 吕便 人、 迦得 人、 玛拿西 半支派的人在 迦南 地对面， 约旦河 一带地方， 以色列 人的境内，筑了一座坛。”
JOSH|22|12|以色列 人一听见，全会众的 以色列 人就聚集在 示罗 ，要上去攻打他们。
JOSH|22|13|以色列 人派 以利亚撒 祭司的儿子 非尼哈 ，往 基列 地，到 吕便 人、 迦得 人和 玛拿西 半支派的人那里。
JOSH|22|14|和他同去的还有十个领袖， 以色列 每个支派在父家中各派一个领袖，这些人每一个在 以色列 族系中都是父家的领袖。
JOSH|22|15|他们来到 基列 地，到 吕便 人、 迦得 人和 玛拿西 半支派的人那里，对他们说：
JOSH|22|16|“耶和华全会众这样说：‘你们今日离弃耶和华不跟从他，干犯 以色列 的上帝，悖逆耶和华，为自己筑了一座坛，你们所犯的是何等的罪！
JOSH|22|17|从前我们在 毗珥 犯的罪孽，导致瘟疫临到耶和华的会众，甚至到今日都还没有洗净，这还算小事吗？
JOSH|22|18|你们今日竟然离弃耶和华不跟从他！你们今日既然悖逆耶和华，明日他必向 以色列 全会众发怒。
JOSH|22|19|若你们认为所得为业之地不洁净，可以过来，到耶和华之地，就是耶和华的帐幕所居住之地，在我们中间得地业。你们却不可悖逆耶和华，也不可背叛我们，在耶和华－我们上帝的坛以外为自己筑坛。
JOSH|22|20|从前 谢拉 的曾孙 亚干 岂不是在那当灭的物上犯了罪，导致愤怒临到 以色列 全会众吗？死在他所犯的罪中的，不只是他一个人而已！’”
JOSH|22|21|于是 吕便 人、 迦得 人、 玛拿西 半支派的人回答 以色列 族系的领袖，说：
JOSH|22|22|“大能者上帝耶和华！大能者上帝耶和华！他已知道，愿 以色列 人也知道，我们若有悖逆的行为，或是干犯耶和华，你今日就不要让我们活着！
JOSH|22|23|若我们为自己筑坛，离弃耶和华不跟从他，或将燔祭、素祭、平安祭献在坛上，愿耶和华亲自追究。
JOSH|22|24|不是这样！我们做这事的原因是惧怕将来你们的子孙对我们的子孙说：‘你们与耶和华－ 以色列 的上帝有什么关系呢？
JOSH|22|25|因为耶和华以 约旦河 作我们和你们 吕便 人、 迦得 人的交界，所以你们在耶和华里无份。’这样，你们的子孙就使我们的子孙不再敬畏耶和华了。
JOSH|22|26|因此我们说：‘不如为自己筑一座坛，不是为献燔祭，也不是为献别样的祭，
JOSH|22|27|而是为你我之间和后代子孙之间作证据，好使我们也在耶和华面前献我们的燔祭、平安祭和别样的祭来事奉他，免得你们的子孙将来对我们的子孙说，你们在耶和华里无份。’
JOSH|22|28|所以我们说：‘将来他们若对我们，或对我们的子孙这样说，我们就可以回答说：你们看，我们列祖所筑的坛是耶和华坛的样式，这并不是为献燔祭，也不是为献别样的祭，而是作为你们和我们之间的证据。’
JOSH|22|29|除了耶和华－我们上帝帐幕前的坛以外，我们绝没有意思要为着献燔祭、素祭和别样的祭而另外筑一座坛，悖逆耶和华，今日离弃不跟从他。”
JOSH|22|30|非尼哈 祭司与会众中的领袖，就是与他同来那些 以色列 族系的领袖，听见 吕便 人、 迦得 人、 玛拿西 人所说的话，就都看为美。
JOSH|22|31|以利亚撒 祭司的儿子 非尼哈 对 吕便 人、 迦得 人、 玛拿西 人说：“今日我们知道耶和华在我们中间，因为你们没有向他犯悖逆的罪。现在你们把 以色列 人从耶和华的手中救出来了。”
JOSH|22|32|以利亚撒 祭司的儿子 非尼哈 与众领袖离开了 吕便 人和 迦得 人，从 基列 地回 迦南 地，到了 以色列 人那里，就把这事向他们回报。
JOSH|22|33|以色列 人看这事为美； 以色列 人就称颂上帝，不再说要上去攻打 吕便 人和 迦得 人，毁坏他们所住的地了。
JOSH|22|34|吕便 人和 迦得 人给这坛起了名，因为这坛在我们之间见证耶和华是上帝。
JOSH|23|1|耶和华使 以色列 人从四围所有的仇敌中得享安宁，已经有很多日子了。 约书亚 年纪老迈，
JOSH|23|2|就召了全 以色列 的众长老、领袖、审判官和官长来，对他们说：“我年纪已经老迈。
JOSH|23|3|耶和华－你们的上帝因你们的缘故向这些国家所做的一切，你们都亲眼看见了，那为你们作战的是耶和华－你们的上帝。
JOSH|23|4|看，我已经把所剩下的列国，连同从 约旦河 起到 大海 日落的方向，我所剪除的列国，都抽签分给你们各支派为业了。
JOSH|23|5|耶和华－你们的上帝必将他们从你们面前赶出去，使他们离开你们，你们就必得他们的地为业，正如耶和华－你们的上帝向你们所应许的。
JOSH|23|6|你们要大大壮胆，谨守遵行写在 摩西 律法书上的一切话，不可偏离左右。
JOSH|23|7|不可与你们中间所剩下的这些国家往来。你们不可提他们神明的名，不可指着它们起誓，不可事奉它们，也不可敬拜它们。
JOSH|23|8|只要紧紧跟随耶和华－你们的上帝，就像你们直到今日所做的。
JOSH|23|9|因为耶和华已经把又大又强的列国从你们面前赶出；直到今日，没有一人能在你们面前站立得住。
JOSH|23|10|你们一人必追赶千人，因为耶和华－你们的上帝照他向你们所应许的，为你们作战。
JOSH|23|11|你们要分外谨慎，爱耶和华－你们的上帝。
JOSH|23|12|你们若断然转离，紧紧跟随你们中间所剩下的这些国家，彼此结亲，互相往来，
JOSH|23|13|就要确实知道，耶和华－你们的上帝必不再将他们从你们面前赶出；他们却要成为你们的罗网、圈套、肋上的鞭、眼中的刺，直到你们在耶和华－你们上帝所赐的这美地上灭亡。
JOSH|23|14|“看哪，我今日要走世人必走的路了。你们要一心一意知道，耶和华－你们上帝所应许要赐给你们的一切福气，没有一件落空，都应验在你们身上了。
JOSH|23|15|耶和华－你们的上帝所应许的一切福气怎样临到你们身上，耶和华也必照样使各样灾祸临到你们身上，直到他把你们从耶和华－你们上帝所赐给你们的这美地上除灭。
JOSH|23|16|你们若违背耶和华－你们上帝吩咐你们所守的约，去事奉别神，敬拜它们，耶和华的怒气必向你们发作，使你们在他所赐给你们的美地上迅速灭亡。”
JOSH|24|1|约书亚 召集 以色列 的众支派到 示剑 ，他召了 以色列 的长老、领袖、审判官和官长来；他们都站在上帝面前。
JOSH|24|2|约书亚 对众百姓说：“耶和华－ 以色列 的上帝如此说：‘古时你们的列祖，就是 亚伯拉罕 和 拿鹤 的父亲 他拉 ，住在 大河 那边事奉别神。
JOSH|24|3|我将你们的祖宗 亚伯拉罕 从 大河 那边带出来，领他走遍 迦南 全地，又使他的子孙众多。我把 以撒 赐给他，
JOSH|24|4|我又把 雅各 和 以扫 赐给 以撒 ，将 西珥山 赐给 以扫 为业。但 雅各 和他的子孙下到 埃及 去了。
JOSH|24|5|我差遣 摩西 和 亚伦 ，照我在 埃及 中间所做的，降灾与 埃及 ，然后把你们领出来。
JOSH|24|6|我领你们的祖宗出 埃及 ，你们就到了 红海 。 埃及 人带领战车骑兵，追赶你们的祖宗到 红海 。
JOSH|24|7|你们的祖宗哀求耶和华，他就用黑暗把你们和 埃及 人隔开了，又使海水冲向 埃及 人，淹没他们。我在 埃及 所做的，你们都亲眼见过。你们在旷野住了很多日子。
JOSH|24|8|我领你们到 约旦河 东 亚摩利 人所住之地。他们与你们争战，我把他们交在你们手中，你们就得了他们的地为业。我也在你们面前灭绝他们。
JOSH|24|9|那时， 摩押 王 西拨 的儿子 巴勒 起来攻击 以色列 人，派人去召 比珥 的儿子 巴兰 来诅咒你们。
JOSH|24|10|但我不愿听 巴兰 ，所以他反而为你们连连祝福。这样，我救了你们脱离他的手。
JOSH|24|11|你们过了 约旦河 ，来到 耶利哥 。 耶利哥 人、 亚摩利 人、 比利洗 人、 迦南 人、 赫 人、 革迦撒 人、 希未 人、 耶布斯 人都与你们争战，我却把他们交在你们手里。
JOSH|24|12|我派遣瘟疫 在你们前面，将 亚摩利 人的两个王从你们面前赶出，并不是用你的刀，也不是用你的弓。
JOSH|24|13|我赐给你们的地，不是你们开垦的；我赐给你们的城镇，不是你们建造的。你们却住在其中，又得吃那不是你们栽植的葡萄园和橄榄园的果子。’
JOSH|24|14|“现在你们要敬畏耶和华，诚心诚意事奉他，除掉你们列祖在 大河 那边和在 埃及 事奉的神明，事奉耶和华。
JOSH|24|15|若你们认为事奉耶和华不好，今日就可以选择所要事奉的：是你们列祖在 大河 那边所事奉的神明，或是你们所住这地 亚摩利 人的神明呢？至于我和我家，我们必定事奉耶和华。”
JOSH|24|16|百姓回答说：“我们绝不离弃耶和华去事奉别神。
JOSH|24|17|因为耶和华－我们的上帝曾领我们和我们的祖宗从 埃及 地为奴之家出来，在我们眼前行了那些大神迹，并在我们所行的一切路上，和所经过的各民族中保护了我们。
JOSH|24|18|耶和华又把各民族和住此地的 亚摩利 人都从我们面前赶出去。所以，我们也必事奉耶和华，因为他是我们的上帝。”
JOSH|24|19|约书亚 对百姓说：“你们不能事奉耶和华，因为他是神圣的上帝，是忌邪 的上帝，必不赦免你们的过犯罪恶。
JOSH|24|20|你们若离弃耶和华去事奉外邦的神明，耶和华在降福之后，必转而降祸给你们，把你们灭绝。”
JOSH|24|21|百姓对 约书亚 说：“不，我们要事奉耶和华。”
JOSH|24|22|约书亚 对百姓说：“你们选择耶和华，要事奉他，你们自己作证吧！”他们说：“我们愿意作证。”
JOSH|24|23|“现在，你们要除掉你们中间外邦的神明，专心归向耶和华－ 以色列 的上帝。”
JOSH|24|24|百姓对 约书亚 说：“我们必事奉耶和华－我们的上帝，听从他的话。”
JOSH|24|25|那日， 约书亚 就与百姓立约，在 示剑 为他们制定律例典章。
JOSH|24|26|约书亚 把这些话写在上帝的律法书上，又拿一块大石头立在橡树下耶和华圣所的旁边。
JOSH|24|27|约书亚 对众百姓说：“看哪，这石头可以向我们作见证，因为它听见了耶和华所吩咐我们的一切话；这石头将向你们作见证，免得你们背叛你们的上帝。”
JOSH|24|28|于是 约书亚 解散百姓，各自回到自己的地业去了。
JOSH|24|29|这些事以后，耶和华的仆人， 嫩 的儿子 约书亚 死了，那时他一百一十岁。
JOSH|24|30|以色列 人把他葬在他自己地业的境内， 以法莲 山区的 亭拿．西拉 ，在 迦实山 的北边。
JOSH|24|31|约书亚 在世的日子和他死了以后，那些知道耶和华为 以色列 所做一切事的长老还在世的时候， 以色列 人事奉耶和华。
JOSH|24|32|以色列 人把从 埃及 所带来 约瑟 的骸骨安葬在 示剑 ，就是 雅各 从前用一百可锡塔 向 示剑 的父亲 哈抹 的众子所买的那块地；这块地就成了 约瑟 子孙的产业。
JOSH|24|33|亚伦 的儿子 以利亚撒 也死了，他们把他葬在他儿子 非尼哈 所得 以法莲 山区的小山上 。
JUDG|1|1|约书亚 死后， 以色列 人求问耶和华说：“我们中间谁当首先上去攻打 迦南 人，与他们争战呢？”
JUDG|1|2|耶和华说：“ 犹大 要先上去。看哪，我已将那地交在他手中。”
JUDG|1|3|犹大 对他哥哥 西缅 说：“请你同我上到我抽签所得之地，与 迦南 人争战；我也同你去你抽签所得之地。”于是 西缅 与他同去。
JUDG|1|4|犹大 就上去，耶和华把 迦南 人和 比利洗 人交在他们手中。他们在 比色 击杀了一万人。
JUDG|1|5|他们在 比色 遇见 亚多尼．比色 ，与他争战，击败了 迦南 人和 比利洗 人。
JUDG|1|6|亚多尼．比色 逃跑，他们追赶他，捉住他，砍断他大拇指和大脚趾。
JUDG|1|7|亚多尼．比色 说：“从前有七十个王，大拇指和大脚趾都被我砍断，在我桌子底下拾取零碎食物。现在上帝照着我所做的报应我了。”他们把 亚多尼．比色 带到 耶路撒冷 ，他就死在那里。
JUDG|1|8|犹大 人攻打 耶路撒冷 ，夺取了它，用刀杀城内的人，并且放火烧城。
JUDG|1|9|后来 犹大 人下去，与住山区、 尼革夫 和低地的 迦南 人争战。
JUDG|1|10|犹大 去攻打住 希伯仑 的 迦南 人，杀了 示筛 、 亚希幔 、 挞买 。 希伯仑 从前名叫 基列．亚巴 。
JUDG|1|11|犹大 从那里去攻击 底壁 的居民。 底壁 从前名叫 基列．西弗 。
JUDG|1|12|迦勒 说：“谁能攻打 基列．西弗 ，夺取那城，我就把我女儿 押撒 嫁给他。”
JUDG|1|13|迦勒 的弟弟 基纳斯 的儿子 俄陀聂 夺取了那城， 迦勒 就把女儿 押撒 嫁给他。
JUDG|1|14|押撒 来的时候，催促丈夫 向她父亲要一块田。 押撒 一下驴， 迦勒 就对她说：“你要什么？”
JUDG|1|15|她对 迦勒 说：“求你赐我福分；你既然把 尼革夫 给了我，求你也给我水泉。” 迦勒 就把上泉和下泉都赐给她。
JUDG|1|16|摩西 的岳父是 基尼 人，他的子孙与 犹大 人一起上到棕树城，往 亚拉得 以南的 犹大 旷野 去，住在百姓当中 。
JUDG|1|17|犹大 和他哥哥 西缅 同去，击杀了住 洗法 的 迦南 人，将城彻底毁灭。因此，那城名叫 何珥玛 。
JUDG|1|18|犹大 攻取了 迦萨 和所属的领土， 亚实基伦 和所属的领土， 以革伦 和所属的领土。
JUDG|1|19|耶和华与 犹大 同在， 犹大 取得了山区，却不能赶出平原的居民，因为他们有铁的战车。
JUDG|1|20|以色列 人照 摩西 所说的，把 希伯仑 给了 迦勒 。 迦勒 从那里赶出 亚衲 的三支后裔。
JUDG|1|21|至于住 耶路撒冷 的 耶布斯 人， 便雅悯 人没有把他们赶出。于是， 耶布斯 人与 便雅悯 人同住在 耶路撒冷 ，直到今日。
JUDG|1|22|约瑟 家也上到 伯特利 去，耶和华与他们同在。
JUDG|1|23|约瑟 家去窥探 伯特利 ，那城起先名叫 路斯 。
JUDG|1|24|探子看见一个人从城里出来，就对他说：“请你把进城的路指示我们，我们会厚待你。”
JUDG|1|25|那人把进城的路指示他们。他们就用刀击杀了城中的居民，却放走那人和他的全家。
JUDG|1|26|那人往 赫 人之地去，建造了一座城，起名叫 路斯 。那城到如今还叫这名。
JUDG|1|27|玛拿西 没有赶出 伯˙善 和所属乡镇 的居民， 他纳 和所属乡镇的居民， 多珥 和所属乡镇的居民， 以伯莲 和所属乡镇的居民， 米吉多 和所属乡镇的居民； 迦南 人仍坚持住在这地。
JUDG|1|28|以色列 强盛的时候，就叫 迦南 人做苦工，没有把他们全然赶走。
JUDG|1|29|以法莲 没有赶出住 基色 的 迦南 人。于是 迦南 人仍住在 基色 ，在 以法莲 中间。
JUDG|1|30|西布伦 没有赶出 基伦 的居民和 拿哈拉 的居民。于是 迦南 人仍住在 西布伦 中间，成了服劳役的人。
JUDG|1|31|亚设 没有赶出 亚柯 的居民和 西顿 的居民，以及 亚黑拉 、 亚革悉 、 黑巴 、 亚弗革 和 利合 的居民。
JUDG|1|32|亚设 人因为没有赶出那地的居民 迦南 人，就住在他们中间。
JUDG|1|33|拿弗他利 没有赶出 伯˙示麦 和 伯˙亚纳 的居民。于是 拿弗他利 就住在那地的居民 迦南 人中，而 伯˙示麦 和 伯˙亚纳 的居民却成了为他们服劳役的人。
JUDG|1|34|亚摩利 人强逼 但 人住在山区，不准他们下到平原。
JUDG|1|35|亚摩利 人仍坚持住在 希烈山 、 亚雅仑 和 沙宾 ；然而 约瑟 家权势强盛的时候，他们成为服劳役的人。
JUDG|1|36|亚摩利 人 的地界是从 亚克拉滨 斜坡，从 西拉 延伸而上。
JUDG|2|1|耶和华的使者从 吉甲 上到 波金 ，说：“我领你们从 埃及 上来，带你们到我向你们列祖起誓应许之地。我曾说：‘我永不废弃我与你们的约。
JUDG|2|2|你们不可与这地的居民立约，要拆毁他们的祭坛。’你们竟没有听从我的话。你们为何这样做呢！
JUDG|2|3|因此我说：‘我必不将他们从你们面前赶出。他们必作你们肋下的荆棘 ，他们的神明必成为你们的圈套。’”
JUDG|2|4|耶和华的使者向 以色列 众人说这些话的时候，百姓放声大哭。
JUDG|2|5|于是他们给那地方起名叫 波金 ，并在那里向耶和华献祭。
JUDG|2|6|约书亚 解散百姓， 以色列 人回到自己的地业，占各自的地。
JUDG|2|7|约书亚 在世的日子和他死了以后，那些见过耶和华为 以色列 所做一切大事的长老还在世的时候，百姓都事奉耶和华。
JUDG|2|8|耶和华的仆人， 嫩 的儿子 约书亚 死了，那时他一百一十岁。
JUDG|2|9|以色列 人把他葬在他自己地业的境内， 以法莲 山区的 亭拿．希烈 ，在 迦实山 的北边。
JUDG|2|10|那世代的人也都归到自己的列祖。后来兴起的另一世代不认识耶和华，也不知道他为 以色列 所做的事。
JUDG|2|11|以色列 人行耶和华眼中看为恶的事，去事奉诸 巴力 。
JUDG|2|12|他们离弃领他们出 埃及 地的耶和华－他们列祖的上帝，去随从别神，就是四围列国的神明，向它们叩拜，惹耶和华发怒。
JUDG|2|13|他们离弃了耶和华，去事奉 巴力 和 亚斯她录 。
JUDG|2|14|耶和华的怒气向 以色列 发作，把他们交在抢夺他们的人手中，又把他们交给四围仇敌的手中 ，以致他们在仇敌面前再也不能站立得住。
JUDG|2|15|他们无论往何处去，耶和华的手都以灾祸攻击他们，正如耶和华所说的，又如耶和华向他们所起的誓；他们就极其困苦。
JUDG|2|16|耶和华兴起士师，士师就拯救他们脱离抢夺他们之人的手。
JUDG|2|17|然而，他们却不听从士师，竟随从别神而行淫，向它们叩拜。他们列祖所行的道，所听从耶和华的命令，他们都速速偏离了，并不照样遵行。
JUDG|2|18|耶和华为他们兴起士师，耶和华与士师同在。士师在世的一切日子，耶和华拯救他们脱离仇敌的手。耶和华因他们受欺压迫害所发出的哀声，就怜悯他们。
JUDG|2|19|但士师一死，他们又转去行恶，比他们祖宗更坏，去随从别神，事奉叩拜它们，总不放弃他们的恶习和顽梗的行为。
JUDG|2|20|于是耶和华的怒气向 以色列 发作，说：“因为这国违背我吩咐他们列祖当守的约，不听从我的话，
JUDG|2|21|约书亚 死的时候所剩下的各国，我必不再从他们面前赶出任何一个，
JUDG|2|22|为要藉此考验 以色列 是否肯谨守遵行耶和华的道，像他们列祖一样地谨守。”
JUDG|2|23|耶和华留下那些国家，不将他们速速赶出，也不把他们交在 约书亚 的手中。
JUDG|3|1|耶和华留下这些国家，为要考验所有未曾经历 迦南 任何战役的 以色列 人，
JUDG|3|2|只是为了要 以色列 人的后代认识战争，教导他们，尤其那些未曾认识这些事的人。
JUDG|3|3|留下的有 非利士 的五个领袖，所有的 迦南 人， 西顿 人，以及从 巴力．黑门山 到 哈马口 ，住 黎巴嫩山 的 希未 人。
JUDG|3|4|他们是为了要考验 以色列 ，好知道他们是否肯听从耶和华藉 摩西 吩咐他们列祖的命令。
JUDG|3|5|以色列 人住在 迦南 人、 赫 人、 亚摩利 人、 比利洗 人、 希未 人、 耶布斯 人中间，
JUDG|3|6|娶他们的女儿，将自己的女儿嫁给他们的儿子，并事奉他们的神明。
JUDG|3|7|以色列 人行耶和华眼中看为恶的事，忘记耶和华－他们的上帝，去事奉诸 巴力 和 亚舍拉 ，
JUDG|3|8|所以耶和华的怒气向 以色列 发作，把他们交给 美索不达米亚 王 古珊．利萨田 的手中。 以色列 人服事 古珊．利萨田 八年。
JUDG|3|9|以色列 人呼求耶和华，耶和华就为 以色列 人兴起一位拯救者来救他们，就是 迦勒 的弟弟 基纳斯 的儿子 俄陀聂 。
JUDG|3|10|耶和华的灵降在他身上，他就作了 以色列 的士师。他出去争战，耶和华将 亚兰 王 古珊．利萨田 交在他手中，他的手战胜了 古珊．利萨田 。
JUDG|3|11|于是这地太平四十年。 基纳斯 的儿子 俄陀聂 死了。
JUDG|3|12|以色列 人又行耶和华眼中看为恶的事。耶和华使 摩押 王 伊矶伦 强大，攻击 以色列 ，因为他们行耶和华眼中看为恶的事。
JUDG|3|13|伊矶伦 召集 亚扪 人和 亚玛力 人到他那里，他就去攻打 以色列 ，占据了棕树城。
JUDG|3|14|于是 以色列 人服事 摩押 王 伊矶伦 十八年。
JUDG|3|15|以色列 人呼求耶和华，耶和华就为他们兴起一位拯救者， 便雅悯 人 基拉 的儿子 以笏 ，他是个惯用左手的人 。 以色列 人托他送礼物给 摩押 王 伊矶伦 。
JUDG|3|16|以笏 打造了一把两刃的剑，长一短肘 ，绑在右腿上衣服里面。
JUDG|3|17|他把礼物献给 摩押 王 伊矶伦 。 伊矶伦 是个很肥胖的人。
JUDG|3|18|以笏 献完礼物的时候，就把抬礼物的人送走。
JUDG|3|19|但他自己却从靠近 吉甲 的雕像那里转回来，说：“王啊，我有一件机密的事要奏告你。”王说：“回避吧！”于是所有侍立在他左右的人都退去了。
JUDG|3|20|以笏 来到王那里，那时他独自一人坐在阴凉的顶楼。 以笏 说：“我有上帝的话向你报告。”王就从座位上站起来。
JUDG|3|21|以笏 伸出左手，从右腿上拔出剑来，刺入王的肚腹。
JUDG|3|22|剑柄连同剑刃都刺进去了，肥肉夹住了剑刃。他没有把剑从王的肚腹拔出来，粪便就流出来了 。
JUDG|3|23|以笏 出到门廊，把王关在楼门里面，就上了锁。
JUDG|3|24|以笏 出来之后，王的仆人就来了。他们观看，看哪，楼门锁住，就说：“他必是在阴凉的房间里大解。”
JUDG|3|25|他们等得不耐烦，看哪，楼门仍然不开，就拿钥匙打开楼门，看哪，他们的主人已经倒在地上死了。
JUDG|3|26|他们耽延的时候， 以笏 就逃跑了。他经过雕像那里，逃到 西伊拉 。
JUDG|3|27|他到了那里，就在 以法莲 山区吹角。 以色列 人跟随他从山区下来，他在他们前面引路，
JUDG|3|28|对他们说：“紧跟着我！因为耶和华已经把你们的仇敌 摩押 交在你们手中。”于是他们跟着他下去，占据了 摩押 对面 约旦河 的渡口，不准一人过去。
JUDG|3|29|那时，他们击杀了约一万 摩押 人，都是强壮的勇士，连一个也没有逃脱。
JUDG|3|30|那日， 摩押 在 以色列 手下制伏了。于是这地太平八十年。
JUDG|3|31|以笏 之后，有 亚拿 的儿子 珊迦 ，他用赶牛的棍子打死六百 非利士 人。他也拯救了 以色列 。
JUDG|4|1|以笏 死后， 以色列 人又行耶和华眼中看为恶的事。
JUDG|4|2|耶和华把他们交给在 夏琐 作王的 迦南 王 耶宾 手中；他的将军是 西西拉 ，住在 夏罗设．哈歌印 。
JUDG|4|3|以色列 人呼求耶和华，因为 耶宾 王有铁的战车九百辆，并且残酷欺压 以色列 人二十年。
JUDG|4|4|有一位女先知 底波拉 ，是 拉比多 的妻子，当时作 以色列 的士师。
JUDG|4|5|她住在 以法莲 山区 拉玛 和 伯特利 的中间，在 底波拉 的棕树下。 以色列 人都上到她那里去听审判。
JUDG|4|6|她派人从 拿弗他利 的 基低斯 把 亚比挪庵 的儿子 巴拉 召来，对他说：“耶和华－ 以色列 的上帝吩咐你：‘你要率领一万 拿弗他利 人和 西布伦 人上 他泊山 去。
JUDG|4|7|我必使 耶宾 的将军 西西拉 率领他的战车和全军往 基顺河 ，到你那里去，我必把他交在你手中。’”
JUDG|4|8|巴拉 对她说：“你若同我去，我就去；你若不同我去，我就不去。”
JUDG|4|9|底波拉 说：“我一定会与你同去，然而你在所行的路上必得不着荣耀，因为耶和华要把 西西拉 交给一个妇人的手里。”于是 底波拉 起来，与 巴拉 一同往 基低斯 去了。
JUDG|4|10|巴拉 召集 西布伦 人和 拿弗他利 人到 基低斯 ，跟他上去的有一万人。 底波拉 也同他上去。
JUDG|4|11|摩西 岳父 何巴 的后裔， 基尼 人 希百 离开了 基尼 族，到靠近 基低斯 的 撒拿音 橡树旁支搭帐棚。
JUDG|4|12|有人告诉 西西拉 ：“ 亚比挪庵 的儿子 巴拉 已经上了 他泊山 。”
JUDG|4|13|西西拉 就召集所有的铁战车九百辆和随从的全军，从 夏罗设．哈歌印 出来，到了 基顺河 。
JUDG|4|14|底波拉 对 巴拉 说：“起来，今日就是耶和华把 西西拉 交在你手中的日子。耶和华岂不在你前面行吗总”于是 巴拉 下了 他泊山 ，跟随他的有一万人。
JUDG|4|15|耶和华使 西西拉 和他一切的战车，以及全军溃乱，在 巴拉 面前倒在刀下。 西西拉 下了车，徒步逃跑。
JUDG|4|16|巴拉 追赶战车、军队，直到 夏罗设．哈歌印 。 西西拉 的全军都倒在刀下，一个也没有留下。
JUDG|4|17|只有 西西拉 徒步逃跑到 基尼 人 希百 之妻 雅亿 的帐棚，因为 夏琐 王 耶宾 与 基尼 人的 希百 家和平共处。
JUDG|4|18|雅亿 出来迎接 西西拉 ，对他说：“请我主进来，进到我这里来，不要怕。” 西西拉 就进了她的帐棚， 雅亿 用被子将他盖住。
JUDG|4|19|西西拉 对 雅亿 说：“我渴了，求你给我一点水喝。” 雅亿 就打开装奶的皮袋，给他喝，再把他盖住。
JUDG|4|20|西西拉 对 雅亿 说：“请你站在帐棚门口，若有人来问你说：‘有人在这里吗？’你就说：‘没有。’”
JUDG|4|21|西西拉 疲乏沉睡了。 希百 的妻 雅亿 取了帐棚的橛子，手拿着锤子，静悄悄地到他那里，将橛子从他的太阳穴钉进去，直钉到地里。 西西拉 就死了。
JUDG|4|22|看哪， 巴拉 追赶 西西拉 ， 雅亿 出来迎接他，对他说：“来，我给你看你要找的人。”他就进入帐棚，看哪， 西西拉 已经倒在地上死了，橛子还在他的太阳穴中。
JUDG|4|23|那日，上帝在 以色列 人面前制伏了 迦南 王 耶宾 。
JUDG|4|24|从此， 以色列 人的手对 迦南 王 耶宾 越来越强硬，直到将 迦南 王 耶宾 剪除。
JUDG|5|1|那日， 底波拉 和 亚比挪庵 的儿子 巴拉 唱歌，说：
JUDG|5|2|“ 以色列 有领袖率领 ， 百姓甘心牺牲自己， 你们当称颂耶和华！
JUDG|5|3|“君王啊，要听！王子啊，要侧耳！ 我要，我要向耶和华歌唱； 我要歌颂耶和华－ 以色列 的上帝。
JUDG|5|4|“耶和华啊，你从 西珥 出来， 从 以东 田野向前行， 地震动 天滴下， 云也滴下雨水。
JUDG|5|5|众山在耶和华面前摇动， 西奈山 在耶和华－ 以色列 上帝面前也摇动。
JUDG|5|6|“在 亚拿 之子 珊迦 的时候， 在 雅亿 的日子， 大道无人行走， 过路人绕道而行。
JUDG|5|7|以色列 农村荒芜， 空无一人， 直到我 底波拉 兴起， 兴起作 以色列 之母！
JUDG|5|8|以色列 人选择新的诸神， 战争就临到城门。 以色列 四万人中， 看得见盾牌枪矛吗？
JUDG|5|9|我心向往 以色列 的领袖， 他们在民中甘心牺牲自己。 你们应当称颂耶和华！
JUDG|5|10|“骑浅色母驴的、 坐绣花毯子的、 行走在路上的， 你们都当思想！
JUDG|5|11|打水的声音胜过弓箭的响声， 那里，人要述说耶和华公义的作为， 他对 以色列 乡民公义的作为。 “那时，耶和华的子民下到城门。
JUDG|5|12|“ 底波拉 啊，兴起！兴起！ 当兴起，兴起，唱歌！ 巴拉 啊，你当兴起！ 亚比挪庵 的儿子啊，当俘掳你的俘虏！
JUDG|5|13|那时，贵族中的幸存者前进， 耶和华的百姓为我前进攻击勇士。
JUDG|5|14|源自 亚玛力 的人从 以法莲 下来 ， 跟着你，你的族人 便雅悯 ； 有领袖从 玛吉 下来， 手握官员权杖的从 西布伦 下来。
JUDG|5|15|以萨迦 的领袖与 底波拉 一起； 巴拉 怎样， 以萨迦 也怎样； 他跟随 巴拉 冲下平原。 吕便 支派 有胸怀大志的人。
JUDG|5|16|你为何坐在羊圈内， 听羊群中吹笛的声音呢？ 吕便 支派具心有大谋的人。
JUDG|5|17|基列 安居在 约旦河 东。 但 为何住在船上呢？ 亚设 在海边居住， 它在港口安居。
JUDG|5|18|西布伦 是拚命敢死的百姓， 拿弗他利 在田野的高处也是如此。 　
JUDG|5|19|“君王都来争战； 那时 迦南 诸王在 米吉多 水旁的 他纳 争战， 却得不到掳掠的银钱。
JUDG|5|20|星宿从天上争战， 从它们的轨道攻击 西西拉 。
JUDG|5|21|基顺 的急流冲走他们， 古老的急流， 基顺 的急流。 我的灵啊，努力前进！
JUDG|5|22|“那时马蹄踢踏， 壮马奔驰飞腾。
JUDG|5|23|“耶和华的使者说：‘要诅咒 米罗斯 ， 重重诅咒其中的居民， 因为他们不来帮助耶和华， 不来帮助耶和华攻击壮士。’
JUDG|5|24|“愿 基尼 人 希百 的妻子 雅亿 比众妇人多得福气， 比帐棚中的妇人更蒙福祉。
JUDG|5|25|西西拉 求水， 雅亿 给他奶， 用贵重的碗装乳酪给他。
JUDG|5|26|雅亿 左手拿着帐棚的橛子， 右手拿着工匠的锤子， 击打 西西拉 ，打碎他的头， 打破穿透他的太阳穴。
JUDG|5|27|西西拉 在她脚下曲身，仆倒，躺卧， 在她脚下曲身，仆倒； 他在哪里曲身，就在哪里仆倒，死亡。
JUDG|5|28|“ 西西拉 的母亲从窗户里往外观看， 她在窗格子中哀号： ‘他的战车为何迟迟未归？ 他的车轮为何走得那么慢呢？’
JUDG|5|29|她聪明的宫女回答她， 她也自言自语说：
JUDG|5|30|‘或许他们得了战利品而分， 每个壮士得了一两个女子？ 西西拉 得了彩衣为掳物， 得了绣花的彩衣为掠物， 这两面绣花的彩衣， 披在颈项上作为战利品。’
JUDG|5|31|“耶和华啊，愿你的仇敌都这样灭亡！ 愿爱你的人如太阳上升，大发光辉！” 于是这地太平四十年。
JUDG|6|1|以色列 人又行耶和华眼中看为恶的事，耶和华就把他们交在 米甸 手里七年。
JUDG|6|2|米甸 的手战胜 以色列 ； 以色列 人躲避 米甸 人，就在山中挖洞穴，挖洞建营寨。
JUDG|6|3|每当 以色列 人撒种之后， 米甸 、 亚玛力 和东边的人都上来攻打他们，
JUDG|6|4|对着他们安营，毁坏那地的农作物，直到 迦萨 ，没有给 以色列 留下食物，牛、羊、驴也没有留下。
JUDG|6|5|因为那些人带着他们的牲畜和帐棚上来，像蝗虫那样多；人和骆驼无数，都进入境内，毁坏全地。
JUDG|6|6|以色列 因 米甸 的缘故极其穷乏， 以色列 人就呼求耶和华。
JUDG|6|7|以色列 人因 米甸 的缘故呼求耶和华的时候，
JUDG|6|8|耶和华就差遣先知到 以色列 人那里，对他们说：“耶和华－ 以色列 的上帝如此说：‘我曾领你们从 埃及 上来，从为奴之家出来，
JUDG|6|9|救你们脱离 埃及 人的手，脱离一切欺压你们之人的手。我从你们面前赶出他们，把他们的地赐给你们。
JUDG|6|10|我对你们说，我是耶和华－你们的上帝。你们住在 亚摩利 人的地，不可敬畏他们的神明，但你们却不听从我的话。’”
JUDG|6|11|耶和华的使者到了 俄弗拉 ，坐在 亚比以谢 族 约阿施 的橡树下。 约阿施 的儿子 基甸 正在醡酒池那里打麦子，为了躲避 米甸 人。
JUDG|6|12|耶和华的使者向 基甸 显现，对他说：“大能的勇士啊，耶和华与你同在！”
JUDG|6|13|基甸 对他说：“主啊，请容许我说，耶和华若与我们同在，我们怎么会遭遇这一切事呢？我们的列祖告诉我们：‘耶和华领我们从 埃及 上来’，他那奇妙的作为在哪里呢？现在耶和华却丢弃了我们，把我们交在 米甸 人的手掌中。”
JUDG|6|14|耶和华转向 基甸 ，说：“去，靠着你这能力拯救 以色列 脱离 米甸 人的手掌。我岂不是已经差遣了你吗？”
JUDG|6|15|基甸 对他说：“主啊，请容许我说，我怎能拯救 以色列 呢？看哪，我这一支在 玛拿西 支派中是最贫寒的，我在我父家又是最微小的。”
JUDG|6|16|耶和华对他说：“我与你同在，你就必击败 米甸 ，如击打一个人。”
JUDG|6|17|基甸 对他说：“我若在你眼前蒙恩，求你给我一个证据，证明是你在跟我说话。
JUDG|6|18|求你不要离开这里，等我回来，将供物带来，供在你面前。”他说：“我必等你回来。”
JUDG|6|19|基甸 去预备一只小山羊，用一伊法细面做了无酵饼，将肉放在篮子里，将汤盛在壶中，带到他那里，在橡树下献上。
JUDG|6|20|上帝的使者对 基甸 说：“将肉和无酵饼放在这磐石上，把汤倒出来。”他就照样做了。
JUDG|6|21|耶和华的使者伸出手里的杖，杖头一碰到肉和无酵饼，就有火从磐石中出来，吞灭了肉和无酵饼。耶和华的使者就从他眼前消失了。
JUDG|6|22|基甸 见他是耶和华的使者，就说：“哎呀！主耶和华啊！因为我真的面对面看见了耶和华的使者。”
JUDG|6|23|耶和华对他说：“安心吧，不要怕，你不会死。”
JUDG|6|24|于是 基甸 在那里为耶和华筑了一座坛，起名叫“耶和华沙龙” 。这坛至今还在 亚比以谢 族的 俄弗拉 。
JUDG|6|25|那夜，耶和华对 基甸 说：“你要把你父亲的公牛，就是 那七岁的第二头公牛取来，并拆毁你父亲为 巴力 筑的坛，砍下坛旁的 亚舍拉 ，
JUDG|6|26|在这堡垒顶上整整齐齐地为耶和华－你的上帝筑一座坛，将第二头公牛献为燔祭，用你所砍下的 亚舍拉 当柴。”
JUDG|6|27|基甸 就从他仆人中选了十个人，照耶和华吩咐他的做了。他因怕父家和本城的人，不敢在白天做这事，就在夜间做。
JUDG|6|28|城里的人清早起来，看哪， 巴力 的坛被拆毁，坛旁的 亚舍拉 被砍下，第二头公牛献在筑好的坛上，
JUDG|6|29|就彼此问：“这是谁做的事呢？”他们寻找查访之后，就说：“这是 约阿施 的儿子 基甸 做的事。”
JUDG|6|30|城里的人对 约阿施 说：“把你的儿子交出来，我们要处死他，因为他拆毁了 巴力 的坛，砍下了坛旁的 亚舍拉 。”
JUDG|6|31|约阿施 对站着敌对他的众人说：“你们是为 巴力 辩护吗？你们要救它吗？谁为它辩护，就在早晨把谁处死吧！ 巴力 如果是上帝，有人拆毁了它的坛，就让它为自己辩护吧！”
JUDG|6|32|所以那日人称 基甸 为 耶路巴力 ，意思是：“他拆毁了 巴力 的坛，让 巴力 与他争辩吧。”
JUDG|6|33|那时，所有的 米甸 人、 亚玛力 人和东边的人都聚集在一起，过了河，在 耶斯列 平原安营。
JUDG|6|34|耶和华的灵降在 基甸 身上；他吹角， 亚比以谢 族都聚集跟随他。
JUDG|6|35|他派使者走遍 玛拿西 ， 玛拿西 人也聚集跟随他。他又派使者到 亚设 、 西布伦 、 拿弗他利 ，他们也都上来会合。
JUDG|6|36|基甸 对上帝说：“你如果真的照你所说的，藉我的手拯救 以色列 ，
JUDG|6|37|看哪，我把一团羊毛放在禾场上，若单是羊毛上有露水，遍地都是干的，我就知道你必照你所说的，藉我的手拯救 以色列 。”
JUDG|6|38|一切果然发生了。次日早晨 基甸 起来，把羊毛拧一拧，从羊毛中挤出露水来，装满一碗的水。
JUDG|6|39|基甸 又对上帝说：“求你不要向我发怒，我再说一次，让我用羊毛再试一次，但愿羊毛是干的，遍地都有露水。”
JUDG|6|40|这夜，上帝也照样做，遍地都有露水，只有羊毛是干的。
JUDG|7|1|耶路巴力 ，就是 基甸 ，和所有跟随他的人早晨起来，在 哈律泉 旁安营。 米甸 营在他北边，靠近 摩利冈 的平原。
JUDG|7|2|耶和华对 基甸 说：“跟随你的人太多，我不能把 米甸 交在他们手中，免得 以色列 向我自夸，说：‘是我自己的手救了我。’
JUDG|7|3|现在你要向这百姓宣告说：‘凡惧怕战兢的，可以离开 基列山 回去。’”于是有二万二千人回去，只剩下一万人。
JUDG|7|4|耶和华对 基甸 说：“人还是太多。你要带他们下到水旁，我好在那里为你试试他们。我指着谁对你说：‘这人可以跟你去’，他就可以跟你去；我指着谁对你说：‘这人不可跟你去’，他就不可跟你去。”
JUDG|7|5|基甸 就带百姓下到水旁。耶和华对 基甸 说：“凡用舌头舔水像狗一样舔的，要使他单独站在一处；那些用双膝跪下喝水的，也要使他单独站在一处。”
JUDG|7|6|用手捧到嘴边舔水的数目有三百人，其余的百姓都用双膝跪下喝水。
JUDG|7|7|耶和华对 基甸 说：“我要用这舔水的三百人拯救你们，把 米甸 交在你手中；其余的百姓都可以各回自己的地方去。”
JUDG|7|8|百姓手里拿着食物和角；其余的 以色列 人， 基甸 都打发他们各自回到自己的帐棚，只留下这三百人。 米甸 营在他下边的平原上。
JUDG|7|9|那夜，耶和华对 基甸 说：“起来，下去攻营，因我已把它交在你手中。
JUDG|7|10|倘若你害怕下去，可以带你的仆人 普拉 下到那营里去，
JUDG|7|11|你必听见他们所说的，这样你的手就有力量下去攻营。”于是 基甸 带着仆人 普拉 下到军营里带着兵器的人边上。
JUDG|7|12|米甸 人、 亚玛力 人和所有东边的人都散布在平原，如同蝗虫那样多。他们的骆驼无数，多如海边的沙。
JUDG|7|13|基甸 到了那里，看哪，有一人把梦告诉同伴说：“看哪，我做了一个梦。看哪，一个大麦饼滚入 米甸 营中，来到帐幕，把帐幕撞倒，帐幕就翻转倒塌了。”
JUDG|7|14|同伴回答说：“这不是别的，而是 以色列 人 约阿施 的儿子 基甸 的刀。上帝已把 米甸 和全军都交在他手中了。”
JUDG|7|15|基甸 听见这梦的叙述和梦的解释，就敬拜上帝。他回到 以色列 营中，说：“起来吧！耶和华已把 米甸 军队交在你们手中了。”
JUDG|7|16|于是 基甸 将三百人分成三队，把角和空瓶交在每个人手中，瓶内有火把。
JUDG|7|17|他对他们说：“看着我，你们要照样做。看哪，我来到营边，我怎样做，你们也要照样做。
JUDG|7|18|我和所有跟随我的人吹角的时候，你们也要在营的四围吹角，喊叫：‘为耶和华！为 基甸 ！’”
JUDG|7|19|基甸 和跟随他的一百人，在半夜之初换岗哨的时候来到营旁。他们就吹角，打破手中的瓶；
JUDG|7|20|三队的人都吹角，打破瓶子。他们左手拿着火把，右手拿着吹的角，喊叫：“耶和华和 基甸 的刀！”
JUDG|7|21|他们围着军营，各人站在自己的地方；全营的人都逃窜，一面喊，一面逃跑。
JUDG|7|22|三百人就吹角，耶和华使全营的人用刀自相击杀。全营的人逃往 西利拉 的 伯．哈示他 ，一直逃到靠近 他巴 的 亚伯．米何拉 。
JUDG|7|23|从 拿弗他利 、 亚设 和 玛拿西 全地来的 以色列 人被召来，追赶 米甸 人。
JUDG|7|24|基甸 也派人走遍 以法莲 山区，说：“你们下来迎击 米甸 人，在他们的前面沿着 约旦河 把守渡口，直到 伯．巴拉 。”于是 以法莲 众人聚集，沿着 约旦河 把守渡口，直到 伯．巴拉 。
JUDG|7|25|他们捉住了 米甸 的两个领袖， 俄立 和 西伊伯 。他们在 俄立 磐石上杀了 俄立 ，在 西伊伯 酒池那里杀了 西伊伯 。他们追赶 米甸 人，把 俄立 和 西伊伯 的首级带到 约旦河 对岸，到 基甸 那里。
JUDG|8|1|以法莲 人对 基甸 说：“你去与 米甸 争战，没有召我们同去，你为什么这样待我们呢？”他们就和 基甸 激烈地争吵。
JUDG|8|2|基甸 对他们说：“我现在所做的怎么与你们所做的相比呢？ 以法莲 拾取剩下的葡萄不强过 亚比以谢 族所摘的葡萄吗？
JUDG|8|3|上帝已把 米甸 的两个领袖 俄立 和 西伊伯 交在你们手中；我所做的怎能与你们所做的相比呢？” 基甸 说了这话，他们对他的怒气就消了。
JUDG|8|4|基甸 和跟随他的三百人来到 约旦河 ，渡了过去；他们虽然疲乏，还是追赶。
JUDG|8|5|基甸 对 疏割 人说：“请你们拿几块饼来给跟随我的百姓，因为他们疲乏了。我正在追击 米甸 王 西巴 和 撒慕拿 。”
JUDG|8|6|疏割 人的领袖回答说：“ 西巴 和 撒慕拿 的手掌现在已经在你手里，因此我们该将饼送给你的军队吗？”
JUDG|8|7|基甸 说：“好吧！耶和华将 西巴 和 撒慕拿 交在我手之后，我必用旷野的荆棘和枳条鞭打你们。”
JUDG|8|8|基甸 从那里上到 毗努伊勒 ，对那里的人也提出同样的请求； 毗努伊勒 人给他的答覆跟 疏割 人的答覆一样。
JUDG|8|9|他也对 毗努伊勒 人说：“我平平安安回来的时候，必拆毁这城楼。”
JUDG|8|10|那时 西巴 和 撒慕拿 ，以及跟随他们的军队都在 加各 ，约有一万五千人，是东边的人全军所剩下的，因为拿刀战死的约有十二万人。
JUDG|8|11|基甸 从 挪巴 和 约比哈 的东边，从住帐棚人 的路上去，趁 米甸 的军兵以为安全的时候攻击他们。
JUDG|8|12|西巴 和 撒慕拿 逃跑； 基甸 追赶他们，捉住 米甸 的两个王 西巴 和 撒慕拿 ，使他们全军溃散。
JUDG|8|13|约阿施 的儿子 基甸 从战场，沿着 希列斯 斜坡回来，
JUDG|8|14|捉住 疏割 人的一个少年，查问他。他就为 基甸 写下 疏割 的领袖和长老的名字，共七十七人。
JUDG|8|15|基甸 到了 疏割 人那里，说：“你们从前讥笑我说：‘ 西巴 和 撒慕拿 的手掌现在已经在你手里，因此我们该将饼送给跟随你的疲乏的人吗？’看哪， 西巴 和 撒慕拿 在这里。”
JUDG|8|16|于是他拿住城内的长老，用旷野的荆棘和枳条责打 疏割 人。
JUDG|8|17|他又拆了 毗努伊勒 的城楼，杀了城里的人。
JUDG|8|18|基甸 对 西巴 和 撒慕拿 说：“你们在 他泊山 所杀的人是什么样子的？”他们说：“他们很像你，个个都有王子的样子。”
JUDG|8|19|基甸 说：“他们都是我的兄弟，我母亲的儿子。我指着永生的耶和华起誓，你们若存留他们的性命，我就不杀你们了。”
JUDG|8|20|他对他的长子 益帖 说：“你起来杀他们！”但是这少年害怕，不敢拔刀，因为他还是个少年。
JUDG|8|21|西巴 和 撒慕拿 说：“你自己起来杀我们吧！因为人如何，力量也如何。” 基甸 就起来，杀了 西巴 和 撒慕拿 ，取了他们骆驼颈项上的月牙圈。
JUDG|8|22|以色列 人对 基甸 说：“你既然救我们脱离 米甸 的手，愿你治理我们，你的儿子孙子也治理我们。”
JUDG|8|23|基甸 对他们说：“我不治理你们，我的儿子也不治理你们，耶和华会治理你们。”
JUDG|8|24|基甸 又对他们说：“我有一件事求你们，请你们各人把所夺的耳环给我。”因敌人都戴金耳环，他们是 以实玛利 人。
JUDG|8|25|以色列 人说：“我们情愿送给你！”他们就铺开一件外衣，各人将所夺的耳环丢在上面。
JUDG|8|26|基甸 所要求的金耳环，重一千七百舍客勒金子。此外还有 米甸 王所戴的月牙圈、耳环，和所穿的紫色衣服，以及骆驼颈项上的链子。
JUDG|8|27|基甸 以此造了一个以弗得，设立在他的本城 俄弗拉 。全 以色列 就在那里拜这以弗得行淫，这就成了 基甸 和他全家的圈套。
JUDG|8|28|这样， 米甸 就被 以色列 人制伏了，再也不能抬头。 基甸 还在的日子，这地太平四十年。
JUDG|8|29|约阿施 的儿子 耶路巴力 回去，住在自己家里。
JUDG|8|30|基甸 有七十个亲生的儿子，因为他有许多妻子。
JUDG|8|31|他在 示剑 的妾也为他生了一个儿子， 基甸 给他起名叫 亚比米勒 。
JUDG|8|32|约阿施 的儿子 基甸 年纪老迈而死，葬在 亚比以谢 族的 俄弗拉 ，他父亲 约阿施 的坟墓里。
JUDG|8|33|基甸 死后， 以色列 人又去随从诸 巴力 而行淫，以 巴力．比利土 为他们的神明。
JUDG|8|34|以色列 人不记得耶和华－他们的上帝，就是那位拯救他们脱离四围仇敌之手的，
JUDG|8|35|也不照着 耶路巴力 ，就是 基甸 向 以色列 所施的恩惠善待他的家。
JUDG|9|1|耶路巴力 的儿子 亚比米勒 到 示剑 他的母舅那里，对他们和他外祖父全家的人说：
JUDG|9|2|“请你们问 示剑 所有的居民：‘是 耶路巴力 的众儿子七十人都治理你们好，还是一人治理你们好呢？’你们要记得，我是你们的骨肉。”
JUDG|9|3|他的母舅们为他把这一切话说给 示剑 所有的居民听，他们的心就倾向 亚比米勒 ，因为他们说：“他是我们的弟兄。”
JUDG|9|4|他们从 巴力．比利土 的庙中取了七十银子给 亚比米勒 ， 亚比米勒 用这些钱雇了一些无赖匪徒跟随他。
JUDG|9|5|他来到 俄弗拉 他父亲的家，在一块磐石上把他的兄弟，就是 耶路巴力 的七十个儿子都杀了，只剩下 耶路巴力 的小儿子 约坦 ，因为他躲了起来。
JUDG|9|6|示剑 所有的居民和全 伯．米罗 都聚集在一起，到 示剑 橡树旁的柱子那里，立 亚比米勒 为王。
JUDG|9|7|有人将这事告诉 约坦 ，他就去站在 基利心山 顶上，高声喊叫，对他们说：“ 示剑 的居民哪，你们要听我，上帝也就会听你们。
JUDG|9|8|有一次，树木要膏一王治理他们，就去对橄榄树说：‘请你来作王治理我们！’
JUDG|9|9|橄榄树对它们说：‘我岂可停止生产使神明和人得尊荣的油，而行走飘摇在众树之上呢？’
JUDG|9|10|树木对无花果树说：‘请你来作王治理我们！’
JUDG|9|11|无花果树对它们说：‘我岂可停止结甜美的果子，而行走飘摇在众树之上呢？’
JUDG|9|12|树木对葡萄树说：‘请你来作王治理我们！’
JUDG|9|13|葡萄树对它们说：‘我岂可停止出产使神明和人欢乐的新酒，而行走飘摇在众树之上呢。’
JUDG|9|14|众树对荆棘说：‘请你来作王治理我们！’
JUDG|9|15|荆棘对众树说：‘你们若真的要膏我作王治理你们，就要来到我的荫下寻求庇护；不然，愿火从荆棘里出来，吞灭 黎巴嫩 的香柏树。’
JUDG|9|16|“现在你们若以诚实正直立 亚比米勒 为王，若善待 耶路巴力 和他的家，若照他手所做的回报他─
JUDG|9|17|从前我父为你们争战，冒生命的危险救你们脱离 米甸 的手，
JUDG|9|18|但是你们如今起来攻击我的父家，在一块磐石上把他的七十个儿子全杀了，又立他使女所生的儿子 亚比米勒 为 示剑 居民的王，因为他是你们的弟兄─
JUDG|9|19|你们如今若以诚实正直对待 耶路巴力 和他的家，就可以因 亚比米勒 欢乐，他也可以因你们欢乐；
JUDG|9|20|不然，愿火从 亚比米勒 发出，吞灭 示剑 居民和 伯．米罗 ，又愿火从 示剑 居民和 伯．米罗 发出，吞灭 亚比米勒 。”
JUDG|9|21|约坦 因躲避他的兄弟 亚比米勒 就逃跑，去到 比珥 ，住在那里。
JUDG|9|22|亚比米勒 治理 以色列 三年。
JUDG|9|23|上帝派邪灵到 亚比米勒 和 示剑 居民中间， 示剑 居民就以诡诈待 亚比米勒 。
JUDG|9|24|这是要使 耶路巴力 七十个儿子受害所流的血，归于他们的兄弟 亚比米勒 ，因他杀害他们，也归于那些出手帮助他杀害兄弟的 示剑 居民。
JUDG|9|25|示剑 居民在山顶上设下埋伏，等候 亚比米勒 。凡沿着那条路，从他们那里经过的人，他们就抢劫。有人把这事告诉 亚比米勒 。
JUDG|9|26|以别 的儿子 迦勒 和他的弟兄经过，来到 示剑 ， 示剑 居民都信任他。
JUDG|9|27|他们出到田间，摘下葡萄，踹酒，作乐。他们进入他们神明的庙中吃喝，诅咒 亚比米勒 。
JUDG|9|28|以别 的儿子 迦勒 说：“ 亚比米勒 是谁，我们 示剑 人是谁，叫我们服事他呢？他不是 耶路巴力 的儿子吗？他的助手不是 西布勒 吗？你们应当服事 示剑 的父亲 哈抹 的后裔！我们为何要服事 亚比米勒 呢？
JUDG|9|29|惟愿这民归到我的手下，我就除掉 亚比米勒 。”他就对 亚比米勒 说：“增加你的军兵，出来吧！”
JUDG|9|30|西布勒 市长听见 以别 的儿子 迦勒 的话，就怒气大发。
JUDG|9|31|他悄悄地派一些使者到 亚比米勒 那里，说：“看哪， 以别 的儿子 迦勒 和他的弟兄到了 示剑 。看哪，他们煽动那城攻击你。
JUDG|9|32|现在，你和跟随你的百姓要夜间起来，在田间埋伏。
JUDG|9|33|早晨太阳一出，你就趁早攻城。看哪， 迦勒 和跟随他的百姓出来攻击你的时候，你就全力对付他们。”
JUDG|9|34|于是， 亚比米勒 和跟随他的众百姓夜间起来，兵分四队，埋伏攻击 示剑 。
JUDG|9|35|以别 的儿子 迦勒 出去，站在城门口。 亚比米勒 和跟随他的百姓从埋伏之处起来。
JUDG|9|36|迦勒 看见百姓，就对 西布勒 说：“看哪，有百姓从山顶上下来。” 西布勒 对他说：“你把山的影子看作是人了。”
JUDG|9|37|迦勒 又继续讲，他说：“看哪，有百姓从地的高处下来，又有一队从 米恶尼尼 橡树 的路前来。”
JUDG|9|38|西布勒 对他说：“你所夸口的在哪里呢？你曾说：‘ 亚比米勒 是谁，叫我们服事他呢？’这不是你所藐视的百姓吗？你现在出去，与他们交战吧！”
JUDG|9|39|于是 迦勒 率领 示剑 居民出去，与 亚比米勒 交战。
JUDG|9|40|亚比米勒 追赶 迦勒 ， 迦勒 在他面前逃跑。有许多人被刺伤仆倒，直到城门口。
JUDG|9|41|亚比米勒 住在 亚鲁玛 。 西布勒 赶出 迦勒 和他的弟兄，不准他们住在 示剑 。
JUDG|9|42|次日，百姓出到田间，有人告诉 亚比米勒 ，
JUDG|9|43|他就带领百姓，把他们分成三队，埋伏在田间窥探。看哪， 示剑 居民从城里出来，他就起来击杀他们。
JUDG|9|44|亚比米勒 和跟随他的一队向前冲，站在城门口；另外两队直冲向田间，击杀了众人。
JUDG|9|45|亚比米勒 攻城一整天，将城夺取，杀了其中的百姓，把城拆毁，撒上了盐。
JUDG|9|46|示剑 城楼里所有的居民听见了，就进入 伊勒．比利土 庙的地窖里。
JUDG|9|47|有人告诉 亚比米勒 ， 示剑 城楼里所有的居民都聚在一起。
JUDG|9|48|亚比米勒 和所有跟随他的百姓都上 撒们山 去。 亚比米勒 手拿斧子，砍下一根树枝，举起来，扛在肩上，对跟随他的百姓说：“你们看我做什么，就赶快照样做。”
JUDG|9|49|众百姓也都各砍一根树枝，跟 亚比米勒 走，把树枝堆在地窖上，放火烧地窖。这样， 示剑 城楼里所有的人都死了，男女约有一千。
JUDG|9|50|亚比米勒 到 提备斯 ，对着 提备斯 安营，攻取了那城。
JUDG|9|51|城中有一座坚固的楼；城里所有的居民，无论男女，都逃到那里，关上门，上了楼顶。
JUDG|9|52|亚比米勒 到了楼前，攻打它。他挨近楼门，要放火焚烧。
JUDG|9|53|有一个妇人把一块上磨石抛在 亚比米勒 的头上，打破了他的头盖骨。
JUDG|9|54|他就急忙叫拿他兵器的青年来，对他说：“拔出你的刀来，杀了我吧！免得有人提到我说：‘他被一个妇人杀了。’”于是那青年把他刺透，他就死了。
JUDG|9|55|以色列 人见 亚比米勒 死了，就各回自己的地方去了。
JUDG|9|56|这样，上帝报应了 亚比米勒 向他父亲所做的恶事，就是杀了自己七十个兄弟。
JUDG|9|57|示剑 人的一切恶事，上帝也都报应在他们头上； 耶路巴力 的儿子 约坦 的诅咒都临到他们身上了。
JUDG|10|1|亚比米勒 以后， 陀拉 兴起，拯救 以色列 ，他是 朵多 的孙子， 普瓦 的儿子， 以萨迦 人，住在 以法莲 山区的 沙密 。
JUDG|10|2|陀拉 作 以色列 的士师二十三年。他死了，葬在 沙密 。
JUDG|10|3|陀拉 以后有 基列 人 睚珥 兴起，作 以色列 的士师二十二年。
JUDG|10|4|他有三十个儿子，骑着三十匹驴驹。他们有三十座城，叫作 哈倭特．睚珥 ，直到如今，都在 基列 地。
JUDG|10|5|睚珥 死了，葬在 加们 。
JUDG|10|6|以色列 人又行耶和华眼中看为恶的事，去事奉诸 巴力 和 亚斯她录 ，以及 亚兰 的神明、 西顿 的神明、 摩押 的神明、 亚扪 人的神明、 非利士 人的神明。他们离弃耶和华，不事奉他。
JUDG|10|7|耶和华的怒气向 以色列 发作，把他们交给 非利士 人和 亚扪 人的手中。
JUDG|10|8|从那年起，他们欺压迫害 以色列 人，在 约旦河 东， 亚摩利 人境内， 基列 一带所有的 以色列 人，长达十八年。
JUDG|10|9|亚扪 人渡过 约旦河 去攻打 犹大 和 便雅悯 ，以及 以法莲 家族。 以色列 的处境非常困苦。
JUDG|10|10|以色列 人哀求耶和华说：“我们得罪了你，因为我们离弃了我们的上帝，去事奉诸 巴力 。”
JUDG|10|11|耶和华对 以色列 人说：“我岂没有救你们脱离 埃及 人、 亚摩利 人、 亚扪 人和 非利士 人吗？
JUDG|10|12|西顿 人、 亚玛力 人和 马云 人 欺压你们，你们哀求我，我也拯救你们脱离他们的手。
JUDG|10|13|你们竟离弃我去事奉别神！所以我不再救你们了。
JUDG|10|14|你们去哀求你们所选择的神明；你们遭遇急难的时候，让它们救你们吧！”
JUDG|10|15|以色列 人对耶和华说：“我们犯罪了，照你看为好的待我们，只求你今日拯救我们吧！”
JUDG|10|16|以色列 人就除掉他们中间的外邦神明，事奉耶和华。耶和华因 以色列 所受的苦难而心里焦急。
JUDG|10|17|亚扪 人被召来，在 基列 安营； 以色列 人也聚集，在 米斯巴 安营。
JUDG|10|18|基列 百姓中的领袖彼此说：“谁领先出去攻打 亚扪 人，谁就作 基列 所有居民的领袖。”
JUDG|11|1|基列 人 耶弗他 是个大能的勇士，是妓女的儿子。 基列 生了 耶弗他 。
JUDG|11|2|基列 的妻子也给他生了几个儿子。他妻子生的儿子长大后，就把 耶弗他 赶出去，说：“你不可在我们父家继承产业，因为你是别的女人生的儿子。”
JUDG|11|3|耶弗他 就逃离他的兄弟，住在 陀伯 地。有些无赖的人聚集在他那里，与他一同出入。
JUDG|11|4|过了些日子， 亚扪 人攻打 以色列 。
JUDG|11|5|亚扪 人攻打 以色列 的时候， 基列 的长老去请 耶弗他 从 陀伯 地回来。
JUDG|11|6|他们对 耶弗他 说：“请你来作我们的指挥官，好让我们跟 亚扪 人打仗。”
JUDG|11|7|耶弗他 对 基列 的长老说：“你们不是恨我，把我赶出父家吗？现在你们遭遇急难，为何到我这里来呢？”
JUDG|11|8|基列 的长老对 耶弗他 说：“现在我们回到你这里，是要请你同我们去跟 亚扪 人打仗，作 基列 所有居民的领袖。”
JUDG|11|9|耶弗他 对 基列 的长老说：“若你们请我回去跟 亚扪 人打仗，耶和华把他们交给我，我就作你们的领袖。”
JUDG|11|10|基列 的长老对 耶弗他 说：“有耶和华在你我之间作证，我们必定照你的话做。”
JUDG|11|11|于是 耶弗他 与 基列 的长老同去，百姓就立 耶弗他 作他们的领袖和指挥官。 耶弗他 在 米斯巴 将他一切的事陈述在耶和华面前。
JUDG|11|12|耶弗他 派使者到 亚扪 人的王那里，说：“你与我有什么相干，竟来到我这里攻打我的地呢？”
JUDG|11|13|亚扪 人的王对 耶弗他 的使者说：“因为 以色列 从 埃及 上来的时候占据我的地，从 亚嫩河 到 雅博河 ，直到 约旦河 。现在你要和平归还这些地方！”
JUDG|11|14|耶弗他 又派使者到 亚扪 人的王那里，
JUDG|11|15|对他说：“ 耶弗他 如此说： 以色列 并没有占据 摩押 地和 亚扪 人的地。
JUDG|11|16|以色列 人从 埃及 上来，是经过旷野到 红海 ，来到 加低斯 。
JUDG|11|17|那时， 以色列 派使者去 以东 王那里，说：‘求你让我穿越你的地。’ 以东 王却不听。 以色列 又照样派使者去 摩押 王那里，他也不肯。于是 以色列 人就住在 加低斯 。
JUDG|11|18|他们又经过旷野，绕过 以东 地和 摩押 地，到 摩押 地的东边 ，在 亚嫩河 边安营，并没有进入 摩押 的境内，因为 亚嫩河 是 摩押 的边界。
JUDG|11|19|以色列 派使者去 亚摩利 王，就是 希实本 王 西宏 那里； 以色列 对他说：‘求你让我们穿越你的地，到我自己的地方去。’
JUDG|11|20|西宏 却不信任 以色列 ，不让他们穿越他的疆界。他召集了他的众百姓在 雅杂 安营，与 以色列 争战。
JUDG|11|21|耶和华－ 以色列 的上帝将 西宏 和他的众百姓都交在 以色列 手中， 以色列 人就击杀他们，占领了那地居民 亚摩利 人的全地。
JUDG|11|22|他们占领了 亚摩利 人所有的疆土，从 亚嫩河 到 雅博河 ，从旷野直到 约旦河 。
JUDG|11|23|耶和华－ 以色列 的上帝如今从他百姓 以色列 面前赶出 亚摩利 人，你竟要占领它吗？
JUDG|11|24|你不是已经得了你的神明 基抹 赐给你的地为业吗？耶和华－我们的上帝在我们面前所赶出的，我们也要得它为业。
JUDG|11|25|现在你比 西拨 的儿子 摩押 王 巴勒 还强吗？他真的曾与 以色列 争执，或是真的与他们争战了吗？
JUDG|11|26|以色列 人住 希实本 和所属的乡镇， 亚罗珥 和所属的乡镇，以及沿着 亚嫩河 的一切城镇，已经有三百年了。在这期间，你们为什么不取回呢？
JUDG|11|27|我并没有得罪你，你却要攻打我，加害于我。愿审判人的耶和华今日在 以色列 人和 亚扪 人之间判断是非。”
JUDG|11|28|但 亚扪 人的王不听 耶弗他 传达给他的话。
JUDG|11|29|耶和华的灵降在 耶弗他 身上，他就经过 基列 和 玛拿西 ，经过 基列 的 米斯巴 ，又从 基列 的 米斯巴 过到 亚扪 人那里。
JUDG|11|30|耶弗他 向耶和华许愿，说：“你若真的将 亚扪 人交在我手中，
JUDG|11|31|我从 亚扪 人那里平平安安回来的时候，无论谁先从我家门出来迎接我，就要归给耶和华，我必将他献上作为燔祭。”
JUDG|11|32|于是 耶弗他 往 亚扪 人那里去，与他们争战。耶和华将他们交在他手中，
JUDG|11|33|他就彻底击败他们，从 亚罗珥 到 米匿 ，直到 亚备勒．基拉明 ，攻取了二十座城。这样， 亚扪 人就在 以色列 人面前被制伏了。
JUDG|11|34|耶弗他 回 米斯巴 去，到了自己的家，看哪，他女儿拿着手鼓跳舞出来迎接他。她是 耶弗他 的独生女，除她以外，没有别的儿女。
JUDG|11|35|耶弗他一看见她，就撕裂衣服，说：“哀哉！我的女儿啊，你使我非常悲痛，叫我十分为难了。因为我已经向耶和华开了口，不能收回。”
JUDG|11|36|他女儿对他说：“我的父亲啊，你既向耶和华开了口，就当照你口中所说的向我行，因为耶和华已经在你的仇敌 亚扪 人身上为你报了仇。”
JUDG|11|37|她又对父亲说：“我只求你这一件事，给我两个月，让我和同伴下到山里，好为我的童贞哀哭。”
JUDG|11|38|耶弗他 说：“你去吧！”他就让她离开两个月。她和同伴去了，在山里为她的童贞哀哭。
JUDG|11|39|过了两个月，她回到父亲那里，父亲就照所许的愿向她行了。她从来没有亲近男人。于是 以色列 中有个风俗，
JUDG|11|40|每年按着日期 以色列 的女子要去为 基列 人 耶弗他 的女儿哀哭四天。
JUDG|12|1|以法莲 人被召来，渡河来到 撒分 。他们对 耶弗他 说：“你去与 亚扪 人争战，为什么没有召我们同去呢？我们必用火将你和你的家烧了。”
JUDG|12|2|耶弗他 对他们说：“我和我的百姓与 亚扪 人有极大的冲突；我曾召你们来，你们却没有来救我脱离他们的手。
JUDG|12|3|我见你们不来救我，就拚了命前去攻打 亚扪 人，耶和华就将他们交在我手中。你们今日为什么上我这里来攻打我呢？”
JUDG|12|4|于是 耶弗他 召集 基列 所有的人，要与 以法莲 人争战。 基列 人击杀 以法莲 人，因 以法莲 人曾说：“你们 基列 人在 以法莲 和 玛拿西 中，不过是 以法莲 逃亡的人而已。”
JUDG|12|5|基列 人把守 约旦河 的渡口，不许 以法莲 人过去。逃跑的 以法莲 人若说：“让我过河。” 基列 人就问他说：“你是不是 以法莲 人？”他若说：“不是”，
JUDG|12|6|基列 人就对他说：“你说‘示播列’。” 以法莲 人因为发音不准，就会说成“西播列”。 基列 人就捉住他，在 约旦河 的渡口把他杀了。那时， 以法莲 人被杀的有四万二千人。
JUDG|12|7|耶弗他 作 以色列 的士师六年。 基列 人 耶弗他 死了，葬在 基列 的城里 。
JUDG|12|8|耶弗他 以后，有 伯利恒 人 以比赞 作 以色列 的士师。
JUDG|12|9|他有三十个儿子。他把三十个女儿都嫁出去了，也为他的儿子从外面娶了三十个媳妇。他作 以色列 的士师七年。
JUDG|12|10|以比赞 死了，葬在 伯利恒 。
JUDG|12|11|以比赞 以后，有 西布伦 人 以伦 作 以色列 的士师，他作 以色列 的士师十年。
JUDG|12|12|西布伦 人 以伦 死了，葬在 西布伦 地的 亚雅仑 。
JUDG|12|13|以伦 以后，有 比拉顿 人 希列 的儿子 押顿 作 以色列 的士师。
JUDG|12|14|他有四十个儿子，三十个孙子，骑着七十匹驴驹。 押顿 作 以色列 的士师八年。
JUDG|12|15|比拉顿 人 希列 的儿子 押顿 死了，葬在 以法莲 地的 比拉顿 ，就在 亚玛力 人的山区。
JUDG|13|1|以色列 人又行耶和华眼中看为恶的事，耶和华将他们交在 非利士 人手中四十年。
JUDG|13|2|那时，有一个 但 支派的 琐拉 人，名叫 玛挪亚 。他的妻子不怀孕，不生育。
JUDG|13|3|耶和华的使者向那妇人显现，对她说：“看哪，以前你不怀孕，不生育，如今你必怀孕生一个儿子。
JUDG|13|4|现在你要谨慎，清酒烈酒都不可喝，任何不洁之物都不可吃，
JUDG|13|5|看哪，你必怀孕，生一个儿子。不可用剃刀剃他的头，因为这孩子一出母胎就归给上帝作拿细耳人。他必开始拯救 以色列 脱离 非利士 人的手。”
JUDG|13|6|那妇人来对丈夫说：“有一个神人到我这里来，他的容貌如上帝使者的容貌，非常可畏。我没有问他从哪里来，他也没有把他的名字告诉我。
JUDG|13|7|他对我说：‘看哪，你要怀孕，生一个儿子 。现在，清酒烈酒都不可喝，任何不洁之物都不可吃，因为这孩子从出母胎一直到死的那一天，要归给上帝作拿细耳人。’”
JUDG|13|8|玛挪亚 祈求耶和华说：“主啊，求你再差遣那神人到我们这里来，指示我们对这将要生的孩子该怎样作。”
JUDG|13|9|上帝垂听了 玛挪亚 的声音。那妇人坐在田间的时候，上帝的使者又到她那里，但是她的丈夫 玛挪亚 没有同她在一起。
JUDG|13|10|妇人急忙跑去告诉丈夫，对他说：“看哪，那日到我这里来的人又向我显现了。”
JUDG|13|11|玛挪亚 起来，跟随他的妻子来到那人那里，对他说：“你就是跟这妇人说话的那个人吗？”他说：“是我。”
JUDG|13|12|玛挪亚 说：“现在，愿你的话应验！这孩子该如何管教呢？他当做什么呢？”
JUDG|13|13|耶和华的使者对 玛挪亚 说：“我告诉这妇人的一切事，她都要遵守。
JUDG|13|14|葡萄树所结的不可吃，清酒烈酒都不可喝，任何不洁之物也不可吃。凡我所吩咐的，她都当遵守。”
JUDG|13|15|玛挪亚 对耶和华的使者说：“请容许我们留你下来，好为你预备一只小山羊。”
JUDG|13|16|耶和华的使者对 玛挪亚 说：“你虽然留我，我却不吃你的食物。你若预备燔祭，就当献给耶和华。”因 玛挪亚 不知道他是耶和华的使者。
JUDG|13|17|玛挪亚 对耶和华的使者说：“请问大名？好让我们在你的话应验的时候尊敬你。”
JUDG|13|18|耶和华的使者对他说：“你何必问我的名字呢？我的名字是奇妙的。”
JUDG|13|19|玛挪亚 取一只小山羊和素祭，在磐石上献给耶和华。他行奇妙的事， 玛挪亚 和他的妻子观看，
JUDG|13|20|火焰从坛上往上升，耶和华的使者也在坛上的火焰中升上去了。 玛挪亚 和他的妻子看见，就脸伏于地。
JUDG|13|21|耶和华的使者不再向 玛挪亚 和他的妻子显现了。那时， 玛挪亚 才知道他是耶和华的使者。
JUDG|13|22|玛挪亚 对他的妻子说：“我们一定会死，因为我们看见了上帝。”
JUDG|13|23|他的妻子却对他说：“耶和华若有意要我们死，就不会从我们手中接受燔祭和素祭，不会将这一切事指示我们，这时也不会让我们听到这话。”
JUDG|13|24|后来妇人生了一个儿子，给他起名叫 参孙 。孩子渐渐长大，耶和华赐福给他。
JUDG|13|25|在 琐拉 和 以实陶 之间的 玛哈尼．但 ，耶和华的灵开始感动 参孙 。
JUDG|14|1|参孙 下到 亭拿 ，在 亭拿 看见一个女子，是 非利士 人的女儿。
JUDG|14|2|他上来告诉他父母说：“我在 亭拿 看见一个女子，是 非利士 人的女儿，现在请你们给我娶她为妻。”
JUDG|14|3|他父母对他说：“在你弟兄的女儿中，或在本族所有的人中，难道没有女子吗？你何必在未受割礼的 非利士 人中去娶妻呢？” 参孙 对他父亲说：“请你给我娶那女子，因为我喜欢她。”
JUDG|14|4|他的父母并不知道这事是出于耶和华，因为他在找机会攻击 非利士 人。那时， 非利士 人辖制 以色列 人。
JUDG|14|5|参孙 跟他父母下 亭拿 去，他们到了 亭拿 的葡萄园。看哪，有一只少壮狮子对着他吼叫。
JUDG|14|6|耶和华的灵大大感动 参孙 ，他就手无寸铁撕裂狮子，如撕裂小山羊一样。他做这事，并没有告诉他的父母亲。
JUDG|14|7|参孙 下去跟那女子说话，看着就喜欢她。
JUDG|14|8|过了些日子，他回来要娶那女子，绕道去看狮子的残骸，看哪，有一群蜜蜂在狮子的尸体内，也有蜜在里面。
JUDG|14|9|他就取了蜜，放在手掌上，边走边吃。他到了父母那里，给他们蜜，他们也吃了。但他没有告诉他们，这蜜是从狮子的尸体内取来的。
JUDG|14|10|他父亲下到女子那里去。 参孙 在那里摆设宴席， 因为这是当时年轻人的习俗。
JUDG|14|11|他们看见 参孙 ，就请了三十个人陪伴他。
JUDG|14|12|参孙 对他们说：“我给你们出个谜语，你们若能在七日宴席之内，猜出谜底告诉我，我就给你们三十件细麻内衣和三十套更换的衣服。
JUDG|14|13|但你们若不能告诉我，你们就给我三十件细麻内衣和三十套更换的衣服。”他们对他说：“请把谜语说给我们听。”
JUDG|14|14|参孙 对他们说： “吃的从吃者出来； 甜的从强者出来”。 三日之久，他们都猜不出谜语来。
JUDG|14|15|第七日 ，他们对 参孙 的妻子说：“你哄骗你的丈夫，为我们探出谜底来，否则我们就用火烧你和你的父家。你们请我们来，是不是要夺走我们所有的呢？”
JUDG|14|16|参孙 的妻子在丈夫面前哭哭啼啼说：“你只是恨我，并不爱我。你给我本族的人出谜语，却不把谜底告诉我。” 参孙 对她说：“看哪，连我的父母我都没有说，我怎么可以告诉你呢？”
JUDG|14|17|在七日宴席中，她一直在丈夫面前哭哭啼啼。第七日， 参孙 因妻子的催逼就把谜底告诉了她。她把谜底告诉了她本族的人。
JUDG|14|18|第七日日落以前，那城里的人对 参孙 说： “有什么比蜜还甜呢？ 有什么比狮子更强呢？” 参孙 对他们说： “你们若不用我的母牛犊耕地， 就无法猜出我的谜底来。”
JUDG|14|19|耶和华的灵大大感动 参孙 ，他就下到 亚实基伦 ，击杀了三十个人，夺了他们身上的衣服，把衣服给了猜出谜语的人。 参孙 怒气大发，就上他父亲的家去了。
JUDG|14|20|参孙 的妻子就归了 参孙 的一个同伴，就是作过他伴郎的。
JUDG|15|1|过了些日子，在割麦子的时候， 参孙 带着一只小山羊去探望他的妻子，说：“我要进内室到我妻子那里。”他岳父不许他进去。
JUDG|15|2|他岳父说：“我以为你极其恨她，因此我把她给了你的同伴。她妹妹不是比她更美丽吗？你可以娶来代替她！”
JUDG|15|3|参孙 对他们说：“这一次我若加害 非利士 人，就不算是我的错了。”
JUDG|15|4|于是 参孙 去捉了三百只狐狸，把它们的尾巴一对一对地绑住，再将火把绑在两条尾巴中间。
JUDG|15|5|他点着火把，把狐狸放进 非利士 人直立的庄稼，把堆积的禾捆和直立的庄稼，葡萄园、橄榄园全都烧了。
JUDG|15|6|非利士 人说：“这事是谁做的呢？”有人说：“是 亭拿 人的女婿 参孙 做的，因为他岳父把他的妻子给了他的同伴。”于是 非利士 人上去，用火烧了女子和她的父亲。
JUDG|15|7|参孙 对他们说：“你们既然这么做，我必向你们报仇才肯罢休。”
JUDG|15|8|参孙 狠狠击杀他们，把他们连腿带腰都砍了。过后，他就下去，住在 以坦岩 的石洞里。
JUDG|15|9|非利士 人上去，安营在 犹大 ，侵犯 利希 。
JUDG|15|10|犹大 人说：“你们为何上来攻击我们呢？”他们说：“我们上来是要捆绑 参孙 ，照他向我们所做的对待他。”
JUDG|15|11|于是，三千 犹大 人下到 以坦岩 的石洞里，对 参孙 说：“ 非利士 人辖制我们，你不知道吗？你向我们做的是什么事呢？”他说：“他们向我怎样做，我也要向他们怎样做。”
JUDG|15|12|犹大 人对他说：“我们下来是要捆绑你，把你交在 非利士 人手中。” 参孙 说：“你们要向我起誓，你们自己不杀害我。”
JUDG|15|13|他们说：“我们绝不杀你，只把你捆绑，交在 非利士 人手中。”于是他们用两条新绳绑住 参孙 ，把他从 以坦岩 带上去。
JUDG|15|14|参孙 到了 利希 ， 非利士 人对着他喊叫。耶和华的灵大大感动 参孙 ，他手臂上的绳子就像着火的麻一样，绑他的绳子从他手上脱落下来。
JUDG|15|15|他找到一块未干的驴腮骨，就伸手拾起来，用它杀了一千人。
JUDG|15|16|参孙 说： “用驴腮骨， 一堆又一堆 ； 用驴腮骨， 我杀了一千人。”
JUDG|15|17|说完这话，就把那腮骨从手里抛出去。因此，那地叫作 拉末．利希 。
JUDG|15|18|参孙 非常口渴，就求告耶和华说：“你既藉仆人的手施行这么大的拯救，现在我要渴死，落在未受割礼的人手中吗？”
JUDG|15|19|上帝就使 利希 的洼地裂开，从中涌出水来。 参孙 喝了，精神恢复。因此那泉名叫 隐．哈歌利 ，直到今日它仍在 利希 。
JUDG|15|20|在 非利士 人辖制的时候， 参孙 作 以色列 的士师二十年。
JUDG|16|1|参孙 到了 迦萨 ，在那里看见一个妓女，就与她亲近。
JUDG|16|2|有人告诉 迦萨 人说：“ 参孙 到这里来了！”他们就包围起来，整夜在城门埋伏等着他。他们整夜静悄悄地，说：“等到天一亮我们就杀他。”
JUDG|16|3|参孙 睡到半夜，在半夜起来，抓住城门的门扇和两个门框，把它们和门闩一起拆下来，扛在肩上，抬到 希伯仑 前面的山顶上。
JUDG|16|4|这事以后， 参孙 在 梭烈谷 爱上了一个女子，名叫 大利拉 。
JUDG|16|5|非利士 人的领袖上去，到那女子那里，对她说：“请你哄骗 参孙 ，探出他为何有这么大的力气，以及我们要用什么方法才能胜他，将他捆绑制伏。我们就每人给你一千一百块银子。”
JUDG|16|6|大利拉 对 参孙 说：“请你告诉我，你为何有这么大的力气，要用什么方法才能捆绑制伏你。”
JUDG|16|7|参孙 对她说：“若用七条未干的新绳子捆绑我，我就像平常人一样软弱。”
JUDG|16|8|于是 非利士 人的领袖拿了七条未干的新绳子来，交给她，她就用绳子捆绑 参孙 。
JUDG|16|9|当时，埋伏的人正在她的内室等着。她对 参孙 说：“ 参孙 ， 非利士 人来捉你了！” 参孙 就挣断绳子，绳子如遇到火的麻线断裂一样。这样，人还是不知道他的力量从哪里来。
JUDG|16|10|大利拉 对 参孙 说：“看哪，你欺骗我，对我说谎。现在请你告诉我，要用什么方法才能捆绑你。”
JUDG|16|11|参孙 对她说：“若用未曾用过的新绳子捆绑我，我就像平常人一样软弱。”
JUDG|16|12|大利拉 就用新绳子捆绑他，对他说：“ 参孙 ， 非利士 人来捉你了！”当时，埋伏的人在内室等着。 参孙 挣断手臂上的绳子，如挣断一条线一样。
JUDG|16|13|大利拉 对 参孙 说：“你到现在还是欺骗我，对我说谎。请你告诉我，要用什么方法才能捆绑你。” 参孙 对她说：“只要用织布的线将我头上的七条发绺编织起来就可以了”。
JUDG|16|14|于是 大利拉 用梭子将他的发绺钉住，对他说：“ 参孙 ， 非利士 人来捉你了！” 参孙 从睡中醒来，将织布机上的梭子和织布的线一齐都拔出来了。
JUDG|16|15|大利拉 对 参孙 说：“你既不与我同心，怎么能说‘我爱你’呢？你这三次欺骗我，不告诉我，你为什么有这么大的力气。”
JUDG|16|16|大利拉 天天用话催逼他，纠缠他，他就心里烦得要死，
JUDG|16|17|终于把心中的一切都告诉她。 参孙 对她说：“从来没有人用剃刀剃我的头，因为我一出母胎就归给上帝作拿细耳人。若有人剃了我的头发，我的力气就会离开我，我就像平常人一样软弱。”
JUDG|16|18|大利拉 见他说出了心中的一切，就派人去召 非利士 人的领袖，说：“请再上来一次，因为他已经说出了心中的一切。”于是 非利士 人的领袖手里拿着银子，上到她那里。
JUDG|16|19|大利拉 哄 参孙 睡在她的膝上，叫一个人来剃掉 参孙 头上的七条发绺。于是 大利拉 开始制伏 参孙 ，他的力气就离开他了。
JUDG|16|20|大利拉 说：“ 参孙 ， 非利士 人来捉你了！” 参孙 从睡中醒来，说：“我要像前几次一样脱身而去。”他却不知道耶和华已经离开他了。
JUDG|16|21|非利士 人逮住他，挖了他的眼睛，带他下到 迦萨 ，用铜链锁住他，叫他在监狱里推磨。
JUDG|16|22|然而他的头发被剃以后，又开始长起来了。
JUDG|16|23|非利士 人的领袖聚集，要向他们的神明 大衮 献大祭，并且庆祝，说：“我们的神明把我们的仇敌 参孙 交在我们手中了。”
JUDG|16|24|众人看见 参孙 ，就赞美他们的神明说：“我们的神明把那毁坏我们的地、杀害我们许多人的仇敌交在我们手中了。”
JUDG|16|25|他们心里高兴的时候，就说：“叫 参孙 来，逗我们欢乐。”于是他们把 参孙 从监狱里提出来，在他们面前戏耍。他们叫他站在两根柱子中间。
JUDG|16|26|参孙 对牵他手的童仆说：“让我摸摸支撑这庙宇的柱子，我要靠一靠。”
JUDG|16|27|那时庙宇内充满男女， 非利士 人的众领袖也都在那里，屋顶上约有三千男女观看 参孙 逗他们欢乐。
JUDG|16|28|参孙 求告耶和华说：“主耶和华啊，求你眷念我。上帝啊，就这一次，求你赐给我力量，使我向 非利士 人报那挖我双眼的仇。”
JUDG|16|29|参孙 抱住中间支撑庙宇的两根柱子，左手抱一根，右手抱一根。
JUDG|16|30|然后他说：“让我与 非利士 人一起死吧！”他尽力弯腰，庙宇就倒塌了，压住领袖和庙宇内的众人。这样， 参孙 死的时候所杀的人比活着所杀的还多。
JUDG|16|31|他的兄弟和他父亲的全家都下去收他的尸首，抬上去，葬在 琐拉 和 以实陶 中间、他父亲 玛挪亚 的坟墓里。 参孙 作 以色列 的士师二十年。
JUDG|17|1|以法莲 山区有一个人，名叫 米迦 。
JUDG|17|2|他对母亲说：“你的一千一百块银子被人拿走了，为此你发咒起誓，也说给我听。看哪，银子在我这里，是我拿的。”他母亲说：“愿我儿蒙耶和华赐福！”
JUDG|17|3|米迦 把这一千一百块银子还他母亲。他母亲说：“我把这银子分别为圣，亲手献给耶和华，为我儿子造一尊雕刻的像，以及一尊铸成的像。现在我把银子交给你。”
JUDG|17|4|米迦 把银子还他母亲，他母亲把二百块银子交给银匠，去造一尊雕刻的像，以及一尊铸成的像，安置在 米迦 的房子里。
JUDG|17|5|米迦 这个人有了神堂，又造了以弗得和家中的神像，派他的一个儿子作祭司。
JUDG|17|6|那时， 以色列 中没有王，各人照自己眼中看为对的去做。
JUDG|17|7|犹大 的 伯利恒 有一个年轻人，是 犹大 族的人。他是 利未 人，寄居在那里。
JUDG|17|8|这人离开 犹大 的 伯利恒城 ，要找一个可住的地方。他来到 以法莲 山区 米迦 的家，还要往前走。
JUDG|17|9|米迦 对他说：“你从哪里来？”他说：“我从 犹大 的 伯利恒 来。我是 利未 人，要找一个可住的地方。”
JUDG|17|10|米迦 说：“你就住在我这里吧！我以你为父为祭司，每年给你十块银子和一套衣服，以及生活所需的食物。” 利未 人就来了。
JUDG|17|11|利未 人愿意和这人同住；他待这年轻人如自己的儿子一样。
JUDG|17|12|米迦 授这年轻的 利未 人祭司的职任，他就住在 米迦 的家里。
JUDG|17|13|米迦 说：“现在我知道耶和华必恩待我，因为我有 利未 人作我的祭司。”
JUDG|18|1|那时， 以色列 中没有王。 但 支派的人还在觅地居住，因为直到那日，他们还没有在 以色列 支派中抽签得地为业。
JUDG|18|2|但 人从 琐拉 和 以实陶 派本族中的五个勇士，去窥探侦察那地，对他们说：“你们去侦察那地。”他们来到 以法莲 山区 米迦 的家中，就在那里住宿。
JUDG|18|3|他们临近 米迦 的家，听出那年轻的 利未 人的口音，就绕到那里，对他说：“谁领你到这里来？你在这里做什么？你在这里得了什么？”
JUDG|18|4|他对他们说：“ 米迦 如此如此待我，他雇用我，我就作了他的祭司。”
JUDG|18|5|他们对他说：“请你求问上帝，使我们知道所走的道路是否通达。”
JUDG|18|6|祭司对他们说：“你们平平安安去吧，你们所行的道路是在耶和华面前的。”
JUDG|18|7|五人就走了，来到 拉亿 ，见那里的人安居，像 西顿 人的生活一样安宁无虑，那地无人羞辱他们，无人夺取侵略。他们离 西顿 人很远，与世无争 。
JUDG|18|8|五人回到 琐拉 和 以实陶 他们的弟兄那里。他们的弟兄对他们说：“你们怎么了？”
JUDG|18|9|他们说：“起来，我们上去攻打他们吧！我们已经窥探了那地，看哪，那地非常好。你们还要待在这里吗？不要再迟延了，立刻出发去得那地为业吧！
JUDG|18|10|你们去，必来到安居的百姓和两边辽阔的地。上帝已将那地方交在你们手中了；那里不缺地上的任何东西。”
JUDG|18|11|于是 但 族的六百人，各带兵器，从 琐拉 和 以实陶 出发，
JUDG|18|12|上到 犹大 的 基列．耶琳 ，在那里安营。因此那地方名叫 玛哈尼．但 ，直到今日。看哪，它在 基列．耶琳 的西边。
JUDG|18|13|他们从那里往 以法莲 山区去，来到 米迦 的家。
JUDG|18|14|先前窥探 拉亿 地的五个人对他们的弟兄说：“你们知道吗？这些屋子里有以弗得和家中的神像，以及一尊雕刻的像与一尊铸成的像。现在你们要知道该怎么做。”
JUDG|18|15|五人转身，进入 米迦 的家，来到那年轻 利未 人的房间，向他问安。
JUDG|18|16|六百 但 人各带兵器，站在门口。
JUDG|18|17|那窥探这地的五个人上前去，进入里面，拿走雕刻的像、以弗得、家中的神像，以及铸成的像。祭司和带兵器的六百人一同站在门口。
JUDG|18|18|当五个人进入 米迦 的家，拿走雕刻的像、以弗得、家中的神像，以及铸成的像，祭司对他们说：“你们做什么呢？”
JUDG|18|19|他们对他说：“不要作声，用手捂口，跟我们去吧！我们必以你为父为祭司。你作一家的祭司好呢？还是作 以色列 一支派一族的祭司好呢？”
JUDG|18|20|祭司心里欢喜，拿着以弗得和家中的神像，以及雕刻的像，跟这些百姓走了。
JUDG|18|21|他们转身离开那里，把孩子、牲畜、财物安排在前头。
JUDG|18|22|他们离了 米迦 的家已远， 米迦 家附近的邻居被召来，追赶 但 人。
JUDG|18|23|他们呼叫 但 人， 但 人回头对 米迦 说：“你召集这许多人来做什么呢？”
JUDG|18|24|米迦 说：“你们把我所造的神像，还有祭司，都带走了，我还有什么呢？你怎么还对我说‘你在做什么’呢？”
JUDG|18|25|但 人对 米迦 说：“你不要让我们再听见你的声音，恐怕这群恼怒成性的人会攻击你们，你和你的全家就会丧命。”
JUDG|18|26|但 人仍走他们的路。 米迦 见他们的势力比自己强，就转身回家去了。
JUDG|18|27|但 人把 米迦 造的神像和他的祭司带走，来到 拉亿 安宁无虑的百姓那里，用刀杀了他们，放火烧了那城。
JUDG|18|28|没有人来搭救，因为这城离 西顿 很远，他们又与世无争；这城在靠近 伯．利合 的平原。 但 人建造这城，在那里居住，
JUDG|18|29|并照着他们祖先 以色列 之子 但 的名字，给这城起名叫 但 。原先这城名叫 拉亿 。
JUDG|18|30|但 人为自己设立了那雕刻的像。 摩西 的孙子， 革舜 的儿子 约拿单 和他的子孙作 但 支派的祭司，直到那地遭掳掠的日子。
JUDG|18|31|上帝的家在 示罗 多少日子， 但 人为自己设立 米迦 所雕刻的像也在 但 多少日子。
JUDG|19|1|当 以色列 中没有王的时候，有一个 利未 人寄居 以法莲 山区的边界，他娶了一个 犹大伯利恒 的女子为妾。
JUDG|19|2|这妾对丈夫生气 ，离开丈夫，回到 犹大伯利恒 的父家，在那里住了四个月。
JUDG|19|3|她的丈夫起来，带着一个仆人、两匹驴跟着她去，要用好话劝她回来。女子就带丈夫进到父亲家里。女子的父亲看见了他，就欢欢喜喜地迎接他。
JUDG|19|4|这岳父，就是女子的父亲，留他住了三天。他们在那里吃喝，住宿。
JUDG|19|5|第四日，他们清早起来， 利未 人起身要走，女子的父亲对女婿说：“先吃点东西，加添心力，然后你们才走。”
JUDG|19|6|于是二人坐下，一同吃喝。女子的父亲对那人说：“请你答应再住一夜，使你的心舒畅。”
JUDG|19|7|那人起身要走，他岳父挽留他，他就留下，在那里又住了一夜。
JUDG|19|8|第五日，他清早起来要走，女子的父亲说：“来，请加添心力，留到太阳偏西吧。”于是二人一同再吃。
JUDG|19|9|那人同他的妾和仆人起身要走，但他岳父，就是女子的父亲，对他说：“看哪，太阳下山，天快晚了，你们再住一夜吧。看哪，太阳偏西了，就在这里住宿，使你的心舒畅，明天你们一早起来上路，回你的帐棚去。”
JUDG|19|10|那人不愿再住一夜，就备上两匹驴，带着他的妾起身走了，来到 耶布斯 的对面， 耶布斯 就是 耶路撒冷 。
JUDG|19|11|将近 耶布斯 的时候，太阳快下山了，仆人对主人说：“来吧，我们进这 耶布斯 人的城，在这里住宿。”
JUDG|19|12|主人对他说：“我们不可进入外邦人的城，那不是 以色列 人的地方，我们越过这里到 基比亚 去吧。”
JUDG|19|13|他又对仆人说：“来，让我们到 基比亚 或 拉玛 的一个地方住宿。”
JUDG|19|14|于是他们越过那里往前走，将到 便雅悯 的 基比亚 的时候，太阳已经下山了。
JUDG|19|15|他们进入 基比亚 要在那里住宿。他来坐在城里的广场上，但没有人接待他们到家里住宿。
JUDG|19|16|看哪，晚上有一个老人从田间做工回来。他是 以法莲 山区的人，寄居在 基比亚 ；那地方的人是 便雅悯 人。
JUDG|19|17|老人举目看见那过路的人在城里的广场上，就说：“你从哪里来？要到哪里去？”
JUDG|19|18|他对他说：“我们从 犹大 的 伯利恒 过来，要到 以法莲 山区的边界去。我是那里的人，去了 犹大 的 伯利恒 ，现在要到耶和华的家去，却没有人接待我到他的家。
JUDG|19|19|其实我有饲料草料可以喂驴，我和你的使女，以及与我们在一起的仆人都有饼有酒，什么都不缺。”
JUDG|19|20|老人说：“愿你平安！你所需用的我都会给你们，只是不可在广场上过夜。”
JUDG|19|21|于是老人领他到家里，喂上驴。他们洗了脚，就吃喝起来。
JUDG|19|22|他们心里欢乐的时候，看哪，城中的无赖围住房子，连连叩门，对老人，这家的主人说：“把那进你家的人带出来，我们要与他交合。”
JUDG|19|23|这家的主人出来对他们说：“弟兄们，不要做这样的恶事。这人既然进了我的家，你们就不要做这样可耻的事。
JUDG|19|24|看哪，我有个女儿还是处女，还有这人的妾，我把她们领出来任由你们污辱她们，就照你们看为好的对待她们吧！但对这人你们不要做这样可耻的事。”
JUDG|19|25|那些人却不肯听从他。那人抓住他的妾，把她拉出去给他们。他们强奸了她，整夜凌辱她，直到早晨，天色快亮才放她走。
JUDG|19|26|到了早晨，妇人回来，仆倒在留她主人住宿的那人的家门前，直到天亮。
JUDG|19|27|早晨，她的主人起来开了门，出去要上路。看哪，那妇人，他的妾倒在屋子门前，双手搭在门槛上。
JUDG|19|28|他对妇人说：“起来，我们走吧！”妇人却没有回应。那人就将她驮在驴上，起身回自己的地方去了。
JUDG|19|29|到了家里，他拿刀，抓住他的妾，把她的尸身切成十二块，分送到 以色列 全境。
JUDG|19|30|凡看见的人都说：“自从 以色列 人离开 埃及 地上来，直到今日，像这样的事还没有发生过，也没有见过。大家应当想一想，商讨一下再说。”
JUDG|20|1|于是 以色列 众人从 但 到 别是巴 ，以及从 基列 地出来，如同一人，聚集在 米斯巴 耶和华那里。
JUDG|20|2|以色列 各支派中众百姓的领袖，都站在上帝百姓的会中。拿刀的步兵共有四十万。
JUDG|20|3|便雅悯 人听见 以色列 人上了 米斯巴 。 以色列 人说：“请说，这恶事是怎么发生的呢？”
JUDG|20|4|那 利未 人，就是被害妇人的丈夫，回答说：“我和我的妾来到 便雅悯 的 基比亚 住宿。
JUDG|20|5|基比亚 人夜间起来攻击我，包围我住的屋子。他们想要杀我，并把我的妾污辱致死。
JUDG|20|6|我把我的妾切成块，分送到 以色列 得为业的全地，因为 基比亚 人在 以色列 中做了邪恶可耻的事。
JUDG|20|7|看哪，你们大家， 以色列 人哪，在此提出你们的建议和对策吧！”
JUDG|20|8|众百姓都起来如同一人，说：“我们谁也不回自己的帐棚，谁也不回自己的家去！
JUDG|20|9|现在，我们要这样对付 基比亚 ，照所抽的签去攻打他们。
JUDG|20|10|我们要在 以色列 各支派中，一百人选十人，一千人选一百人，一万人选一千人，为那到 便雅悯 的 迦巴 去的士兵运粮；因为 基比亚 在 以色列 中行了可耻的事。”
JUDG|20|11|于是 以色列 众人彼此联合如同一人，聚集攻击那城。
JUDG|20|12|以色列 众支派派人去，问 便雅悯 支派的各家说：“你们中间怎么做了这样的恶事呢？
JUDG|20|13|现在你们要把 基比亚 的那些无赖交出来，我们好处死他们，从 以色列 中除掉这恶。” 便雅悯 人却不肯听从他们弟兄 以色列 人的话。
JUDG|20|14|便雅悯 人从各城聚集到 基比亚 ，出来要与 以色列 人打仗。
JUDG|20|15|那日， 便雅悯 人从各城里征召了拿刀的士兵，共有二万六千，另外还从 基比亚 居民中征召七百个精兵。
JUDG|20|16|全军中有特选的七百个精兵，都是惯用左手的，个个能用机弦甩石，毫发不差。
JUDG|20|17|以色列 人，除了 便雅悯 之外，共征召了四十万拿刀的，个个都是战士。
JUDG|20|18|以色列 人起来，上到 伯特利 去求问上帝说：“我们中间谁当首先上去与 便雅悯 人争战呢？”耶和华说：“ 犹大 先上去。”
JUDG|20|19|以色列 人早晨起来，对着 基比亚 安营。
JUDG|20|20|以色列 人出来与 便雅悯 人打仗， 以色列 人在 基比亚 对着他们摆阵。
JUDG|20|21|便雅悯 人从 基比亚 出来，当日把 以色列 中二万二千人杀倒在地。
JUDG|20|22|以色列 人的士兵鼓起勇气，在第一日摆阵的地方又摆阵。
JUDG|20|23|因 以色列 人上去，在耶和华面前哀哭，直到晚上。他们求问耶和华说：“我可以再出兵与我弟兄 便雅悯 人打仗吗？”耶和华说：“可以上去攻打他们。”
JUDG|20|24|第二日， 以色列 人就上前攻击 便雅悯 人。
JUDG|20|25|便雅悯 人也在第二日从 基比亚 出来与他们交战，又把 以色列 人一万八千个拿刀的士兵杀倒在地。
JUDG|20|26|以色列 众人和全体士兵上到 伯特利 ，坐在耶和华面前哭泣。那日，他们禁食直到晚上，又在耶和华面前献燔祭和平安祭。
JUDG|20|27|以色列 人去求问耶和华；那时，上帝的约柜在那里。
JUDG|20|28|那时， 亚伦 的孙子， 以利亚撒 的儿子 非尼哈 侍立在约柜前。他们说：“我可以再出去与我弟兄 便雅悯 人打仗吗？还是停战呢？”耶和华说：“你们可以上去，因为明日我必把他交在你手中。”
JUDG|20|29|以色列 在 基比亚 的四围设下埋伏。
JUDG|20|30|第三日， 以色列 人又上去攻击 便雅悯 人，在 基比亚 前摆阵，与前两次一样。
JUDG|20|31|便雅悯 人也出来迎敌，就被引诱出城外。在田间的两条路上，一条通往 伯特利 ，一条通往 基比亚 ，他们像前两次一样，动手杀了约三十个 以色列 人。
JUDG|20|32|便雅悯 人说：“他们仍像以前一样败在我们面前。”但 以色列 人说：“让我们逃跑，引诱他们离开城到路上来。”
JUDG|20|33|以色列 众人都起来，在 巴力．他玛 摆阵， 以色列 的伏兵从 马利．迦巴 埋伏的地方冲上前去。
JUDG|20|34|全 以色列 中的一万精兵来到 基比亚 前，战争十分激烈。 便雅悯 人却不知道灾祸临近了。
JUDG|20|35|耶和华在 以色列 面前击打 便雅悯 。那日， 以色列 人歼灭二万五千一百个 便雅悯 人，都是拿刀的士兵。
JUDG|20|36|便雅悯 人看到自己战败了。 以色列 人因为信任在 基比亚 前所设的伏兵，就在 便雅悯 人面前假装撤退。
JUDG|20|37|伏兵迅速闯进 基比亚 ；他们继续前进，用刀杀死全城的人。
JUDG|20|38|以色列 人预先与伏兵约定在城内放火，以上腾的烟为信号。
JUDG|20|39|以色列 人从阵上撤退， 便雅悯 人动手杀死 以色列 人，约有三十个，就说：“他们仍像以前一样败在我们面前。”
JUDG|20|40|当烟如柱一般从城中上腾的时候， 便雅悯 人回头，看哪，全城已经浓烟冲天了。
JUDG|20|41|以色列 人又转身回来， 便雅悯 人就很惊惶，因为看见灾祸临到自己了。
JUDG|20|42|他们在 以色列 人面前转身往旷野逃跑，战况对他们不利，那从城里出来的也去夹攻，杀灭他们。
JUDG|20|43|以色列 人围攻 便雅悯 人，追赶他们，在他们歇脚之处，直到向日出方向的 基比亚 的对面，践踏他们。
JUDG|20|44|便雅悯 人倒下的有一万八千名，这些全都是勇士。
JUDG|20|45|其余的人转身往旷野逃跑，到 临门岩 去。 以色列 人在路上杀了五千人，如拾穗一样，紧追他们直到 基顿 ，又杀了二千人。
JUDG|20|46|那日 便雅悯 人倒下的有二万五千名，这些全都是拿刀的勇士。
JUDG|20|47|有六百人转身往旷野逃跑，到了 临门岩 ，在 临门岩 住了四个月。
JUDG|20|48|以色列 人又转回去攻击 便雅悯 人，凡经过的各城，其中的人和牲畜都用刀杀了，又放火烧了所经过的一切城镇。
JUDG|21|1|以色列 人在 米斯巴 曾起誓说：“我们中谁都不把女儿嫁给 便雅悯 人。”
JUDG|21|2|以色列 人来到 伯特利 ，坐在那里直到晚上，在上帝面前放声大哭，
JUDG|21|3|说：“耶和华－ 以色列 的上帝啊，为何 以色列 中会发生这样的事，使 以色列 今日缺了一个支派呢？”
JUDG|21|4|次日，百姓清早起来，在那里筑了一座坛，献燔祭和平安祭。
JUDG|21|5|以色列 人说：“ 以色列 各支派中，谁没有同会众一起上到耶和华那里呢？”因为 以色列 人曾起重誓说：“凡不上 米斯巴 到耶和华那里的，必被处死。”
JUDG|21|6|以色列 人怜悯他们的弟兄 便雅悯 ，说：“如今 以色列 中断绝一个支派了。
JUDG|21|7|我们既然向耶和华起誓说，必不把我们的女儿嫁给 便雅悯 人，现在我们该怎么办，使他们剩下的人可以娶妻呢？”
JUDG|21|8|他们又说：“ 以色列 支派中谁没有上 米斯巴 到耶和华那里呢？”看哪， 基列 的 雅比 没有一人进营到会众那里，
JUDG|21|9|百姓被数点的时候，看哪， 基列 的 雅比 居民没有一人在那里。
JUDG|21|10|会众就派一万二千名大勇士，吩咐他们说：“你们去用刀把 基列 的 雅比 居民连妇女带孩子都杀了。
JUDG|21|11|这是你们当做的事：要把所有男人和曾与男人同房共寝的女人全都杀了。”
JUDG|21|12|他们在 基列 的 雅比 居民中，找到四百个未曾与男人同房共寝的处女，就带她们到 迦南 地的 示罗 营里。
JUDG|21|13|全会众派人到 临门岩 的 便雅悯 人那里，与他们讲和。
JUDG|21|14|当时 便雅悯 人回来了， 以色列 人就把所留下， 基列 的 雅比 活着的女子嫁给他们，可是还是不够。
JUDG|21|15|百姓怜悯 便雅悯 人，因为耶和华使 以色列 支派中有一个缺口。
JUDG|21|16|会众中的长老说：“ 便雅悯 中的女子既然都除灭了，我们该怎么办，使剩下的人可以娶妻呢？”
JUDG|21|17|他们又说：“ 便雅悯 逃脱的人应当有地业，免得 以色列 中的一个支派被涂去。
JUDG|21|18|只是我们不能把自己的女儿嫁给他们。”因为 以色列 人曾起誓说：“把女儿嫁给 便雅悯 人的必受诅咒。”
JUDG|21|19|他们又说：“看哪，一年一度耶和华的节期正在 示罗 举行。” 示罗 位于 利波拿 的南边， 伯特利 的北边，从 伯特利 往 示剑 大路的东边。
JUDG|21|20|他们吩咐 便雅悯 人说：“你们去，躲在葡萄园中，
JUDG|21|21|观看；看哪，若 示罗 的女子出来跳舞，你们就从葡萄园出来，各人从 示罗 的女子中抢一个为妻，然后到 便雅悯 地去。
JUDG|21|22|他们的父亲或兄弟若来与我们争论，我们就对他们说：‘请看我们的情面恩待这些人吧！因为我们在战争的时候没有给他们任何人留下女子为妻。这次也不是你们给他们的，若是你们给的，就算有罪了。’”
JUDG|21|23|于是 便雅悯 人就照样做了，按照他们的人数，把从跳舞女子中抢来的娶为妻子，带回自己的地业，重建城镇，居住在其中。
JUDG|21|24|那时 以色列 人离开那里，各自回到自己的支派、宗族；他们从那里起行，各自回到自己的地业去了。
JUDG|21|25|那时， 以色列 中没有王，各人照自己眼中看为对的去做。
RUTH|1|1|士师统治的时候，国中有饥荒。在 犹大 的 伯利恒 ，有一个人带着妻子和两个儿子往 摩押 地去寄居。
RUTH|1|2|这人名叫 以利米勒 ，他的妻子名叫 拿娥米 ；他两个儿子，一个名叫 玛伦 ，一个名叫 基连 ，都是 犹大伯利恒 的 以法他 人。他们到了 摩押 地，就住在那里。
RUTH|1|3|后来 拿娥米 的丈夫 以利米勒 死了，剩下她和两个儿子。
RUTH|1|4|两个儿子娶了 摩押 女子，一个名叫 俄珥巴 ，第二个名叫 路得 ，在那里住了约有十年。
RUTH|1|5|玛伦 和 基连 二人也死了，剩下 拿娥米 ，没有丈夫，也没有儿子。
RUTH|1|6|拿娥米 与两个媳妇起身，要从 摩押 地回去，因为她在 摩押 地听见耶和华眷顾自己的百姓，赐粮食给他们。
RUTH|1|7|她和两个媳妇就起行，离开所住的地方，上路回 犹大 地去。
RUTH|1|8|拿娥米 对两个媳妇说：“你们各自回娘家去吧！愿耶和华恩待你们，像你们待已故的人和我一样。
RUTH|1|9|愿耶和华使你们各自在新的丈夫家中得归宿！”于是 拿娥米 与她们亲吻，她们就放声大哭，
RUTH|1|10|对她说：“不，我们要与你一同回你的百姓那里去。”
RUTH|1|11|拿娥米 说：“我的女儿啊，回去吧！为何要跟我去呢？我还能生儿子作你们的丈夫吗？
RUTH|1|12|我的女儿啊，回去吧！我年纪老了，不能再有丈夫。就算我还有希望，今夜有丈夫，而且也生了儿子，
RUTH|1|13|你们岂能等着他们长大呢？你们能守住自己不嫁人吗？我的女儿啊，不要这样。我比你们更苦，因为耶和华伸手击打我。”
RUTH|1|14|两个媳妇又放声大哭， 俄珥巴 与婆婆吻别，但是 路得 却紧跟着 拿娥米 。
RUTH|1|15|拿娥米 说：“看哪，你嫂嫂已经回她的百姓和她的神明那里去了，你也跟你嫂嫂回去吧！”
RUTH|1|16|路得 说： “不要劝我离开你， 转去不跟随你。 你往哪里去， 我也往哪里去； 你在哪里住， 我也在哪里住； 你的百姓就是我的百姓； 你的上帝就是我的上帝。
RUTH|1|17|你死在哪里， 我也死在哪里，葬在哪里。 只有死能使你我分离； 不然，愿耶和华重重惩罚我！”
RUTH|1|18|拿娥米 见 路得 决意要跟自己去，就不再对她说什么了。
RUTH|1|19|于是二人同行，来到 伯利恒 。她们到了 伯利恒 ，全城因她们骚动起来。妇女们说：“这是 拿娥米 吗？”
RUTH|1|20|拿娥米 对她们说： “不要叫我 拿娥米 ， 要叫我 玛拉 ， 因为全能者使我受尽了苦。
RUTH|1|21|我满满地出去， 耶和华使我空空地回来。 耶和华使我受苦， 全能者降祸于我。 你们为何还叫我 拿娥米 呢？”
RUTH|1|22|拿娥米 从 摩押 地回来了，她的媳妇 摩押 女子 路得 跟她在一起。她们到了 伯利恒 ，正是开始收割大麦的时候。
RUTH|2|1|拿娥米 有一个亲戚，是她丈夫 以利米勒 本族的人，名叫 波阿斯 ，是个大财主。
RUTH|2|2|摩押 女子 路得 对 拿娥米 说：“让我到田里去拾取麦穗，我在谁的眼中蒙恩，就跟在谁的身后。” 拿娥米 说：“女儿啊，你去吧。”
RUTH|2|3|路得 就去了。她来到田间，在收割的人身后拾取麦穗。她恰巧来到 以利米勒 本族的人 波阿斯 那块田里。
RUTH|2|4|看哪， 波阿斯 正从 伯利恒 来，对收割的人说：“愿耶和华与你们同在！”他们对他说：“愿耶和华赐福给你！”
RUTH|2|5|波阿斯 对监督收割的仆人说：“那是谁家的女子？”
RUTH|2|6|监督收割的仆人回答说：“她是 摩押 女子，跟随 拿娥米 从 摩押 地回来的。
RUTH|2|7|她说：‘请你容许我拾取麦穗，在收割的人身后捡禾捆中掉落的麦穗。’她就来了，从早晨直到如今，除了在屋子里坐一会儿，她都留在这里。”
RUTH|2|8|波阿斯 对 路得 说：“女儿啊，听我说，不要到别人田里去拾取麦穗，也不要离开这里，要紧跟着我的女仆们。
RUTH|2|9|你要看好我的仆人正在哪块田收割，就跟着女仆们去。我已经吩咐仆人不可侵犯你。你渴了，可以到水缸那里喝仆人打来的水。”　
RUTH|2|10|路得 就脸伏于地叩拜，对他说：“我既是外邦女子，怎么会在你眼中蒙恩，使你这样照顾我呢？”
RUTH|2|11|波阿斯 回答她说：“自从你丈夫死后，凡你向婆婆所行的，以及你离开父母和你的出生地，到素不相识的百姓中，这些事人都告诉我了。
RUTH|2|12|愿耶和华照你所行的报偿你。你来投靠在耶和华－ 以色列 上帝的翅膀下，愿你满得他的报偿。”
RUTH|2|13|路得 说：“我主啊，愿我在你眼前蒙恩。我虽然不及你的一个婢女，你还安慰我，对你的婢女说关心的话。”
RUTH|2|14|吃饭的时候， 波阿斯 对 路得 说：“你到这里来吃些饼，把你的一块蘸在醋里。” 路得 就在收割的人旁边坐下。 波阿斯 把烘了的穗子递给她。她吃饱了，还有剩余的。
RUTH|2|15|她又起来拾取麦穗， 波阿斯 吩咐仆人说：“她即使在禾捆中拾取麦穗，也不可羞辱她。
RUTH|2|16|你们还要从捆里抽一些出来，留给她拾取，不可责备她。”
RUTH|2|17|这样， 路得 在田间拾取麦穗，直到晚上。她把所拾取的麦穗打了约有一伊法的大麦。
RUTH|2|18|路得 把所拾取的带进城去给婆婆看，又把她吃饱所剩的拿出来，给了婆婆。
RUTH|2|19|婆婆问她说：“你今日在哪里拾取麦穗？在哪里做工呢？愿那照顾你的得福。” 路得 告诉婆婆，她在谁那里做工，说：“我今日在一个名叫 波阿斯 的人那里做工。”
RUTH|2|20|拿娥米 对媳妇说：“愿那人蒙耶和华赐福，因为他不断地恩待活人死人。” 拿娥米 又对她说：“那人是我们本族的人，是一个可以赎我们产业的至亲。”
RUTH|2|21|摩押 女子 路得 说：“他还对我说：‘你要紧跟着我的仆人拾取麦穗，直到他们把我所有的庄稼收割完毕。’”
RUTH|2|22|拿娥米 对媳妇 路得 说：“女儿啊，你要跟着他的女仆出去，免得你在别人的田间受人骚扰。”
RUTH|2|23|于是 路得 紧跟着 波阿斯 的女仆拾取麦穗，直到大麦和小麦收割完毕。 路得 仍与婆婆同住。
RUTH|3|1|路得 的婆婆 拿娥米 对她说：“女儿啊，我不该为你找个归宿，使你享福吗？
RUTH|3|2|你与 波阿斯 的女仆常在一处，现在， 波阿斯 不是我们的亲人吗？看哪，他今夜将在禾场簸大麦。
RUTH|3|3|你要沐浴抹膏，穿上外衣，下到禾场，一直到那人吃喝完了，都不要让他认出你来。
RUTH|3|4|他躺下的时候，你看准他躺卧的地方，就进去掀露他的脚，躺卧在那里，他必告诉你所当做的事。”
RUTH|3|5|路得 说：“凡你所吩咐我的，我必遵行。”
RUTH|3|6|路得 就下到禾场，照她婆婆吩咐她的一切去做。
RUTH|3|7|波阿斯 吃喝完了，心情畅快，就去躺卧在麦堆旁边。 路得 悄悄走来，掀露他的脚，躺卧在那里。
RUTH|3|8|到了半夜，那人惊醒，翻过身来，看哪，有个女子躺在他的脚旁。
RUTH|3|9|他就说：“你是谁？” 路得 说：“我是你的使女 路得 。请你用你衣服的边来遮盖你的使女，因为你是可以赎我产业的至亲。”
RUTH|3|10|波阿斯 说：“女儿啊，愿你蒙耶和华赐福。你后来的忠诚比先前的更美，因为无论贫富的年轻人，你都没有跟从。
RUTH|3|11|女儿啊，现在不要惧怕，凡你所说的，我必为你做，因为我城里的百姓都知道你是个贤德的女子。
RUTH|3|12|现在，我的确是一个可以赎你产业的至亲，可是还有一个人比我更亲。
RUTH|3|13|你今夜在这里住宿，明早他若肯为你尽至亲的本分，很好，就由他吧！倘若他不肯，我指着永生的耶和华起誓，我必为你尽上至亲的本分。你只管躺到早晨。”
RUTH|3|14|路得 就在他脚旁躺到早晨，在人还无法彼此辨认的时候就起来了。 波阿斯 说：“不可让人知道有女子到禾场来。”　
RUTH|3|15|他又对 路得 说：“把你所披的外衣拿来，握紧它。”她就握紧外衣， 波阿斯 量了六簸箕的大麦，帮 路得 扛上，他就进城去了 。”
RUTH|3|16|路得 回到婆婆那里，婆婆说：“女儿啊，怎么样了 ？” 路得 就把那人向她所做的一切都告诉了婆婆，
RUTH|3|17|又说：“那人给了我这六簸箕的大麦，对我说：‘你不可空手回去见婆婆。’”
RUTH|3|18|婆婆说：“女儿啊，等着吧，看这事结果如何，因为那人今日不办妥这事，必不罢休。”
RUTH|4|1|波阿斯 上到城门，坐在那里，看哪， 波阿斯 所说那个可以赎产业的至亲经过。 波阿斯 说：“某某先生，请你转回来，坐在这里。”他就转回来坐下。
RUTH|4|2|波阿斯 又请了本城的十个长老来，对他们说：“请你们坐在这里。”他们就都坐下。
RUTH|4|3|波阿斯 对那至亲说：“从 摩押 地回来的 拿娥米 ，现在要卖我们弟兄 以利米勒 的那块地。
RUTH|4|4|我想我应该向你说清楚：你可以买那块地，当着在座的众人和我百姓的长老面前，你若要赎就赎吧！倘若你不赎 就告诉我，让我知道，因为除了你以外，没有人可以先赎，在你之后才轮到我。”那人说：“我要赎。”
RUTH|4|5|波阿斯 说：“你从 拿娥米 和 摩押 女子 路得 手中买这地的时候，也当买死人的妻子，使死人在产业上留名。”
RUTH|4|6|那至亲说：“这样我就不能赎了，免得对我的产业有损。你尽管去赎我所当赎的吧，我不能赎了！”
RUTH|4|7|从前，在 以色列 中要确认任何交易，无论是赎业或买卖，一方必须脱鞋给另一方。 以色列 中都以此为证。
RUTH|4|8|那至亲对 波阿斯 说：“你自己买吧！”于是把鞋脱了下来。
RUTH|4|9|波阿斯 对长老和所有在场的百姓说：“你们今日都是证人；凡属 以利米勒 ，以及 基连 和 玛伦 的，我都从 拿娥米 手中买下来了。
RUTH|4|10|我也娶 玛伦 的妻子 摩押 女子 路得 ，好让死人可以在产业上留名，免得他的名在本族本乡的城门中消失了。你们今日都是证人。”
RUTH|4|11|在城门坐着的所有百姓和长老说：“我们都是证人。愿耶和华使进你家的这女子，像建立 以色列 家的 拉结 和 利亚 二人一样。又愿你在 以法他 得亨通，在 伯利恒 有名声。
RUTH|4|12|愿耶和华从这年轻女子赐你后裔，使你的家像 她玛 从 犹大 所生 法勒斯 的家一样。”
RUTH|4|13|于是， 波阿斯 娶了 路得 为妻，与她同房。耶和华使她怀孕生了一个儿子。
RUTH|4|14|妇女们对 拿娥米 说：“耶和华是应当称颂的！因为他今日没有使你断绝可以赎产业的至亲。愿这孩子在 以色列 中得名声。
RUTH|4|15|他必振奋你的精神，奉养你的晚年，因为他是爱慕你的媳妇所生的。有这样的媳妇，比有七个儿子更好！”
RUTH|4|16|拿娥米 接过孩子来，抱在怀中抚养他。
RUTH|4|17|邻居的妇人给孩子起名，说：“ 拿娥米 得了一个孩子了！”她们就给他起名叫 俄备得 。 俄备得 是 耶西 的父亲，是 大卫 的祖父。
RUTH|4|18|这是 法勒斯 的后代： 法勒斯 生 希斯仑 ；
RUTH|4|19|希斯仑 生 兰 ； 兰 生 亚米拿达 ；
RUTH|4|20|亚米拿达 生 拿顺 ； 拿顺 生 撒门 ；
RUTH|4|21|撒门 生 波阿斯 ； 波阿斯 生 俄备得 ；
RUTH|4|22|俄备得 生 耶西 ； 耶西 生 大卫 。
1SAM|1|1|以法莲 山区有一个 拉玛 的 琐非 人 ，名叫 以利加拿 ，他是 苏弗 的玄孙， 托户 的曾孙， 以利户 的孙子， 耶罗罕 的儿子，是 以法莲 人。
1SAM|1|2|他有两个妻子：一个名叫 哈拿 ，另一个名叫 毗尼拿 。 毗尼拿 有孩子， 哈拿 却没有孩子。
1SAM|1|3|这人每年从本城上到 示罗 ，敬拜万军之耶和华，向他献祭。在那里有 以利 的两个儿子 何弗尼 和 非尼哈 当耶和华的祭司。
1SAM|1|4|每逢献祭的日子， 以利加拿 把祭肉分给他的妻子 毗尼拿 和 毗尼拿 所生的儿女。
1SAM|1|5|他给 哈拿 的却是双分，因为他爱 哈拿 。耶和华却不使 哈拿 生育。
1SAM|1|6|她的对头 毗尼拿 因耶和华不使 哈拿 生育，就常常惹她发怒，要使她生气。
1SAM|1|7|年年都是如此。每当她上到耶和华殿的时候， 毗尼拿 就这样惹她发怒，以致她哭泣不吃饭。
1SAM|1|8|她丈夫 以利加拿 对她说：“ 哈拿 ，你为何哭泣？为何不吃饭？为何伤心难过呢？有我不比有十个儿子更好吗？”
1SAM|1|9|他们在 示罗 吃喝完了， 哈拿 就站起来。祭司 以利 坐在耶和华殿门框旁边的位子上。
1SAM|1|10|哈拿 心里愁苦，就痛痛哭泣，向耶和华祈祷。
1SAM|1|11|她许愿说：“万军之耶和华啊，你若垂顾你使女的苦情，眷念不忘你的使女，赐你的使女一个子嗣，我必使他终生归给耶和华，不用剃刀剃他的头。”
1SAM|1|12|哈拿 在耶和华面前不住地祈祷， 以利 注意她的嘴。
1SAM|1|13|哈拿 心中默祷，只动嘴唇，听不到她的声音，因此 以利 以为她喝醉了。
1SAM|1|14|以利 对她说：“你要醉到几时呢？不要再喝酒了！”
1SAM|1|15|哈拿 回答说：“我主啊，不是这样。我是心里愁苦的妇人，清酒烈酒都没有喝，只在耶和华面前倾心吐意。
1SAM|1|16|不要将你的使女看作不正经的女子。我因极其难过和生气，所以一直祷告到如今。”
1SAM|1|17|以利 回答说：“平平安安地回去吧。愿 以色列 的上帝允准你向他所求的！”
1SAM|1|18|哈拿 说：“愿你的婢女在你眼前蒙恩。”于是妇人上路，去吃饭，脸上不再带愁容了。
1SAM|1|19|他们清早起来，在耶和华面前敬拜，就回去，往 拉玛 自己的家里。 以利加拿 和妻子 哈拿 同房，耶和华顾念 哈拿 。
1SAM|1|20|时候到了， 哈拿 怀孕生了一个儿子， 哈拿 给他起名叫 撒母耳 ，说：“这是我从耶和华那里求来的。”
1SAM|1|21|以利加拿 和他全家都上去，要向耶和华献年祭和还愿祭。
1SAM|1|22|哈拿 却没有上去，因为她对丈夫说：“等孩子断了奶，我就带他上去朝见耶和华，让他永远住在那里。”
1SAM|1|23|她丈夫 以利加拿 对她说：“就照你看为好的去做吧！可以留到儿子断了奶，愿耶和华应验他的话。”于是妇人留在家里乳养儿子，直到断了奶。
1SAM|1|24|断奶之后，她就带着孩子，连同一头三岁的公牛 ，一伊法细面 ，一皮袋酒，上 示罗 耶和华的殿去。那时，孩子还小。
1SAM|1|25|他们宰了公牛，就领孩子到 以利 面前。
1SAM|1|26|妇人说：“我主啊，请容许我说，我向你，我的主起誓，从前在你这里站着祈求耶和华的那妇人就是我。
1SAM|1|27|我祈求为要得这孩子，耶和华已将我向他所求的赐给我了。
1SAM|1|28|所以，我将这孩子献给耶和华，使他终生归给耶和华。” 他就在那里敬拜耶和华。
1SAM|2|1|哈拿 祷告说： “我的心因耶和华快乐， 我的角因耶和华高举。 我的口向仇敌张开； 我因你的救恩欢欣。
1SAM|2|2|“没有一位圣者像耶和华， 除你以外没有别的了， 也没有磐石像我们的上帝。
1SAM|2|3|不要夸口说骄傲的话， 也不要口出狂妄的言语， 因耶和华是有知识的上帝， 人的行为被他衡量。
1SAM|2|4|勇士的弓折断， 跌倒的人以力量束腰。
1SAM|2|5|饱足的人作雇工求食； 饥饿的人也不再饥饿。 不生育的生了七个； 儿女多的反倒孤独。
1SAM|2|6|耶和华使人死，也使人活， 使人下阴间，也使人往上升。
1SAM|2|7|耶和华使人贫穷，也使人富足； 使人降卑，也使人升高。
1SAM|2|8|他从灰尘里抬举贫寒人， 从粪堆中提拔贫穷人， 使他们与贵族同坐， 继承荣耀的座位。 地的柱子属耶和华， 他将世界立在其上。
1SAM|2|9|“他必保护他圣民的脚步， 但恶人却在黑暗中毁灭， 因为人不是靠力量得胜。
1SAM|2|10|与耶和华相争的，必被打碎； 他必从天上打雷攻击他们。 耶和华审判地极的人， 将力量赐给所立的王， 高举受膏者的角。”
1SAM|2|11|以利加拿 往 拉玛 回自己的家去了。那孩子在 以利 祭司面前事奉耶和华。
1SAM|2|12|以利 的两个儿子是无赖，不认识耶和华。
1SAM|2|13|这二祭司对待百姓的规矩是这样：凡有人献祭，正煮肉的时候，祭司的仆人就手拿三齿的叉子来，
1SAM|2|14|将叉子往盆里，或锅里，或釜里，或壶里一插，插上来的肉，祭司都拿了去。他们对所有上到 示罗 的 以色列 人都这样做。
1SAM|2|15|甚至在未烧脂肪之前，祭司的仆人就来对献祭的人说：“把肉给祭司，让他烤吧。他不要拿你煮过的肉，要生的。”
1SAM|2|16|献祭的人若说：“他们必须先烧脂肪，然后你才可以随意拿。”仆人就说：“不，你立刻给我，不然我就要抢了。”
1SAM|2|17|这些年轻人的罪在耶和华面前非常严重，因为这些人藐视耶和华的祭物。
1SAM|2|18|那时， 撒母耳 还是孩子，穿着细麻布的以弗得，侍立在耶和华面前。
1SAM|2|19|他母亲每年为他做一件小外袍，同丈夫上来献年祭的时候带来给他。
1SAM|2|20|以利 为 以利加拿 和他妻子祝福，说：“愿耶和华由这妇人再赐你后裔，代替从耶和华求来的孩子。”他们就回自己的地方去了。
1SAM|2|21|耶和华眷顾 哈拿 ，她就怀孕生了三个儿子，两个女儿。那孩子 撒母耳 在耶和华面前渐渐长大。
1SAM|2|22|以利 年纪老迈，听见他两个儿子对 以色列 众人所做一切的事，又听见他们与会幕门前伺候的妇人同寝，
1SAM|2|23|就对他们说：“你们为何做这样的事呢？我从这众百姓听见了你们的恶行。
1SAM|2|24|我儿啊，不可这样！我听到耶和华的百姓传出你们不好的名声 。
1SAM|2|25|人若得罪人，有上帝 可以裁决；人若得罪耶和华，谁能为他代求呢？”然而他们还是不听父亲的话，因为耶和华想要他们死。
1SAM|2|26|撒母耳 这孩子渐渐长大，耶和华与人越发喜爱他。
1SAM|2|27|有神人来见 以利 ，对他说：“耶和华如此说：‘你祖宗的家在 埃及 法老家 的时候，我不是向他们显现吗？
1SAM|2|28|在 以色列 众支派中，我不是拣选他作我的祭司，上我的祭坛，烧香，在我面前穿以弗得吗？我不是将 以色列 人所献的火祭都赐给你祖宗的家吗？
1SAM|2|29|你们为何践踏我所吩咐献在我居所的祭物和供物呢 ？你为何尊重你的儿子过于尊重我，将我百姓 以色列 所献美好的祭物都拿去养肥你们自己呢？’
1SAM|2|30|因此，耶和华－ 以色列 的上帝说：‘我确实说过，你和你祖宗的家必永远行在我面前，但现在耶和华却说，我绝不会这样做。因为尊重我的，我必尊重他；藐视我的，他必被轻视。
1SAM|2|31|看哪，日子将到，我要折断你的膀臂和你祖宗家的膀臂，使你家中没有一个老年人。
1SAM|2|32|你在 以色列 人享福的时候必看见我居所的衰败 ，你家中必永远没有一个老年人。
1SAM|2|33|你家中的人，我没有从我坛前剪除的，必使你眼睛失明，心中忧伤。你家中所添的人口都必夭折。
1SAM|2|34|你的两个儿子 何弗尼 、 非尼哈 所遭遇的事是给你的预兆：他们二人必在同一日死亡。
1SAM|2|35|我要为自己立一个忠心的祭司，他行事必照我的心、如我的意。我要为他建立坚固的家，他必天天行走在我受膏者的面前。
1SAM|2|36|你家所剩下的人都必来叩拜他，求一块银子，一个饼，说：求你给我一个祭司的职分，好使我得点饼吃。’”
1SAM|3|1|那孩子 撒母耳 在 以利 面前事奉耶和华。在那些日子，耶和华的言语稀少，不常有异象。
1SAM|3|2|那时， 以利 在自己的地方睡觉；他眼目开始昏花，不能看见。
1SAM|3|3|上帝的灯还没有熄灭， 撒母耳 睡在耶和华的殿内，上帝的约柜就在那里。
1SAM|3|4|耶和华呼唤 撒母耳 ， 撒母耳 说：“我在这里！”
1SAM|3|5|他跑到 以利 那里，说：“你叫我吗？我在这里。” 以利 说：“我没有叫你，回去睡吧。”他就回去睡了。
1SAM|3|6|耶和华又呼唤 撒母耳 。 撒母耳 起来，到 以利 那里，说：“你叫我吗？我在这里。” 以利 说：“我儿，我没有叫你，回去睡吧。”
1SAM|3|7|那时 撒母耳 还未认识耶和华，耶和华的话也未曾向他启示。
1SAM|3|8|耶和华第三次再呼唤 撒母耳 。 撒母耳 起来，到 以利 那里，说：“你叫我吗？我在这里。” 以利 才明白是耶和华呼唤这小孩。
1SAM|3|9|以利 对 撒母耳 说：“你回去睡吧。他若再叫你，你就说：‘耶和华啊，请说，仆人敬听！’” 撒母耳 就回去，仍睡在原处。
1SAM|3|10|耶和华来站着，像前几次呼唤：“ 撒母耳 ！ 撒母耳 ！” 撒母耳 说：“请说，仆人敬听！”
1SAM|3|11|耶和华对 撒母耳 说：“看哪，我在 以色列 中必行一件事，凡听见的人都必双耳齐鸣。
1SAM|3|12|我指着 以利 家所说的话，到了时候，必从头到尾应验在 以利 身上。
1SAM|3|13|我曾告诉他，我必永远惩罚他的家，因为他知道自己的儿子作恶，亵渎上帝 ，却不禁止他们。
1SAM|3|14|所以我向 以利 家起誓：‘ 以利 家的罪孽，就是献祭物和供物，也永不得赎。’”
1SAM|3|15|撒母耳 睡到天亮，就开了耶和华殿的门。 撒母耳 害怕，不敢将异象告诉 以利 。
1SAM|3|16|以利 呼唤 撒母耳 说：“我儿 撒母耳 ！” 撒母耳 说：“我在这里！”
1SAM|3|17|以利 说：“他对你说了什么话，你不要向我隐瞒。你若将他对你所说的话向我隐瞒一句，愿上帝重重惩罚你。”
1SAM|3|18|撒母耳 就把一切话都告诉 以利 ，并没有隐瞒。 以利 说：“他是耶和华，愿他照他看为好的去做。”
1SAM|3|19|撒母耳 长大了，耶和华与他同在，使他所说的话一句都不落空。
1SAM|3|20|从 但 到 别是巴 ，所有的 以色列 人都知道耶和华立 撒母耳 为先知。
1SAM|3|21|耶和华又在 示罗 显现，因为耶和华在 示罗 藉他的话向 撒母耳 启示他自己。
1SAM|4|1|撒母耳 的话传遍了全 以色列 。 以色列 人出去与 非利士 人打仗，安营在 以便．以谢 ， 非利士 人安营在 亚弗 。
1SAM|4|2|非利士 人向 以色列 人摆阵。两军交战的时候， 以色列 人败在 非利士 人面前； 非利士 人在战场上杀了他们约四千人。
1SAM|4|3|百姓回到营里， 以色列 的长老说：“耶和华今日为何使我们败在 非利士 人面前呢？我们要将耶和华的约柜从 示罗 抬到我们这里来，好让他来到我们中间，救我们脱离敌人的手掌。”
1SAM|4|4|于是百姓派人到 示罗 ，从那里将坐在二基路伯上万军之耶和华的约柜抬来。 以利 的两个儿子 何弗尼 、 非尼哈 也与上帝的约柜同来。
1SAM|4|5|耶和华的约柜到了营中，全 以色列 就大声欢呼，连地都震动。
1SAM|4|6|非利士 人听见欢呼的声音，就说：“为何 希伯来 人在营里这么大声欢呼呢？”他们知道耶和华的约柜到了营中。
1SAM|4|7|非利士 人就惧怕，说：“有神明到了他们营中。”又说：“我们有祸了！从来不曾有这样的事。
1SAM|4|8|我们有祸了！谁能救我们脱离这些大能之神明的手呢？从前在旷野用各样灾祸击打 埃及 人的，就是这些神明。
1SAM|4|9|非利士 人哪，要刚强，要作大丈夫，免得作 希伯来 人的奴仆，如同他们作你们的奴仆一样。你们要作大丈夫，与他们争战。”
1SAM|4|10|非利士 人进攻， 以色列 人败了，各往自己的家逃跑。被杀的人很多， 以色列 倒下的步兵有三万。
1SAM|4|11|上帝的约柜被掳去， 以利 的两个儿子 何弗尼 、 非尼哈 也都被杀了。
1SAM|4|12|有一个 便雅悯 人从战场上逃跑，衣服撕裂，头蒙灰尘，当日来到 示罗 。
1SAM|4|13|他到了的时候，看哪， 以利 正坐在路旁的位子上观望，为上帝的约柜心里担忧。那人进城报信，全城的人就都呼喊起来。
1SAM|4|14|以利 听见呼喊的声音就说：“这喧嚷的声音是什么呢？”那人急忙来报信给 以利 。
1SAM|4|15|那时 以利 九十八岁了，两眼发直，不能看见。
1SAM|4|16|那人对 以利 说：“我是从战场上来的，今日刚从战场上逃回来。” 以利 说：“我儿，事情怎样了？”
1SAM|4|17|报信的回答说：“ 以色列 人在 非利士 人面前逃跑，百姓中被杀的很多！你的两个儿子 何弗尼 和 非尼哈 也都死了，并且上帝的约柜已经被掳去了。”
1SAM|4|18|他一提到上帝的约柜， 以利 就从城门旁自己的位子上往后跌倒，折断颈项而死，因为他年纪老迈，身体沉重。 以利 作 以色列 的士师四十年。
1SAM|4|19|以利 的媳妇， 非尼哈 的妻子怀孕将到产期，她听见上帝的约柜被掳，公公和丈夫都死了，就曲身生产，极其疼痛。
1SAM|4|20|她将要死的时候，旁边站着的妇人们对她说：“不要怕！你生了男孩了。”她不回答，也不放在心上。
1SAM|4|21|她给孩子起名叫 以迦博 ，说：“荣耀离开 以色列 了！”这是因为上帝的约柜被掳去，又因为她公公和丈夫都死了。
1SAM|4|22|她又说：“荣耀离开 以色列 ，因为上帝的约柜被掳去了。”
1SAM|5|1|非利士 人掳去上帝的约柜，从 以便．以谢 带到 亚实突 。
1SAM|5|2|非利士 人掳了上帝的约柜，带进 大衮 庙，放在 大衮 的旁边。
1SAM|5|3|次日， 亚实突 人清早起来，看哪， 大衮 仆倒在耶和华的约柜前，脸伏于地，他们就扶起 大衮 ，把它放回原处。
1SAM|5|4|又次日，他们清早起来，看哪， 大衮 仆倒在耶和华的约柜前，脸伏于地，并且 大衮 的头和两手都在门槛上折断，只剩下 大衮 的躯干。
1SAM|5|5|因此， 大衮 的祭司和所有进 大衮 庙的人，都不踏 亚实突 的 大衮 庙的门槛，直到今日。
1SAM|5|6|耶和华的手重重击打 亚实突 人，使他们恐惧，使 亚实突 和 亚实突 周围的人都生痔疮。
1SAM|5|7|亚实突 人见这情况，就说：“ 以色列 上帝的约柜不可留在我们这里，因为他的手重重击打我们和我们的神明 大衮 ”。
1SAM|5|8|他们就派人去请 非利士 的众领袖来聚集，对他们说：“我们向 以色列 上帝的约柜应当怎样做呢？”他们说：“可以把 以色列 上帝的约柜运到 迦特 去。”于是他们把 以色列 上帝的约柜运到那里。
1SAM|5|9|运到之后，耶和华的手击打那城，使那城的人非常惊慌，无论大小都生痔疮。
1SAM|5|10|他们就把上帝的约柜送到 以革伦 。上帝的约柜到了 以革伦 ， 以革伦 人就呼喊说：“他们把 以色列 上帝的约柜运到我这里，要害我和我的百姓！”
1SAM|5|11|于是他们派人去请 非利士 的众领袖来，说：“请你们把 以色列 上帝的约柜送回原处，免得害死我和我的百姓！”原来上帝的手重重攻击那城，死亡的恐惧弥漫全城，
1SAM|5|12|没有死的人都受痔疮的折磨。城里的哀声上达于天。
1SAM|6|1|耶和华的约柜在 非利士 人之地七个月。
1SAM|6|2|非利士 人召了祭司和占卜的来，说：“我们向耶和华的约柜应当怎样做呢？请指示我们要用什么方法把约柜送回原处。”
1SAM|6|3|他们说：“若要将 以色列 上帝的约柜送回去，不可空手送回，一定要给他献赔罪的礼物，然后你们才可以得痊愈，并且知道他的手为何不离开你们。”
1SAM|6|4|非利士 人说：“应当用什么献为赔罪的礼物呢？”他们说：“当按照 非利士 领袖的数目，献五个金痔疮和五个金老鼠，因为你们众人和领袖所遭遇的都是一样的灾祸。
1SAM|6|5|当制造你们痔疮的像和毁坏田地老鼠的像，并要将荣耀归给 以色列 的上帝，或者他向你们和你们的神明，以及你们的田地，把手放轻些。
1SAM|6|6|你们为何硬着心，像 埃及 人和法老硬着心一样呢？上帝岂不是严厉对付 埃及 ，使 埃及 人释放 以色列 人，他们就走了吗？
1SAM|6|7|现在你们应当造一辆新车，把两头未曾负轭，还在哺乳的母牛套在车上，赶牛犊离开母牛，回家去。
1SAM|6|8|你们要把耶和华的约柜放在车上，把所献赔罪的金器装在匣子里，放在柜旁，送走柜子，让它去。
1SAM|6|9|你们要观察：车若直行过 以色列 的边界，上到 伯．示麦 去，这大灾祸就是耶和华降在我们身上的；若不然，我们就知道，这不是他的手击打我们，而是我们偶然遭遇的。”
1SAM|6|10|非利士 人就照样做了。他们取了两头哺乳的母牛套在车上，把牛犊关在家里，
1SAM|6|11|把耶和华的约柜和装金老鼠以及金痔疮像的匣子都放在车上。
1SAM|6|12|牛直行大路，在往 伯．示麦 的一条大道上，一面走一面叫，不偏左右。 非利士 的领袖跟在后面，直到 伯．示麦 的地界。
1SAM|6|13|那时， 伯．示麦 人正在平原收割麦子，举目看见约柜，就欢欢喜喜地迎见它。
1SAM|6|14|车到了 伯．示麦 人 约书亚 的田间，就在那里停了。在那里有一块大磐石，他们把车的木头劈了，把两头母牛献给耶和华为燔祭。
1SAM|6|15|利未 人将耶和华的约柜和柜子旁边装金器的匣子拿下来，放在大磐石上。当日 伯．示麦 人献上燔祭，又献其他祭物给耶和华。
1SAM|6|16|非利士 人的五个领袖看见了，当日就回 以革伦 去。
1SAM|6|17|非利士 人献给耶和华作赔罪的金痔疮像如下：一个为 亚实突 ，一个为 迦萨 ，一个为 亚实基伦 ，一个为 迦特 ，一个为 以革伦 。
1SAM|6|18|金老鼠的数目是按照 非利士 五个领袖的城镇，就是坚固的城镇和乡村，以及大磐石。这磐石是安放耶和华约柜的，到今日还在 伯．示麦 人 约书亚 的田间。
1SAM|6|19|耶和华击杀 伯．示麦 人，因为他们观看他的约柜。他击杀了百姓七十人 。百姓因耶和华大大击杀他们，就哀哭了。
1SAM|6|20|伯．示麦 人说：“谁能在耶和华这位圣洁的上帝面前侍立呢？这约柜可以从我们这里上到谁那里去呢？”
1SAM|6|21|于是他们派使者到 基列．耶琳 的居民那里，说：“ 非利士 人将耶和华的约柜送回来了，你们下来将约柜接了，上到你们那里去吧！”
1SAM|7|1|基列．耶琳 人就来了，将耶和华的约柜接上去，抬到山上 亚比拿达 的家中，将他儿子 以利亚撒 分别为圣，看守耶和华的约柜。
1SAM|7|2|从约柜留在 基列．耶琳 的那天起，经过了许多日子，有二十年； 以色列 全家都哀哭归向耶和华。
1SAM|7|3|撒母耳 对 以色列 全家说：“你们若全心回转归向耶和华，就要从你们中间除掉外邦的神明和 亚斯她录 ，预备你们的心归向耶和华，单单事奉他，他必救你们脱离 非利士 人的手。”
1SAM|7|4|以色列 人就除掉诸 巴力 和 亚斯她录 ，单单事奉耶和华。
1SAM|7|5|撒母耳 说：“要召集 以色列 众人到 米斯巴 去，我好为你们向耶和华祷告。”
1SAM|7|6|他们就聚集在 米斯巴 ，打水浇在耶和华面前。当日他们禁食，说：“我们得罪了耶和华。” 撒母耳 在 米斯巴 作 以色列 人的士师。
1SAM|7|7|非利士 人听见 以色列 人聚集在 米斯巴 ， 非利士 的领袖就上来要攻击 以色列 。 以色列 人听见，就惧怕 非利士 人。
1SAM|7|8|以色列 人对 撒母耳 说：“愿你不住为我们呼求耶和华－我们的上帝，救我们脱离 非利士 人的手。”
1SAM|7|9|撒母耳 就把一只吃奶的羔羊献给耶和华作全牲的燔祭，为 以色列 人呼求耶和华，耶和华就应允他。
1SAM|7|10|撒母耳 正献燔祭的时候， 非利士 人前来要与 以色列 争战。当日，耶和华打雷，发出极大的声音，使 非利士 人溃乱，他们就败在 以色列 面前。
1SAM|7|11|以色列 人从 米斯巴 出来，追赶 非利士 人，击杀他们，直到 伯．甲 的下边。
1SAM|7|12|撒母耳 拿一块石头立在 米斯巴 和 善 的中间，给石头起名叫 以便．以谢 ，说：“到如今耶和华都帮助我们。”
1SAM|7|13|因此， 非利士 人被制伏了，不再入侵 以色列 境内。 撒母耳 有生之年，耶和华的手攻击 非利士 人。
1SAM|7|14|非利士 人所夺取 以色列 的城镇，从 以革伦 直到 迦特 ，都归回 以色列 了。 以色列 也从 非利士 人手中收回这些城所属的地界。那时 以色列 与 亚摩利 人和平相处。
1SAM|7|15|撒母耳 一生作 以色列 的士师。
1SAM|7|16|他每年巡行到 伯特利 、 吉甲 、 米斯巴 ，在这些地方审判 以色列 人。
1SAM|7|17|随后他回到 拉玛 ，因为他的家在那里；他在那里审判 以色列 人，并且在那里为耶和华筑了一座坛。
1SAM|8|1|撒母耳 年纪老迈，就立他的儿子作 以色列 的士师。
1SAM|8|2|他的长子名叫 约珥 ，次子名叫 亚比亚 ；他们在 别是巴 作士师。
1SAM|8|3|他的儿子不行他的道，贪图财利，收取贿赂，屈枉正直。
1SAM|8|4|以色列 的长老都聚集在 拉玛 ，来到 撒母耳 那里，
1SAM|8|5|对他说：“看哪，你年纪老了，你的儿子又不行你的道。现在请你为我们立一个王治理我们，像列国一样。”
1SAM|8|6|撒母耳 不喜悦他们说“立一个王治理我们”，他就向耶和华祷告。
1SAM|8|7|耶和华对 撒母耳 说：“你只管听从百姓向你说的一切话，因为他们不是厌弃你，而是厌弃我，不要我作他们的王。
1SAM|8|8|自从我领他们出 埃及 的日子到如今，他们离弃我，事奉别神；正像他们从前所做的一切事，现在他们也照样向你做了。
1SAM|8|9|现在你只管听从他们的话，不过要严厉警告他们，告诉他们将来王会用什么方式管辖他们。”
1SAM|8|10|撒母耳 将耶和华一切的话转告求他立王的百姓。
1SAM|8|11|他说：“管辖你们的王必用这样的方式：他必派你们的儿子为他驾车，赶马，在他的战车前奔跑。
1SAM|8|12|他要为自己立千夫长、五十夫长；耕种他的田地，收割他的庄稼；打造他的兵器和车上的器械。
1SAM|8|13|他必叫你们的女儿为他制造香膏，作厨师与烤饼的，
1SAM|8|14|也必取你们最好的田地、葡萄园、橄榄园，赐给他的臣仆。
1SAM|8|15|你们的粮食和葡萄园所出产的，他必征收十分之一给他的官员和臣仆，
1SAM|8|16|又必叫你们的仆人婢女，健壮的青年和你们的驴为他做工。
1SAM|8|17|你们的羊群，他必征收十分之一，你们自己也必作他的仆人。
1SAM|8|18|那日，你们必因自己所选的王哀求耶和华，但那日耶和华却不应允你们。”
1SAM|8|19|百姓却不肯听 撒母耳 的话，说：“不！我们一定要一个王治理我们，
1SAM|8|20|使我们像列国一样，有王治理我们，率领我们，为我们争战。”
1SAM|8|21|撒母耳 听见百姓这一切话，就禀告给耶和华听。
1SAM|8|22|耶和华对 撒母耳 说：“你只管听从他们的话，为他们立一个王。” 撒母耳 对 以色列 人说：“去，你们各归各城吧！”
1SAM|9|1|有一个 便雅悯 人名叫 基士 ，是 便雅悯 人 亚斐亚 的玄孙， 比歌拉 的曾孙， 洗罗 的孙子， 亚别 的儿子，是个大能的勇士 。
1SAM|9|2|他有一个儿子名叫 扫罗 ，又健壮、又英俊，在 以色列 人中没有一个可以与他相比；他比众百姓高出一个头 。
1SAM|9|3|扫罗 的父亲 基士 丢失了几匹母驴，他就吩咐儿子 扫罗 说：“起来，带一个仆人去寻找驴子。”
1SAM|9|4|扫罗 走过 以法莲 山区，又过 沙利沙 地，都没有找着。他们走过 沙琳 地，驴不在那里，又走过 便雅悯 地，也没有找到。
1SAM|9|5|到了 苏弗 地， 扫罗 对跟随他的仆人说：“我们不如回去，免得我父亲不为驴挂虑，反为我们担忧。”
1SAM|9|6|仆人对他说：“看哪，这城里有一位神人，受人敬重，凡他所说的全都应验。现在让我们到他那里去，或者他能指示我们当走的路。”
1SAM|9|7|扫罗 对仆人说：“看哪，我们若去，送什么给那人呢？我们袋子里的食物都吃完了，也没有礼物可以送给神人，我们还有些什么呢？”
1SAM|9|8|仆人又回答 扫罗 说：“看哪，我手里还有四分之一舍客勒的银子，可以送给神人，请他指示我们当走的路。”
1SAM|9|9|从前 以色列 中，若有人去求问上帝，就这么说：“来，我们到先见那里去吧！”因现在的先知，从前称为先见。
1SAM|9|10|扫罗 对仆人说：“好主意！来，我们去吧。”于是他们往神人所住的城里去了。
1SAM|9|11|他们上坡要进城，遇见几个少女出来打水，就问她们说：“先见有没有在这里呢？”
1SAM|9|12|她们回答说：“有的，看哪，他就在你们前面。快！他今日正来到城里，因为今日百姓要在丘坛献祭。
1SAM|9|13|你们一进城，他还没有上丘坛吃祭物之前，就会遇见他。因为他没有到，百姓不能吃，必须等他先为祭物祝谢，然后受邀的人才可以吃。现在就上去吧，因为这时候你们会遇见他。”
1SAM|9|14|他们就上到那城，进入城中的时候，看哪， 撒母耳 正迎着他们来，要上丘坛去。
1SAM|9|15|扫罗 还没有到的前一日，耶和华已经对 撒母耳 启示说：
1SAM|9|16|“明日这时候，我必使一个人从 便雅悯 地到你这里来，你要膏他作我百姓 以色列 的君王。他必救我的百姓脱离 非利士 人的手，因为我眷顾我的百姓 ，他们的哀声已上达于我。”
1SAM|9|17|撒母耳 看见 扫罗 的时候，耶和华对他说：“看哪，这就是我对你所说的人，他必治理我的百姓。”
1SAM|9|18|扫罗 在城门中走到 撒母耳 跟前，说：“请告诉我，先见的家在哪里？”
1SAM|9|19|撒母耳 回答扫罗说：“我就是先见。你在我前面先上丘坛去，因为你们今日必跟我同席。明日早晨我送你走，会把你心里一切的事都告诉你。
1SAM|9|20|至于你前三日所丢失的几匹母驴，你心里不必挂虑，都已经找到了。 以色列 众人所仰慕的是谁呢？不是仰慕你和你父的全家吗？”
1SAM|9|21|扫罗 回答说：“我不是 以色列 支派中最小的 便雅悯 人吗？我的家族不是 便雅悯 支派中最小的家族吗？你为何对我说这样的话呢？”
1SAM|9|22|撒母耳 领 扫罗 和他的仆人进了大厅，使他们在受邀的人中坐首位；受邀者约有三十个。
1SAM|9|23|撒母耳 对厨师说：“我交给你的那一份祭肉，吩咐你收存的，现在可以拿来。”
1SAM|9|24|厨师就举起祭肉的腿和腿上的部分 ，摆在 扫罗 面前。 撒母耳 说：“看哪，所存留的摆在你面前了。吃吧！因为这是为你保留到这特定的时候的，好让你说，是我请了这百姓来，” 当日， 扫罗 就与 撒母耳 同席。
1SAM|9|25|他们从丘坛下来进城， 撒母耳 和 扫罗 在房顶上说话。
1SAM|9|26|次日他们清早起来。黎明的时候， 撒母耳 呼叫在房顶上的 扫罗 ，说：“起来，我好送你回去。” 扫罗 就起来，和 撒母耳 二人一同到外面去。
1SAM|9|27|二人下到城边， 撒母耳 对 扫罗 说：“你要吩咐仆人先走，仆人走了以后， 你要留在这里，这时候我要将上帝的话传给你听。”
1SAM|10|1|撒母耳 拿一瓶膏油倒在 扫罗 的头上，亲吻他，说：“耶和华岂不是膏你作他产业的君王吗？
1SAM|10|2|你今日离开我之后，会在 便雅悯 境内的 谢撒 ，靠近 拉结 的坟墓，遇见两个人。他们会对你说：‘你要找的几匹母驴已经找到了。看哪，你父亲不为驴子的事挂虑，反为你担忧，说：我为儿子该做些什么呢？’
1SAM|10|3|你从那里往前走，到了 他泊 的橡树那里，会遇见三个往 伯特利 去敬拜上帝的人：一个带着三只小山羊，一个带着三个饼，一个带着一皮袋酒。
1SAM|10|4|他们会向你问安，给你两个饼，你就从他们手中接过来。
1SAM|10|5|然后你要到上帝的山去，在那里有 非利士 的驻军。你到了城里的时候，会遇见一队先知从丘坛下来，前面有鼓瑟的、击鼓的、吹笛的、弹琴的，他们都受感说话。
1SAM|10|6|耶和华的灵必大大感动你，你就与他们一同受感说话，转变成另一个人。
1SAM|10|7|这征兆临到你，你就要趁机做该做的事，因为上帝与你同在。
1SAM|10|8|你要在我以先下到 吉甲 。看哪，我必下到你那里献燔祭和平安祭。你要等候七日，等我到你那里指示你当做的事。”
1SAM|10|9|扫罗 转身离开 撒母耳 ，上帝就改变他，赐给他另一颗心。当日这一切征兆都应验了。
1SAM|10|10|他们来到那座山，看哪，有一队先知遇见 扫罗 。上帝的灵大大感动他，他就在先知中受感说话。
1SAM|10|11|所有先前认识 扫罗 的人看见了，看哪，他和先知一同受感说话，百姓就彼此说：“ 基士 的儿子遇见了什么呢？ 扫罗 也在先知中吗？”
1SAM|10|12|那地方有一个人说：“这些人的父亲是谁呢？”因此就有一句俗语说：“ 扫罗 也在先知中吗？”
1SAM|10|13|扫罗 受感说完了话，就上丘坛去了。
1SAM|10|14|扫罗 的叔叔问 扫罗 和他的仆人说：“你们到哪里去了？”他说：“我们找驴子去了。但我们找不到，就去了 撒母耳 那里。”
1SAM|10|15|扫罗 的叔叔说：“告诉我 撒母耳 对你们说了些什么。”
1SAM|10|16|扫罗 对他的叔叔说：“他明明告诉我们，驴子已经找到了。”至于 撒母耳 所说君王的事， 扫罗 没有告诉叔叔。
1SAM|10|17|撒母耳 召集百姓到 米斯巴 耶和华那里。
1SAM|10|18|他对 以色列 众人说：“耶和华－ 以色列 的上帝如此说：‘我领 以色列 出 埃及 ，救你们脱离 埃及 人的手，以及脱离欺压你们各国之人的手。’
1SAM|10|19|你们今日却厌弃救你们脱离一切灾祸和患难的上帝，对他说：‘求你立一个王治理我们。’现在你们应当按支派和宗族站在耶和华面前。”
1SAM|10|20|于是， 撒母耳 叫 以色列 众支派近前来抽签，抽到了 便雅悯 支派。
1SAM|10|21|然后，他叫 便雅悯 支派按宗族近前来，抽到了 玛特利 族，接着又抽到了 基士 的儿子 扫罗 。众人寻找他却找不到，
1SAM|10|22|就再问耶和华说：“那人来到这里了没有？”耶和华说：“看哪，他藏在物品堆中。”
1SAM|10|23|众人就跑去从那里领他出来。他站在百姓中间，比众百姓高出一个头。
1SAM|10|24|撒母耳 对众百姓说：“你们看到了耶和华所拣选的人吗？众百姓中没有人可以与他相比。”众百姓就欢呼说：“愿王万岁！”
1SAM|10|25|撒母耳 将君王的典章对百姓说明，又记在书上，放在耶和华面前，然后 撒母耳 遣散众百姓，各回自己的家去了。
1SAM|10|26|扫罗 也往 基比亚 自己的家去，有一群心中被上帝感动的勇士跟随他。
1SAM|10|27|但有些无赖之辈说：“这人怎么能救我们呢？”他们就藐视他，不送礼物给他。 扫罗 却保持沉默。
1SAM|11|1|亚扪 人 拿辖 上来，对着 基列 的 雅比 安营。 雅比 众人对 拿辖 说：“你与我们立约，我们就服事你。”
1SAM|11|2|亚扪 人 拿辖 对他们说：“你们若由我挖出你们各人的右眼，以此凌辱 以色列 众人，我就与你们立约。”
1SAM|11|3|雅比 的长老对他说：“求你宽容我们七日，等我们派人到 以色列 的全境去。若没有人来救我们，我们就出来归顺你。”
1SAM|11|4|使者到了 扫罗 住的 基比亚 ，把这事说给百姓听，众百姓就都放声大哭。
1SAM|11|5|看哪， 扫罗 正从田间赶牛回来，说：“百姓为什么哭呢？”众人把 雅比 人的话告诉他。
1SAM|11|6|扫罗 听见这些话，就被上帝的灵催逼，大发怒气。
1SAM|11|7|他把一对牛切成小块，吩咐使者传送到 以色列 全境，说：“凡不出来跟随 扫罗 和 撒母耳 的，就必这样待他的牛。”耶和华使百姓惧怕，他们就都出来如同一人。
1SAM|11|8|扫罗 在 比色 数点他们： 以色列 人有三十万， 犹大 人有三万。
1SAM|11|9|他们对那些来的使者说：“你们要对 基列 的 雅比 人这样说，明天太阳快到中午的时候，你们必得解救。”使者回去告诉 雅比 人，他们就欢喜了。
1SAM|11|10|于是 雅比 人对 亚扪 人说：“明日我们出来归顺你们，可以照你们看为好的待我们。”
1SAM|11|11|第二日， 扫罗 把百姓分为三队，在清晨换岗哨的时候入侵 亚扪 人的军营，击杀他们直到中午的时候。逃脱的人都分散了，甚至没有两个人同在一起。
1SAM|11|12|百姓对 撒母耳 说：“那说‘ 扫罗 岂能作我们的王’的是谁呢？把他们交出来，我们好处死他们。”
1SAM|11|13|扫罗 说：“今日耶和华在 以色列 中施行拯救，所以今日不可处死人。”
1SAM|11|14|撒母耳 对百姓说：“来，我们到 吉甲 去，在那里开始新的王国。”
1SAM|11|15|众百姓到了 吉甲 那里，在耶和华面前拥立 扫罗 为王，又在耶和华面前献平安祭。 扫罗 和 以色列 众人在那里都非常欢喜。
1SAM|12|1|撒母耳 对 以色列 众人说：“看哪，我已听了你们对我所说一切的话，为你们立了一个王。
1SAM|12|2|现在，看哪，有这王行走在你们前面。我已年老发白，看哪，我的儿子都在你们这里。我从幼年直到今日都行走在你们前面。
1SAM|12|3|我在这里，你们要在耶和华和他的受膏者面前为我作证，我夺过谁的牛，抢过谁的驴，欺负过谁，虐待过谁，从谁手里收过贿赂而蒙蔽自己的眼目呢？若有，我必偿还。”
1SAM|12|4|众人说：“你未曾欺负我们，虐待我们，也未曾从任何人手里收过任何东西。”
1SAM|12|5|撒母耳 对他们说：“你们在我手里没有找着什么，有耶和华在你们中间作证，也有他的受膏者今日作证。”他们说 ：“愿耶和华作证。”
1SAM|12|6|撒母耳 对百姓说：“从前立 摩西 和 亚伦 ，又领你们祖先出 埃及 地的是耶和华。
1SAM|12|7|现在你们要站住，让我在耶和华面前，以耶和华向你们和你们祖先所行一切公义的事来和你们争辩。
1SAM|12|8|从前 雅各 到了 埃及 ，后来你们的祖先呼求耶和华，耶和华就差遣 摩西 和 亚伦 领你们的祖先出 埃及 ，来到这地方居住。
1SAM|12|9|他们却忘记耶和华－他们的上帝，他就把他们交给 夏琐 将军 西西拉 的手中，以及 非利士 人和 摩押 王的手中 。于是这些人常来攻击他们。
1SAM|12|10|他们呼求耶和华说：‘我们离弃了耶和华去事奉诸 巴力 和 亚斯她录 ，我们有罪了。现在求你救我们脱离仇敌的手，我们必事奉你。’
1SAM|12|11|耶和华就差遣 耶路巴力 、 比但 、 耶弗他 、 撒母耳 救你们脱离四围仇敌的手，你们才安然居住。
1SAM|12|12|你们见 亚扪 人的王 拿辖 来攻击你们，就对我说：‘不，要有一个王治理我们。’其实耶和华－你们的上帝是你们的王。
1SAM|12|13|现在，看哪，这就是你们所选的、你们所求的王。看哪，耶和华已经为你们立王了。
1SAM|12|14|你们若敬畏耶和华，事奉他，听从他的话，不违背耶和华的命令，你们和治理你们的王也都跟从耶和华－你们的上帝就好了。
1SAM|12|15|倘若不听从耶和华的话，违背他的命令，耶和华的手必攻击你们，像从前攻击你们祖先一样。
1SAM|12|16|现在你们要站住，看耶和华在你们眼前要行的一件大事。
1SAM|12|17|这不是割麦子的时候吗？我求告耶和华，他必打雷降雨，让你们知道并且看出，你们为自己求立王的事在耶和华眼前是犯大罪了。”
1SAM|12|18|于是 撒母耳 求告耶和华，耶和华就在这日打雷降雨，众百姓就非常惧怕耶和华和 撒母耳 。
1SAM|12|19|众百姓对 撒母耳 说：“请你为仆人向耶和华－你的上帝祷告，免得我们死亡，因为我们求立王的事，正是罪上加罪了。”
1SAM|12|20|撒母耳 对百姓说：“不要惧怕！你们虽然行了这恶，却不要偏离耶和华，只要尽心事奉他。
1SAM|12|21|不可偏离去随从那没有益处、不能救人的虚无的神明 ，因为它们是虚无的。
1SAM|12|22|耶和华必因他大名的缘故不撇弃他的子民，因为耶和华喜悦你们作他的子民。
1SAM|12|23|至于我，我如果停止为你们祷告，就得罪耶和华了，我绝不会这样做。我必以善道正路指教你们。
1SAM|12|24|但你们要敬畏耶和华，诚诚实实地尽心事奉他，因你们要留意，他向你们所行的事何等大。
1SAM|12|25|你们若不断作恶，你们和你们的王必一同灭亡。”
1SAM|13|1|扫罗 登基的时候年三十 岁，作 以色列 王二年 。
1SAM|13|2|扫罗 从 以色列 中选出三千人：二千跟随 扫罗 在 密抹 和 伯特利 山区，一千跟随 约拿单 在 便雅悯 的 基比亚 。其余的百姓， 扫罗 打发他们各自回自己的帐棚去了。
1SAM|13|3|约拿单 攻击 非利士 人在 迦巴 的驻军， 非利士 人听见了这事。 扫罗 就在遍地吹角，说：“让 希伯来 人都听见。”
1SAM|13|4|以色列 众人听见 扫罗 攻击 非利士 的驻军，又听见 以色列 为 非利士 人所憎恶，百姓就跟随 扫罗 ，在 吉甲 集合。
1SAM|13|5|非利士 人集合，要与 以色列 人作战。他们有战车三万辆，骑兵六千，士兵像海边的沙那样多。他们上来，在 伯．亚文 东边的 密抹 安营。
1SAM|13|6|以色列 人见自己危急，军队被围攻，百姓就藏在山洞、丛林、岩隙、地窖和深坑中。
1SAM|13|7|有些 希伯来 人过了 约旦河 ，逃到 迦得 和 基列 地。 扫罗 还在 吉甲 ，所有的人都战战兢兢地跟随他。
1SAM|13|8|扫罗 照着 撒母耳 所定的日期等了七日。但是， 撒母耳 还没有来到 吉甲 ，百姓就离开 扫罗 散去了。
1SAM|13|9|于是 扫罗 说：“把燔祭和平安祭带到我这里来。” 扫罗 就献上燔祭。
1SAM|13|10|他刚献完燔祭，看哪， 撒母耳 就到了。 扫罗 出去迎接他，向他问安。
1SAM|13|11|撒母耳 说：“你做了什么事啊？” 扫罗 说：“因为我见百姓离开我散去，你又不照所定的日期来到，而且 非利士 人已在 密抹 集合；
1SAM|13|12|我说：‘现在 非利士 人已经下到 吉甲 来攻击我，可是我还没有向耶和华祷告。’所以我就勉强献上燔祭。”
1SAM|13|13|撒母耳 对 扫罗 说：“你做了糊涂事了，没有遵守耶和华－你上帝吩咐你的命令。不然，耶和华会在 以色列 中坚立你的国度，直到永远。
1SAM|13|14|现在你的国度必不长久。耶和华已经寻着一个合他心意的人，立他作百姓的君王，因为你没有遵守耶和华所吩咐你的。”
1SAM|13|15|撒母耳 就起来，从 吉甲 上到 便雅悯 的 基比亚 。 扫罗 数点跟随他的百姓，约有六百人。
1SAM|13|16|扫罗 和他儿子 约拿单 ，以及跟随他们的百姓，都住在 便雅悯 的 迦巴 ， 非利士 人却在 密抹 安营。
1SAM|13|17|有突击队从 非利士 营中出来，分成三队：一队往 俄弗拉 到 书亚 地去，
1SAM|13|18|一队往 伯．和仑 去，一队往边界，下望朝着旷野的 洗波音谷 。
1SAM|13|19|那时， 以色列 全地找不到一个铁匠，因为 非利士 人说：“恐怕 希伯来 人制造刀枪。”
1SAM|13|20|以色列 众人要磨锄、犁、斧、铲，就各自下到 非利士 人那里去磨。
1SAM|13|21|磨锄或犁的价钱是三分之二舍客勒，磨斧或修整刺棒的价钱是三分之一舍客勒。
1SAM|13|22|所以到了战争的日子，所有跟随 扫罗 和 约拿单 的百姓找不到一个手里有刀有枪的，惟 扫罗 和他儿子 约拿单 有。
1SAM|13|23|非利士 人的一队驻军出来，到 密抹 的隘口。
1SAM|14|1|有一日， 扫罗 的儿子 约拿单 对拿他兵器的青年说：“来，我们过去到 非利士 的驻军那里。”但他没有告诉父亲。
1SAM|14|2|扫罗 在 基比亚 的郊外，坐在 米矶仑 的石榴树下，跟随他的百姓约有六百人。
1SAM|14|3|在那里有 亚希突 的儿子 亚希亚 ，穿着以弗得。 亚希突 是 以迦博 的哥哥， 非尼哈 的儿子， 以利 的孙子。 以利 从前在 示罗 作耶和华的祭司。 约拿单 去了，百姓却不知道。
1SAM|14|4|约拿单 要从隘口过到 非利士 驻军那里去。这隘口两边各有一座齿状峭壁：一座名叫 播薛 ，另一座名叫 西尼 ；
1SAM|14|5|一座向北，对着 密抹 ，一座向南，对着 迦巴 。
1SAM|14|6|约拿单 对拿兵器的青年说：“来，我们过去到那些未受割礼之人的驻军那里，或者耶和华为我们施展能力，因为耶和华使人得胜，不在乎人多人少 。”
1SAM|14|7|拿兵器的对他说：“随你的心意做吧。你上去，看哪，我一定跟随你，与你同心。”
1SAM|14|8|约拿单 说：“看哪，我们要过去到那些人那里，在他们那里展现我们自己。
1SAM|14|9|他们若对我们这么说：‘站住，等我们到你们那里去’，我们就站在原地，不上他们那里去；
1SAM|14|10|但他们若这么说：‘上到我们这里来吧’，我们就上去，因为耶和华把他们交在我们手里了。这就是我们的凭据。”
1SAM|14|11|二人就让 非利士 的驻军看见。 非利士 人说：“看哪， 希伯来 人从躲藏的洞穴里出来了！”
1SAM|14|12|站岗的士兵对 约拿单 和拿兵器的人说：“上到这里来，我们有一件事要告诉你们。” 约拿单 就对拿兵器的人说：“跟我上去，因为耶和华把他们交在 以色列 人手里了。”
1SAM|14|13|约拿单 手脚并用爬上去，拿兵器的人跟随他。 非利士 人仆倒在 约拿单 面前，拿兵器的人跟着他，杀死他们。
1SAM|14|14|约拿单 和拿兵器的人第一次击杀的约有二十人，都在一亩 地的半犁沟之内。
1SAM|14|15|于是在军营、在田野、在众百姓中，人心惶惶，驻军和突击队都战兢；地也震动，这是从上帝那里来的惊恐 。
1SAM|14|16|在 便雅悯 的 基比亚 ， 扫罗 的哨兵观看，看哪， 非利士 全军溃乱，四处乱窜。
1SAM|14|17|扫罗 就对跟随他的百姓说：“你们去数点人数，看是谁从我们这里出去。”他们一数点，看哪， 约拿单 和拿兵器的人不在其中。
1SAM|14|18|那时上帝的约柜 在 以色列 人那里。 扫罗 对 亚希亚 说：“你把上帝的约柜请到这里来。”
1SAM|14|19|扫罗 正与祭司说话的时候， 非利士 营中的骚乱越来越剧烈； 扫罗 就对祭司说：“停手吧！”
1SAM|14|20|扫罗 和所有跟随他的百姓都集合，来到战场，看哪， 非利士 人用刀互相击杀，大大混乱。
1SAM|14|21|那先前由四方来跟随 非利士 人、在他们营中的 希伯来 人，现在也转过来帮助跟随 扫罗 和 约拿单 的 以色列 人了。
1SAM|14|22|那藏在 以法莲 山区的 以色列 众人听说 非利士 人逃跑，就出来紧紧地追击他们。
1SAM|14|23|那日，耶和华使 以色列 人得胜，战争一直打到 伯．亚文 。
1SAM|14|24|那日， 以色列 人非常困惫，因为 扫罗 叫百姓起誓说：“凡不等到晚上我向敌人报完了仇就吃东西的，必受诅咒。”因此所有的百姓都没有尝食物。
1SAM|14|25|所有的百姓 进入树林，见地面上有蜜。
1SAM|14|26|百姓进了树林，看哪，有蜜流出来，却没有人敢用手取蜜入口，因为百姓怕那誓言。
1SAM|14|27|约拿单 没有听见他父亲叫百姓起誓，所以他伸出手中的杖，以杖头蘸在蜂房里，用手取回送入口内，他的眼睛就明亮了。
1SAM|14|28|百姓中有一人对他说：“你父亲曾叫百姓严严地起誓说，今日吃东西的人必受诅咒；因此百姓就疲乏了。”
1SAM|14|29|约拿单 说：“我父亲给这地添麻烦了。你们看，我尝了这一点蜜，眼睛就明亮了。
1SAM|14|30|今日百姓若随意吃了从仇敌夺来的东西，现在击杀的 非利士 人岂不更多吗？”
1SAM|14|31|这日， 以色列 人击杀 非利士 人，从 密抹 直到 亚雅仑 。但百姓非常疲乏，
1SAM|14|32|就急着扑向掠物，夺取牛羊和牛犊，宰于地上，连肉带血吃了。
1SAM|14|33|有人告诉 扫罗 说：“看哪，百姓吃带血的肉，得罪耶和华了。” 扫罗 说：“你们行了诡诈，今日把一块大石头滚到我这里来吧。”
1SAM|14|34|扫罗 又说：“你们分散到百姓中，对他们说，你们各人把牛羊牵到我这里来宰了吃，不可吃带血的肉得罪耶和华。”那夜，所有的百姓把自己手中的牛 牵到那里宰了。
1SAM|14|35|扫罗 为耶和华筑了一座坛，这是他开始为耶和华筑的坛。
1SAM|14|36|扫罗 说：“我们要在夜里下去追赶 非利士 人，抢掠他们，直到天亮，不给他们留下一人。”众百姓说：“你看怎样好就做吧！”祭司说：“我们要先在这里亲近上帝。”
1SAM|14|37|扫罗 求问上帝说：“我可以下去追赶 非利士 人吗？你把他们交在 以色列 人手里吗？”这日上帝没有回答他。
1SAM|14|38|扫罗 说：“百姓中的众领袖，你们都要近前来到这里，查明今日这罪是怎样发生的。
1SAM|14|39|我指着拯救 以色列 的永生的耶和华起誓，就是我儿子 约拿单 犯了罪，他也必被处死。”但众百姓中无人回答他。
1SAM|14|40|扫罗 对 以色列 众人说：“你们站在一边，我与我儿子 约拿单 也站在一边。”百姓对 扫罗 说：“你看怎样好就做吧！”
1SAM|14|41|扫罗 向耶和华－ 以色列 的上帝祷告说：“求你指示正确的答案。”抽中的是 扫罗 和 约拿单 ，百姓尽都无事。
1SAM|14|42|扫罗 说：“你们再抽签，看是我，还是我儿子 约拿单 。”抽中的是 约拿单 。
1SAM|14|43|扫罗 对 约拿单 说：“你告诉我，你做了什么事？” 约拿单 说：“我只是用手中的杖，以杖头蘸了一点蜜尝尝，看哪，我就要死吗？”
1SAM|14|44|扫罗 说：“ 约拿单 哪，你一定要死！若不然，愿上帝重重惩罚我。”
1SAM|14|45|百姓对 扫罗 说：“ 约拿单 在 以色列 中大行拯救，岂可死呢？绝对不可！我们指着永生的耶和华起誓，连他的一根头发也不可落地，因为他今日与上帝一同做事。”于是百姓救 约拿单 免了死亡。
1SAM|14|46|扫罗 上去，不追赶 非利士 人， 非利士 人也回本地去了。
1SAM|14|47|扫罗 执掌 以色列 的国权，攻打他四围所有的仇敌，就是 摩押 人、 亚扪 人、 以东 人和 琐巴 诸王，以及 非利士 人。他无论往何处去，都打败他们。
1SAM|14|48|扫罗 奋勇作战，击败 亚玛力 人，救了 以色列 脱离抢掠他们之人的手。
1SAM|14|49|扫罗 的儿子是 约拿单 、 亦施韦 、 麦基．舒亚 。他的两个女儿：长女名叫 米拉 ，次女名叫 米甲 。
1SAM|14|50|扫罗 的妻子名叫 亚希暖 ，是 亚希玛斯 的女儿。 扫罗 军队的元帅名叫 押尼珥 ，是 扫罗 的叔叔 尼珥 的儿子。
1SAM|14|51|扫罗 的父亲 基士 ， 押尼珥 的父亲 尼珥 ，都是 亚别 的儿子。
1SAM|14|52|扫罗 有生之年常与 非利士 人激烈争战，他看到任何有能力的人或勇士，都招募来跟随他。
1SAM|15|1|撒母耳 对 扫罗 说：“耶和华差遣我膏你为王，治理他的百姓 以色列 ，现在你要听从耶和华的话。
1SAM|15|2|万军之耶和华如此说：‘ 以色列 人从 埃及 上来的时候，在路上 亚玛力 人怎样待他们，怎样抵挡他们，我都要惩罚。
1SAM|15|3|现在你要去攻打 亚玛力 人，灭尽他们所有的，不可怜惜他们，将男女、孩童、吃奶的，以及牛、羊、骆驼和驴全都杀死。’”
1SAM|15|4|于是 扫罗 在 提拉因 召集百姓，数点他们，共有二十万步兵和一万 犹大 人。
1SAM|15|5|扫罗 到了 亚玛力 的京城，在谷中设下埋伏。
1SAM|15|6|扫罗 对 基尼 人说：“你们离开 亚玛力 人下去吧，免得我把你们和 亚玛力 人一同杀灭，因为 以色列 众人从 埃及 上来的时候，你们曾恩待他们。”于是 基尼 人离开了 亚玛力 人。
1SAM|15|7|扫罗 攻打 亚玛力 人，从 哈腓拉 直到 埃及 东边的 书珥 ，
1SAM|15|8|生擒了 亚玛力 王 亚甲 ，用刀杀尽 亚玛力 的众百姓。
1SAM|15|9|扫罗 和百姓却怜惜 亚甲 ，爱惜上好的牛、羊、牛犊、羔羊，以及一切美物，不肯灭绝。但是凡看不上眼和没有价值的，他们尽都杀了。
1SAM|15|10|耶和华的话临到 撒母耳 说：
1SAM|15|11|“我立 扫罗 为王，我感到遗憾，因为他转去不跟从我，不遵守我的命令。” 撒母耳 就很生气，终夜哀求耶和华。
1SAM|15|12|撒母耳 清早起来，去见 扫罗 。有人告诉 撒母耳 说：“ 扫罗 到了 迦密 ，看哪，他在那里为自己立了纪念碑，又转身下到 吉甲 。”
1SAM|15|13|撒母耳 到了 扫罗 那里， 扫罗 对他说：“愿耶和华赐福给你，耶和华的命令我已遵守了。”
1SAM|15|14|撒母耳 说：“我耳中听见有羊叫、牛鸣的声音，又是什么呢？”
1SAM|15|15|扫罗 说：“这是百姓从 亚玛力 人那里带来的，因为他们爱惜上好的牛羊，要献给耶和华－你的上帝。其余的，我们都灭尽了。”
1SAM|15|16|撒母耳 对 扫罗 说：“住口吧！等我把耶和华昨夜向我所说的话告诉你。” 扫罗 说：“请说。”
1SAM|15|17|撒母耳 说：“你虽然看自己为小，你岂不是作了 以色列 诸支派的元首吗？耶和华膏你作了 以色列 的王。
1SAM|15|18|耶和华差遣你，吩咐你说：‘你去除灭那些犯罪的 亚玛力 人，攻打他们，直到把他们完全灭尽。’
1SAM|15|19|你为何没有听从耶和华的话呢？你为何急着扑向掠物，行耶和华眼中看为恶的事呢？”
1SAM|15|20|扫罗 对 撒母耳 说：“我听从了耶和华的话，行了耶和华派我行的路，擒了 亚玛力 王 亚甲 来，灭尽了 亚玛力 人。
1SAM|15|21|百姓却从掠物中取了牛羊，是当灭之物中最好的，要在 吉甲 献给耶和华－你的上帝。”
1SAM|15|22|撒母耳 说： “耶和华喜爱燔祭和祭物， 岂如喜爱人听从他的话呢？ 看哪，听命胜于献祭， 顺从胜于公羊的脂肪。
1SAM|15|23|悖逆与占卜的罪相等， 顽梗与拜偶像的罪孽相同。 因为你厌弃耶和华的命令， 耶和华也厌弃你作王。”
1SAM|15|24|扫罗 对 撒母耳 说：“我有罪了！我违背了耶和华的指示和你的命令；因为我惧怕百姓，听从了他们的话。
1SAM|15|25|现在求你赦免我的罪，同我回去，我好敬拜耶和华。”
1SAM|15|26|撒母耳 对 扫罗 说：“我不同你回去，因为你厌弃耶和华的命令，耶和华也厌弃你作 以色列 的王。”
1SAM|15|27|撒母耳 转身要走， 扫罗 抓住他外袍的衣角，外袍就断裂了。
1SAM|15|28|撒母耳 对他说：“今日耶和华使 以色列 国与你断绝，把这国赐给另一个比你更好的人。
1SAM|15|29|以色列 的大能者必不说谎，也不后悔，因为他不是世人，绝不后悔。”
1SAM|15|30|扫罗 说：“我有罪了。现在求你在我百姓的长老和 以色列 人面前尊重我，同我回去，我好敬拜耶和华－你的上帝。”
1SAM|15|31|于是 撒母耳 转身跟随 扫罗 回去， 扫罗 就敬拜耶和华。
1SAM|15|32|撒母耳 说：“把 亚玛力 王 亚甲 带到我这里来。” 亚甲 就欢欢喜喜地来到他面前，说：“死亡的苦难必定过去了。”
1SAM|15|33|撒母耳 说：“你既用刀使妇人丧子，你母亲在妇人中也必照样丧子。”于是， 撒母耳 在 吉甲 耶和华面前把 亚甲 砍碎了。
1SAM|15|34|撒母耳 回了 拉玛 。 扫罗 上他所住的 基比亚 ，回自己的家去了。
1SAM|15|35|撒母耳 直到死的日子，再没有见 扫罗 。但 撒母耳 为 扫罗 悲伤，因为耶和华遗憾立 扫罗 为 以色列 的王。
1SAM|16|1|耶和华对 撒母耳 说：“我既厌弃 扫罗 作 以色列 的王，你为他悲伤要到几时呢？你将膏油盛满了角；来，我差遣你到 伯利恒 人 耶西 那里去，因为我在他儿子中已看中了一个为我作王的。”
1SAM|16|2|撒母耳 说：“我怎么能去呢？ 扫罗 一听见，就会杀我。”耶和华说：“你可以手里牵一头小母牛去，说：‘我来是要向耶和华献祭。’
1SAM|16|3|你要请 耶西 来一同献祭，我会指示你当做的事。我对你说的那个人，你要为我膏他。”
1SAM|16|4|撒母耳 遵照耶和华的话去做，来到 伯利恒 ，城里的长老都战战兢兢出来迎接他，有人问他说：“你是为平安来的吗？”
1SAM|16|5|他说：“为平安来的，我来是要向耶和华献祭。你们要使自己分别为圣，来跟我一同献祭。” 撒母耳 把 耶西 和他众儿子分别为圣，请他们来一同献祭。
1SAM|16|6|他们来的时候， 撒母耳 看见 以利押 ，就心里说，耶和华的受膏者一定在耶和华面前了。
1SAM|16|7|耶和华却对 撒母耳 说：“不要只看他的外貌和他身材高大，我不拣选他。因为耶和华不像人看人，人是看外貌 ，耶和华是看内心。”
1SAM|16|8|耶西 叫 亚比拿达 从 撒母耳 面前经过， 撒母耳 说：“耶和华也不拣选他。”
1SAM|16|9|耶西 又叫 沙玛 经过， 撒母耳 说：“耶和华也不拣选他。”
1SAM|16|10|耶西 叫他七个儿子都从 撒母耳 面前经过， 撒母耳 对 耶西 说：“这些都不是耶和华所拣选的。”
1SAM|16|11|撒母耳 对 耶西 说：“你的儿子都在这里了吗？”他说：“还有一个最小的，看哪，他正在放羊。” 撒母耳 对 耶西 说：“你派人去叫他来；他若不来这里，我们必不坐席。”
1SAM|16|12|耶西 就派人去叫他来。他面色红润，双目清秀，容貌俊美。耶和华说：“起来，膏他，因为这就是他了。”
1SAM|16|13|撒母耳 就用角里的膏油，在他的兄长中膏了他。从这日起，耶和华的灵就大大感动 大卫 。 撒母耳 起身回 拉玛 去了。
1SAM|16|14|耶和华的灵离开 扫罗 ，有邪灵从耶和华那里来扰乱他。
1SAM|16|15|扫罗 的臣仆对他说：“看哪，有邪灵从上帝那里来扰乱你。
1SAM|16|16|我们的主可以吩咐你面前的臣仆，去找一个善于弹琴的来。上帝那里来的邪灵临到你身上的时候，他用手弹琴，你就会感觉爽快。”
1SAM|16|17|扫罗 对臣仆说：“你们给我找一个善于弹琴的，带到我这里来。”
1SAM|16|18|仆人中有一个回答说：“看哪，我曾见 伯利恒 人 耶西 的一个儿子善于弹琴，是大能的勇士，说话合宜，容貌俊美，耶和华也与他同在。”
1SAM|16|19|于是 扫罗 差遣使者到 耶西 那里，说：“叫你放羊的儿子 大卫 到我这里来。”
1SAM|16|20|耶西 把几个饼和一皮袋酒，以及一只小山羊，驮在驴上，由儿子 大卫 的手送给 扫罗 。
1SAM|16|21|大卫 到了 扫罗 那里，就侍立在 扫罗 面前。 扫罗 很喜欢他，他就作了 扫罗 拿兵器的人。
1SAM|16|22|扫罗 派人到 耶西 那里，说：“让 大卫 侍立在我面前，因为他在我眼前蒙了恩宠。”
1SAM|16|23|从上帝那里来的邪灵临到 扫罗 身上的时候， 大卫 就拿琴，用手弹奏，使 扫罗 舒畅，感觉爽快，那邪灵就离开他了。
1SAM|17|1|非利士 人召集他们的军队来争战。他们聚集在 犹大 的 梭哥 ，在 梭哥 和 亚西加 中间的 以弗．大悯 安营。
1SAM|17|2|扫罗 和 以色列 人也聚集，在 以拉谷 安营，摆阵迎战，要与 非利士 人打仗。
1SAM|17|3|非利士 人站在这边的山上， 以色列 人站在那边的山上，当中有谷。
1SAM|17|4|从 非利士 营中出来一个挑战的人，名叫 歌利亚 ，是 迦特 人，身高六肘一虎口。
1SAM|17|5|他头戴铜盔，身穿铠甲，甲重五千舍客勒铜。
1SAM|17|6|他腿上有铜护膝，两肩之中背负铜矛。
1SAM|17|7|他的枪杆粗如织布机的轴，枪头的铁重六百舍客勒。有一个拿盾牌的人走在他前面。
1SAM|17|8|歌利亚 站着，对 以色列 的军队喊叫，对他们说：“你们出来摆阵作战是为了什么呢？我不是 非利士 人吗？你们不是 扫罗 的仆人吗？你们选一个人出来，叫他下来到我这里吧。
1SAM|17|9|他若能与我决斗，把我杀死，我们就作你们的奴隶；我若胜了他，把他杀死，你们就作我们的奴隶，服事我们。”
1SAM|17|10|那 非利士 人又说：“我今日向 以色列 的军队骂阵。你们叫一个人出来，跟我决斗吧。”
1SAM|17|11|扫罗 和 以色列 众人听见 非利士 人这些话就惊惶，非常害怕。
1SAM|17|12|大卫 是 犹大 伯利恒 的 以法他 人 耶西 的儿子， 耶西 有八个儿子。在 扫罗 的时候，这人年老，在众人中受敬重 。
1SAM|17|13|耶西 最大的三个儿子跟随 扫罗 出征。出征的三个儿子名字是：长子 以利押 ，次子 亚比拿达 ，三子 沙玛 。
1SAM|17|14|大卫 是最小的，最大的三个儿子跟随 扫罗 。
1SAM|17|15|大卫 有时离开 扫罗 ，回 伯利恒 为他父亲放羊。
1SAM|17|16|那 非利士 人早晚都出来站着，共四十日。
1SAM|17|17|耶西 对他儿子 大卫 说：“你拿一伊法烘了的穗子和十个饼，跑到营里去，交给你的哥哥，
1SAM|17|18|再拿这十块奶饼，送给他们的千夫长，并要问你哥哥好，向他们要个凭据回来。”
1SAM|17|19|扫罗 和 大卫 的三个哥哥，以及 以色列 众人，都在 以拉谷 与 非利士 人打仗。
1SAM|17|20|大卫 早晨起来，把羊交托一个看守的人，照 耶西 所吩咐的带着食物去了。到了军营，军队刚出到战场，呐喊叫阵。
1SAM|17|21|以色列 人和 非利士 人都摆列阵势，彼此相对。
1SAM|17|22|大卫 把东西留在看守物件的人手中，跑到战场，问他哥哥好。
1SAM|17|23|他与他们说话的时候，看哪，那挑战的人，就是 迦特 的 非利士 人 歌利亚 ，从 非利士 队伍中上来，说了同样的话， 大卫 听见了。
1SAM|17|24|以色列 众人看见那人就非常害怕，从他面前逃跑。
1SAM|17|25|以色列 人说：“这上来的人你看见了吗？他上来是要向 以色列 人骂阵。若有人能杀他，王必赏赐他大财，将自己的女儿嫁给他，并在 以色列 人中免除他父家纳粮服役。”
1SAM|17|26|大卫 对站在旁边的人说：“若有人杀这 非利士 人，除掉 以色列 人的羞辱，他会怎样呢？这未受割礼的 非利士 人是谁，竟敢向永生上帝的军队骂阵！”
1SAM|17|27|百姓照同样的话对他说：“若有人杀了那人，必这样待他。”
1SAM|17|28|大卫 的长兄 以利押 听见 大卫 与他们所说的话，就向他发怒，说：“你下来做什么呢？在旷野的那几只羊，你交托谁了呢？我知道你的骄傲和你心里的恶意，你下来只是为了看战争！”
1SAM|17|29|大卫 说：“我现在做了什么呢？只是问一句话也不可以吗？”
1SAM|17|30|大卫 离开他转向别人，问了同样的事，百姓也照先前的话回答他。
1SAM|17|31|有人听见 大卫 所说的话，就在 扫罗 面前报告； 扫罗 就派人叫他来。
1SAM|17|32|大卫 对 扫罗 说：“人不必因那 非利士 人灰心。你的仆人要去与他决斗。”
1SAM|17|33|扫罗 对 大卫 说：“你不能去与那 非利士 人决斗，因为你年纪太轻，他从小就是战士。”
1SAM|17|34|大卫 对 扫罗 说：“你仆人为父亲放羊，有时狮子来了，有时熊来了，从群中抓走一只羔羊。
1SAM|17|35|我就追赶它，击打它，把羔羊从它口中救出来。它起来攻击我，我就揪它的胡子，打死它。
1SAM|17|36|你仆人曾打死狮子和熊，这未受割礼的 非利士 人必像狮子和熊一样，因为他向永生上帝的军队骂阵。”
1SAM|17|37|大卫 又说：“耶和华救我脱离狮子和熊的爪，他必救我脱离这 非利士 人的手。” 扫罗 对 大卫 说：“你去吧！耶和华必与你同在。”
1SAM|17|38|扫罗 把自己的战衣给 大卫 穿上，将铜盔戴在他头上，又给他穿上铠甲。
1SAM|17|39|大卫 佩刀在战衣上，试着走走看。因 大卫 没有试过，就对 扫罗 说：“我穿戴这些不能走路，因为我没有试过。”于是他脱下身上的这些军装。
1SAM|17|40|他手中拿杖，又在溪中挑选了五块光滑的石子，放在袋里，就是牧人带的囊里，手里拿着甩石的机弦，迎向那 非利士 人。
1SAM|17|41|那 非利士 人渐渐走近 大卫 ，拿盾牌的人在他前面。
1SAM|17|42|非利士 人观看，见了 大卫 ，就藐视他，因为他年轻，面色红润，容貌俊美。
1SAM|17|43|非利士 人对 大卫 说：“你拿着杖到我这里来，我岂是狗吗？” 非利士 人就指着自己的神明诅咒 大卫 。
1SAM|17|44|非利士 人又对 大卫 说：“来吧！我要把你的肉给空中的飞鸟和田野的走兽。”
1SAM|17|45|大卫 对 非利士 人说：“你来攻击我，是靠着刀枪和铜矛，但我来攻击你，是靠着万军之耶和华的名，就是你所辱骂、带领 以色列 军队的上帝。
1SAM|17|46|今日耶和华必将你交在我手里。我必杀你，砍下你的头，今日我要把 非利士 军兵的尸体给空中的飞鸟和地上的野兽，使全地的人都知道以色列中有上帝，
1SAM|17|47|又使这里的全会众知道，耶和华使人得胜，不是用刀用枪，因为战争全在乎耶和华。他必将你们交在我们手里。”
1SAM|17|48|那 非利士 人起来，迎向 大卫 ，走近前来。 大卫 急忙往战场，迎向 非利士 人跑去。
1SAM|17|49|大卫 伸手入囊中，从里面掏出一块石子来，用机弦甩去，击中 非利士 人的前额，石子进入额内，他就仆倒，面伏于地。
1SAM|17|50|这样， 大卫 用机弦和石子胜了那 非利士 人，击中了他，把他杀死； 大卫 手中没有刀。
1SAM|17|51|大卫 跑去，站在那 非利士 人身旁，把他的刀从鞘中拔出来，杀死他，用刀割下他的头。 非利士 众人看见他们的勇士死了，就都逃跑。
1SAM|17|52|以色列 人和 犹大 人就起来呐喊，追赶 非利士 人，直到 该 和 以革伦 的城门。被杀的 非利士 人倒在路上，从 沙拉音 直到 迦特 和 以革伦 。
1SAM|17|53|以色列 人追赶 非利士 人回来，抢夺了他们的军营。
1SAM|17|54|大卫 拿着那 非利士 人的头带到 耶路撒冷 ，却把那 非利士 人的军装放在自己的帐棚里。
1SAM|17|55|扫罗 看见 大卫 去迎战 非利士 人，就问 押尼珥 元帅说：“ 押尼珥 ，那年轻人是谁的儿子？” 押尼珥 说：“王啊，我在你面前起誓，我不知道。”
1SAM|17|56|王说：“你可以问问那孩子是谁的儿子。”
1SAM|17|57|大卫 打死那 非利士 人回来， 押尼珥 领他到 扫罗 面前， 大卫 手中拿着 非利士 人的头。
1SAM|17|58|扫罗 问他说：“年轻人，你是谁的儿子？” 大卫 说：“我是你仆人 伯利恒 人 耶西 的儿子。”
1SAM|18|1|大卫 对 扫罗 说完了话， 约拿单 的心与 大卫 的心深相契合。 约拿单 爱 大卫 ，如同爱自己的性命。
1SAM|18|2|那日 扫罗 留住 大卫 ，不让他回父家。
1SAM|18|3|约拿单 爱 大卫 如同爱自己的性命，就与他立约。
1SAM|18|4|约拿单 从身上脱下外袍，给了 大卫 ，又把战衣、刀、弓、腰带都给了他。
1SAM|18|5|扫罗 无论差遣 大卫 往何处去，他都做事精明。 扫罗 立他作军队的指挥官，众百姓和 扫罗 的臣仆都看为美。
1SAM|18|6|大卫 打死了那 非利士 人，同众人回来的时候，妇女们从 以色列 各城里出来，欢欢喜喜，打鼓奏乐，唱歌跳舞，迎接 扫罗 王。
1SAM|18|7|众妇女欢乐唱和，说： “ 扫罗 杀死千千， 大卫 杀死万万。”
1SAM|18|8|扫罗 非常愤怒，不喜欢这话。他说：“将万万归给 大卫 ，千千归给我，只剩下王国没有给他！”
1SAM|18|9|从这日起， 扫罗 就敌视 大卫 。
1SAM|18|10|次日，从上帝来的邪灵紧抓住 扫罗 ，他就在家中胡言乱语。 大卫 照常弹琴， 扫罗 手里拿着枪。
1SAM|18|11|扫罗 把枪一掷，心里说：“我要将 大卫 刺透，钉在墙上。” 大卫 闪避了他两次。
1SAM|18|12|扫罗 惧怕 大卫 ，因为耶和华离开自己，与 大卫 同在。
1SAM|18|13|所以 扫罗 叫 大卫 离开自己，立他为千夫长，他就领兵出入。
1SAM|18|14|大卫 所做的每一件事都精明，耶和华也与他同在。
1SAM|18|15|扫罗 见 大卫 做事精明，就更怕他。
1SAM|18|16|但 以色列 和 犹大 众人都爱 大卫 ，因为他领他们出入。
1SAM|18|17|扫罗 对 大卫 说：“看哪，我将大女儿 米拉 嫁给你，只要你作我的勇士，为耶和华争战。” 扫罗 心里说：“我不好亲手害他，要藉 非利士 人的手害他。”
1SAM|18|18|大卫 对 扫罗 说：“我是谁，我是什么出身，我父家在 以色列 中算什么，岂敢作王的女婿呢？”
1SAM|18|19|扫罗 的女儿 米拉 到了当嫁给 大卫 的时候， 扫罗 却将她嫁给了 米何拉 人 亚得列 。
1SAM|18|20|扫罗 的女儿 米甲 爱 大卫 。有人告诉 扫罗 ，这件事在 扫罗 眼中看为合宜。
1SAM|18|21|扫罗 心里说：“我把这女儿嫁给 大卫 ，作他的圈套，好藉 非利士 人的手害他。”所以 扫罗 第二次对 大卫 说：“你今日可以作我的女婿。”
1SAM|18|22|扫罗 吩咐臣仆：“你们暗中对 大卫 说：‘看哪，王喜欢你，王的臣仆也都爱戴你，现在你就作王的女婿吧。’”
1SAM|18|23|扫罗 的臣仆照这话说给 大卫 听。 大卫 说：“你们把作王的女婿看为小事吗？我是贫穷卑微的人。”
1SAM|18|24|扫罗 的臣仆回奏说， 大卫 说了这样的话。
1SAM|18|25|扫罗 说：“你们要对 大卫 这样说：‘王不要什么聘礼，只要一百 非利士 人的包皮，好在王的仇敌身上报仇。’” 扫罗 的意图是要 大卫 落在 非利士 人的手中。
1SAM|18|26|扫罗 的臣仆把这话告诉 大卫 ， 大卫 就欢喜作王的女婿。日期还没有到，
1SAM|18|27|大卫 和跟随他的人起来前往，杀了二百 非利士 人，将包皮足数交给王，为要作王的女婿。于是 扫罗 将女儿 米甲 嫁给 大卫 。
1SAM|18|28|扫罗 见耶和华与 大卫 同在，女儿 米甲 又爱 大卫 ，
1SAM|18|29|就更怕 大卫 ，常常与 大卫 为敌。
1SAM|18|30|每逢 非利士 的军官出来打仗， 大卫 做事比 扫罗 任何臣仆更精明，因此他的名极受尊重。
1SAM|19|1|扫罗 吩咐他儿子 约拿单 和众臣仆要杀 大卫 ，但 扫罗 的儿子 约拿单 却很喜爱 大卫 。
1SAM|19|2|约拿单 告诉 大卫 说：“我父 扫罗 想要杀你，现在你要小心，明日早晨留在一个僻静的地方藏起来。
1SAM|19|3|我会出去，到你所藏的田里，站在我父亲旁边，与父亲谈论到你。我看情形怎样，会告诉你。”
1SAM|19|4|约拿单 向他父亲 扫罗 说 大卫 的好话，对他说：“王不可得罪王的仆人 大卫 ，因为他未曾得罪你，他所行的对你都很有益处。
1SAM|19|5|他拚了命杀那 非利士 人，并且耶和华为全 以色列 大施拯救。那时你看见，也很欢喜，现在为何要犯罪，流无辜人的血，无缘无故杀 大卫 呢？”
1SAM|19|6|扫罗 听了 约拿单 的话，就指着永生的耶和华起誓：“我绝不杀他。”
1SAM|19|7|约拿单 叫 大卫 来，把这一切事告诉他。 约拿单 带他去见 扫罗 ，他就像以前一样侍立在 扫罗 面前。
1SAM|19|8|此后又有战争， 大卫 出去与 非利士 人打仗。他大大击败他们，他们就在他面前逃跑。
1SAM|19|9|从耶和华来的邪灵又降在 扫罗 身上， 扫罗 手里拿枪坐在屋里， 大卫 正用手弹琴。
1SAM|19|10|扫罗 想要用枪刺透 大卫 ，把他钉在墙上，他却躲开 扫罗 ， 扫罗 的枪刺入墙内。当夜 大卫 逃走，躲起来了。
1SAM|19|11|扫罗 派一些使者到 大卫 的房屋那里守着他，等到天亮要杀他。 大卫 的妻子 米甲 对 大卫 说：“你今夜若不逃命，明日就要被杀。”
1SAM|19|12|于是 米甲 将 大卫 从窗户缒下去，让他走； 大卫 就逃走，躲起来了。
1SAM|19|13|米甲 把家中的神像放在床上，头枕在山羊毛的枕头上，用衣服盖起来。
1SAM|19|14|扫罗 派一些使者去捉拿 大卫 ， 米甲 说：“他病了。”
1SAM|19|15|扫罗 又派一些使者去看 大卫 ，说：“把他连床一起抬到我这里，我好杀他。”
1SAM|19|16|使者进去，看哪，神像在床上，头枕在山羊毛的枕头上。
1SAM|19|17|扫罗 对 米甲 说：“你为什么这样欺骗我，放我仇敌逃走呢？” 米甲 对 扫罗 说：“他对我说：‘你放我走吧，我何必要杀你呢？’”
1SAM|19|18|大卫 逃跑躲避，来到 拉玛 的 撒母耳 那里，把 扫罗 向他所行的事全告诉他。他和 撒母耳 就去，住在 拿约 。
1SAM|19|19|有人告诉 扫罗 说：“看哪， 大卫 在 拉玛 的 拿约 ”。
1SAM|19|20|扫罗 派一些使者去捉拿 大卫 。去的人见一队先知受感说话， 撒母耳 站在当中领导他们， 扫罗 派去的使者也受上帝的灵感动说话。
1SAM|19|21|有人把这事告诉 扫罗 ，他又派另一些使者去，他们也受感说话。 扫罗 第三次派使者去，他们也受感说话。
1SAM|19|22|然后 扫罗 亲自往 拉玛 去，到了 西沽 的大井，问人说：“ 撒母耳 和 大卫 在哪里？”有人说：“看哪，在 拉玛 的 拿约 。”
1SAM|19|23|他就往那里去，到了 拉玛 的 拿约 。上帝的灵也临到他，他一面走一面受感说话，直到 拉玛 的 拿约 。
1SAM|19|24|他也脱了衣服，也在 撒母耳 面前受感说话，一日一夜赤身躺卧。因此有人说：“ 扫罗 也在先知中吗？”
1SAM|20|1|大卫 从 拉玛 的 拿约 逃跑，来到 约拿单 面前，对他说：“我做了什么，有什么罪孽，在你父亲面前犯了什么罪，他竟要寻索我的性命呢？”
1SAM|20|2|约拿单 对他说：“绝无此事！你必不至于死。看哪，我父做事，无论大小，没有不告诉我的。我父亲为什么要隐瞒我这件事呢？不会这样的！”
1SAM|20|3|大卫 又起誓说：“你父亲确实知道我在你眼前蒙恩。所以他说，‘这事不要让 约拿单 知道，免得他愁烦。’我指着永生的耶和华起誓，又指着你的性命起誓，我离死只差一步而已。”
1SAM|20|4|约拿单 对 大卫 说：“你心里所求的，我必为你成就。”
1SAM|20|5|大卫 对 约拿单 说：“看哪，明日是初一，我必须与王同席用餐，求你让我去藏在田野，直到第三日傍晚。
1SAM|20|6|你父亲若见我不在席上，你就说：‘ 大卫 恳求我允许他赶回本城 伯利恒 去，因为他全家在那里献年祭。’
1SAM|20|7|你父亲若说好，你的仆人就平安了；他若大怒，你就知道他决意行恶。
1SAM|20|8|求你施恩于仆人，因你在耶和华面前曾与仆人立约。我若有罪孽，你就亲自杀死我，何必把我交给你父亲呢？”
1SAM|20|9|约拿单 说：“绝无此事！我若确实知道我父亲决意害你，怎么会不告诉你呢？”
1SAM|20|10|大卫 对 约拿单 说：“你父亲若严厉回答你，谁来告诉我呢？”
1SAM|20|11|约拿单 对 大卫 说：“来，让我们到田野去。”二人就往田野去了。
1SAM|20|12|约拿单 对 大卫 说：“愿耶和华－ 以色列 的上帝作证。明日约在这时候，或第三日，我一探出我父亲的心意，看哪，若对 大卫 是好意，我怎么会不派人来告诉你呢？
1SAM|20|13|我父亲若有意害你，而我不告诉你，送你平安地离开，愿耶和华重重惩罚 约拿单 。愿耶和华与你同在，如同从前与我父亲同在一样。
1SAM|20|14|你要照耶和华的慈爱恩待我，不但我活着的时候免我死亡，
1SAM|20|15|就是耶和华从地面逐一剪除 大卫 仇敌的时候，你也永不可向我家断绝恩惠。”
1SAM|20|16|于是 约拿单 与 大卫 家立约：“愿耶和华从 大卫 仇敌 的手来追讨。”
1SAM|20|17|约拿单 因爱 大卫 如同爱自己的性命，就叫他再起誓。
1SAM|20|18|约拿单 对他说：“明日是初一，你的座位空着，人必察觉你不在。
1SAM|20|19|到第三日，就要走一段长路下去 ，去到你遇事那天所藏的地方，在 以色 磐石 的旁边等候。
1SAM|20|20|我会向磐石旁边射三箭，如同射箭靶一样。
1SAM|20|21|看哪，我会派僮仆，说：‘去把箭找来。’我若对僮仆喊说：‘看哪，箭在你的这边，把箭拿来’，你就可以平安回来；我指着永生的耶和华起誓，你一定没有事。
1SAM|20|22|我若对孩子说：‘看哪，箭在你的前方’，你就要离开，因为是耶和华差你去的。
1SAM|20|23|至于你和我，我们所说的话，看哪，耶和华在你我中间作证，直到永远。”
1SAM|20|24|大卫 就去藏在田野。到了初一，王要坐席用餐。
1SAM|20|25|王照常坐在靠墙的位子上， 约拿单 在对面 ， 押尼珥 坐在 扫罗 旁边， 大卫 的座位却是空的。
1SAM|20|26|这日 扫罗 没有说什么，因为他说：“ 大卫 或许有事，偶染不洁，还未得洁净。”
1SAM|20|27|初二， 大卫 的座位还空着。 扫罗 对他儿子 约拿单 说：“ 耶西 的儿子为何昨日、今日都没有来用餐呢？”
1SAM|20|28|约拿单 回答 扫罗 说：“ 大卫 恳求我允许他回 伯利恒 去，
1SAM|20|29|说：‘求你让我去，因为我家在城里有献祭的事，我哥哥吩咐我去。如今我若在你眼前蒙恩，求你让我去见我的兄弟。’所以 大卫 没有来赴王的筵席。”
1SAM|20|30|扫罗 向 约拿单 怒气大发，对他说：“你这顽梗悖逆之妇人所生的，我怎么会不知道你选择 耶西 的儿子 ，自取羞辱，也使你母亲露体蒙羞呢？
1SAM|20|31|只要 耶西 的儿子还活在世上一天，你和你的国必保不住。现在你要派人去，把他带到我这里来，因为他是该死的。”
1SAM|20|32|约拿单 回答父亲 扫罗 说：“他为什么该死呢？他做了什么呢？”
1SAM|20|33|扫罗 向 约拿单 掷枪要刺他， 约拿单 就知道他父亲决意要杀死 大卫 。
1SAM|20|34|于是 约拿单 气愤愤地从席上起来。他在初二这天没有吃饭，因为他为 大卫 愁烦，又因为他父亲羞辱了他。
1SAM|20|35|次日早晨， 约拿单 按着与 大卫 约定的时候到田野去，有一个小僮仆跟随他。
1SAM|20|36|约拿单 对僮仆说：“你跑去把我所射的箭找来。”僮仆跑去， 约拿单 就把箭射在僮仆的前方。
1SAM|20|37|僮仆到了 约拿单 落箭之地， 约拿单 呼叫僮仆说：“箭不是在你的前方吗？”
1SAM|20|38|约拿单 又呼叫僮仆说：“快去，不要站在那里！”僮仆就捡起箭来，回到主人那里。
1SAM|20|39|僮仆不知道这是什么意思，只有 约拿单 和 大卫 知道这事。
1SAM|20|40|约拿单 把他的弓箭交给僮仆，吩咐他说：“你拿到城里去。”
1SAM|20|41|僮仆一去， 大卫 就从南边 出来，俯伏在地，拜了三拜。他们彼此亲吻，一起哭泣， 大卫 哭得更悲哀。
1SAM|20|42|约拿单 对 大卫 说：“你平平安安地去吧！因为我们二人曾指着耶和华的名起誓说：‘愿耶和华在你我中间，以及你我后裔中间作证，直到永远。’” 大卫 就起身走了， 约拿单 也回城里去了。
1SAM|21|1|大卫 到了 挪伯 的 亚希米勒 祭司那里， 亚希米勒 战战兢兢地出来迎接他，对他说：“你为什么独自一人，没有人跟随你呢？”
1SAM|21|2|大卫 对 亚希米勒 祭司说：“王吩咐我一件事，对我说：‘我差遣你，吩咐你的这件事，不可让任何人知道。’因此我已告诉一些仆人到某处去 。
1SAM|21|3|现在你手中有什么？请你给我五个饼或是可以找到的食物。”
1SAM|21|4|祭司对 大卫 说：“我手中没有普通的饼，只有圣饼，只能给没有亲近妇人的年轻人。”
1SAM|21|5|大卫 回答祭司说：“我们确实没有亲近妇人，如同往常我出征的时候一样。平常行路，仆人的身体 都还分别为圣，何况今日岂不更使自己分别为圣吗？”
1SAM|21|6|祭司拿圣饼给他，因为在那里没有别的饼，只有那从耶和华面前撤下的供饼，就是换上热饼的日子取下来的。
1SAM|21|7|当日，有 扫罗 的一个臣仆在那里，他留在耶和华的面前，名叫 多益 ，是 以东 人，作 扫罗 的畜牧长。
1SAM|21|8|大卫 对 亚希米勒 说：“你手中有没有枪或刀？因为王的事紧急，连刀剑兵器我都没有带。”
1SAM|21|9|祭司说：“你在 以拉谷 所杀的 非利士 人 歌利亚 的那刀，看哪，裹在布中，放在以弗得后边。你若要可以拿去，除此以外，再没有别的了。” 大卫 说：“没有什么可以跟它比的了！请你给我。”
1SAM|21|10|那日 大卫 起来，躲避 扫罗 ，逃到 迦特 王 亚吉 那里。
1SAM|21|11|亚吉 的臣仆对他说：“这不是那地的国王 大卫 吗？那里的人跳舞唱和： ‘ 扫罗 杀死千千， 大卫 杀死万万’， 不是指着他说的吗？”
1SAM|21|12|大卫 把这些话放在心里，就很惧怕 迦特 王 亚吉 。
1SAM|21|13|于是他在众人眼前一反常态，在他们中间 装疯作癫，在城门的门扇上胡写乱画，任由唾沫流在胡子上。
1SAM|21|14|亚吉 对臣仆说：“看哪，你们看这人疯了，为什么带他到我这里来呢？
1SAM|21|15|我岂缺少疯子，你们竟然带这人到我面前疯癫吗？这个人可以进我的家吗？”
1SAM|22|1|大卫 离开那里，逃到 亚杜兰 洞。他的兄弟和他父亲全家听见了，都下到他那里去。
1SAM|22|2|凡生活窘迫的、欠债的、心里苦恼的都聚集到 大卫 那里，他就作他们的领袖，跟随他的约有四百人。
1SAM|22|3|大卫 从那里往 摩押 的 米斯巴 去，对 摩押 王说：“请你让我父母搬来，跟你们在一起，等我知道上帝要为我怎样做。”
1SAM|22|4|大卫 领他父母到 摩押 王面前。 大卫 住山寨一切的日子，他父母也都住在 摩押 王那里。
1SAM|22|5|先知 迦得 对 大卫 说：“你不要住在山寨，要到 犹大 地去。” 大卫 就去，来到 哈列 的树林。
1SAM|22|6|扫罗 听见 大卫 和跟随他之人的下落， 扫罗 正在 基比亚 ，坐在山顶 的柳树下，手里拿着枪，众臣仆侍立在左右。
1SAM|22|7|扫罗 对左右侍立的臣仆说：“ 便雅悯 人哪，听着！ 耶西 的儿子也能把田地和葡萄园赐给你们各人吗？他能立你们各人作千夫长和百夫长吗？
1SAM|22|8|你们竟都结党害我！我儿子与 耶西 的儿子立约的时候，无人告诉我；我儿子挑唆我的臣仆谋害我，像今日这样，也无人告诉我，为我忧虑。”
1SAM|22|9|那时 以东 人 多益 站在 扫罗 的臣仆中，回答说：“我曾看见 耶西 的儿子往 挪伯 去，到了 亚希突 的儿子 亚希米勒 那里。
1SAM|22|10|亚希米勒 为他求问耶和华，给他食物，又把 非利士 人 歌利亚 的刀给了他。”
1SAM|22|11|王就派人把 亚希突 的儿子 亚希米勒 祭司和他父亲的全家，就是在 挪伯 的祭司都召了来，他们都来到王那里。
1SAM|22|12|扫罗 说：“ 亚希突 的儿子，听着！”他说：“我主，我在这里。”
1SAM|22|13|扫罗 对他说：“你为什么与 耶西 的儿子结党害我，把食物和刀给他，又为他求问上帝，使他起来谋害我，像今日这样？”
1SAM|22|14|亚希米勒 回答王说：“王的众臣仆中有谁比 大卫 忠心呢？他是王的女婿，又是你的侍卫长 ，并且是你宫中受敬重的人。
1SAM|22|15|我今日才开始为他求问上帝吗？绝非如此！王不要归罪于我和我父全家，因为这事，无论大小，仆人都不知情。”
1SAM|22|16|王说：“ 亚希米勒 ，你和你父全家都是该死的！”
1SAM|22|17|王吩咐左右的侍卫说：“你们转身去杀耶和华的祭司吧！因为他们帮助 大卫 ，知道 大卫 逃跑却不告诉我。”但王的臣仆都不愿动手杀耶和华的祭司。
1SAM|22|18|王吩咐 多益 说：“你转身去杀祭司吧！” 以东 人 多益 就转身去杀祭司，那日杀了穿细麻布以弗得的，共八十五人，
1SAM|22|19|又用刀把祭司城 挪伯 中的男女、孩童和吃奶的都杀了，又用刀杀了牛、羊和驴子。
1SAM|22|20|亚希突 的儿子 亚希米勒 有一个儿子逃脱了；他名叫 亚比亚他 ，逃到 大卫 那里。
1SAM|22|21|亚比亚他 把 扫罗 杀耶和华祭司的事告诉 大卫 。
1SAM|22|22|大卫 对 亚比亚他 说：“那日我见 以东 人 多益 在那里，就知道他一定会告诉 扫罗 。你父的全家丧命，都是因我的缘故。
1SAM|22|23|你可以住在我这里，不要惧怕。因为寻索你命的也要寻索我的命，你在我这里可得保护。”
1SAM|23|1|有人告诉 大卫 说：“看哪， 非利士 人攻击 基伊拉 ，抢夺禾场。”
1SAM|23|2|大卫 求问耶和华说：“我可以去吗？我可以去攻打那些 非利士 人吗？”耶和华对 大卫 说：“你可以去攻打 非利士 人，拯救 基伊拉 。”
1SAM|23|3|大卫 的人对他说：“看哪，我们在 犹大 这里尚且惧怕，何况到 基伊拉 去攻打 非利士 人的军队呢？”
1SAM|23|4|大卫 又再求问耶和华，耶和华回答说：“你起身下 基伊拉 去，我必将 非利士 人交在你手里。”
1SAM|23|5|于是 大卫 和他的人往 基伊拉 去，与 非利士 人打仗，大大击败他们，夺取他们的牲畜。这样， 大卫 救了 基伊拉 的居民。
1SAM|23|6|亚希米勒 的儿子 亚比亚他 逃往 基伊拉 到 大卫 那里的时候，手里拿着以弗得。
1SAM|23|7|有人告诉 扫罗 ， 大卫 到了 基伊拉 。 扫罗 说：“上帝将他交在我手里了，因为他进了有门有闩的城，把自己关起来了。”
1SAM|23|8|于是 扫罗 召集众百姓，要下去攻打 基伊拉 ，围困 大卫 和他的人。
1SAM|23|9|大卫 知道 扫罗 设计陷害他，就对 亚比亚他 祭司说：“把以弗得拿过来。”
1SAM|23|10|大卫 说：“耶和华－ 以色列 的上帝啊，你仆人确实听见 扫罗 设法要到 基伊拉 来，为我的缘故毁灭这城。
1SAM|23|11|基伊拉 人会把我交在 扫罗 手里吗？ 扫罗 会下来，正如你仆人所听见的吗？耶和华－ 以色列 的上帝啊，求你指示仆人！”耶和华说：“他会下来。”
1SAM|23|12|大卫 又说：“ 基伊拉 人会把我和我的人交在 扫罗 手里吗？”耶和华说：“他们会交出来。”
1SAM|23|13|于是 大卫 和他的人约有六百名起身离开 基伊拉 ，往他们所能去的地方去。有人告诉 扫罗 ， 大卫 离开 基伊拉 逃走了， 扫罗 就停止出发了。
1SAM|23|14|大卫 住在旷野的山寨里，在 西弗 旷野的山区。 扫罗 天天寻索 大卫 ，上帝却不将 大卫 交在他手里。
1SAM|23|15|大卫 看到 扫罗 出来寻索他的命。那时，他住在 西弗 旷野的树林里 ；
1SAM|23|16|扫罗 的儿子 约拿单 起身，到树林里去见 大卫 ，使他的手倚靠上帝得以坚固，
1SAM|23|17|对他说：“不要惧怕！我父 扫罗 的手无法害你 ，你必作 以色列 的王，我必作你的宰相。我父 扫罗 也知道这事。”
1SAM|23|18|于是二人在耶和华面前立约。 大卫 仍住在树林里， 约拿单 就回家去了。
1SAM|23|19|西弗 人上 基比亚 到 扫罗 那里，说：“ 大卫 不是在我们那里，在树林里的山寨中，在荒野 南边的 哈基拉山 藏着吗？
1SAM|23|20|现在，王啊，请随你的心愿要下来，就请下来；至于我们，一定会把他交在王的手里。”
1SAM|23|21|扫罗 说：“愿耶和华赐福给你们，因为你们体恤我。
1SAM|23|22|请你们回去，再确定一下，调查并看清楚他落脚的地方，是谁看见他在那里 ，因为有人告诉我他很狡猾。
1SAM|23|23|你们要看清楚，调查他藏匿的每一个地方，回来给我确实的报告，我就与你们同去。他若在境内，我必从 犹大 的千门万户中搜出他来。”
1SAM|23|24|西弗 人动身，在 扫罗 以先往 西弗 去。 大卫 和他的人却在 玛云 旷野，在荒野南边的 亚拉巴 。
1SAM|23|25|扫罗 和他的人去寻索 大卫 。有人告诉 大卫 ，他就下到岩石那里，留在 玛云 的旷野。 扫罗 听见了，就在 玛云 的旷野追赶 大卫 。
1SAM|23|26|扫罗 在山的这一边走， 大卫 和他的人在山的那一边。 大卫 急忙躲避 扫罗 ， 扫罗 和他的人正四面围住 大卫 和他的人，要捉拿他们。
1SAM|23|27|有使者来对 扫罗 说：“ 非利士 人入境抢掠，请快快回去！”
1SAM|23|28|于是 扫罗 不再追赶 大卫 ，回去迎击 非利士 人。因此那地方名叫 西拉．哈玛希罗结 。
1SAM|23|29|大卫 从那里上去，住在 隐．基底 的山寨里。
1SAM|24|1|扫罗 追赶 非利士 人回来，有人告诉他说：“看哪， 大卫 在 隐．基底 的旷野。”
1SAM|24|2|扫罗 就从全 以色列 中挑选三千精兵，往 野山羊磐石 的东边 去，寻索 大卫 和他的人。
1SAM|24|3|到了路旁的羊圈，在那里有个洞， 扫罗 进去大解。 大卫 和他的人正藏在洞里的深处。
1SAM|24|4|大卫 的人对 大卫 说：“看哪，这日子到了！耶和华曾对你说：‘看哪，我要将你的仇敌交在你手里，你可以照你看为好的对待他。’” 大卫 就起来，悄悄地割下 扫罗 外袍的衣角。
1SAM|24|5|随后 大卫 心中自责，因为他割下了 扫罗 的衣角。
1SAM|24|6|他对他的人说：“耶和华绝不允许我对我的主，耶和华的受膏者做这事，伸手害他，因为他是耶和华的受膏者。”
1SAM|24|7|大卫 用这话劝阻他的人，不许他们起来害 扫罗 。 扫罗 起来，从洞里出去，预备上路。
1SAM|24|8|然后 大卫 也起来，从洞里出去，呼唤 扫罗 说：“我主，我王！” 扫罗 回头观看， 大卫 就屈身，脸伏于地下拜。
1SAM|24|9|大卫 对 扫罗 说：“你为何听信人的谗言，说‘看哪， 大卫 想要害你’呢？
1SAM|24|10|看哪，今日你亲眼看见，在洞中耶和华将你交在我手里。有人要我杀你，我却爱惜你，说：‘我不敢伸手害我的主，因为他是耶和华的受膏者。’
1SAM|24|11|我父啊，请看，看你外袍的衣角在我手中。我割下你外袍的衣角，却没有杀你。你知道，并且看见我没有恶意要悖逆你。你虽然要猎取我的命，我却没有得罪你。
1SAM|24|12|愿耶和华在你我中间判断，愿耶和华在你身上为我伸冤，我却不亲手加害于你。
1SAM|24|13|古人有句俗语说：‘恶事出于恶人。’我却不亲手加害于你。
1SAM|24|14|以色列 王出来要寻找谁呢？你要追赶谁呢？不过是一条死狗，一只跳蚤而已。
1SAM|24|15|愿耶和华作仲裁者，在你我中间判断。愿他鉴察，为我伸冤，救我脱离你的手。”
1SAM|24|16|大卫 向 扫罗 说完了这些话， 扫罗 说：“我儿 大卫 ，这是你的声音吗？”于是 扫罗 放声大哭，
1SAM|24|17|对 大卫 说：“你比我公义，因为你以善待我，我却以恶待你。
1SAM|24|18|今日你已显明是以善待我，因为耶和华将我交在你手里，你却没有杀我。
1SAM|24|19|人若遇见仇敌，岂肯放他平安上路呢？愿耶和华因你今日向我所做的，以善回报你。
1SAM|24|20|现在，看哪，我知道你一定会作王， 以色列 的国必要坚立在你手里。
1SAM|24|21|现在你要指着耶和华向我起誓，你必不剪除我的后裔，必不从我父家除去我的名。”
1SAM|24|22|于是 大卫 向 扫罗 起誓， 扫罗 就回家去， 大卫 和他的人也上山寨去了。
1SAM|25|1|撒母耳 死了， 以色列 众人聚集，为他哀哭，把他葬在 拉玛 他的家里。 大卫 动身，下到 巴兰 的旷野。
1SAM|25|2|在 玛云 有一个人，他的产业在 迦密 。这人是一个大富翁，有三千只绵羊，一千只山羊；他正在 迦密 剪羊毛。
1SAM|25|3|这人名叫 拿八 ，他的妻子名叫 亚比该 。 拿八 的妻子有美好的见识，又有美丽的容貌，但 拿八 为人刚愎凶恶，是 迦勒 族的人。
1SAM|25|4|大卫 在旷野听见 拿八 正在剪羊毛，
1SAM|25|5|就派十个仆人，对他们说：“你们上 迦密 到 拿八 那里，提我的名向他问安。
1SAM|25|6|你们要如此说：‘愿你来年平安 ，愿你家平安，愿你一切所有的都平安。
1SAM|25|7|现在我听说你有剪羊毛的人，你的牧人和我们在一起，他们在 迦密 一切的日子，我们没有欺负过他们，他们也未曾失去什么。
1SAM|25|8|你问你的仆人，他们会告诉你。愿我的仆人在你眼前得欢心，因为我们是在好日子来的。请你随手分点食物给仆人和你儿子 大卫 。’”
1SAM|25|9|大卫 的仆人到了，就提 大卫 的名，把这一切话告诉 拿八 ，他们就停顿下来。
1SAM|25|10|拿八 回答 大卫 的仆人说：“ 大卫 是谁？ 耶西 的儿子是谁？今日悖逆主人奔逃的仆人很多。
1SAM|25|11|我岂可把饮食，以及我为剪羊毛的人所宰的肉给那些我不知道从哪里来的人呢？”
1SAM|25|12|大卫 的仆人转身从原路回去，照这一切的话告诉 大卫 。
1SAM|25|13|大卫 对他的人说：“你们各人都要佩上刀！”各人就都佩上刀， 大卫 也佩上刀。跟随 大卫 上去的约有四百人，留下二百人看守物件。
1SAM|25|14|拿八 的一个仆人告诉 拿八 的妻子 亚比该 说：“看哪， 大卫 从旷野派使者来向我主人问安，主人却辱骂他们。
1SAM|25|15|但是那些人待我们真好；我们在田野与他们一切来往的日子，没有受他们欺负，也未曾失去什么。
1SAM|25|16|我们在他们那里牧羊，一切的日子他们昼夜保护我们 。
1SAM|25|17|现在，你当知道，看怎样做才好。不然，祸患必定临到我主人和他全家。他性情凶暴，无人敢与他说话。”
1SAM|25|18|亚比该 急忙将二百个饼，两皮袋酒，五只宰好的羊，五细亚烘熟的穗子，一百个葡萄干饼，二百个无花果饼，都驮在驴上，
1SAM|25|19|对仆人说：“你们在我前面走，看哪，我跟着你们去。”她却没有告诉丈夫 拿八 。
1SAM|25|20|亚比该 骑着驴，正下山坡，看哪， 大卫 和他的人正迎着 亚比该 下来，她就去迎接他们。
1SAM|25|21|大卫 曾说：“我在旷野为那人看守他一切所有的，以致他未失去任何一样东西，实在是徒然了！他竟然向我以恶报善。
1SAM|25|22|凡属 拿八 的男丁，我若留一个到明日早晨，愿上帝重重惩罚 大卫 ！”
1SAM|25|23|亚比该 看见 大卫 ，就急忙下驴，在 大卫 面前脸伏于地叩拜。
1SAM|25|24|她俯伏在 大卫 的脚前，说：“我主啊，愿这罪归于我！求你容许使女向你进言，更求你听使女的话。
1SAM|25|25|我主不必理会 拿八 这性情凶暴的人，他就像他的名字一样；他名叫 拿八 ，为人也真是愚顽。至于我，你的使女并没有看见我主所派来的仆人。
1SAM|25|26|现在，我主啊，耶和华既然阻止你亲手报仇，避免流人的血，我指着永生的耶和华起誓，又指着你的性命起誓：‘现在，愿你的仇敌和谋害我主的人都像 拿八 一样。’
1SAM|25|27|现在求我主把婢女送来的礼物给跟随我主的仆人。
1SAM|25|28|求你原谅使女的冒犯。耶和华必为我主建立坚固的家，因为我主为耶和华争战，并且你一生的日子查不出有什么恶来。
1SAM|25|29|虽有人起来追逼你，要寻索你的性命，我主的性命在耶和华－你的上帝那里，如同藏在生命的宝藏中。至于你仇敌的性命，耶和华必甩去，如用机弦甩石一样。
1SAM|25|30|耶和华照所应许你的福气赐给我主，立你作 以色列 王的时候，
1SAM|25|31|我主就不至于因为亲手报仇，流了无辜人的血，而心里不安，良心有亏了。耶和华赐福给我主的时候，求你记得你的使女。”
1SAM|25|32|大卫 对 亚比该 说：“耶和华－ 以色列 的上帝是应当称颂的，因为他今日派你来迎接我。
1SAM|25|33|你和你的见识也配得称赞，因为你今日拦阻我亲手报仇、流人的血。
1SAM|25|34|我指着阻止我加害于你的耶和华－ 以色列 永生的上帝起誓，若不是你很快地来迎接我，到早晨天亮的时候，凡属 拿八 的男丁，必定一个也不留。”
1SAM|25|35|大卫 从 亚比该 手中收了她带来的礼物，对她说：“平平安安上你的家去吧！你看，我看了你的情面，听了你的话。”
1SAM|25|36|亚比该 到 拿八 那里，看哪，他在家里摆设宴席，如同王的宴席。 拿八 心情舒畅，酩酊大醉。所以 亚比该 大小事都没有告诉他，直等到早晨天亮的时候。
1SAM|25|37|到了早晨， 拿八 酒醒了，他的妻子把这些事都告诉他，他就发心脏病快死了，僵如石头。
1SAM|25|38|过了十天，耶和华击打 拿八 ，他就死了。
1SAM|25|39|大卫 听见 拿八 死了，就说：“耶和华是应当称颂的，因为我从 拿八 手中受了羞辱，他为我伸冤，又阻止他的仆人行恶；耶和华使 拿八 的恶归到他自己头上。”于是 大卫 派人去向 亚比该 说，要娶她为妻。
1SAM|25|40|大卫 的仆人来到 迦密 ，到 亚比该 那里，对她说：“ 大卫 派我们到你这里，要娶你作他的妻子。”
1SAM|25|41|亚比该 起来叩拜，俯伏在地，说：“看哪，你的使女情愿作婢女，为我主的仆人洗脚。”
1SAM|25|42|亚比该 立刻起身，骑上驴，五个女仆跟着她走。她跟从 大卫 的使者去，就作了 大卫 的妻子。
1SAM|25|43|大卫 先前娶了 耶斯列 人 亚希暖 ，她们二人都作了他的妻子。
1SAM|25|44|扫罗 已把他的女儿 米甲 ，就是 大卫 的妻子，给了 迦琳 人 拉亿 的儿子 帕提 为妻。
1SAM|26|1|西弗 人来到 基比亚 ，到 扫罗 那里，说：“ 大卫 不是在荒野 东边 的 哈基拉山 藏着吗？”
1SAM|26|2|扫罗 动身，带领 以色列 人中挑选的三千精兵下到 西弗 的旷野，要在那里寻索 大卫 。
1SAM|26|3|扫罗 在荒野东边的 哈基拉山 ，在路旁安营。那时 大卫 住在旷野，看见 扫罗 到旷野来追赶他，
1SAM|26|4|大卫 就派人去探听，知道 扫罗 果然来了。
1SAM|26|5|大卫 起来，到 扫罗 安营的地方，看见 扫罗 和 尼珥 的儿子 押尼珥 元帅躺卧之处； 扫罗 睡在军营里，士兵安营在他周围。
1SAM|26|6|大卫 对 赫 人 亚希米勒 和 洗鲁雅 的儿子 约押 的兄弟 亚比筛 说：“谁同我下到 扫罗 营里去？” 亚比筛 说：“我同你下去。”
1SAM|26|7|于是 大卫 和 亚比筛 夜间到了士兵那里；看哪， 扫罗 睡在军营里，他的枪在头旁，插在地上。 押尼珥 和士兵睡在他周围。
1SAM|26|8|亚比筛 对 大卫 说：“上帝将你的仇敌交在你手里，现在让我拿枪把他刺透在地上，一刺就成，不用再刺他了。”
1SAM|26|9|大卫 对 亚比筛 说：“不可杀害他！有谁伸手害耶和华的受膏者而无罪呢？”
1SAM|26|10|大卫 又说：“我指着永生的耶和华起誓，他或被耶和华击杀，或死期到了，或出战阵亡，
1SAM|26|11|耶和华绝不允许我伸手害耶和华的受膏者。现在你可以把他头旁的枪和水壶拿来，我们就走。”
1SAM|26|12|大卫 从 扫罗 的头旁拿了枪和水壶，他们就走了。没有人看见，没有人知道，也没有人醒过来。他们都睡着了，因为耶和华使他们沉睡了。
1SAM|26|13|大卫 过到另一边去，远远地站在山顶上，与他们相离很远。
1SAM|26|14|大卫 呼叫百姓和 尼珥 的儿子 押尼珥 说：“ 押尼珥 ，你为何不回答呢？” 押尼珥 回答说：“你是谁？竟敢呼唤王呢？”
1SAM|26|15|大卫 对 押尼珥 说：“你不是个大丈夫吗？ 以色列 中谁能比你呢？百姓中有一个人进来要害死你主你王，你为何没有保护你主你王呢？
1SAM|26|16|你做的这件事不好！我指着永生的耶和华起誓，你们都是该死的，因为你们没有保护你们的主，就是耶和华的受膏者。现在你看，王头旁的枪和水壶在哪里？”
1SAM|26|17|扫罗 认出 大卫 的声音，就说：“我儿 大卫 ，这是你的声音吗？” 大卫 说：“我主我王啊，是我的声音。”
1SAM|26|18|又说：“我主为何要追赶仆人呢？我做了什么？我手做了什么恶事呢？
1SAM|26|19|现在求我主我王听仆人的话：若是耶和华激发你来攻击我，愿耶和华悦纳供物；若是出于人，愿他们在耶和华面前受诅咒，因为他们今日赶逐我，不让我在耶和华的产业中有分，说：‘你去事奉别神吧！’
1SAM|26|20|现在不要使我的血流在远离耶和华面的地上。因为 以色列 王出来，只不过是寻找一只跳蚤，如同人在山上猎取一只鹧鸪。”
1SAM|26|21|扫罗 说：“我有罪了！我儿 大卫 ，回来吧！我必不再加害于你，因为你今日看我的性命为宝贵。看哪，我是个糊涂人，大大错了。”
1SAM|26|22|大卫 回答说：“看哪，这是王的枪，可以吩咐一个仆人过来拿去。
1SAM|26|23|今日耶和华将王交在我手里，我却不肯伸手害耶和华的受膏者。耶和华必照各人的公义诚实报应他。
1SAM|26|24|看哪，我今日看重你的性命，愿耶和华也照样看重我的性命，并且拯救我脱离一切患难。”
1SAM|26|25|扫罗 对 大卫 说：“我儿 大卫 ，愿你得福！你必做大事，也必得胜。”于是 大卫 上路， 扫罗 也回自己的地方去了。
1SAM|27|1|大卫 心里说：“总有一天我会死在 扫罗 手里，现在我最好逃到 非利士 人的地去， 扫罗 就会绝望，不会继续在 以色列 全境内寻索我了。这样，我才可以脱离他的手。”
1SAM|27|2|于是 大卫 动身，和跟随他的六百人投奔 玛俄 的儿子 迦特 王 亚吉 去了。
1SAM|27|3|大卫 和他的两个妻子，就是 耶斯列 人 亚希暖 和作过 拿八 妻子的 迦密 人 亚比该 ，以及他的人，连同各人的眷属，都住在 迦特 的 亚吉 那里。
1SAM|27|4|有人告诉 扫罗 ：“ 大卫 逃到 迦特 。” 扫罗 就不再寻索他了。
1SAM|27|5|大卫 对 亚吉 说：“我若蒙你看得起，求你在郊外的城镇中赐我一个地方，让我住在那里。仆人何必与王同住京城呢？”
1SAM|27|6|当日 亚吉 把 洗革拉 赐给他，因此 洗革拉 属于 犹大 王，直到今日。
1SAM|27|7|大卫 在 非利士 人的地，住的期间有一年四个月。
1SAM|27|8|大卫 和他的人上去，侵夺 基述 人、 基色 人、 亚玛力 人，这些是从 帖兰 经过 书珥 直到 埃及 地的居民 。
1SAM|27|9|大卫 攻击那地，无论男女没有留下一个活口，又夺获牛、羊、驴、骆驼和衣服，回来到 亚吉 那里。
1SAM|27|10|亚吉 说：“今日你们没有去抢夺什么地方吧 ？” 大卫 说：“侵夺了 犹大 、 耶拉篾 、 基尼 等地的南方。”
1SAM|27|11|无论男女， 大卫 没有留下一个活口带到 迦特 来。他说：“恐怕他们把我们的事告诉人，说：‘ 大卫 如此做了。’”这是他住在 非利士 人之地一切日子的惯例。
1SAM|27|12|亚吉 信了 大卫 ，说：“ 大卫 已经使本族 以色列 人憎恶他，所以他必永远作我的仆人了。”
1SAM|28|1|那时， 非利士 人召集军队，要与 以色列 打仗。 亚吉 对 大卫 说：“你当知道，你和你的人都要随我出征。”
1SAM|28|2|大卫 对 亚吉 说：“好，仆人所能做的事，王都知道。” 亚吉 对 大卫 说：“好，我立你终生作我 的侍卫。”
1SAM|28|3|那时 撒母耳 已经死了， 以色列 众人为他哀哭，把他葬在他的本城 拉玛 。 扫罗 曾在国内驱除招魂的和行巫术的人。
1SAM|28|4|非利士 人集合，来到 书念 安营； 扫罗 集合 以色列 众人在 基利波 安营。
1SAM|28|5|扫罗 看见 非利士 的军队，就惧怕，心中大大战兢。
1SAM|28|6|扫罗 求问耶和华，耶和华却不藉梦，或乌陵，或先知回答他。
1SAM|28|7|扫罗 吩咐臣仆说：“为我找一个招魂的妇人，我好去问她。”臣仆对他说：“看哪，在 隐．多珥 有一个招魂的妇人。”
1SAM|28|8|于是 扫罗 改了装，穿上别的衣服，带着两个人，夜里去见那妇人。 扫罗 说：“请你用招魂的法术，把我所告诉你的死人，为我招上来。”
1SAM|28|9|妇人对他说：“看哪，你知道 扫罗 所做的，他从国中剪除招魂的和行巫术的。你为何为我的性命设下罗网，要害死我呢？”
1SAM|28|10|扫罗 向妇人指着耶和华起誓说：“我指着永生的耶和华起誓，你必不因这事受罚。”
1SAM|28|11|妇人说：“我为你招谁上来呢？”他说：“为我招 撒母耳 上来。”
1SAM|28|12|妇人看见 撒母耳 ，就大声喊叫。妇人对 扫罗 说：“你是 扫罗 ，为什么欺骗我呢？”
1SAM|28|13|王对妇人说：“不要惧怕，你看见什么呢？”妇人对 扫罗 说：“我看见有神明从地里上来。”
1SAM|28|14|扫罗 说：“他是怎样的形状？”妇人说：“有一个老人上来，身穿长袍。” 扫罗 知道是 撒母耳 ，就屈身，脸伏于地下拜。
1SAM|28|15|撒母耳 对 扫罗 说：“你为什么搅扰我，招我上来呢？” 扫罗 说：“我十分为难，因为 非利士 人攻击我，上帝离开我，不再藉先知或梦回答我。因此请你上来，好指示我应当怎样做。”
1SAM|28|16|撒母耳 说：“耶和华已经离开你，与你为敌，你何必问我呢？
1SAM|28|17|耶和华照他藉我所说的话为他自己 实现了。耶和华已经从你手里夺去国权，赐给别人，就是 大卫 。
1SAM|28|18|因为你没有听从耶和华的话，没有执行他对 亚玛力 人的恼怒，所以今日耶和华向你做这事。
1SAM|28|19|耶和华也必将你和 以色列 交在 非利士 人手里。明日你和你儿子们必与我在一处了；耶和华也必将 以色列 的军兵交在 非利士 人手里。”
1SAM|28|20|扫罗 突然全身仆倒在地，因为 撒母耳 的话令他十分惧怕。他毫无气力，因为他一日一夜都没有吃什么。
1SAM|28|21|妇人到 扫罗 面前，见他极其惊恐，对他说：“看哪，婢女听从了你，不顾惜自己的性命，遵从你吩咐我的话。
1SAM|28|22|现在求你也听婢女的话，让我在你面前摆上一点食物，你吃了才有气力上路。”
1SAM|28|23|扫罗 不肯，说：“我不吃。”但他的仆人和那妇人再三劝他，他才听他们的话，从地上起来，坐在床上。
1SAM|28|24|妇人急忙把家里的一只肥牛犊宰了，又拿面来揉，烤成无酵饼，
1SAM|28|25|摆在 扫罗 和他仆人面前。他们吃了，当夜就起身走了。
1SAM|29|1|非利士 人聚集他们所有的军队到 亚弗 ； 以色列 人在 耶斯列 的泉旁安营。
1SAM|29|2|非利士 人的领袖各率队伍，或百或千的前进； 大卫 和他的人同 亚吉 跟在后边前进。
1SAM|29|3|非利士 人的领袖说：“这些 希伯来 人在这里做什么呢？” 亚吉 对 非利士 人的领袖说：“这不是 以色列 王 扫罗 的臣仆 大卫 吗？他在我这里有些年日了。自从他投降直到今日，我未曾见他有什么过错。”
1SAM|29|4|非利士 人的领袖向 亚吉 发怒，对他说：“叫这人回去！叫他回到你指派他的地方去，不可让他同我们出征，免得他在阵上反成为我们的敌人。他用什么与他主人复和呢？岂不是用我们这些人的首级吗？
1SAM|29|5|有人跳舞唱和说： ‘ 扫罗 杀死千千， 大卫 杀死万万’， 不就是这个 大卫 吗？”
1SAM|29|6|亚吉 叫 大卫 来，对他说：“我指着永生的耶和华起誓，你是个正直人。你随我在军中出入，我也很满意。自从你投奔我到如今，我未曾看见你有什么过失，但是众领袖看你不顺眼。
1SAM|29|7|现在你平平安安地回去，不要做 非利士 人领袖眼中看为恶的事。”
1SAM|29|8|大卫 对 亚吉 说：“但我做了什么呢？自从仆人到你面前，直到今日，你查出我有什么过错，使我不去攻击我主我王的仇敌呢？”
1SAM|29|9|亚吉 回答 大卫 说：“我知道你在我眼中是好人，如同上帝的使者一样，只是 非利士 人的领袖说：‘这人不可同我们上战场。’
1SAM|29|10|现在，你和跟随你来的，就是你主人的仆人，清晨要早早起来，回到我所指派你的地方去，不要把中伤的话放在心上，因为你在我面前很好 。你们清晨早早起来，天一亮就回去吧！”
1SAM|29|11|于是 大卫 和他的人清晨早早起来，回到 非利士 人的地去。 非利士 人也上 耶斯列 去了。
1SAM|30|1|第三日， 大卫 和他的人到了 洗革拉 。 亚玛力 人已经侵夺 尼革夫 和 洗革拉 。他们攻破 洗革拉 ，用火焚烧。
1SAM|30|2|他们掳去城内的妇女和城中的大小人口，一个都没有杀，全都带走，他们就上路去了。
1SAM|30|3|大卫 和他的人到了那城，看哪，城已被火烧毁，他们的妻子儿女都被掳去了。
1SAM|30|4|大卫 和跟随他的百姓就放声大哭，直到没有气力再哭。
1SAM|30|5|大卫 的两个妻子， 耶斯列 人 亚希暖 和作过 拿八 妻子的 迦密 人 亚比该 ，也被掳去了。
1SAM|30|6|大卫 非常焦急，因为众百姓为自己的儿女痛心，说要用石头打死他。 大卫 却倚靠耶和华－他的上帝，坚定自己。
1SAM|30|7|大卫 对 亚希米勒 的儿子 亚比亚他 祭司说：“请你把以弗得拿来给我。” 亚比亚他 就把以弗得拿给 大卫 。
1SAM|30|8|大卫 求问耶和华说：“我追赶这群人，是否追得上呢？”耶和华对他说：“你可以追，一定追得上，也一定救得回来。”
1SAM|30|9|于是， 大卫 出发，他和跟随他的六百人来到 比梭溪 ，那些不能前去的就留在那里。
1SAM|30|10|大卫 带着四百人往前追赶；有二百人疲乏，不能过 比梭溪 ，留在那里。
1SAM|30|11|这四百人在田野遇见一个 埃及 人，就带他到 大卫 面前，给他饼吃，给他水喝，
1SAM|30|12|又给他一块无花果饼，两个葡萄干饼。他吃了，精神就恢复了，因为他三日三夜没有吃饼，没有喝水。
1SAM|30|13|大卫 对他说：“你是谁的人？你从哪里来？”他说：“我是 埃及 的青年，是 亚玛力 人的奴仆。因为我三天前生病，我主人就把我撇弃了。
1SAM|30|14|我们侵夺了 基利提 的南方和属 犹大 的地，以及 迦勒 地的南方，又用火烧了 洗革拉 。”
1SAM|30|15|大卫 对他说：“你肯领我们下到那群人那里吗？”他说：“你要向我指着上帝起誓，你不杀我，也不把我交在我主人手里，我就领你下到那群人那里。”
1SAM|30|16|那人领 大卫 下去，看哪，他们分散在全地面，吃喝跳舞，因为他们从 非利士 人的地和 犹大 地掳来的财物非常多。
1SAM|30|17|大卫 击杀他们，从黎明直到次日晚上，除了四百个骑骆驼逃走的青年之外，一个也没有逃脱。
1SAM|30|18|亚玛力 人所掳去的财物， 大卫 全都夺回，并救回他的两个妻子。
1SAM|30|19|凡 亚玛力 人所掳去的，无论大小、儿女、掠物和一切被掳去的， 大卫 全都夺回来。
1SAM|30|20|大卫 所夺来的牛群羊群，有人赶在群畜前面，说：“这是 大卫 的掠物。”
1SAM|30|21|大卫 到了那疲乏不能跟随、留在 比梭溪 的二百人那里。他们出来迎接 大卫 和跟随他的百姓。 大卫 上前向他们问安。
1SAM|30|22|跟随 大卫 去的人中，每一个恶人和无赖都说：“这些人既然没有和我同去，我们所夺的财物就不分给他们，只把他们各人的妻子儿女给他们，让他们带回去就好了。”
1SAM|30|23|大卫 说：“我的弟兄，耶和华所赐给我们的，你们不可这么做，因为他保佑了我们，把那群来攻击我们的人交在我们手里。
1SAM|30|24|谁肯在这事上听你们呢？上阵的分得多少，留下看守物件的也分得多少，大家应当平分。”
1SAM|30|25|从那日起， 大卫 定此为 以色列 的律例典章，直到今日。
1SAM|30|26|大卫 到了 洗革拉 ，从掠物中取些送给他的朋友，就是 犹大 的长老，说：“看哪，这是从耶和华仇敌那里夺来的，送给你们作礼物。”
1SAM|30|27|有在 伯特利 的， 尼革夫 之 拉末 的， 雅提珥 的，
1SAM|30|28|有在 亚罗珥 的， 息末 的， 以实提莫 的，
1SAM|30|29|有在 拉哈勒 的， 耶拉篾 各城的， 基尼 各城的，
1SAM|30|30|有在 何珥玛 的， 坡拉珊 的， 亚挞 的，
1SAM|30|31|有在 希伯仑 的，以及 大卫 和跟随他的人经常进出之处的。
1SAM|31|1|非利士 人攻打 以色列 。 以色列 人在 非利士 人面前逃跑，很多人 在 基利波山 被杀仆倒。
1SAM|31|2|非利士 人紧追 扫罗 和他的儿子，杀了 扫罗 的儿子 约拿单 、 亚比拿达 、 麦基．舒亚 。
1SAM|31|3|攻击 扫罗 的战事激烈，弓箭手追上他，他被弓箭手射中，伤势很重 。
1SAM|31|4|扫罗 吩咐拿他兵器的人说：“你拔出刀来，把我刺死，免得那些未受割礼的人来刺我，凌辱我。”但拿兵器的人不肯，因为他非常惧怕。于是 扫罗 拿起刀来，伏在刀上。
1SAM|31|5|拿兵器的人见 扫罗 已死，也伏在刀上跟他一起死。
1SAM|31|6|这样， 扫罗 和他三个儿子，与拿他兵器的人，以及他所有的人 ，都在那日一起死了。
1SAM|31|7|住平原那边和 约旦河 那边的 以色列 人，见 以色列 军兵逃跑， 扫罗 和他儿子都死了，就弃城逃跑。 非利士 人前来住在其中。
1SAM|31|8|次日， 非利士 人来剥那些被杀之人的衣服，看见 扫罗 和他三个儿子仆倒在 基利波山 。
1SAM|31|9|他们割下他的首级，剥了他的盔甲，派人到 非利士 人之地的四境，报信给他们庙里的偶像和百姓。
1SAM|31|10|他们将 扫罗 的盔甲放在 亚斯她录 庙里，把他的尸身钉在 伯．珊 的城墙上。
1SAM|31|11|基列 的 雅比 居民听见 非利士 人向 扫罗 所行的事，
1SAM|31|12|他们所有的勇士就起身，走了一夜，把 扫罗 和他儿子的尸身从 伯．珊 城墙上取下来，送到 雅比 ，在那里用火烧了，
1SAM|31|13|把骸骨葬在 雅比 的柳树下，并且禁食七日。
2SAM|1|1|扫罗 死后， 大卫 击杀 亚玛力 人回来，在 洗革拉 住了两天。
2SAM|1|2|第三天，看哪，有一人从 扫罗 的营里出来，衣服撕裂，头蒙灰尘，到 大卫 面前伏地叩拜。
2SAM|1|3|大卫 对他说：“你从哪里来？”他说：“我从 以色列 的营里逃来。”
2SAM|1|4|大卫 又对他说：“事情怎么样？请你告诉我。”他说：“士兵从阵上逃跑，也有许多士兵仆倒死亡， 扫罗 和他儿子 约拿单 也死了。”
2SAM|1|5|大卫 问报信的青年说：“你怎么知道 扫罗 和他儿子 约拿单 死了呢？”
2SAM|1|6|报信的青年说：“我恰巧到 基利波山 ，看哪， 扫罗 靠在自己的枪上，看哪，有战车、骑兵紧紧地追他。
2SAM|1|7|他回头看见我，就呼叫我。我说：‘我在这里。’
2SAM|1|8|他问我说：‘你是什么人？’我说：‘我是 亚玛力 人。’
2SAM|1|9|他对我说：‘请你站到我这里来，把我杀死，因为我非常痛苦，只剩下一口气。’
2SAM|1|10|我就站到他那里，杀了他，因为我知道他一倒下就活不了。然后，我把他头上的冠冕和臂上的镯子拿到我主这里来。”
2SAM|1|11|大卫 就抓着自己的衣服，把衣服撕裂，所有跟随他的人也都如此。
2SAM|1|12|他们为 扫罗 和他儿子 约拿单 ，以及耶和华的百姓和 以色列 家的人悲哀哭泣，禁食到晚上，因为他们都倒在刀下。
2SAM|1|13|大卫 问报信的青年说：“你是哪里人？”他说：“我是一个寄居者的儿子，是 亚玛力 人。”
2SAM|1|14|大卫 对他说：“你动手杀害耶和华的受膏者，怎么不畏惧呢？”
2SAM|1|15|大卫 叫了一个仆人来，说：“来，杀了他！”仆人击杀他，他就死了。
2SAM|1|16|大卫 对他说：“你的血归到你自己头上，因为你亲口作证控诉自己，说：‘我杀了耶和华的受膏者。’”
2SAM|1|17|大卫 作了这首哀歌，哀悼 扫罗 和他儿子 约拿单 ，
2SAM|1|18|并吩咐人把这首“弓歌”教导 犹大 人，看哪，它写在《雅煞珥书》上：
2SAM|1|19|以色列 啊，尊荣者在你的高处被杀！ 大英雄竟然仆倒！
2SAM|1|20|不要在 迦特 报告， 不要在 亚实基伦 街上传扬， 免得 非利士 的女子欢喜， 免得未受割礼之人的女子欢乐。
2SAM|1|21|基利波山 哪，愿你那里没有雨，没有露！ 愿你的田地无土产可作供物！ 因为英雄的盾牌在那里受辱， 扫罗 的盾牌没有抹油。
2SAM|1|22|在被杀者的血前， 在勇士的脂肪前， 约拿单 的弓绝不退缩， 扫罗 的刀断不虚回。
2SAM|1|23|扫罗 和 约拿单 生时相悦相爱， 死时也不分离。 他们比鹰更快， 比狮子还强。
2SAM|1|24|以色列 的女子啊，当为 扫罗 哭泣！ 他曾使你们穿朱红色的美衣， 使你们衣服有黄金的妆饰。
2SAM|1|25|英雄竟然在阵上仆倒！ 约拿单 竟然在你的高处被杀！
2SAM|1|26|我兄 约拿单 哪，我为你悲伤！ 我甚喜爱你！ 你对我的爱何等奇妙， 过于妇女的爱情。
2SAM|1|27|英雄竟然仆倒！ 兵器竟然废弃！
2SAM|2|1|此后， 大卫 求问耶和华说：“我可以上 犹大 的一个城去吗？”耶和华对他说：“可以上去。” 大卫 说：“我上哪一个城去呢？”耶和华说：“ 希伯仑 。”
2SAM|2|2|于是 大卫 和他的两个妻子，一个是 耶斯列 人 亚希暖 ，一个是作过 迦密 人 拿八 妻子的 亚比该 ，都上那里去了。
2SAM|2|3|大卫 也把跟随他的人和他们各人的眷属一同带上去，住在 希伯仑 的城镇中。
2SAM|2|4|犹大 人来，在那里膏 大卫 作 犹大 家的王。 有人告诉 大卫 说：“埋葬 扫罗 的是 基列 的 雅比 人。”
2SAM|2|5|大卫 就派使者到 基列 的 雅比 人那里，对他们说：“愿耶和华赐福给你们！因为你们忠心对待你们的主 扫罗 ，埋葬了他。
2SAM|2|6|你们既做了这事，愿耶和华以慈爱和信实待你们，我也要为此厚待你们。
2SAM|2|7|现在，你们的主 扫罗 死了， 犹大 家也已经膏我作他们的王，你们的手要坚强，要作英勇的人。”
2SAM|2|8|扫罗 军队的元帅， 尼珥 的儿子 押尼珥 ，曾将 扫罗 的儿子 伊施．波设 带过河，到 玛哈念 ，
2SAM|2|9|立他作王，治理 基列 、 亚书利 、 耶斯列 、 以法莲 、 便雅悯 和 以色列 众人。
2SAM|2|10|扫罗 的儿子 伊施．波设 登基的时候年四十岁，作 以色列 王二年，但是 犹大 家却随从 大卫 。
2SAM|2|11|大卫 在 希伯仑 作 犹大 家的王，共七年六个月。
2SAM|2|12|尼珥 的儿子 押尼珥 和 扫罗 的儿子 伊施．波设 的仆人从 玛哈念 出来，往 基遍 去。
2SAM|2|13|洗鲁雅 的儿子 约押 和 大卫 的仆人也出来，在 基遍 池旁与他们相遇；一队坐在池的这边，一队坐在池的那边。
2SAM|2|14|押尼珥 对 约押 说：“让年轻人起来，在我们面前较量一下吧！” 约押 说：“让他们起来吧。”
2SAM|2|15|他们就起来，点了人数过来：属 扫罗 儿子 伊施．波设 的有 便雅悯 人十二名， 大卫 的仆人也有十二名。
2SAM|2|16|每人抓住对方的头，用刀刺对方的肋旁，一同仆倒。所以，那地叫做 希利甲．哈素林 ，就在 基遍 。
2SAM|2|17|那日战况激烈， 押尼珥 和 以色列 人败在 大卫 的仆人面前。
2SAM|2|18|在那里有 洗鲁雅 的三个儿子： 约押 、 亚比筛 、 亚撒黑 。 亚撒黑 的脚快如野地里的羚羊；
2SAM|2|19|亚撒黑 追赶 押尼珥 ，直追赶他不偏左右。
2SAM|2|20|押尼珥 回头说：“ 亚撒黑 ，是你吗？”他说：“是我。”
2SAM|2|21|押尼珥 对他说：“你转左或转右，去抓一个年轻人，剥去他的战衣吧。” 亚撒黑 却不肯转开而不追赶他。
2SAM|2|22|押尼珥 又对 亚撒黑 说：“转开，不要再追我了！我何必把你击杀在地上呢？我若杀了你，怎么有脸见你哥哥 约押 呢？”
2SAM|2|23|亚撒黑 仍不肯转开， 押尼珥 就用回马枪 刺入他的肚腹，甚至枪从背后穿出， 亚撒黑 就仆倒在那里，当场死了。众人赶到 亚撒黑 仆倒而死的地方，就都站住。
2SAM|2|24|约押 和 亚比筛 追赶 押尼珥 。日落的时候，他们到了通往 基遍 旷野的路旁， 基亚 对面的 亚玛山 。
2SAM|2|25|便雅悯 人聚集在 押尼珥 后面，成为一队，站在一座山顶上。
2SAM|2|26|押尼珥 呼叫 约押 说：“刀剑岂可永远吞噬呢？你岂不知，结局必是痛苦的吗？你要等到何时才叫百姓回去，不追赶他们的弟兄呢？”
2SAM|2|27|约押 说：“我指着永生的上帝起誓：你若没有这么说，百姓就必继续追赶弟兄，直到早晨 。”
2SAM|2|28|于是 约押 吹角，众百姓就站住，不再追赶 以色列 人，也不再打仗了。
2SAM|2|29|押尼珥 和他的人整夜行过 亚拉巴 。他们过了 约旦河 ，走过 毕伦 ，到了 玛哈念 。
2SAM|2|30|约押 追赶 押尼珥 回来，聚集众百姓， 大卫 的仆人中缺少了十九个人和 亚撒黑 。
2SAM|2|31|但 大卫 的仆人杀了 押尼珥 的人， 便雅悯 人三百六十名。
2SAM|2|32|他们把 亚撒黑 送到 伯利恒 ，葬在他父亲的坟墓里。 约押 和他的人走了一整夜，天亮的时候他们才到 希伯仑 。
2SAM|3|1|扫罗 家和 大卫 家争战许久。 大卫 家日见强盛， 扫罗 家却日见衰弱。
2SAM|3|2|大卫 在 希伯仑 生了几个儿子：长子 暗嫩 是 耶斯列 人 亚希暖 所生的；
2SAM|3|3|次子 基利押 是作过 迦密 人 拿八 的妻子 亚比该 所生的；三子 押沙龙 是 基述 王 达买 的女儿 玛迦 所生的；
2SAM|3|4|四子 亚多尼雅 是 哈及 所生的；五子 示法提雅 是 亚比她 所生的；
2SAM|3|5|六子 以特念 是 大卫 的妻子 以格拉 所生的。 大卫 这六个儿子都是在 希伯仑 生的。
2SAM|3|6|扫罗 家和 大卫 家争战的时候， 押尼珥 在 扫罗 家大有权势。
2SAM|3|7|扫罗 有一妃子，名叫 利斯巴 ，是 爱亚 的女儿。一日， 伊施．波设 对 押尼珥 说：“你为什么与我父的妃子同寝呢？”
2SAM|3|8|押尼珥 因 伊施．波设 的话非常生气，说：“我岂是狗的头，向着 犹大 呢？我今日忠心对待你父 扫罗 的家和他的弟兄、朋友，不将你交在 大卫 手里，今日你竟为这妇人责备我吗？
2SAM|3|9|愿上帝重重惩罚 押尼珥 ！我要照着耶和华起誓应许 大卫 的话为他成就，
2SAM|3|10|废去 扫罗 家的国度，建立 大卫 的王位，使他治理 以色列 和 犹大 ，从 但 直到 别是巴 。”
2SAM|3|11|伊施．波设 惧怕 押尼珥 ，一句话也不能回答。
2SAM|3|12|押尼珥 派使者到 大卫 所在的地方 ，说：“这地归谁呢？”又说：“你与我立约，看哪，我必帮助你，使全 以色列 都拥护你。”
2SAM|3|13|大卫 说：“好！我与你立约。但有一件事我要求你，你来见我面的时候，除非把 扫罗 的女儿 米甲 带来，就不必来见我的面了。”
2SAM|3|14|大卫 派使者到 扫罗 的儿子 伊施．波设 那里，说：“你要把我的妻子 米甲 归还我；她是我从前用一百 非利士 人的包皮所聘定的。”
2SAM|3|15|伊施．波设 就派人去，把 米甲 从 拉亿 的儿子，她丈夫 帕铁 那里带来。
2SAM|3|16|米甲 的丈夫跟着她，一面走一面哭，直跟到 巴户琳 。 押尼珥 对他说：“你回去吧！” 帕铁 就回去了。
2SAM|3|17|押尼珥 与 以色列 长老商议，说：“从前你们企盼 大卫 作王治理你们，
2SAM|3|18|现在你们可以这样做了。因为耶和华曾论到 大卫 说：‘我必藉我仆人 大卫 的手，救我民 以色列 脱离 非利士 人和众仇敌的手。’”
2SAM|3|19|押尼珥 也说给 便雅悯 人听。 押尼珥 又到 希伯仑 ，把 以色列 人和 便雅悯 全家所看为好的，说给 大卫 听。
2SAM|3|20|押尼珥 带着二十个人来到 希伯仑大卫 那里， 大卫 就为 押尼珥 和他带来的人摆设宴席。
2SAM|3|21|押尼珥 对 大卫 说：“我要起身去召集全 以色列 ，来到我主我王这里，与你立约，你就可以照你的心愿作王，统治一切。”于是 大卫 送走 押尼珥 ，他就平安地去了。
2SAM|3|22|看哪， 大卫 的仆人和 约押 突击回来，带回许多掠物。那时 押尼珥 不在 希伯仑大卫 那里，因 大卫 已经送他走，他也平安地去了。
2SAM|3|23|约押 和跟随他的全军到了，有人告诉 约押 说：“ 尼珥 的儿子 押尼珥 来到王这里，王送走他，他也平安地去了。”
2SAM|3|24|约押 到王那里，说：“你这是做什么呢？看哪， 押尼珥 来到你这里，你为何送他走，让他去了呢？
2SAM|3|25|你知道， 尼珥 的儿子 押尼珥 来，是要骗你，要打听你的出入，知道你一切所行的事。”
2SAM|3|26|约押 从 大卫 那里出来，派些使者去追 押尼珥 ，从 西拉井 那里带他回来， 大卫 却不知道。
2SAM|3|27|押尼珥 回到 希伯仑 ， 约押 领他到城门中间，要与他私下交谈，就在那里刺穿了他的肚腹。他就死了，因为他流了 约押 兄弟 亚撒黑 的血。
2SAM|3|28|这事以后， 大卫 听见了，说：“流 尼珥 儿子 押尼珥 的血，我和我的国在耶和华面前永远是无辜的。
2SAM|3|29|愿这血归到 约押 头上和他父的全家；又愿 约押 家不断有患漏症的，长痲疯 的，架柺杖而行的 ，仆倒在刀下的，缺乏食物的。”
2SAM|3|30|约押 和他弟弟 亚比筛 杀了 押尼珥 ，是因为在 基遍 战争的时候， 押尼珥 杀了他们的弟弟 亚撒黑 。
2SAM|3|31|大卫 对 约押 和跟随他的众百姓说：“你们当撕裂衣服，腰束麻布，在 押尼珥 前面哀哭。” 大卫 王也跟在棺木后面。
2SAM|3|32|他们把 押尼珥 葬在 希伯仑 。王在 押尼珥 的墓旁放声大哭，众百姓也都哭了。
2SAM|3|33|王为 押尼珥 举哀，说： 押尼珥 怎么会像愚顽人一样地死呢？
2SAM|3|34|你手未曾被捆绑，脚未曾被脚镣锁住。 你仆倒，如仆倒在凶恶之子手下一样。 于是众百姓又为 押尼珥 哀哭。
2SAM|3|35|白天的时候，众百姓来劝 大卫 吃饭，但 大卫 起誓说：“我若在太阳未下山以前吃饭，或吃任何东西，愿上帝重重惩罚我！”
2SAM|3|36|众百姓知道了就看为好。凡王所做的，众百姓都看为好。
2SAM|3|37|那日， 以色列 众百姓才知道杀 尼珥 的儿子 押尼珥 并非出于王意。
2SAM|3|38|王对臣仆说：“你们岂不知今日在 以色列 中倒了一个作元帅的大人物吗？
2SAM|3|39|我虽然受膏为王，今日还是软弱。 洗鲁雅 的两个儿子，这些人比我强硬。愿耶和华照着恶人所行的恶报应他。”
2SAM|4|1|扫罗 的儿子 伊施．波设 听见 押尼珥 死在 希伯仑 ，手就发软，全 以色列 也都惊惶。
2SAM|4|2|扫罗 的儿子 伊施．波设 有两个军官，一个叫 巴拿 ，第二个叫 利甲 ，都是 便雅悯 支派 比录 人 临门 的儿子；因为 比录 也算是属于 便雅悯 的。
2SAM|4|3|比录 人先前逃到 基他音 ，在那里寄居，直到今日。
2SAM|4|4|扫罗 的儿子 约拿单 有一个儿子，名叫 米非波设 ，是瘸腿的。 扫罗 和 约拿单 的消息从 耶斯列 传来的时候，他才五岁。他的奶妈抱着他逃跑；因为跑得太急，孩子掉在地上，腿就瘸了。
2SAM|4|5|比录 人 临门 的两个儿子 利甲 和 巴拿 出去，天正热的时候到了 伊施．波设 的家。那时， 伊施．波设 在睡午觉。
2SAM|4|6|妇人进到房子中间，要取麦子。 利甲 和他的哥哥 巴拿 刺穿了 伊施．波设 的肚腹，然后逃跑了。
2SAM|4|7|他们进到房子的时候， 伊施．波设 正躺在卧房的床上，他们就把他杀死，割了他的首级，拿着首级在 亚拉巴 的路上走了一整夜。
2SAM|4|8|他们把 伊施．波设 的首级拿到 希伯仑 大卫 那里，对王说：“王的仇敌 扫罗 曾寻索你的性命。看哪，这是他儿子 伊施．波设 的首级；耶和华今日为我主我王在 扫罗 和他后裔身上报了仇。”
2SAM|4|9|大卫 回答 比录 人 临门 的儿子 利甲 和他哥哥 巴拿 说：“我指着救我性命脱离一切苦难、永生的耶和华起誓：
2SAM|4|10|从前有人告诉我说：‘看哪， 扫罗 死了。’他自以为报好消息，我就拿住他，把他杀在 洗革拉 ，作为他报消息的赏赐。
2SAM|4|11|更何况恶人把义人杀在他家的床上，我岂不从你们手中追讨他的血，从地上除灭你们吗？”
2SAM|4|12|于是 大卫 吩咐仆人把他们杀了，砍断他们的手脚，挂在 希伯仑 的池旁。然后，他们把 伊施．波设 的首级葬在 希伯仑押尼珥 的坟墓里。
2SAM|5|1|以色列 众支派来到 希伯仑 见 大卫 ，说：“看哪，我们是你的骨肉。
2SAM|5|2|从前 扫罗 作我们王的时候，率领 以色列 人出入的是你。耶和华也曾对你说：‘你必牧养我的百姓 以色列 ，你必作 以色列 的君王。’”
2SAM|5|3|于是 以色列 的众长老都来到 希伯仑 见王 。 大卫 在 希伯仑 ，在耶和华面前与他们立约，他们就膏 大卫 作 以色列 的王。
2SAM|5|4|大卫 登基的时候年三十岁，作王四十年。
2SAM|5|5|他在 希伯仑 作 犹大 王七年六个月，在 耶路撒冷 作 以色列 和 犹大 王三十三年。
2SAM|5|6|王和他的人到了 耶路撒冷 ，要攻打住那地方的 耶布斯 人。 耶布斯 人对 大卫 说：“你必不能进到这里，就是盲人、瘸子都可以把你击退。”就是说：“ 大卫 绝不能进到这里。”
2SAM|5|7|然而 大卫 攻取了 锡安 的堡垒，就是 大卫 的城。
2SAM|5|8|当日， 大卫 说：“谁攻打 耶布斯 人，就要从水道上去，攻打我心里所恨恶的 瘸子、盲人。”因此有人说：“盲人和瘸子不得进殿里去。”
2SAM|5|9|大卫 住在堡垒里，给它起名叫 大卫城 。 大卫 又从 米罗 往内，周围建筑。
2SAM|5|10|大卫 日见强大，耶和华－万军之上帝与他同在。
2SAM|5|11|推罗 王 希兰 派使者把香柏木运到 大卫 那里，又派木匠和石匠给 大卫 建造宫殿。
2SAM|5|12|大卫 知道耶和华坚立他作 以色列 王，又为自己百姓 以色列 的缘故，使他的国兴盛。
2SAM|5|13|大卫 离开 希伯仑 之后，在 耶路撒冷 又立后妃，又生儿女。
2SAM|5|14|在 耶路撒冷 所生的孩子的名字是 沙母亚 、 朔罢 、 拿单 、 所罗门 、
2SAM|5|15|益辖 、 以利书亚 、 尼斐 、 雅非亚 、
2SAM|5|16|以利沙玛 、 以利雅大 、 以利法列 。
2SAM|5|17|非利士 人听见 大卫 受膏作 以色列 王， 非利士 众人就上来寻索 大卫 。 大卫 听见了，就下到堡垒去。
2SAM|5|18|非利士 人来了，散布在 利乏音谷 。
2SAM|5|19|大卫 求问耶和华说：“我可以上去攻打 非利士 人吗？你将他们交在我手里吗？”耶和华对 大卫 说：“你可以上去，我必将 非利士 人交在你手里。”
2SAM|5|20|大卫 来到 巴力．毗拉心 ，在那里击败了 非利士 人。他说：“耶和华在我面前冲破敌人，如水冲破一样。”因此他称那地方为 巴力．毗拉心 。
2SAM|5|21|非利士 人把偶像抛弃在那里， 大卫 和他的人拿去了。
2SAM|5|22|非利士 人又上来，散布在 利乏音谷 。
2SAM|5|23|大卫 求问耶和华；耶和华说：“不要直上，要绕到他们后头，从桑树林对面攻打他们。
2SAM|5|24|你听见桑树梢上有脚步的声音，就要急速前去，因为那时耶和华已经出去，在你前头攻打 非利士 人的军队了。”
2SAM|5|25|大卫 就遵照耶和华所吩咐的去做，攻打 非利士 人，从 迦巴 直到 基色 。
2SAM|6|1|大卫 又聚集 以色列 中所有挑选的人，共三万名。
2SAM|6|2|大卫 起身，和跟随他的众百姓前往，要从 巴拉．犹大 那里将上帝的约柜接上来；这约柜是以坐在二基路伯上万军之耶和华的名所命名的。
2SAM|6|3|他们将上帝的约柜从山冈上 亚比拿达 的家里抬出来，放在新车上； 亚比拿达 的儿子 乌撒 和 亚希约 赶这新车。
2SAM|6|4|他们将上帝的约柜从山冈上 亚比拿达 家里抬出来 ， 亚希约 在约柜前行走。
2SAM|6|5|大卫 和 以色列 全家在耶和华面前，随着松木制造的各样乐器 和琴、瑟、鼓、钹、锣跳舞。
2SAM|6|6|到了 拿艮 的禾场，因为牛失前蹄 ， 乌撒 就伸手扶住上帝的约柜。
2SAM|6|7|耶和华的怒气向 乌撒 发作；上帝因这冒犯在那里击打他，他就死在那里，在上帝的约柜旁。
2SAM|6|8|大卫 因耶和华突然冲出撞死 乌撒 就生气，称那地方为 毗列斯．乌撒 ，直到今日。
2SAM|6|9|那日， 大卫 惧怕耶和华，说：“耶和华的约柜怎可到我这里来呢？”
2SAM|6|10|于是 大卫 不愿将耶和华的约柜接进 大卫城 他自己的地方，却转送到 迦特 人 俄别．以东 的家中。
2SAM|6|11|耶和华的约柜停在 迦特 人 俄别．以东 家中三个月，耶和华赐福给 俄别．以东 和他的全家。
2SAM|6|12|有人告诉 大卫 王说：“耶和华因约柜的缘故赐福给 俄别．以东 的家和一切属他的。” 大卫 就去，欢欢喜喜地将上帝的约柜从 俄别．以东 家中接上来，到 大卫城 里。
2SAM|6|13|抬耶和华约柜的人走了六步， 大卫 就献牛与肥畜为祭。
2SAM|6|14|大卫 穿着细麻布以弗得，在耶和华面前极力跳舞。
2SAM|6|15|这样， 大卫 和 以色列 全家欢呼吹角，将耶和华的约柜接了上来。
2SAM|6|16|耶和华的约柜进 大卫城 的时候， 扫罗 的女儿 米甲 从窗户里往外观看，见 大卫 王在耶和华面前踊跃跳舞，心里就轻视他。
2SAM|6|17|众人将耶和华的约柜请进去，安放在所预备的地方，就是 大卫 为它搭的帐幕中。 大卫 在耶和华面前献燔祭和平安祭。
2SAM|6|18|大卫 献完了燔祭和平安祭，就奉万军之耶和华的名祝福百姓，
2SAM|6|19|并且分给 以色列 众人，所有的百姓，无论男女，每人一个饼，一个枣子饼 ，一个葡萄饼。众人就各自回家去了。
2SAM|6|20|大卫 回去要为家里的人祝福， 扫罗 的女儿 米甲 出来迎接他，说：“ 以色列 王今日有好大的荣耀啊！他今日在臣仆的使女眼前露体，如同一个无赖赤身露体一样，”
2SAM|6|21|大卫 对 米甲 说：“这是在耶和华面前的。耶和华已拣选我，在你父和你父的全家之上，立我作耶和华百姓 以色列 的君王，所以我在耶和华面前跳舞，
2SAM|6|22|我也必更加卑微，自己看为低贱 。至于你所说的那些使女，她们反而尊重我。”
2SAM|6|23|扫罗 的女儿 米甲 ，直到死的那日没有孩子。
2SAM|7|1|王住在自己宫中，耶和华使他平静，不被四围的仇敌扰乱。
2SAM|7|2|王对 拿单 先知说：“你看，我住在香柏木的宫中，上帝的约柜却停在幔子里。”
2SAM|7|3|拿单 对王说：“你可以完全照你的心意去做，因为耶和华与你同在。”
2SAM|7|4|当夜耶和华的话临到 拿单 ，说：
2SAM|7|5|“你去对我仆人 大卫 说：‘耶和华如此说：你要建造殿宇给我居住吗？
2SAM|7|6|自从我领 以色列 人从 埃及 上来，直到今日，我未曾住过殿宇，却在会幕和帐幕中行走。
2SAM|7|7|凡我同 以色列 人所走的地方，我何曾向 以色列 任何一个领袖 ，就是我吩咐牧养我百姓 以色列 的，说过这话：你们为何不给我建造香柏木的殿宇呢？’
2SAM|7|8|现在，你要对我仆人 大卫这样 说：‘万军之耶和华如此说：我从羊圈中将你召来，叫你不再牧放羊群，立你作我百姓 以色列 的君王。
2SAM|7|9|你无论往哪里去，我都与你同在，剪除你所有的仇敌。我必使你得大名，好像世上伟人的名一样。
2SAM|7|10|我必为我百姓 以色列 选定一个地方，栽植他们，使他们住自己的地方，不再受搅扰；凶恶之子也不像从前那样苦待他们，
2SAM|7|11|并不像我命令士师治理我百姓 以色列 的日子。我必使你平静，不受任何仇敌搅扰，并且耶和华应许你，耶和华必为你建立家室。
2SAM|7|12|当你寿数满足、与你祖先同睡的时候，我必使你身所生的后裔接续你；我也必坚定他的国。
2SAM|7|13|他必为我的名建造殿宇，我必坚定他国度的王位，直到永远。
2SAM|7|14|我要作他的父，他要作我的子；他若犯了罪，我必用人的杖，用世人的鞭责罚他。
2SAM|7|15|但我的慈爱仍不离开他，像离开在你面前所废的 扫罗 一样。
2SAM|7|16|你的家和你的国必在你 面前永远坚立，你的王位也必坚定，直到永远。’”
2SAM|7|17|拿单 就按这一切话，照这一切异象告诉 大卫 。
2SAM|7|18|于是 大卫 王进去，坐在耶和华面前，说：“主耶和华啊，我是谁，我的家算什么，你竟带领我到这地步呢？
2SAM|7|19|主耶和华啊，这在你眼中还看为小，你又说到你仆人的家将来的情况。主耶和华啊，这岂是人的常理吗？
2SAM|7|20|大卫 还有什么可以对你说呢？主耶和华啊，你是知道你仆人的。
2SAM|7|21|你行这一切大事，使你的仆人明白，是因你应许的缘故，也照着你的心意。
2SAM|7|22|因此，主耶和华啊，你本为大；照我们耳中一切所听见的，没有可比你的，除你以外再没有上帝。
2SAM|7|23|谁像你的百姓 以色列 呢？上帝亲自去救赎世上的一国 ，作自己的子民，显出他的大名；为了你的地，从列国和他们的神明中，在你亲自从埃及赎出来的子民面前，为自己行了大而可畏的事 。
2SAM|7|24|你曾坚立你的百姓 以色列 作你的子民，直到永远；你－耶和华也作他们的上帝。
2SAM|7|25|现在，耶和华上帝啊，你所应许仆人和仆人家的话，求你坚定，直到永远；求你照你所说的而行。
2SAM|7|26|愿人永远尊你的名为大，说：‘万军之耶和华是治理 以色列 的上帝。’这样，你仆人 大卫 的家必在你面前坚立。
2SAM|7|27|万军之耶和华－ 以色列 的上帝啊，因你启示你的仆人说：‘我必为你建立家室’，所以仆人大胆向你如此祈祷。
2SAM|7|28|现在，主耶和华啊，惟有你是上帝！你的话是真实的，你也应许将这福气赐给仆人。
2SAM|7|29|现在，求你赐福给你仆人的家，可以永存在你面前。主耶和华啊，因为这是你所应许的。愿你的福分永远赐给你仆人的家，使之蒙福！”
2SAM|8|1|此后， 大卫 攻打 非利士 人，制伏了他们。 大卫 从 非利士 人手中夺取了京城的治理权 。
2SAM|8|2|他又攻打 摩押 人，使他们躺卧在地上，用绳来量，量二绳的杀了，量一绳的活着。 摩押 人就臣服 大卫 ，向他进贡。
2SAM|8|3|利合 的儿子 琐巴 王 哈大底谢 往 幼发拉底河 去，要夺回他的国权， 大卫 就攻打他，
2SAM|8|4|俘掳了他的骑兵一千七百人，步兵二万人。 大卫 把所有战马的蹄筋砍断，只留下一百辆战车。
2SAM|8|5|大马士革 的 亚兰 人来帮助 琐巴 王 哈大底谢 ， 大卫 杀了 亚兰 人二万二千。
2SAM|8|6|于是 大卫 在 大马士革 的 亚兰 设立军营， 亚兰 人就臣服 大卫 ，向他进贡。 大卫 无论往哪里去，耶和华都使他得胜。
2SAM|8|7|大卫夺了 哈大底谢 臣仆拥有的金盾牌，带到 耶路撒冷 。
2SAM|8|8|大卫 王又从 哈大底谢 的 比他 和 比罗他 二城夺取了许多的铜。
2SAM|8|9|哈马 王 陀以 听见 大卫 击败 哈大底谢 的全军，
2SAM|8|10|就派他儿子 约兰 到 大卫 王那里，向他请安，为他祝福，因他与 哈大底谢 争战，并且击败了他；原来 哈大底谢 与 陀以 常常争战。 约兰 手里带了金银铜的器皿来。
2SAM|8|11|大卫 王把这些器皿分别为圣，连同他制伏各国所分别为圣的金银，献给耶和华，
2SAM|8|12|就是从 亚兰 、 摩押 、 亚扪 人、 非利士 人、 亚玛力 人，以及从 利合 的儿子 琐巴 王 哈大底谢 所掠之物。
2SAM|8|13|大卫 得了名声。当他回来的时候，在 盐谷 击杀了一万八千 以东 人。
2SAM|8|14|大卫 在 以东 设立军营；他在全 以东 设立军营， 以东 人就都臣服他。 大卫 无论往哪里去，耶和华都使他得胜。
2SAM|8|15|大卫 作全 以色列 的王，又向众百姓秉公行义。
2SAM|8|16|洗鲁雅 的儿子 约押 作元帅； 亚希律 的儿子 约沙法 作史官；
2SAM|8|17|亚希突 的儿子 撒督 和 亚比亚他 的儿子 亚希米勒 作祭司； 西莱雅 作书记；
2SAM|8|18|耶何耶大 的儿子 比拿雅 管辖 基利提 人和 比利提 人。 大卫 的众子都作祭司。
2SAM|9|1|大卫 说：“ 扫罗 家还有剩下的人没有？我要因 约拿单 的缘故向他施恩。”
2SAM|9|2|扫罗 家有一个仆人名叫 洗巴 ，有人叫他来到 大卫 那里。王对他说：“你是 洗巴 吗？”他说：“仆人是。”
2SAM|9|3|王说：“ 扫罗 家还有没有剩下的人？我要照上帝的慈爱恩待他。” 洗巴 对王说：“还有 约拿单 的一个儿子，双腿是瘸的。”
2SAM|9|4|王对他说：“他在哪里？” 洗巴 对王说：“看哪，他在 罗．底巴 ， 亚米利 的儿子 玛吉 家里。”
2SAM|9|5|于是 大卫 王派人去，从 罗．底巴 ， 亚米利 的儿子 玛吉 家里召了他来。
2SAM|9|6|扫罗 的孙子， 约拿单 的儿子 米非波设 来到 大卫 那里，脸伏于地叩拜。 大卫 说：“ 米非波设 ！” 米非波设 说：“看哪，仆人在此。”
2SAM|9|7|大卫 对他说：“你不要惧怕，我必因你父亲 约拿单 的缘故向你施恩，把你祖父 扫罗 的一切田地都归还你，你也可以常与我同席吃饭。”
2SAM|9|8|米非波设 叩拜，说：“你的仆人算什么，不过如死狗一般，竟蒙你这样眷顾！”
2SAM|9|9|王召了 扫罗 的仆人 洗巴 来，对他说：“我已把属 扫罗 和他的一切家产都赐给你主人的儿子了。
2SAM|9|10|你，你的众子和仆人要为你主人的儿子耕种田地，把所收获的拿来供他食用；你主人的儿子 米非波设 却要常与我同席吃饭。” 洗巴 有十五个儿子和二十个仆人。
2SAM|9|11|洗巴 对王说：“凡我主我王吩咐仆人的，仆人都必遵行。”于是 米非波设 与王 同席吃饭，如王的儿子一样。
2SAM|9|12|米非波设 有一个小儿子，名叫 米迦 。凡住在 洗巴 家里的人都作了 米非波设 的仆人。
2SAM|9|13|米非波设 住在 耶路撒冷 ，常与王同席吃饭。他两腿都是瘸的。
2SAM|10|1|此后， 亚扪 人的王死了，他儿子 哈嫩 接续他作王。
2SAM|10|2|大卫 说：“ 哈嫩 的父亲 拿辖 怎样向我施恩，我也要怎样向 哈嫩 施恩。”于是 大卫 派臣仆为他的父亲安慰他。当 大卫 的臣仆到了 亚扪 人的境内，
2SAM|10|3|亚扪 人的领袖对他们的主 哈嫩 说：“ 大卫 派人来安慰你，你看他是要尊敬你父亲吗？ 大卫 派臣仆到你这里，不是为了要窥探侦察，而倾覆这城吗？”
2SAM|10|4|哈嫩 就抓住 大卫 的臣仆，把他们的胡须剃去一半，又割断他们下半截的袍子，露出下体，然后放了他们。
2SAM|10|5|有人告诉 大卫 ，他就派人去迎接他们，因为这些人觉得很羞耻。王说：“可以住在 耶利哥 ，等到胡须长出来再回来。”
2SAM|10|6|亚扪 人看到 大卫 憎恶他们，就派人去雇用 伯．利合 的 亚兰 人和 琐巴 的 亚兰 人，步兵二万，以及 玛迦 王的人一千、 陀伯 人一万二千。
2SAM|10|7|大卫 听见了，就派 约押 和所有勇猛的军队出去。
2SAM|10|8|亚扪 人出来，在城门前摆阵； 琐巴 与 利合 的 亚兰 人、 陀伯 人，以及 玛迦 人另外在郊野摆阵。
2SAM|10|9|约押 看见战阵对着他前后摆列，就把从 以色列 所有精兵中挑选出来的，摆阵迎战 亚兰 人。
2SAM|10|10|他把其余的兵交在他兄弟 亚比筛 手里， 亚比筛 就摆阵迎战 亚扪 人。
2SAM|10|11|约押 对 亚比筛说：“ 亚兰 人若强过我，你就来帮助我； 亚扪 人若强过你，我就去帮助你。
2SAM|10|12|你要刚强，我们要为自己的百姓，为我们上帝的城镇奋勇。愿耶和华照他所看为好的去做！”
2SAM|10|13|于是， 约押 和跟随他的士兵前进攻打 亚兰 人； 亚兰 人在他面前逃跑。
2SAM|10|14|亚扪 人见 亚兰 人逃跑，他们也在 亚比筛 面前逃跑进城。 约押 就离开 亚扪 人，回 耶路撒冷 去了。
2SAM|10|15|亚兰 人见自己被 以色列 打败，就集合起来。
2SAM|10|16|哈大底谢 派人去，把 大河 那边的 亚兰 人调来；他们到了 希兰 ，由 哈大底谢 的将军 朔法 在他们前面率领。
2SAM|10|17|有人告诉 大卫 ，他就聚集 以色列 众人过 约旦河 ，来到 希兰 。 亚兰 人迎着 大卫 摆阵，与他打仗。
2SAM|10|18|亚兰 人在 以色列 人面前逃跑。 大卫 杀了 亚兰 七百辆战车的士兵，四万骑兵 ，又击杀 亚兰 的将军 朔法 ，他就死在那里。
2SAM|10|19|哈大底谢 属下的诸王见自己被 以色列 打败，就与 以色列 讲和，臣服他们。于是 亚兰 人害怕，不再帮助 亚扪 人了。
2SAM|11|1|过了一年，正是诸王出战的时候， 大卫 派 约押 率领臣仆和 以色列 众人出去。他们打败 亚扪 人，围攻 拉巴 。 大卫 仍然留在 耶路撒冷 。
2SAM|11|2|黄昏的时候， 大卫 从床上起来，在王宫的平顶上散步。他从平顶上看见一个妇人沐浴，这妇人容貌非常美丽。
2SAM|11|3|大卫 派人打听那妇人是谁。有人说：“她不是 以连 的女儿， 赫 人 乌利亚 的妻子 拔示巴 吗？”
2SAM|11|4|大卫 派使者去把妇人接来；她来到大卫那里，那时她的月经刚洁净， 大卫 与她同寝。她就回家去了。
2SAM|11|5|那妇人怀了孕，派人去告诉 大卫 说：“我怀孕了。”
2SAM|11|6|大卫 派人告诉 约押 ：“你派 赫 人 乌利亚 到我这里来。” 约押 就派 乌利亚 到 大卫 那里。
2SAM|11|7|乌利亚 来到 大卫那里， 大卫 问 约押 好，也问士兵好，又问战争的情况。
2SAM|11|8|大卫 对 乌利亚 说：“下到你家去，洗洗脚吧！” 乌利亚 出了王宫，随后王送他一份礼物。
2SAM|11|9|乌利亚 却和他主人所有的仆人一同睡在王宫门口，没有下到他家去。
2SAM|11|10|有人告诉 大卫 说：“ 乌利亚 没有下到他的家。” 大卫 就对 乌利亚 说：“你不是从远路上来吗？为什么不下到你家去呢？”
2SAM|11|11|乌利亚 对 大卫 说：“约柜， 以色列 和 犹大 都留在棚里，我主 约押 和我主的仆人都在田野安营，我岂可回家吃喝，与妻子同房呢？我指着王和王的性命起誓：‘我绝不做这事！’”
2SAM|11|12|大卫 对 乌利亚 说：“你今日仍留在这里，明日我打发你去。”于是 乌利亚 那日留在 耶路撒冷 。次日，
2SAM|11|13|大卫 召了 乌利亚 来，叫他在自己面前吃喝，使他喝醉。黄昏的时候， 乌利亚 出去，躺卧在自己的床上；与他主的仆人在一起，并没有下到他的家去。
2SAM|11|14|早晨， 大卫 写信给 约押 ，交 乌利亚 亲手带去。
2SAM|11|15|他在信内写着说：“要派 乌利亚 到战争激烈的前线去，然后你们撤退离开他，使他被击杀而死。”
2SAM|11|16|约押 侦察城的时候，知道敌人哪里有勇士，就派 乌利亚 到那地方。
2SAM|11|17|城里的人出来和 约押 打仗， 大卫 的仆人中有几个士兵被杀， 赫 人 乌利亚 也死了。
2SAM|11|18|于是， 约押 派人去将战争的一切事奏告 大卫 ，
2SAM|11|19|又吩咐使者说：“你把战争的一切事对王说完了，
2SAM|11|20|王若发怒，对你说：‘你们打仗为什么挨近城呢？岂不知敌人会从城墙上射箭吗？
2SAM|11|21|从前击杀 耶路比设 的儿子 亚比米勒 的是谁呢？岂不是一个妇人从城墙上抛下一块上磨石来，打在他身上，他就死在 提备斯 吗？你们为什么挨近城墙呢？’你就说：‘你的仆人 赫 人 乌利亚 也死了。’”
2SAM|11|22|使者就去，照着 约押 所吩咐的一切话来奏告 大卫 。
2SAM|11|23|使者对 大卫 说：“敌人强过我们，出到郊外攻打我们，我们把他们赶回到城门口。
2SAM|11|24|弓箭手从城墙上射你的仆人，射死几个王的仆人，你的仆人 赫 人 乌利亚 也死了。”
2SAM|11|25|大卫 向使者说：“你对 约押 这样说：‘不要为这事难过，因为刀剑可能吞灭这人或那人。你只管竭力攻城，将城倾覆。’你要勉励 约押 。”
2SAM|11|26|乌利亚 的妻听见丈夫 乌利亚 死了，就为丈夫哀哭。
2SAM|11|27|居丧的日子过了， 大卫 派人把她接到宫里，她就作了 大卫 的妻子，给 大卫 生了一个儿子。但 大卫 做的这事，耶和华的眼中看为恶。
2SAM|12|1|耶和华差遣 拿单 到 大卫 那里。 拿单 到了他那里，对他说：“在一座城里有两个人，一个是富翁，一个是穷人。
2SAM|12|2|富翁有极多的牛群羊群；
2SAM|12|3|穷人除了所买来养活的一只小母羊之外，一无所有。小羊在他家里和他儿女一同长大，吃他所吃的，喝他所喝的，睡在他怀中，在他看来如同女儿一样。
2SAM|12|4|有一客人来到这富翁那里，富翁舍不得从自己的牛群羊群中取一只招待来到他那里的旅客，却取了穷人的小母羊，招待来到他那里的人。”
2SAM|12|5|大卫 就非常恼怒那人，对 拿单 说：“我指着永生的耶和华起誓，做这事的人该死！
2SAM|12|6|他必须偿还小母羊四倍，因为他做这事，没有怜悯的心。”
2SAM|12|7|拿单 对 大卫 说：“你就是那人！耶和华－ 以色列 的上帝如此说：‘我膏你作 以色列 的王，我救你脱离 扫罗 的手；
2SAM|12|8|我将你主人的家业赐给你，将你主人的妃嫔交在你怀里，又将 以色列 和 犹大 家赐给你；若还嫌少，我也会如此这般加倍赐给你。
2SAM|12|9|你为什么藐视耶和华的命令，做他眼中看为恶的事呢？你用刀击杀 赫 人 乌利亚 ，又娶了他的妻子为妻，借 亚扪 人的刀杀死他。
2SAM|12|10|现在刀剑必永不离开你的家，因你藐视我，娶了 赫 人 乌利亚 的妻子为妻。’
2SAM|12|11|耶和华如此说：‘看哪，我必从你家中兴起灾祸攻击你；我必在你眼前把你的妃嫔赐给你身边的人，他要在光天化日下与你的妃嫔同寝。
2SAM|12|12|你在暗中做那事，我却要在 以色列 众人面前，在日光之下做这事。’”
2SAM|12|13|大卫 对 拿单 说：“我得罪耶和华了！” 拿单 说：“耶和华已经除去你的罪，你必不至于死。
2SAM|12|14|只是在这事上，你大大藐视耶和华 ，因此，你生的孩子必定要死。”
2SAM|12|15|拿单 就回家去了。 耶和华击打 乌利亚 的妻子为 大卫 生的孩子，他就得了重病。
2SAM|12|16|大卫 为这孩子恳求上帝。 大卫 刻苦禁食，到里面去，躺在地上过夜。
2SAM|12|17|他家中的老臣来到他旁边，要把他从地上扶起来，他却不肯，也不同他们吃饭。
2SAM|12|18|到第七日，孩子死了。 大卫 的臣仆不敢告诉他孩子死了，因他们说：“看哪，孩子还活着的时候，我们劝他，他尚且不听我们的话，我们怎么能告诉他孩子死了，让他做出不好的事呢？”
2SAM|12|19|大卫 见臣仆彼此低声说话，就知道孩子死了。他问臣仆说：“孩子死了吗？”他们说：“死了。”
2SAM|12|20|大卫 就从地上起来，沐浴，抹膏，换了衣服，进耶和华的殿敬拜。然后他回宫，吩咐人为他摆饭，他就吃了。
2SAM|12|21|臣仆对他说：“你所做的是什么事呢？孩子活着的时候，你为他禁食哭泣；孩子死了，你却起来吃饭。”
2SAM|12|22|大卫 说：“孩子还活着，我禁食哭泣，因为我想，或许耶和华怜悯我，会让孩子活下来。
2SAM|12|23|现在孩子死了，我何必禁食呢？我能使他回来吗？我必往他那里去，他却不能回到我这里来。”
2SAM|12|24|大卫 安慰他的妻子 拔示巴 ，与她同房，她就生了儿子，给他起名叫 所罗门 。耶和华喜爱他，
2SAM|12|25|就藉 拿单 先知赐他一个名字，叫 耶底底亚 ；这是为了耶和华的缘故。
2SAM|12|26|约押 攻打 亚扪 人的 拉巴 ，攻占了京城。
2SAM|12|27|约押 派使者到 大卫 那里，说：“我攻打 拉巴 ， 也攻占了水城。
2SAM|12|28|现在你要召集其余的军兵，安营围攻这城，攻占它，免得我攻占这城，人就以我的名叫这城。”
2SAM|12|29|于是 大卫 召集全军，往 拉巴 去攻城，就攻占了它。
2SAM|12|30|他也夺了 米勒公 头上所戴的冠冕，其上的金子重一他连得，又嵌着宝石。这冠冕就戴在 大卫 头上。 大卫 又从城里夺了许多财物，
2SAM|12|31|把城里的百姓拉出来，叫他们用锯，用铁耙，用铁斧做工，派他们在砖窑中服役； 大卫 待 亚扪 各城的居民都是如此。于是， 大卫 和全军都回 耶路撒冷 去了。
2SAM|13|1|后来发生了一件事。 大卫 的儿子 押沙龙 有一个美貌的妹妹，名叫 她玛 。 大卫 的儿子 暗嫩 爱上了她。
2SAM|13|2|暗嫩 为他妹妹 她玛 苦恋成疾，因为 她玛 还是处女， 暗嫩 眼看难以向她行事。
2SAM|13|3|暗嫩 有一个密友，名叫 约拿达 ，是 大卫 长兄 示米亚 的儿子。这 约拿达 为人极其狡猾。
2SAM|13|4|他对 暗嫩 说：“王的儿子啊，你何不告诉我，为何你一天比一天憔悴呢？” 暗嫩 对他说：“我爱上了我兄弟 押沙龙 的妹妹 她玛 。”
2SAM|13|5|约拿达 对他说：“你躺在床上装病，等你父亲来看你，就对他说：‘请让我妹妹 她玛 来，给我东西吃，在我眼前预备食物，使我可以看见，好从她手里接过来吃。’”
2SAM|13|6|于是 暗嫩 躺着装病，王来看他。 暗嫩 对王说：“请让我妹妹 她玛 来，在我眼前为我做两个饼，我好从她手里接过来吃。”
2SAM|13|7|大卫 就派人去宫里，到 她玛 那里，说：“你到你哥哥 暗嫩 的屋里去，为他预备食物。”
2SAM|13|8|她玛 就到她哥哥 暗嫩 的屋里，那时 暗嫩 正躺着。 她玛 拿了面团揉面，在他眼前做饼，把饼烤熟了。
2SAM|13|9|她玛 拿了锅子，在他面前把饼倒出来，他却不肯吃。 暗嫩 说：“每一个人都离开我，出去吧！”众人就都离开他，出去了。
2SAM|13|10|暗嫩 对 她玛 说：“你把食物拿进卧房，我好从你手里接过来吃。” 她玛 就把所做的饼拿进卧房，到她哥哥 暗嫩 那里。
2SAM|13|11|她玛 上前去给他吃，他就拉住 她玛 ，对她说：“我妹妹，你来与我同寝。”
2SAM|13|12|她玛 对他说：“哥哥，不可以！不要玷辱我！ 以色列 中不可以这样做，你不要做这丑事！
2SAM|13|13|我蒙受耻辱，该往那里去呢？至于你，你在 以色列 中也成了一个愚顽人。现在你可以求王，他必不禁止我归你。”
2SAM|13|14|但 暗嫩 不肯听她的话，因他比她更有力，就玷辱她，与她同寝。
2SAM|13|15|随后， 暗嫩 极其恨她，恨她的心比先前爱她的心更甚，就对她说：“你起来，去吧！”
2SAM|13|16|她玛 对 暗嫩 说：“不要这样！你赶我出去的这恶比你刚才向我所做的更严重！”但 暗嫩 不肯听她，
2SAM|13|17|就叫伺候自己的仆人来，说：“把这女子从我这里赶出去！她一出去，你就闩上门。”
2SAM|13|18|那时 她玛 穿着彩衣，因为没有出嫁的公主都穿这样的外袍。 暗嫩 的仆人把她赶出去，她一出去，仆人就闩上门。
2SAM|13|19|她玛 把灰尘撒在头上，撕裂所穿的彩衣，以手抱头，一面走一面哭喊。
2SAM|13|20|她胞兄 押沙龙 对她说：“你哥哥 暗嫩 与你亲近了吗？妹妹，现在暂且不要作声，他是你的哥哥，不要把这事放在心上。” 她玛 就孤孤单单地住在她胞兄 押沙龙 的家里。
2SAM|13|21|大卫 王听见这一切的事，就非常愤怒。
2SAM|13|22|押沙龙 却不和 暗嫩 说好说歹；因为 暗嫩 玷辱他妹妹 她玛 ，所以 押沙龙 恨恶他。
2SAM|13|23|过了二年，有人在靠近 以法莲 的 巴力．夏琐 为 押沙龙 剪羊毛。 押沙龙 请了王所有的儿子来。
2SAM|13|24|押沙龙 来到王那里，说：“看哪，有人正为你的仆人剪羊毛，请王和王的臣仆与你的仆人同去。”
2SAM|13|25|王对 押沙龙 说：“不，我儿，我们不必都去，免得成了你的负担。” 押沙龙 再三请王，王仍是不肯去，只为他祝福。
2SAM|13|26|押沙龙 说：“王若不去，请让我哥哥 暗嫩 与我们同去。”王对他说：“为何要他与你同去呢？”
2SAM|13|27|押沙龙 再三求王，王就派 暗嫩 和王所有的儿子与他同去。
2SAM|13|28|押沙龙 吩咐仆人说：“你们注意， 暗嫩 开怀畅饮的时候，我对你们说击杀 暗嫩 ，你们就杀他。不要惧怕，这不是我吩咐你们的吗？你们要刚强，作勇士！”
2SAM|13|29|押沙龙 的仆人就照 押沙龙 所吩咐的，向 暗嫩 行了。王所有的儿子都起来，各人骑上骡子逃跑了。
2SAM|13|30|他们还在路上，就有风声传到 大卫 那里，说：“ 押沙龙 击杀了王所有的儿子，没有留下一个。”
2SAM|13|31|王就起来，撕裂衣服，躺在地上。王的臣仆全都撕裂衣服，站在旁边。
2SAM|13|32|大卫 的长兄 示米亚 的儿子 约拿达 说：“我主，不要以为他们把所有的年轻人，就是王的儿子都杀了，只有 暗嫩 一个人死了。自从 暗嫩 玷辱了 押沙龙 的妹妹 她玛 那日， 押沙龙 已经决定这事了。
2SAM|13|33|现在，我主我王，不要把这事放在心上，以为王所有的儿子都死了。其实，只有 暗嫩 一人死了。”
2SAM|13|34|押沙龙 逃跑了。守望的年轻人举目观看，看哪，有许多人从 何罗念 山坡的路上来。
2SAM|13|35|约拿达 对王说：“看哪，王的儿子都来了，正如你仆人所说的，事情就这样发生了。”
2SAM|13|36|话刚说完，看哪，王的儿子都到了，放声大哭。王和他的众臣仆也都号啕痛哭。
2SAM|13|37|押沙龙 逃到 亚米忽 的儿子 基述 王 达买 那里去了。 大卫 天天为他儿子悲哀。
2SAM|13|38|押沙龙 逃到 基述 去了，在那里住了三年。
2SAM|13|39|王想要出去对付 押沙龙 的心化解了 ，因为王对 暗嫩 之死这事已经得了安慰。
2SAM|14|1|洗鲁雅 的儿子 约押 知道王心里想念 押沙龙 。
2SAM|14|2|他派人往 提哥亚 去，从那里叫了一个有智慧的妇人来，对她说：“请你装作居丧的人，穿上丧服，不用膏抹身，装作为死者悲哀多日的妇人。
2SAM|14|3|你到王那里，对王如此如此说。”于是 约押 把当说的话放在她口中。
2SAM|14|4|提哥亚 妇人到王面前 ，脸伏于地叩拜，说：“王啊，求你拯救！”
2SAM|14|5|王对她说：“你有什么事呢？”她说：“我实在是个寡妇，我丈夫死了。
2SAM|14|6|婢女有两个儿子，二人在田间打架，没有人从中劝解，一个击杀另一个，把他打死了。
2SAM|14|7|看哪，全家族都起来攻击婢女，说：‘把那打死兄弟的交出来，我们好处死他，为他所打死的兄弟偿命，灭绝那承受家业的。’这样，他们要把我剩下的炭火灭尽，不给我丈夫留名或留后在地面上。”
2SAM|14|8|王对妇人说：“你回家去吧！我必为你下个命令。”
2SAM|14|9|提哥亚 妇人又对王说：“我主我王，愿这罪孽归我和我的父家，与王和王的位无关。”
2SAM|14|10|王说：“有人说话难为你，你就带他到我这里来，他必不再搅扰你。”
2SAM|14|11|妇人说：“愿王对耶和华－你的上帝发誓，不许报血仇的人施行毁灭，免得他们灭绝我的儿子。”王说：“我指着永生的耶和华起誓：你的儿子连一根头发也不致落在地上。”
2SAM|14|12|妇人说：“求我主我王容许婢女再说一句话。”王说：“你说吧！”
2SAM|14|13|妇人说：“王为何起意做这事，要害上帝的百姓呢？王不使那逃亡的人回来，王说这话就证实自己错了！
2SAM|14|14|我们都必死，如同水泼在地上，不能收回。上帝不会让人不死，但仍设法 使逃亡的人不致成为赶出、回不来的人。
2SAM|14|15|现在我来将这话告诉我主我王，是因百姓使我惧怕。婢女想：‘不如告诉王，或者王会成就使女所求的。
2SAM|14|16|人要把我和我儿子从上帝的地业上一同除灭，王必应允救使女脱离他的手。’
2SAM|14|17|婢女想：‘我主我王的话必安慰我’；因为我主我王能辨别是非，如同上帝的使者一样。惟愿耶和华－你的上帝与你同在！”
2SAM|14|18|王回答妇人说：“我问你一句话，你一点也不可瞒我。”妇人说：“我主我王，请说。”
2SAM|14|19|王说：“这一切莫非是 约押 的手指使你的吗？”妇人回答说：“我敢在我主我王面前起誓：我主我王所说的一切不偏左右，这是王的仆人 约押 吩咐我的，这一切话是他放在婢女口中的。
2SAM|14|20|王的仆人 约押 做这事，为要扭转局面。我主的智慧却如上帝使者的智慧，能知地上一切的事。”
2SAM|14|21|王对 约押 说：“看哪，我应允这事。你去，把那年轻人 押沙龙 带回来。”
2SAM|14|22|约押 脸伏于地叩拜，为王祝福，说：“王既应允仆人这件事，仆人今日知道在我主我王眼前蒙恩宠了。”
2SAM|14|23|于是 约押 起身往 基述 去，把 押沙龙 带回 耶路撒冷 。
2SAM|14|24|王说：“让他回自己的家去，不要来见我的面。” 押沙龙 就回自己的家去，没有见王的面。
2SAM|14|25|全 以色列 中，无人像 押沙龙 那样俊美，得人称赞，从脚底到头顶毫无瑕疵。
2SAM|14|26|他的头发很重，每到年底剪发一次，所剪下来的，按王的秤称一称，重二百舍客勒。
2SAM|14|27|押沙龙 生了三个儿子，一个女儿。女儿名叫 她玛 ，是个容貌美丽的女子。
2SAM|14|28|押沙龙 住在 耶路撒冷 ，足足有二年没有见王的面。
2SAM|14|29|押沙龙 派人去叫 约押 来，要托他到王那里去， 约押 却不肯来。 押沙龙 第二次派人去叫他，他仍不肯来。
2SAM|14|30|于是 押沙龙 对仆人说：“你们看， 约押 有一块田靠近我的田，其中有大麦，你们去放火把它烧了。” 押沙龙 的仆人就去放火烧了那田。
2SAM|14|31|于是 约押 起来，到了 押沙龙 家里，对他说：“你的仆人为何放火烧我的田呢？”
2SAM|14|32|押沙龙 对 约押 说：“看哪，我派人去请你来，好托你到王那里去，说：‘我为何从 基述 回来呢？我仍在那里比较好。’现在让我去见王的面；我若有罪孽，就任凭王杀了我吧。”
2SAM|14|33|于是 约押 到王那里，奏告王，王就叫 押沙龙 来。 押沙龙 到王那里，在王面前脸伏于地，王就亲吻 押沙龙 。
2SAM|15|1|此后， 押沙龙 为自己预备车马，又派五十人在他前头奔跑。
2SAM|15|2|押沙龙 常常早晨起来，站在城门的路旁，任何人有争讼要去求王判决， 押沙龙 就叫他过来，说：“你是哪一城的人？”他说：“仆人是 以色列 某支派的人。”
2SAM|15|3|押沙龙 就对他说：“看，你的案件合情合理，无奈王没有委派人听你申诉。”
2SAM|15|4|押沙龙 又说：“恨不得我作这地的审判官！ 凡有争讼的人可以到我这里来，我必秉公判断。”
2SAM|15|5|若有人近前来要拜 押沙龙 ， 押沙龙 就伸手拉住他，亲吻他。
2SAM|15|6|以色列 中，凡到王那里求判决的， 押沙龙 都这么做。这样， 押沙龙 暗中赢得了 以色列 人的心。
2SAM|15|7|过了四年 ， 押沙龙 对王说：“求你准我往 希伯仑 去，还我向耶和华所许的愿。
2SAM|15|8|因为仆人住在 亚兰 的 基述 时，曾许愿说：‘耶和华若使我再回 耶路撒冷 ，我必事奉他 。’”
2SAM|15|9|王对他说：“你平安地去吧！” 押沙龙 就动身，往 希伯仑 去了。
2SAM|15|10|押沙龙 派密使走遍 以色列 各支派，说：“你们一听见角声就说：‘ 押沙龙 在 希伯仑 作王了！’”
2SAM|15|11|押沙龙 在 耶路撒冷 请了二百人与他同去，都是诚心诚意去的，一点也不知道实情。
2SAM|15|12|押沙龙 献祭的时候，派人去把 大卫 的谋士， 基罗 人 亚希多弗 从他本城 基罗 请来 。于是叛乱越发强大，因为随从 押沙龙 的百姓日渐增多。
2SAM|15|13|报信的人来到 大卫 那里，说：“ 以色列 人的心都归向 押沙龙 了！”
2SAM|15|14|大卫 就对 耶路撒冷 所有跟随他的臣仆说：“起来，我们逃吧！否则，我们来不及逃避 押沙龙 。要快点离开，免得他很快追上我们，加害于我们，用刀击杀城里的人。”
2SAM|15|15|王的臣仆对王说：“我主我王所决定的一切，看哪，仆人都愿遵行。”
2SAM|15|16|于是王出去了，他的全家都跟随他，但留下十个妃嫔看守宫殿。
2SAM|15|17|王出去，众百姓都跟随他；到了最后一座屋子 ，他们就停下来。
2SAM|15|18|王的众臣仆都在他旁边过去。 基利提 人、 比利提 人，和从 迦特 跟随王来的六百个 迦特 人，也都在王面前过去。
2SAM|15|19|王对 迦特 人 以太 说：“你是外邦人，从你本地逃来的，为什么与我们同去呢？你回去留在新王那里吧！
2SAM|15|20|你昨天才到，我今日怎好叫你与我们一同流亡，而我却要到处飘流呢？回去吧，你带你的弟兄回去吧！愿主用慈爱信实待你 。”
2SAM|15|21|以太 回答王说：“我指着永生的耶和华起誓，又敢在王面前起誓：无论生死，王在哪里，你的仆人也必在哪里。”
2SAM|15|22|大卫 对 以太 说：“去，过去吧！”于是 迦特 人 以太 带着所有跟随他的人和孩子过去了。
2SAM|15|23|众百姓过去时，当地的人全都放声大哭。王过了 汲沦溪 ，众百姓就往旷野的路上去了。
2SAM|15|24|看哪， 撒督 和所有抬上帝约柜的 利未 人也一同来了。他们将上帝的约柜放下， 亚比亚他 上来 ，直到众百姓从城里出来走过去为止。
2SAM|15|25|王对 撒督 说：“你将上帝的约柜请回城去。我若在耶和华眼前蒙恩，他必使我回来，再见到约柜和他的居所。
2SAM|15|26|倘若他说：‘我不喜爱你’；我在这里，就照他眼中看为好的待我！”
2SAM|15|27|王对 撒督 祭司说：“你不是先见吗？你可以平安地回城，你儿子 亚希玛斯 和 亚比亚他 的儿子 约拿单 ，你们二人的儿子可以与你们同去。
2SAM|15|28|看，我在旷野的渡口那里等，直到你们来报信给我。”
2SAM|15|29|于是 撒督 和 亚比亚他 将上帝的约柜请回 耶路撒冷 ，他们就留在那里。
2SAM|15|30|大卫 蒙头赤脚走上 橄榄山 的斜坡，一面上一面哭。所有跟随他的百姓也都各自蒙头哭着上去；
2SAM|15|31|有人告诉 大卫 说 ：“ 亚希多弗 也在叛党之中，随从 押沙龙 。” 大卫 说：“耶和华啊，求你使 亚希多弗 的计谋变为愚拙！”
2SAM|15|32|大卫 到了山顶，敬拜上帝的地方，看哪， 亚基 人 户筛 衣服撕裂，头蒙灰尘来迎见他。
2SAM|15|33|大卫 对他说：“你若与我一同过去，必拖累我；
2SAM|15|34|你若回城去，对 押沙龙 说：‘王啊，我愿作你的仆人。我向来作你父亲的仆人，现在我也愿意作你的仆人。’你就可以为我破坏 亚希多弗 的计谋。
2SAM|15|35|撒督 和 亚比亚他 二位祭司岂不都在你那里吗？你在王宫里听见什么，就要告诉 撒督 和 亚比亚他 二位祭司。
2SAM|15|36|看哪， 撒督 的儿子 亚希玛斯 ， 亚比亚他 的儿子 约拿单 ，也跟二位祭司在那里。凡你们所听见的事，可以托这二人来向我报告。”
2SAM|15|37|于是， 大卫 的朋友 户筛 进了城， 押沙龙 也进了 耶路撒冷 。
2SAM|16|1|大卫 刚过山顶，看哪， 米非波设 的仆人 洗巴 拉着装好鞍子的两匹驴，驴上驮着二百个面饼，一百个葡萄饼，一百个夏天的果饼，一皮袋酒来迎接他。
2SAM|16|2|王对 洗巴 说：“你的这些东西是什么意思呢？” 洗巴 说：“驴是给王的家眷骑的，面饼和夏天的果饼是给年轻人吃的，酒是给在旷野疲乏的人喝的。”
2SAM|16|3|王说：“你主人的儿子在哪里呢？” 洗巴 对王说：“看哪，他留在 耶路撒冷 ，因他说：‘ 以色列 家今日必将我父的国归还我。’”
2SAM|16|4|王对 洗巴 说：“看哪，凡属 米非波设 的都是你的了。” 洗巴 说：“我叩拜我主我王，愿我在你眼前蒙恩宠。”
2SAM|16|5|大卫 王到了 巴户琳 ，看哪，有一个人从那里出来，是 扫罗 家族中 基拉 的儿子，名叫 示每 。他一面走一面咒骂，
2SAM|16|6|又向 大卫 王和王的众臣仆扔石头；众百姓和勇士都在王的左右。
2SAM|16|7|示每 这样咒骂说：“你这好流人血的，你这无赖，滚吧！滚吧！
2SAM|16|8|你流了 扫罗 全家的血，接续他作王，耶和华把这罪归在你身上。耶和华将这国交在你儿子 押沙龙 的手中。看哪，你咎由自取，因为你是好流人血的人。”
2SAM|16|9|洗鲁雅 的儿子 亚比筛 对王说：“这死狗为何咒骂我主我王呢？让我过去，割下他的头来。”
2SAM|16|10|王说：“ 洗鲁雅 的儿子，我与你们有何相干呢？他这样咒骂是因耶和华吩咐他：‘你要咒骂 大卫 。’如此，谁敢说：‘你为什么这样做呢？’”
2SAM|16|11|大卫 又对 亚比筛 和众臣仆说：“看哪，我亲生的儿子尚且寻索我的性命，何况现在这 便雅悯 人呢？由他咒骂吧！因为这是耶和华吩咐他的。
2SAM|16|12|或者耶和华见我遭难 ，因我今日被这人咒骂而向我施恩。”
2SAM|16|13|于是 大卫 和他的人在路上走。 示每 走在 大卫 对面的山坡，一面走一面咒骂，又向他扔石头，扬起尘土。
2SAM|16|14|王和跟随他的众百姓来了，非常疲乏，就在那里歇息。
2SAM|16|15|押沙龙 和 以色列 众百姓来到 耶路撒冷 ， 亚希多弗 也与他同来。
2SAM|16|16|大卫 的朋友 亚基 人 户筛 来到 押沙龙 那里，对他说：“愿王万岁！愿王万岁！”
2SAM|16|17|押沙龙 对 户筛 说：“你这样做是忠诚对待你的朋友吗？为什么不与你的朋友同去呢？”
2SAM|16|18|户筛 对 押沙龙 说：“不，谁是耶和华和这百姓，以及 以色列 众人所拣选的，我必归顺他，留在他那里。
2SAM|16|19|再者，我当服事谁呢？岂不是前王的儿子吗？我怎样服事你父亲，也必照样服事你。”
2SAM|16|20|押沙龙 对 亚希多弗 说：“你们出个主意，我们该怎么做？”
2SAM|16|21|亚希多弗 对 押沙龙 说：“你父亲所留下看守宫殿的妃嫔，你可以与她们亲近。 以色列 众人听见你敢惹你父亲憎恶你，凡归顺你人的手就更坚强了。”
2SAM|16|22|于是他们为 押沙龙 在屋顶上支搭帐棚， 押沙龙 就在 以色列 众人眼前，与他父亲的妃嫔亲近。
2SAM|16|23|那时 亚希多弗 所出的主意好像人从上帝求问得来的话一样；他给 大卫 ，给 押沙龙 所出的一切主意，都是这样。
2SAM|17|1|亚希多弗 对 押沙龙 说：“请让我挑选一万二千人，今夜起身追赶 大卫 。
2SAM|17|2|我必趁他疲乏手软的时候追上他，使他惊惶。跟随他的众百姓必都逃跑，我就只杀王一个人。
2SAM|17|3|我必使众百姓都归顺你，正如众人归顺你所追杀的人一样 ，众百姓就都平安无事了。”
2SAM|17|4|这话在 押沙龙 和 以色列 众长老的眼中都看为好。
2SAM|17|5|押沙龙 说：“把 亚基 人 户筛 也召来，我们也要听他怎么说。”
2SAM|17|6|户筛 到了 押沙龙 那里， 押沙龙 向他说：“ 亚希多弗 说了这样的话，我们要照他的话做吗？若不可，你就说吧！”
2SAM|17|7|户筛 对 押沙龙 说：“ 亚希多弗 这次所出的主意不好。”
2SAM|17|8|户筛 又说：“你知道，你父亲和他的人都是勇士，他们心里恼怒，如同田野中失去小熊的母熊一样；而且你父亲是个战士，必不和百姓一同住宿。
2SAM|17|9|看哪，他现今或藏在一个坑中或在别处，若我们 有人首先被杀，听见的必说：‘跟随 押沙龙 的百姓被杀了。’
2SAM|17|10|虽有勇士胆大如狮子，他的心也必定融化，因为全 以色列 都知道你父亲是英雄，跟随他的人都是勇士。
2SAM|17|11|依我之计，要把如同海边的沙那样多的 以色列 众人，从 但 直到 别是巴 ，聚集到你这里来，由你亲自率领他们出战。
2SAM|17|12|我们到他那里，在任何地方遇见他，就突然临到他，如同露水滴在泥土上。这样，他和所有跟随他的人，一个也不留。
2SAM|17|13|他若撤退到一座城， 以色列 众人必带绳子去那城，把城拉到河里，甚至连一块小石子也找不到。”
2SAM|17|14|押沙龙 和 以色列 众人都说：“ 亚基 人 户筛 的计谋比 亚希多弗 的更好！”这是因为耶和华定意破坏 亚希多弗 的良谋，为的是耶和华要降祸给 押沙龙 。
2SAM|17|15|户筛 对 撒督 和 亚比亚他 二位祭司说：“ 亚希多弗 为 押沙龙 和 以色列 的长老出的主意是如此如此，我出的主意是如此如此。
2SAM|17|16|现在你们要急速派人去告诉 大卫 说：‘今夜不可在旷野的渡口住宿，务要过河，免得王和所有跟随他的百姓都被吞灭。’”
2SAM|17|17|约拿单 和 亚希玛斯 在 隐．罗结 等候，不敢进城，恐怕被人看见。有一个婢女出来，把这话告诉他们，他们就去报信给 大卫 王。
2SAM|17|18|然而有一个僮仆看见他们，就去告诉 押沙龙 。他们二人急忙离开，跑到 巴户琳 一个人的家里。那人院中有一口井，他们就下到那里。
2SAM|17|19|那家的妇人用盖盖上井口，又在上头铺上碎麦，事情就没有泄漏。
2SAM|17|20|押沙龙 的仆人来到妇人的家，说：“ 亚希玛斯 和 约拿单 在哪里？”妇人对他们说：“他们过了河了。”仆人搜寻，却找不着，就回 耶路撒冷 去了。
2SAM|17|21|他们走后，二人从井里上来，去告诉 大卫 王。他们对 大卫 说：“ 亚希多弗 出这样的主意要害你，你们起来，快快过河。”
2SAM|17|22|于是 大卫 和所有跟随他的百姓都起来，过 约旦河 。到了天亮，无一人不过 约旦河 的。
2SAM|17|23|亚希多弗 见他的计谋不被接纳，就备上驴，动身归回本城，到了自己的家。他留下遗嘱给他的家，就上吊死了，葬在他父亲的坟墓里。
2SAM|17|24|大卫 到了 玛哈念 ， 押沙龙 和跟随他的 以色列 众人也都过了 约旦河 。
2SAM|17|25|押沙龙 立 亚玛撒 作元帅，取代 约押 。 亚玛撒 是 以实玛利 人 以特拉 的儿子。 以特拉 曾与 拿辖 的女儿 亚比该 亲近；这 亚比该 与 约押 的母亲 洗鲁雅 是姊妹。
2SAM|17|26|押沙龙 和 以色列 人安营在 基列 地。
2SAM|17|27|大卫 到了 玛哈念 ， 亚扪 族的 拉巴 人 拿辖 的儿子 朔比 ， 罗．底巴 人 亚米利 的儿子 玛吉 ，来自 罗基琳 的 基列 人 巴西莱 ，
2SAM|17|28|带着被褥、盆、瓦器，还有小麦、大麦、麦面、烤熟的谷穗、豆子、红豆、炒豆、
2SAM|17|29|蜂蜜、奶油、绵羊、奶饼，供给 大卫 和跟随他的人吃，因为他们想：“百姓在旷野中，必定又饥渴又疲乏。”
2SAM|18|1|大卫 数点跟随他的百姓，立千夫长、百夫长率领他们。
2SAM|18|2|大卫 把军兵分为三队 ：三分之一在 约押 手下，三分之一在 洗鲁雅 的儿子 约押 弟弟 亚比筛 手下，三分之一在 迦特 人 以太 手下。王对军兵说：“我必与你们一同出战。”
2SAM|18|3|军兵却说：“你不可出战。若是我们逃跑，敌人不会把心放在我们身上；我们阵亡一半，敌人也不会把心放在我们身上。但现在你一人抵过我们万人，所以你最好留在城里支援我们。”
2SAM|18|4|王对他们说：“你们看怎样好，我就怎样做。”于是王站在城门旁，所有的军兵成百成千地挨次出战去了。
2SAM|18|5|王嘱咐 约押 、 亚比筛 、 以太 说：“你们要为我的缘故宽待那年轻人 押沙龙 。”王为 押沙龙 的事嘱咐众将领的话，所有的军兵都听见了。
2SAM|18|6|军兵出到田野迎战 以色列 ，在 以法莲 的树林里交战。
2SAM|18|7|在那里， 以色列 百姓败在 大卫 的臣仆面前。那日在那里阵亡的很多，共有二万人。
2SAM|18|8|战争蔓延到整个地面，那日被树林吞噬的军兵比被刀剑吞噬的更多。
2SAM|18|9|押沙龙 刚好遇见了 大卫 的臣仆。 押沙龙 骑着骡子，从大橡树密枝底下经过，他的头被橡树夹住，悬挂在空中 ，所骑的骡子就离他去了。
2SAM|18|10|有个人看见，就告诉 约押 说：“看哪，我看见 押沙龙 挂在橡树上了。”
2SAM|18|11|约押 对报信的人说：“看哪，你既看见了，为什么不当场把他击杀在地呢？我必赏你十个银子和一条带子。”
2SAM|18|12|那人对 约押 说：“即使我手里得了一千银子，也不敢伸手害王的儿子，因为我们听见王嘱咐你、 亚比筛 、 以太 说：‘你们要谨慎，不可害那年轻人 押沙龙 。’
2SAM|18|13|我若冒着生命危险做这傻事 ，无论何事都瞒不过王，你自己也必远远站在一旁。”
2SAM|18|14|约押 说：“我不能在你面前这样耗下去！” 约押 手拿三枝短枪，趁 押沙龙 在橡树上 还活着，就刺透他的心。
2SAM|18|15|给 约押 拿兵器的十个青年围着 押沙龙 ，击杀他，将他杀死。
2SAM|18|16|约押 吹角，军兵就回来，不去追赶 以色列 人，因为 约押 制止了军兵。
2SAM|18|17|他们拿下 押沙龙 ，把他丢在树林中一个大坑里，上头堆起一大堆石头。 以色列 众人都逃跑，各回自己的帐棚去了。
2SAM|18|18|押沙龙 活着的时候，曾在 王谷 立了一根柱子，因他说：“我没有儿子为我留名。”他就以自己的名字称那柱子为 押沙龙碑 ，直到今日。
2SAM|18|19|撒督 的儿子 亚希玛斯 说：“让我跑去报信给王，耶和华已经为王伸冤，使他脱离仇敌的手了。”
2SAM|18|20|约押 对他说：“你今日不可作报信的人，改日再去报信；因为今日王的儿子死了，所以你不可去报信。”
2SAM|18|21|约押 对 古实 人说：“你去把你所看见的告诉王。” 古实 人向 约押 叩拜后，就跑去了。
2SAM|18|22|撒督 的儿子 亚希玛斯 又对 约押 说：“无论怎样，让我随着 古实 人跑去吧！” 约押 说：“我儿，你报这信息，既不得赏赐，何必要跑去呢？”
2SAM|18|23|他说：“无论怎样，我要跑去。” 约押 对他说：“你跑去吧！” 亚希玛斯 就从平原的路往前跑，越过了 古实 人。
2SAM|18|24|大卫 正坐在内外城门之间。守望的人上到城墙，在城门的顶上举目观看，看哪，有一个人独自跑来。
2SAM|18|25|守望的人就大声告诉王。王说：“他若独自来，必是报口信的。”那人跑得越来越近了。
2SAM|18|26|守望的人又见一人跑来，就对守城门的人喊说：“看哪，又有一人独自跑来。”王说：“这也是报信的。”
2SAM|18|27|守望的人说：“我看前面那人的跑法，好像 撒督 的儿子 亚希玛斯 的跑法。”王说：“他是个好人，是来报好消息的。”
2SAM|18|28|亚希玛斯 向王呼叫说：“平安了！”他就脸伏于地向王叩拜，说：“耶和华－你的上帝是应当称颂的，他已把些那举手攻击我主我王的人交出来了。”
2SAM|18|29|王说：“年轻人 押沙龙 平安吗？” 亚希玛斯 说：“ 约押 派王的仆人，就是你的仆人时，我看见一阵大骚动，却不知道是什么事。”
2SAM|18|30|王说：“你退去，站在这里。”他就退去，站着。
2SAM|18|31|看哪， 古实 人也来到，说：“有信息报给我主我王！耶和华今日为你伸冤，使你脱离一切起来攻击你之人的手。”
2SAM|18|32|王对 古实 人说：“年轻人 押沙龙 平安吗？” 古实 人说：“愿我主我王的仇敌，和一切起来恶意要害你的人，都像那年轻人一样。”
2SAM|18|33|王战抖，就上城门的楼房去痛哭，一面走一面说：“我儿 押沙龙 啊！我儿，我儿 押沙龙 啊！我恨不得替你死， 押沙龙 啊，我儿！我儿！”
2SAM|19|1|有人告诉 约押 ：“看哪，王为 押沙龙 悲哀哭泣。”
2SAM|19|2|那日众军兵听说王为他儿子悲伤，他们得胜的日子变成悲哀了。
2SAM|19|3|那日军兵暗暗地进城，如同战场上逃跑、羞愧的士兵一般。
2SAM|19|4|王蒙着脸，大声哭号说：“我儿 押沙龙 啊！ 押沙龙 ，我儿，我儿啊！”
2SAM|19|5|约押 进了宫到王那里，说：“你今日使你众臣仆的脸面羞愧了！他们今日救了你的性命和你儿女妻妾的性命，
2SAM|19|6|你却爱那些恨你的人，恨那些爱你的人。今日你摆明了不以将帅、臣仆为念。我今日看得出，若 押沙龙 活着，我们今日全都死了，你就高兴了。
2SAM|19|7|现在你要起来，出去安慰你臣仆的心。我指着耶和华起誓：你若不出去，今夜必没有一人跟你在一起了。这祸患比你从幼年到如今所遭受的更严重！”
2SAM|19|8|于是王起来，坐在城门口。有人告诉众军兵说：“看哪，王坐在城门口。”众军兵就都到王的面前。 那时， 以色列 人已经逃跑，各回自己的帐棚去了。
2SAM|19|9|以色列 众支派的百姓都议论纷纷，说：“王曾救我们脱离仇敌的手，又救我们脱离 非利士 人的手，现在他为了 押沙龙 逃离这地了。
2SAM|19|10|我们所膏治理我们的 押沙龙 已经阵亡。现在你们为什么沉默，不请王回来呢？”
2SAM|19|11|大卫 王派人到 撒督 和 亚比亚他 二位祭司那里，说：“你们当向 犹大 长老说：‘ 以色列 众人已经有话到了王那里 ，你们为什么最后才请王回宫呢？
2SAM|19|12|你们是我的弟兄，是我的骨肉，为什么最后才请王回来呢？’
2SAM|19|13|你们要对 亚玛撒 说：‘你不是我的骨肉吗？我若不立你在我面前取代 约押 永久作元帅，愿上帝重重惩罚我！’”
2SAM|19|14|这样，他挽回了 犹大 众人的心，如同一人。他们就派人到王那里，说：“请王和王的众臣仆回来。”
2SAM|19|15|王回来了，到 约旦河 。 犹大 人来到 吉甲 ，去迎接王，请王过 约旦河 。
2SAM|19|16|来自 巴户琳 的 便雅悯 人 基拉 的儿子 示每 急忙与 犹大 人一同下去迎接 大卫 王。
2SAM|19|17|跟从 示每 的有一千个 便雅悯 人，还有 扫罗 家的仆人 洗巴 和他十五个儿子、二十个随从仆人，他们都赶紧过 约旦河 到王的面前。
2SAM|19|18|渡船就渡王的家眷过河 ，照王看为好的去做。 王过 约旦河 的时候， 基拉 的儿子 示每 俯伏在王面前，
2SAM|19|19|对王说：“我主我王离开 耶路撒冷 的那日，仆人行了悖逆的事，现在求我主不要因此加罪于仆人，不要记得，也不要放在心上。
2SAM|19|20|仆人明知自己有罪，看哪， 约瑟 全家之中，今日我首先下来迎接我主我王。”
2SAM|19|21|洗鲁雅 的儿子 亚比筛 回答说：“ 示每 既然咒骂耶和华的受膏者，不应当为这缘故处死他吗？”
2SAM|19|22|大卫 说：“ 洗鲁雅 的儿子，我与你们有何相干，你们今日要跟我作对吗？今日在 以色列 中岂可把任何人处死呢？我岂不知今日我是 以色列 的王吗？”
2SAM|19|23|于是王对 示每 说：“你必不死。”王就向他起誓。
2SAM|19|24|扫罗 的孙子 米非波设 也下去迎接王。他自从王离开的那一日，直到王平安回 耶路撒冷 的日子，没有修脚，没有剃胡须，也没有洗衣服。
2SAM|19|25|他来迎接王的时候 ，王对他说：“ 米非波设 ，你为什么没有与我同去呢？”
2SAM|19|26|他说：“我主我王啊，我的仆人欺骗了我。那日仆人想要备驴骑上，与王同去，因为仆人是瘸腿的。
2SAM|19|27|他却在我主我王面前毁谤仆人。然而我主我王如同上帝的使者一样，你看怎样好，就怎样做吧！
2SAM|19|28|因为我祖全家的人，在我主我王面前不过是该死的人，王却使仆人列在王的席上吃饭的人当中，我现在还有什么权利能向王请求呢？”
2SAM|19|29|王对他说：“你何必再提你的事呢？我说，你与 洗巴 要平分土地。”
2SAM|19|30|米非波设 对王说：“我主我王既然平安地回宫，甚至让 洗巴 全都拿去也没关系。”
2SAM|19|31|基列 人 巴西莱 从 罗基琳 下来，要护送王过 约旦河 ，就跟王一同过 约旦河 。
2SAM|19|32|巴西莱 年纪老迈，已经八十岁了。王住在 玛哈念 的时候，他拿食物来供给王，因他是个大富翁。
2SAM|19|33|王对 巴西莱 说：“你与我一同渡过去，我要在 耶路撒冷 我的身边奉养你。”
2SAM|19|34|巴西莱 对王说：“我还能活多少年日，可以与王一同上 耶路撒冷 呢？
2SAM|19|35|今日我已八十岁了，还能辨别美丑吗？仆人还能尝出饮食的滋味吗？还能听男女歌唱的声音吗？仆人何必拖累我主我王呢？
2SAM|19|36|仆人护送王过 约旦河 只是一件小事，王何必用这样的赏赐来报答我呢？
2SAM|19|37|请让我回去，死在我本城，葬在我父母的墓旁。看哪，这里有 金罕 作王的仆人，让他同我主我王过去，你看怎样好，就怎样对待他吧。”
2SAM|19|38|王说：“ 金罕 可以与我一同过去，我必照你看为好的待他。你要我做的，我都会为你做。”
2SAM|19|39|于是众百姓过了 约旦河 ，王也过去了。王亲吻 巴西莱 ，为他祝福， 巴西莱 就回自己的地方去了。
2SAM|19|40|王渡过去 ，到了 吉甲 ， 金罕 也跟他过去。 犹大 众百姓和 以色列 百姓的一半也都送王过去。
2SAM|19|41|看哪， 以色列 众人来到王那里，对王说：“我们的弟兄 犹大 人为什么暗暗地送王和王的家眷，以及所有跟随王的人，过 约旦河 呢？”
2SAM|19|42|犹大 众人回答 以色列 人说：“因为王与我们是亲属，你们为何因这事发怒呢？我们靠王吃了什么呢？王真正给了我们什么赏赐呢？”
2SAM|19|43|以色列 人回答 犹大 人说：“我们与王有十倍的关系，就是在 大卫 身上，我们也比你们更有权利 。你们为何藐视我们呢？我们不是最先提议请王回来的吗？”但 犹大 人的话比 以色列 人的话更强硬。
2SAM|20|1|在那里恰巧有一个无赖，名叫 示巴 ，是 便雅悯 人 比基利 的儿子。他吹角，说： “我们与 大卫 无份， 与 耶西 的儿子无关。 以色列 啊，各回自己的帐棚去吧！”
2SAM|20|2|于是 以色列 众人都离弃 大卫 去跟随 比基利 的儿子 示巴 ，但 犹大 人从 约旦河 直到 耶路撒冷 ，都紧紧跟随他们的王。
2SAM|20|3|大卫 王来到 耶路撒冷 ，进了宫，就把从前留下看守宫殿的十个妃嫔软禁在冷宫，养活她们，却不与她们亲近。她们被关起来，活着如同寡妇，直到死的日子。
2SAM|20|4|王对 亚玛撒 说：“你要在三日之内召集 犹大 人到我这里来，你自己也要留在这里。”
2SAM|20|5|亚玛撒 就去召集 犹大 人，不过他却耽延，过了王所定的期限。
2SAM|20|6|大卫 对 亚比筛 说：“现在 比基利 的儿子 示巴 对我们的危害恐怕比 押沙龙 更大。你要带领你主的一些仆人追赶他，免得他得了坚固的城镇，在我们眼前逃脱 。”
2SAM|20|7|约押 的人和 基利提 人、 比利提 人，以及所有的勇士都跟着 亚比筛 ，从 耶路撒冷 出去追赶 比基利 的儿子 示巴 。
2SAM|20|8|他们到了 基遍 的大石头那里， 亚玛撒 来迎接他们。那时 约押 穿着战衣，腰束佩刀的带子，刀在鞘内。 约押 前行时，刀从鞘内掉出来。
2SAM|20|9|约押 对 亚玛撒 说：“我的弟兄，你平安吗？”他就用右手抓住 亚玛撒 的胡子，要亲吻他。
2SAM|20|10|亚玛撒 没有防备 约押 手里拿着的刀； 约押 用刀刺入他的肚腹，他的肠子流在地上， 约押 没有再刺，他就死了。 约押 和他弟弟 亚比筛 往前追赶 比基利 的儿子 示巴 。
2SAM|20|11|有 约押 的一个仆人站在 亚玛撒 尸体的旁边，说：“谁喜爱 约押 ，谁归顺 大卫 ，就当跟随 约押 。”
2SAM|20|12|亚玛撒 浑身是血，躺在路中间。那人见众百姓都站住，就把 亚玛撒 的尸体从路上移到田间，把衣服盖在他身上，因为他看见众人经过时都站住。
2SAM|20|13|尸体从路上移走之后，众人就都跟随 约押 去追赶 比基利 的儿子 示巴 。
2SAM|20|14|示巴 走遍 以色列 各支派，直到 伯．玛迦 的 亚比拉 ；所有精选的人 都聚集跟随他。
2SAM|20|15|跟随 约押 的众百姓到了 伯．玛迦 的 亚比拉 ，围困 示巴 ，对着城建土堆，与城郭相对。他们猛撞城墙，要使城倒塌。
2SAM|20|16|一个有智慧的妇人从城上呼叫：“听啊，听啊，请你们告诉 约押 ：‘近前来到这里，我好与你说话。’”
2SAM|20|17|约押 就近前到她那里，妇人对他说：“你是 约押 吗？”他说：“我是。”妇人对他说：“请你听使女的话。” 约押 说：“我正在听。”
2SAM|20|18|妇人说：“古时有话说，当在 亚比拉 求问，事情就可以解决。
2SAM|20|19|我在 以色列 中是和平、忠诚的。你现在想要毁坏这城， 以色列 的根源 ，为何你要吞灭耶和华的产业呢？”
2SAM|20|20|约押 回答说：“不，我绝不吞灭和毁坏！
2SAM|20|21|话不是这么说的，只是因为有一个 以法莲 山区的人，就是 比基利 的儿子名叫 示巴 ，他举手攻击 大卫 王；你们只要把他一人交出来，我就离城而去。”妇人对 约押 说：“看哪，他的首级必从城墙上丢给你。”
2SAM|20|22|妇人凭她的智慧去劝众百姓，他们就割下 比基利 的儿子 示巴 的首级，丢给 约押 。 约押 吹角，众人就离城散开，各回自己的帐棚去了。 约押 回 耶路撒冷 ，到王那里。
2SAM|20|23|约押 统管 以色列 全军； 耶何耶大 的儿子 比拿雅 统管 基利提 人和 比利提 人；
2SAM|20|24|亚多兰 管理劳役的人； 亚希律 的儿子 约沙法 作史官；
2SAM|20|25|示法 作书记； 撒督 和 亚比亚他 作祭司；
2SAM|20|26|睚珥 人 以拉 也作 大卫 的祭司。
2SAM|21|1|大卫 在位年间有饥荒，一连三年， 大卫 求问耶和华，耶和华说：“ 扫罗 和他家犯了流人血之罪，因为他杀死了 基遍 人。”
2SAM|21|2|大卫 王召了 基遍 人来，跟他们说话。 基遍 人不是 以色列 人，而是 亚摩利 人中所剩下的人。 以色列 人曾向他们起誓， 扫罗 却为 以色列 人和 犹大 人大发热心，追杀他们，为了要消灭他们。
2SAM|21|3|大卫 对 基遍 人说：“我当为你们做什么呢？要用什么赎这罪，使你们为耶和华的产业祝福呢？”
2SAM|21|4|基遍 人对他说：“我们和 扫罗 以及他家的事与金银无关，也不要因我们的缘故杀任何 以色列 人。” 大卫 说：“你们怎样说，我就为你们怎样做。”
2SAM|21|5|他们对王说：“那谋害我们、要消灭我们、使我们不得住 以色列 境内的人，
2SAM|21|6|请把他的子孙七人交给我们，我们好在耶和华面前，把他们悬挂在 基比亚 ，就是耶和华拣选 扫罗 的地方。”王说：“我必交给你们。”
2SAM|21|7|王顾惜 扫罗 的孙子， 约拿单 的儿子 米非波设 ，因为在 大卫 和 扫罗 的儿子 约拿单 之间，有指着耶和华的誓言。
2SAM|21|8|王却把 爱亚 的女儿 利斯巴 为 扫罗 所生的两个儿子 亚摩尼 和 米非波设 ，以及 扫罗 的女儿 米拉 为 米何拉 人 巴西莱 儿子 亚得列 所生的五个儿子
2SAM|21|9|交在 基遍 人的手里。 基遍 人在耶和华面前把他们悬挂在山上，这七人就一起死了。他们被杀的时候正是收割的头几天，就是开始收割大麦的时候。
2SAM|21|10|爱亚 的女儿 利斯巴 用麻布铺在磐石上搭棚，从收割的开始直到天降雨在尸体上，她白日不许空中的飞鸟落在尸体上，夜间不让田野的走兽前来。
2SAM|21|11|有人把 扫罗 的妃子 爱亚 女儿 利斯巴 所做的事告诉 大卫 。
2SAM|21|12|大卫 就去，从 基列 的 雅比 人那里把 扫罗 和他儿子 约拿单 的骸骨搬来。先前 非利士 人在 基利波 杀了 扫罗 ，把尸体悬挂在 伯．珊 的广场上，后来 基列 的 雅比 人把尸体偷走。
2SAM|21|13|大卫 把 扫罗 和他儿子 约拿单 的骸骨从那里搬上来，又收殓了被悬挂的那些人的骸骨。
2SAM|21|14|他们将 扫罗 和他儿子 约拿单 的骸骨葬在 便雅悯 的 洗拉 ，在 扫罗 父亲 基士 的坟墓里。他们遵照王所吩咐的一切做了。此后上帝垂听了为那地的祈求。
2SAM|21|15|非利士 人与 以色列 人打仗。 大卫 带领仆人下去，与 非利士 人交战， 大卫 就疲乏了。
2SAM|21|16|巨人族的后裔 以实．比诺 说要杀 大卫 ；他的铜枪重三百舍客勒，腰间又佩着新刀 。
2SAM|21|17|但 洗鲁雅 的儿子 亚比筛 帮助 大卫 攻击 非利士 人，杀死了他。当日， 大卫 的人向 大卫 起誓说：“你不可再与我们一同出战，免得 以色列 的灯熄灭了。”
2SAM|21|18|后来，在 歌伯 又与 非利士 人打仗，那时 户沙 人 西比该 杀了巨人族的后裔 撒弗 。
2SAM|21|19|他们又在 歌伯 与 非利士 人打仗， 伯利恒 人 雅雷 的儿子 伊勒哈难 杀了 迦特 人 歌利亚 ；这人的枪杆粗如织布机的轴。
2SAM|21|20|又有一次，他们在 迦特 打仗。那里有一个身材高大的人，双手各有六根手指，双脚各有六根脚趾，共有二十四根；他也是巨人族的后裔。
2SAM|21|21|他向 以色列 骂阵， 大卫 的哥哥 示米亚 的儿子 约拿单 就杀了他。
2SAM|21|22|这四个人是 迦特 巨人族的后裔，都仆倒在 大卫 和他仆人的手下。
2SAM|22|1|当耶和华救 大卫 脱离所有仇敌和 扫罗 之手的日子，他用这诗的歌词向耶和华说话。
2SAM|22|2|他说： 耶和华是我的岩石、我的山寨、我的救主、
2SAM|22|3|我的上帝、我的磐石、我所投靠的。 他是我的盾牌，是拯救我的角， 是我的碉堡，是我的避难所， 是我的救主，救我脱离凶暴的。
2SAM|22|4|我要求告当赞美的耶和华， 我必从仇敌手中被救出来。
2SAM|22|5|死亡的波浪环绕我， 毁灭的急流惊吓我，
2SAM|22|6|阴间的绳索缠绕我， 死亡的圈套临到我。
2SAM|22|7|我在急难中求告耶和华， 向我的上帝呼求。 他从殿中听了我的声音； 我的呼求进入他的耳中。
2SAM|22|8|那时，因他发怒地就摇撼震动； 天的根基也战抖摇撼。
2SAM|22|9|他的鼻孔冒烟上腾； 他的口发火焚烧，连煤炭也烧着了。
2SAM|22|10|他使天下垂，亲自降临； 黑云在他脚下。
2SAM|22|11|他乘坐基路伯飞行， 在风的翅膀上显现。
2SAM|22|12|他以黑暗和聚集的水、 天空的密云为四围的行宫。
2SAM|22|13|因他发出光辉， 火炭都烧着了。
2SAM|22|14|耶和华在天上打雷； 至高者发出声音。
2SAM|22|15|他射出箭来，使仇敌四散； 发出闪电，击溃他们。
2SAM|22|16|耶和华的斥责一发，鼻孔的气一出， 海底就显现，大地的根基也暴露。
2SAM|22|17|他从高天伸手抓住我， 把我从大水中拉上来。
2SAM|22|18|他救我脱离我的强敌， 脱离那些恨我的人， 因为他们比我强盛。
2SAM|22|19|我遭遇灾难的日子，他们来攻击我； 但耶和华是我的倚靠。
2SAM|22|20|他领我到宽阔之处， 他救拔我，因他喜爱我。
2SAM|22|21|耶和华必按我的公义报答我， 按我手中的清洁赏赐我。
2SAM|22|22|因为我遵守耶和华的道， 未曾作恶离开我的上帝。
2SAM|22|23|他的一切典章在我面前， 他的律例我也未曾丢弃。
2SAM|22|24|我在他面前作了完全人， 我也持守自己远离罪孽。
2SAM|22|25|所以耶和华按我的公义， 在他眼前按我的清洁赏赐我。
2SAM|22|26|慈爱的人，你以慈爱待他； 完全的人，你以完善待他；
2SAM|22|27|清洁的人，你以清洁待他； 歪曲的人，你以弯曲待他。
2SAM|22|28|困苦的百姓，你必拯救； 但你的眼目察看高傲的人，使他们降卑。
2SAM|22|29|耶和华啊，你是我的灯； 耶和华必照明我的黑暗。
2SAM|22|30|我藉着你冲入敌军， 藉着我的上帝跳过城墙。
2SAM|22|31|至于上帝，他的道是完全的； 耶和华的话是纯净的。 凡投靠他的，他就作他们的盾牌。
2SAM|22|32|除了耶和华，谁是上帝呢？ 除了我们的上帝，谁是磐石呢？
2SAM|22|33|上帝是我坚固的保障， 他为我开完全的路。
2SAM|22|34|他使我的脚快如母鹿， 使我站稳在高处。
2SAM|22|35|他教导我的手能争战， 我的膀臂能开铜造的弓。
2SAM|22|36|你赐救恩给我作盾牌， 你的庇护 使我为大。
2SAM|22|37|你使我脚步宽阔， 我的脚踝未曾滑跌。
2SAM|22|38|我追赶我的仇敌，消灭他们； 若不将他们灭绝，我总不归回。
2SAM|22|39|我灭绝了他们， 打伤了他们，使他们站不起来； 他们都倒在我的脚下。
2SAM|22|40|你曾以力量束我的腰，使我能争战； 也曾使那起来攻击我的，都服在我以下。
2SAM|22|41|你又使我的仇敌在我面前转身逃跑， 使我能歼灭那恨我的人。
2SAM|22|42|他们仰望，却无人拯救； 就是呼求耶和华，他也不应允。
2SAM|22|43|我捣碎他们，如同地上的灰尘； 践踏压碎他们，如同街上的泥土。
2SAM|22|44|你救我脱离我百姓 的纷争， 保护我作列国的元首； 我素不认识的百姓必事奉我。
2SAM|22|45|外邦人要向我投降， 一听见我的名声就必顺从我。
2SAM|22|46|外邦人要丧胆， 战战兢兢地出营寨。
2SAM|22|47|耶和华永远活着。 愿我的磐石被称颂， 愿上帝－救我的磐石受尊崇。
2SAM|22|48|这位上帝为我伸冤， 使万民服在我以下。
2SAM|22|49|他救我脱离仇敌， 又把我举起，高过那些起来攻击我的人， 救我脱离残暴的人。
2SAM|22|50|耶和华啊，因此我要在列国中称谢你， 歌颂你的名。
2SAM|22|51|耶和华赐极大的救恩给他所立的王， 施慈爱给他的受膏者， 就是给 大卫 和他的后裔，直到永远！
2SAM|23|1|以下是 大卫 末了的话： “ 耶西 的儿子 大卫 的话， 得居高位的， 雅各 的上帝所膏的， 以色列 所喜爱的诗人的话。
2SAM|23|2|耶和华的灵藉着我说话， 他的言语在我的舌头上。
2SAM|23|3|以色列 的上帝说， 以色列 的磐石向我说： ‘那以公义治理人， 以敬畏上帝来治理的，
2SAM|23|4|他必像晨光， 如无云清晨的日出， 如雨后的光辉， 在嫩草地上。’
2SAM|23|5|我的家在上帝面前不是如此吗？ 上帝与我立永远的约， 这约既全备又稳妥。 我的一切救恩和我一切所想望的， 他岂不成全吗？
2SAM|23|6|但无赖全都像被丢弃的荆棘； 它们不能用手去拿；
2SAM|23|7|碰它们的人必须用铁器和枪杆， 它们必在那里被火烧尽。”
2SAM|23|8|大卫 勇士的名字如下： 哈革摩尼 人 约设．巴设 ，他是三勇士之首；他又名叫 伊斯尼 人 亚底挪 ，曾一次就杀了八百人 。
2SAM|23|9|跟随 大卫 的三勇士中，其次是 亚何亚 人 朵多 的儿子 以利亚撒 。从前 非利士 人聚集要打仗，他们向 非利士 人骂阵。 以色列 人上去的时候，
2SAM|23|10|他起来击杀 非利士 人，直到手臂疲乏，手粘住刀把。那日耶和华大获全胜，百姓跟在 以利亚撒 后面只顾夺取掠物。
2SAM|23|11|再其次是 哈拉 人 亚基 的儿子 沙玛 。一次， 非利士 人聚集在 利希 ，在一块长满红豆的田里，百姓在 非利士 人面前逃跑。
2SAM|23|12|沙玛 却站在那田的中间，防守那田，击败了 非利士 人。耶和华大获全胜。
2SAM|23|13|开始收割的时候，三个 侍卫 下到 亚杜兰洞 ，到 大卫 那里。 非利士 的军兵在 利乏音谷 安营。
2SAM|23|14|那时 大卫 在山寨， 非利士 人的驻军在 伯利恒 。
2SAM|23|15|大卫 渴想着说：“但愿有人从 伯利恒 城门旁的井里打水来给我喝！”
2SAM|23|16|这三个勇士就闯过 非利士 人的军营，从 伯利恒 城门旁的井里打水，拿来给 大卫 喝。他却不肯喝，将水浇在耶和华面前，
2SAM|23|17|说：“耶和华啊，我绝不做这事！这三个人冒生命的危险，这不是他们的血吗？” 大卫 不肯喝这水。这是三个勇士所做的事。
2SAM|23|18|洗鲁雅 的儿子， 约押 的兄弟 亚比筛 是这三个勇士的领袖；他曾举枪杀了三百人，就在三个勇士中得了名。
2SAM|23|19|他在这三个 勇士中是最有名望的，所以作他们的领袖，只是不及前三个勇士。
2SAM|23|20|耶何耶大 的儿子 比拿雅 是来自 甲薛 的勇士，曾行了大事。他杀了 摩押 人 亚利伊勒 的两个儿子，又在下雪的时候下到坑里去，杀了一只狮子。
2SAM|23|21|他又杀了一个魁梧的 埃及 人； 埃及 人手里拿着枪。 比拿雅 只拿着棍子下到他那里去，从 埃及 人手里夺过枪来，用那枪杀死了他。
2SAM|23|22|这些是 耶何耶大 的儿子 比拿雅 所做的事，就在三个勇士里得了名。
2SAM|23|23|他比那三十个勇士 更有名望，只是不及前三个勇士。 大卫 立他作护卫长。
2SAM|23|24|三十个勇士中有 约押 的兄弟 亚撒黑 ， 伯利恒 人 朵多 的儿子 伊勒哈难 ，
2SAM|23|25|哈律 人 沙玛 ， 哈律 人 以利加 ，
2SAM|23|26|帕勒提 人 希利斯 ， 提哥亚 人 益吉 的儿子 以拉 ，
2SAM|23|27|亚拿突 人 亚比以谢 ， 户沙 人 米本乃 ，
2SAM|23|28|亚何亚 人 撒们 ， 尼陀法 人 玛哈莱 ，
2SAM|23|29|尼陀法 人 巴拿 的儿子 希立 ， 便雅悯 族 基比亚 人 利拜 的儿子 以太 ，
2SAM|23|30|比拉顿 人 比拿雅 ， 迦实溪 人 希太 ，
2SAM|23|31|亚拉巴 人 亚比．亚本 ， 巴鲁米 人 押斯玛弗 ，
2SAM|23|32|沙本 人 以利雅哈巴 ， 雅善 儿子中的 约拿单 ，
2SAM|23|33|哈拉 人 沙玛 ， 哈拉 人 沙拉 的儿子 亚希暗 ，
2SAM|23|34|玛迦 人 亚哈拜 的儿子 以利法列 ， 基罗 人 亚希多弗 的儿子 以连 ，
2SAM|23|35|迦密 人 希斯莱 ， 亚巴 人 帕莱 ，
2SAM|23|36|琐巴 人 拿单 的儿子 以甲 ， 迦得 人 巴尼 ，
2SAM|23|37|亚扪 人 洗勒 ， 比录 人 拿哈莱 ，是给 洗鲁雅 的儿子 约押 拿兵器的，
2SAM|23|38|以帖 人 以拉 ， 以帖 人 迦立 ，
2SAM|23|39|赫 人 乌利亚 ，共三十七人。
2SAM|24|1|耶和华的怒气又向 以色列 发作，激起 大卫 来对付他们，说：“去，数点 以色列 人和 犹大 人。”
2SAM|24|2|大卫 对跟随他的 约押 元帅说：“你来回走遍 以色列 众支派，从 但 直到 别是巴 ，数点百姓，我好知道百姓的数目。”
2SAM|24|3|约押 对王说：“愿耶和华－你的上帝使百姓的数目增加百倍，使我主我王亲眼得见。我主我王何必要做这事呢？”
2SAM|24|4|但王坚持他对 约押 和众军官的命令。 约押 和众军官就从王面前出去，数点 以色列 的百姓。
2SAM|24|5|他们过 约旦河 ，在 迦得谷 中、城的右边 亚罗珥 安营，与 雅谢 相对。
2SAM|24|6|他们来到 基列 ，到了 他停．合示 地 ，又来到 但．雅安 ，绕到 西顿 。
2SAM|24|7|他们来到 推罗 的堡垒，以及 希未 人和 迦南 人的各城，又出来，到 犹大尼革夫 的 别是巴 。
2SAM|24|8|他们来回走遍全地，过了九个月又二十天，就回到 耶路撒冷 。
2SAM|24|9|约押 向王报告百姓的总数： 以色列 拿刀的勇士有八十万； 犹大 有五十万人。
2SAM|24|10|大卫 数点百姓以后，心中自责。大卫向耶和华说：“我做这事大大有罪了。耶和华啊，现在求你除掉仆人的罪孽，因我所做的非常愚昧。”
2SAM|24|11|大卫 早晨起来，耶和华的话临到 迦得 先知，就是 大卫 的先见，说：
2SAM|24|12|“你去告诉 大卫 ：‘耶和华如此说：我向你提出三样，随你选择一样，我好降给你。’”
2SAM|24|13|于是 迦得 来到 大卫 那里告诉他，问他：“你要国中有七 年的饥荒呢？或是你在敌人面前逃跑，被追赶三个月呢？或是在你国中有三日的瘟疫呢？现在你要考虑思量，我怎样去回覆那差我来的。”
2SAM|24|14|大卫 对 迦得 说：“我很为难。我们宁愿落在耶和华的手里，因为他有丰盛的怜悯；我不愿落在人的手里。”
2SAM|24|15|于是，耶和华降瘟疫给 以色列 。自早晨到所定的时候，从 但 直到 别是巴 ，百姓中死了七万人。
2SAM|24|16|天使向 耶路撒冷 伸手要毁灭这城的时候，耶和华改变心意，不降那灾难，就对那在百姓中施行毁灭的天使说：“够了！住手吧！”耶和华的使者正在 耶布斯 人 亚劳拿 的禾场那里。
2SAM|24|17|大卫 看见那在百姓中施行毁灭的天使，就向耶和华说：“看哪，我犯了罪，行了恶，但这群羊做了什么呢？愿你的手攻击我和我的父家。”
2SAM|24|18|当日， 迦得 来到 大卫 那里，对他说：“你上去，在 耶布斯 人 亚劳拿 的禾场上为耶和华立一座坛。”
2SAM|24|19|大卫 就照着 迦得 的话，照着耶和华所吩咐的上去了。
2SAM|24|20|亚劳拿 观看，看见王和臣仆向他走过来。 亚劳拿 就出去，脸伏于地，向王下拜。
2SAM|24|21|亚劳拿 说：“我主我王为何来到仆人这里呢？” 大卫 说：“我要买你这禾场，为耶和华筑一座坛，使瘟疫在百姓中停止。”
2SAM|24|22|亚劳拿 对 大卫 说：“我主我王，你眼中看为好，就拿去献祭。看，这里有牛可以作燔祭，有打粮的器具和套牛的轭可以当作柴。
2SAM|24|23|王啊，这一切， 亚劳拿 都献给王。” 亚劳拿 又对王说：“愿耶和华－你的上帝悦纳你。”
2SAM|24|24|王对 亚劳拿 说：“不，我一定要按价钱向你买；我不能用白白得来的东西作燔祭献给耶和华－我的上帝。” 大卫 就用五十舍客勒银子买了那禾场与牛。
2SAM|24|25|大卫 在那里为耶和华筑了一座坛，献燔祭和平安祭。耶和华垂听了为那地的祈求，瘟疫就在 以色列 中停止了。
1KGS|1|1|大卫 王年纪老迈，虽然盖着外袍，仍不够暖和。
1KGS|1|2|臣仆对他说：“不如为我主我王找一个年轻的少女，侍立在王面前，照顾王，睡在王的怀中，好使我主我王得暖。”
1KGS|1|3|于是他们在 以色列 全境寻找美貌的少女，找到了一个 书念 女子 亚比煞 ，带到王那里。
1KGS|1|4|这少女极其美貌，她照顾王，伺候王，王却没有与她亲近。
1KGS|1|5|那时， 哈及 的儿子 亚多尼雅 妄自尊大，说：“我要作王”，就为自己预备座车、骑兵，又派五十人在他前头奔跑。
1KGS|1|6|他父亲从来没有责怪他，说：“你为何这么做？”他非常俊美，生在 押沙龙 之后。
1KGS|1|7|亚多尼雅 与 洗鲁雅 的儿子 约押 和 亚比亚他 祭司商议；他们就顺从 亚多尼雅 ，帮助他。
1KGS|1|8|但 撒督 祭司、 耶何耶大 的儿子 比拿雅 、 拿单 先知、 示每 、 利以 ，以及 大卫 自己的勇士 都不顺从 亚多尼雅 。
1KGS|1|9|亚多尼雅 在 隐．罗结 旁 琐希列 磐石那里献牛羊、肥犊为祭，请了他的众兄弟，就是王的众儿子，以及所有作王臣仆的 犹大 人。
1KGS|1|10|但他没有邀请 拿单 先知、 比拿雅 和勇士们，以及他的弟弟 所罗门 。
1KGS|1|11|拿单 对 所罗门 的母亲 拔示巴 说：“ 哈及 的儿子 亚多尼雅 作王了，你没有听见吗？我们的主 大卫 却不知道。
1KGS|1|12|现在，来，我给你出个主意，好保全你和你儿子 所罗门 的性命。
1KGS|1|13|你去，进到 大卫 王那里，对他说：‘我主我王啊，你不是曾向使女起誓说：你儿子 所罗门 必接续我作王，他必坐在我的王位上吗？ 亚多尼雅 怎么作了王呢？’
1KGS|1|14|看哪，你还在那里与王说话的时候，我会随后进去，证实你的话。”
1KGS|1|15|拔示巴 进入内室，到王那里。那时，王很老了， 书念 女子 亚比煞 正伺候着王。
1KGS|1|16|拔示巴 向王屈身下拜，王说：“你要什么？”
1KGS|1|17|她对王说：“我主啊，你曾向使女指着耶和华－你的上帝起誓：‘你儿子 所罗门 必接续我作王，他必坐在我的王位上。’
1KGS|1|18|现在，看哪， 亚多尼雅 作王了，你 ，我主我王却不知道。
1KGS|1|19|他献许多牛羊、肥犊为祭，请了王的众儿子和 亚比亚他 祭司，以及 约押 元帅，他却没有请王的仆人 所罗门 。
1KGS|1|20|但你 ，我主我王啊， 以色列 众人的眼目都仰望你，等你告诉他们，在我主我王之后谁坐你的王位。
1KGS|1|21|若不然，我主我王与祖先同睡的时候，我和我儿子 所罗门 必列为罪犯了。”
1KGS|1|22|看哪， 拔示巴 还与王说话的时候， 拿单 先知也进来了。
1KGS|1|23|有人奏告王说：“看哪， 拿单 先知来了。” 拿单 进到王面前，脸伏于地，向王叩拜。
1KGS|1|24|拿单 说：“我主我王，你果真说过‘ 亚多尼雅 必接续我作王，他要坐在我的王位上’吗？
1KGS|1|25|他今日下去，献了许多牛羊、肥犊为祭，请了王的众儿子和军官们，以及 亚比亚他 祭司；看哪，他们正在 亚多尼雅 面前吃喝，说：‘ 亚多尼雅 王万岁！’
1KGS|1|26|至于我，就是你的仆人，和 撒督 祭司、 耶何耶大 的儿子 比拿雅 、王的仆人 所罗门 ，他都没有请。
1KGS|1|27|这事果真出于我主我王吗？王却没有告诉仆人们，在我主我王之后谁坐你的王位。”
1KGS|1|28|大卫 王回答说：“召 拔示巴 到我这里来。” 拔示巴 就来，站在王面前。
1KGS|1|29|王起誓说：“我指着救我性命脱离一切苦难的永生的耶和华起誓。
1KGS|1|30|我既然指着耶和华－ 以色列 的上帝向你起誓说：你儿子 所罗门 必接续我作王，他必继承我坐在我的王位上，我今日必这样做。”
1KGS|1|31|于是， 拔示巴 屈身，脸伏于地，向王叩拜，说：“我主 大卫 王万岁！”
1KGS|1|32|大卫 王又说：“召 撒督 祭司、 拿单 先知、 耶何耶大 的儿子 比拿雅 到我这里来！”他们就都来到王面前。
1KGS|1|33|王对他们说：“要带领你们主的仆人，让我儿子 所罗门 骑我自己的骡子，送他下到 基训 。
1KGS|1|34|在那里， 撒督 祭司和 拿单 先知要膏他作 以色列 的王；你们也要吹角，说：‘ 所罗门 王万岁！’
1KGS|1|35|你们要跟随他上来，使他坐在我的王位上，他要接续我作王。我已立他作 以色列 和 犹大 的君王。”
1KGS|1|36|耶何耶大 的儿子 比拿雅 回应王说：“阿们！愿耶和华－我主我王的上帝这样说。
1KGS|1|37|耶和华怎样与我主我王同在，愿他照样与 所罗门 同在，使他的王位比我主 大卫 王的王位更大。”
1KGS|1|38|于是， 撒督 祭司、 拿单 先知、 耶何耶大 的儿子 比拿雅 ，以及 基利提 人和 比利提 人都下去，让 所罗门 骑上 大卫 王的骡子，送他到 基训 。
1KGS|1|39|撒督 祭司从帐幕中取了盛膏油的角来，膏 所罗门 。他们就吹角，众百姓都说：“ 所罗门 王万岁！”
1KGS|1|40|众百姓跟随他上来，吹着笛，大大欢呼，地被他们的声音震裂。
1KGS|1|41|亚多尼雅 和所有的宾客刚吃完，听见这声音； 约押 听见角声就说：“城中为何有这响声呢？”
1KGS|1|42|他正说话的时候，看哪， 亚比亚他 祭司的儿子 约拿单 来了。 亚多尼雅 说：“进来吧！你是个贤明的人，必是来报好消息的。”
1KGS|1|43|约拿单 回答 亚多尼雅 说：“我们的主 大卫 王已经立 所罗门 为王了！
1KGS|1|44|王派 撒督 祭司、 拿单 先知、 耶何耶大 的儿子 比拿雅 ，以及 基利提 人和 比利提 人和 所罗门 一起去，叫他骑上王的骡子。
1KGS|1|45|撒督 祭司和 拿单 先知已经在 基训 膏他作王了。他们从那里欢呼着上来，城都震动，这就是你们所听见的声音。
1KGS|1|46|所罗门 也已经登上国度的王位了。
1KGS|1|47|王的臣仆也来为我们的主 大卫 王祝福，说：‘愿上帝使 所罗门 的名比你的名更尊荣，使他的王位比你的王位更大。’王在床上屈身敬拜，
1KGS|1|48|王也这样说：‘耶和华－ 以色列 的上帝是应当称颂的，因他今日赏赐一个人坐在我的王位上，我也亲眼看见了。’”
1KGS|1|49|亚多尼雅 所有的宾客都战兢，起来，各走各路去了。
1KGS|1|50|亚多尼雅 惧怕 所罗门 ，就起来，去抓住祭坛的翘角。
1KGS|1|51|有人告诉 所罗门 说：“看哪， 亚多尼雅 惧怕 所罗门 王。看哪，他抓住祭坛的翘角，说：‘愿 所罗门 王先向我起誓，必不用刀杀死仆人。’”
1KGS|1|52|所罗门 说：“他若作贤明的人，连一根头发也不致落在地上；他若作恶，必要死亡。”
1KGS|1|53|于是 所罗门 王派人叫 亚多尼雅 从坛上下来，他就来向 所罗门 王下拜。 所罗门 对他说：“你回家去吧！”
1KGS|2|1|大卫 的死期临近了，就吩咐他儿子 所罗门 说：
1KGS|2|2|“我要走世人必走的路了。你当刚强，作大丈夫，
1KGS|2|3|遵守耶和华－你上帝所吩咐的，照着 摩西 律法上所写的行耶和华的道，谨守他的律例、诫命、典章、法度，好让你无论做什么，不拘往何处去，尽都亨通。
1KGS|2|4|耶和华必成就他所说关于我的话，说：‘你的子孙若谨慎自己的行为，尽心尽意凭信实行在我面前，就不断有人坐 以色列 的王位。’
1KGS|2|5|你也知道 洗鲁雅 的儿子 约押 向我所做的事，他对付 以色列 的两个元帅， 尼珥 的儿子 押尼珥 和 益帖 的儿子 亚玛撒 ，杀了他们。他在太平之时，如同战争一般，流这二人的血，把这战争的血染了他腰间束的带和脚上穿的鞋。
1KGS|2|6|所以你要照你的智慧去做，不让他白发安然下阴间。
1KGS|2|7|你当恩待 基列 人 巴西莱 的众儿子，请他们常与你同席吃饭，因为我躲避你哥哥 押沙龙 的时候，他们亲近我。
1KGS|2|8|看哪，在你这里有来自 巴户琳 的 便雅悯 人， 基拉 的儿子 示每 。我到 玛哈念 去的那日，他用狠毒的言语咒骂我。后来他却下 约旦河 迎接我，我就指着耶和华向他起誓说：‘我必不用刀杀死你。’
1KGS|2|9|但现在你不要以他为无罪。你是有智慧的人，必知道怎样待他，使他白发流血下阴间。”
1KGS|2|10|大卫 与他祖先同睡，葬在 大卫城 。
1KGS|2|11|大卫 作 以色列 王四十年：在 希伯仑 作王七年，在 耶路撒冷 作王三十三年。
1KGS|2|12|所罗门 坐他父亲 大卫 的王位，他的国度非常稳固。
1KGS|2|13|哈及 的儿子 亚多尼雅 到 所罗门 的母亲 拔示巴 那里， 拔示巴 问他说：“你是为平安来的吗？”他说：“为平安来的。”
1KGS|2|14|他又说：“我有话对你说。” 拔示巴 说：“你说吧。”
1KGS|2|15|亚多尼雅 说：“你知道这国原是归我的，全 以色列 也都期望我作王。然而，这国反归了我兄弟，因这国归了他是出乎耶和华。
1KGS|2|16|现在我有一件事求你，请你不要推辞。” 拔示巴 对他说：“你说吧。”
1KGS|2|17|他说：“求你请 所罗门 王把 书念 女子 亚比煞 赐我为妻，因他必不拒绝你。”
1KGS|2|18|拔示巴 说：“好，我必为你对王提说。”
1KGS|2|19|于是， 拔示巴 来到 所罗门 王那里，要为 亚多尼雅 说话。王起来迎接，向她下拜，然后坐在自己的位上，又为王的母亲设一座位，她就坐在王的右边。
1KGS|2|20|拔示巴 说：“我要向你提出一个小小的请求，请你不要回绝我。”王对她说：“母亲，请提出来，我必不回绝你。”
1KGS|2|21|拔示巴 说：“请你把 书念 女子 亚比煞 赐给你哥哥 亚多尼雅 为妻。”
1KGS|2|22|所罗门 王回答母亲说：“为何替 亚多尼雅 求 书念 女子 亚比煞 呢？可以为他求王国吧！他是我的兄长，不但为他，也为 亚比亚他 祭司和 洗鲁雅 的儿子 约押 求吧！ ”
1KGS|2|23|所罗门 王指着耶和华起誓说：“ 亚多尼雅 讲这话是自己送命，不然，愿上帝重重惩罚我。
1KGS|2|24|耶和华坚立我，使我坐在父亲 大卫 的王位上，照着他所应许的为我建立家室；现在我指着永生的耶和华起誓， 亚多尼雅 今日必被处死。”
1KGS|2|25|于是 所罗门 王派 耶何耶大 的儿子 比拿雅 去击杀 亚多尼雅 ，他就死了。
1KGS|2|26|王对 亚比亚他 祭司说：“你回 亚拿突 归自己的田地去吧！你本是该死的，但因你在我父亲 大卫 面前抬过主耶和华的约柜，又与我父亲同受一切苦难，所以我今日不杀死你。”
1KGS|2|27|所罗门 就革除 亚比亚他 ，不让他作耶和华的祭司。这就应验了耶和华在 示罗 论 以利 家所说的话。
1KGS|2|28|虽然 约押 没有拥护 押沙龙 ，却拥护了 亚多尼雅 ；这消息传到 约押 那里，他就逃到耶和华的帐幕，抓住祭坛的翘角。
1KGS|2|29|有人告诉 所罗门 王：“ 约押 逃到耶和华的帐幕，看哪，他在祭坛的旁边。” 所罗门 就派 耶何耶大 的儿子 比拿雅 ，说：“去，杀了他。”
1KGS|2|30|比拿雅 来到耶和华的帐幕，对 约押 说：“王这样吩咐：‘你出来吧！’”他说：“不，我要死在这里。” 比拿雅 就去回覆王，说：“ 约押 这样说，他这样回答我。”
1KGS|2|31|王对他说：“你可以照着他的话去做，杀了他，把他葬了，好叫 约押 流无辜人血的罪不归在我和我的父家。
1KGS|2|32|耶和华必使 约押 的血归到他自己头上，因为他击杀两个比他又公义又良善的人，就是 尼珥 的儿子 以色列 的元帅 押尼珥 和 益帖 的儿子 犹大 的元帅 亚玛撒 ，用刀杀了他们，我父亲 大卫 却不知道。
1KGS|2|33|这二人的血必归到 约押 和他后裔头上，直到永远；惟有 大卫 和他的后裔，以及他的家与王位，必从耶和华那里得平安，直到永远。”
1KGS|2|34|于是 耶何耶大 的儿子 比拿雅 上去，击杀 约押 ，杀死他，把他葬在旷野 约押 自己的家里。
1KGS|2|35|王就立 耶何耶大 的儿子 比拿雅 作元帅，代替 约押 ，又使 撒督 祭司代替 亚比亚他 。
1KGS|2|36|王派人召 示每 来，对他说：“你要在 耶路撒冷 为自己建造房屋，住在那里，不可从那里出来到任何地方去。
1KGS|2|37|你当确实知道，你何日出来过 汲沦溪 ，就必定死！你的血必归到自己头上。”
1KGS|2|38|示每 对王说：“这话很好！我主我王怎样说，仆人必照样做。”于是 示每 住在 耶路撒冷 许多日子。
1KGS|2|39|过了三年， 示每 的两个奴仆逃到 玛迦 的儿子 迦特 王 亚吉 那里去。有人告诉 示每 说：“看哪，你的奴仆在 迦特 。”
1KGS|2|40|示每 起来，备上驴，往 迦特 到 亚吉 那里去找他的奴仆，从 迦特 带他的奴仆回来。
1KGS|2|41|有人告诉 所罗门 ：“ 示每 出 耶路撒冷 到 迦特 去，又回来了。”
1KGS|2|42|王就派人召 示每 来，对他说：“我岂不是叫你指着耶和华起誓，并且警告你说‘你当确实知道，你何日出来到任何地方去，就必定死’吗？你也对我说：‘这话很好，我必听从。’
1KGS|2|43|你为何不遵守你对耶和华的誓言和我吩咐你的命令呢？”
1KGS|2|44|王又对 示每 说：“你向我父亲 大卫 所做的一切恶事，你自己心里都知道，耶和华必使你的罪恶归到你自己的头上。
1KGS|2|45|但 所罗门 王必蒙福， 大卫 的王位必在耶和华面前坚立，直到永远。”
1KGS|2|46|于是王吩咐 耶何耶大 的儿子 比拿雅 ，他就出去，击杀 示每 ， 示每 就死了。这样，国度在 所罗门 的手中巩固了。
1KGS|3|1|所罗门 与 埃及 王法老结亲，娶了法老的女儿，接她进入 大卫城 ，直等到建完了自己的宫和耶和华的殿，以及 耶路撒冷 周围的城墙。
1KGS|3|2|当那些日子，百姓仍在丘坛献祭，因为还没有为耶和华的名建殿。
1KGS|3|3|所罗门 爱耶和华，遵行他父亲 大卫 的律例，只是还在丘坛献祭烧香。
1KGS|3|4|所罗门 王到 基遍 ，在那里献祭，因为 基遍 有极大的丘坛。 所罗门 在那坛上献了一千祭牲为燔祭。
1KGS|3|5|在 基遍 ，耶和华夜间在梦中向 所罗门 显现；上帝说：“你愿我赐你什么，你可以求。”
1KGS|3|6|所罗门 说：“你曾向你仆人我父亲 大卫 大施慈爱，因为他用忠信、公义、正直的心行在你面前。你又为他存留大慈爱，赐他一个儿子坐在他的王位上，正如今日一样。
1KGS|3|7|现在，耶和华－我的上帝啊，你使仆人接续我父亲 大卫 作王；但我是幼小的孩子，不知道应当怎样出入。
1KGS|3|8|仆人住在你拣选的百姓中，这百姓之多，多得不可点，不可算。
1KGS|3|9|所以求你赐仆人善于了解的心，可以判断你的百姓，辨别是非。不然，谁能判断你这么多的百姓呢？”
1KGS|3|10|所罗门 因为求这事，就蒙主喜悦。
1KGS|3|11|上帝对他说：“你既然求这事，不为自己求寿、求富，也不求灭绝你仇敌的性命，只求能明辨，可以听讼，
1KGS|3|12|看哪，我会照你的话去做，看哪，我会赐你智慧和明辨的心，在你以前没有像你的，在你以后也没有兴起像你的。
1KGS|3|13|你没有求的，我也赐给你，就是富足、尊荣，使你在世一切的日子，列王中没有一个能比你的。
1KGS|3|14|你若遵行我的道，谨守我的律例、诫命，正如你父亲 大卫 所行的，我必使你长寿。”
1KGS|3|15|所罗门 醒了，看哪，是个梦。他就来到 耶路撒冷 ，站在耶和华的约柜前，献燔祭和平安祭，又为众臣仆摆设宴席。
1KGS|3|16|那时，有两个妓女来，站在王面前。
1KGS|3|17|一个妇人说：“我主啊，我和这妇人同住一屋。她在屋子里的时候，我生了一个孩子。
1KGS|3|18|我生了以后第三天，这妇人也生了。我们是一起的，屋子里除了我们二人之外，再没有别人在屋子里。
1KGS|3|19|夜间，这妇人的儿子死了，因为她压在她的儿子身上。
1KGS|3|20|她半夜起来，趁你使女睡着的时候，从我旁边把我儿子抱走，放在她怀里，又把她死的儿子放在我怀里。
1KGS|3|21|清早，我起来要给我的儿子吃奶，看哪，他死了；早晨我仔细察看他，看哪，他不是我所生的儿子。”
1KGS|3|22|另一个妇人说：“不！我的儿子是活的，你的儿子是死的。”但这一个说：“不！你的儿子是死的，我的儿子是活的。”她们就在王面前争吵。
1KGS|3|23|王说：“这妇人说：‘这是我的儿子，他是活的，你的儿子是死的。’那妇人说：‘不！你的儿子是死的，我的儿子是活的。’”
1KGS|3|24|王就说：“给我拿刀来！”人就把刀拿到王面前来。
1KGS|3|25|王说：“把活孩子劈成两半，一半给这妇人，一半给那妇人。”
1KGS|3|26|活孩子的母亲为自己的儿子心急如焚，对王说：“求我主把活孩子给那妇人吧，万不可杀死他！”那妇人说：“这孩子也不归我，也不归你，你们就劈了吧！”
1KGS|3|27|王回应说：“把活孩子给这妇人，万不可杀死他，因为这妇人是他的母亲。”
1KGS|3|28|全 以色列 听见王这样判断，就都敬畏王，因为他们看见他心中有上帝的智慧，能够断案。
1KGS|4|1|所罗门 作全 以色列 的王。
1KGS|4|2|这些是他的官员： 撒督 的儿子 亚撒利雅 作祭司，
1KGS|4|3|示沙 的两个儿子 以利何烈 、 亚希亚 作书记， 亚希律 的儿子 约沙法 作史官，
1KGS|4|4|耶何耶大 的儿子 比拿雅 作元帅， 撒督 和 亚比亚他 作祭司，
1KGS|4|5|拿单 的儿子 亚撒利雅 作宰相， 拿单 的儿子 撒布得 作祭司和王的顾问，
1KGS|4|6|亚希煞 作管家， 亚比大 的儿子 亚多尼兰 掌管服劳役的工人。
1KGS|4|7|所罗门 在全 以色列 有十二个官员，供给王和王室的食物，每年各人供给一个月。
1KGS|4|8|这些是他们的名字：在 以法莲 山区有 便．户珥 ；
1KGS|4|9|在 玛迦斯 、 沙宾 、 伯．示麦 、 以伦．伯．哈南 有 便．底甲 ；
1KGS|4|10|在 亚鲁泊 有 便．希悉 ，他管理 梭哥 和 希弗 全地；
1KGS|4|11|在 多珥 山冈 有 便．亚比拿达 ，他娶了 所罗门 的女儿 她法 为妻；
1KGS|4|12|在 他纳 和 米吉多 ，以及靠近 撒拉他拿 、 耶斯列 下边的 伯．善 全地，从 伯．善 到 亚伯．米何拉 直到 约缅 的另一边有 亚希律 的儿子 巴拿 ；
1KGS|4|13|在 基列 的 拉末 有 便．基别 ，他管理在 基列 的 玛拿西 子孙 睚珥 的城镇， 巴珊 的 亚珥歌伯 地的六十座大城，各有城墙和铜闩；
1KGS|4|14|在 玛哈念 有 易多 的儿子 亚希拿达 ；
1KGS|4|15|在 拿弗他利 有 亚希玛斯 ，他也娶了 所罗门 的一个女儿 巴实抹 为妻；
1KGS|4|16|在 亚设 和 亚禄 有 户筛 的儿子 巴拿 ；
1KGS|4|17|在 以萨迦 有 帕路亚 的儿子 约沙法 ；
1KGS|4|18|在 便雅悯 有 以拉 的儿子 示每 ；
1KGS|4|19|在 基列 地，就是 亚摩利 王 西宏 和 巴珊 王 噩 之地，有 乌利 的儿子 基别 ，他一个官员管理这地 。
1KGS|4|20|犹大 人和 以色列 人如同海边的沙那样多，都吃喝快乐。
1KGS|4|21|所罗门 统治诸国，从 大河 到 非利士 地，直到 埃及 的边界。 所罗门 在世的日子，这些国都向他进贡，服事他。
1KGS|4|22|所罗门 每日所用的食物：三十歌珥细面，六十歌珥粗面，
1KGS|4|23|十头肥牛，二十头草场的牛，一百只羊，还有鹿、羚羊、麃子，以及肥禽。
1KGS|4|24|所罗门 管理整个 大河 西边，从 提弗萨 直到 迦萨 ，以及 大河 西边的诸王，属他的四境尽都平安。
1KGS|4|25|所罗门 在世的日子，从 但 到 别是巴 ， 犹大 和 以色列 各人都在自己的葡萄树下和无花果树下安然居住。
1KGS|4|26|所罗门 拥有给战车用的四万个 马棚，还有一万二千名骑兵。
1KGS|4|27|这些官员各按自己的月份供给 所罗门 王，以及一切与他同席之人的食物，一无所缺。
1KGS|4|28|他们各按其分，把给马与快马吃的大麦和干草送到指定的地方去。
1KGS|4|29|上帝赐给 所罗门 极大的智慧和聪明，以及宽阔的心，如同海边的沙。
1KGS|4|30|所罗门 的智慧超过所有东方人的智慧，和 埃及 人一切的智慧。
1KGS|4|31|他的智慧胜过万人，胜过 以斯拉 人 以探 ，以及 玛曷 的儿子 希幔 、 甲各 、 达大 。他的名声传遍四围的列国。
1KGS|4|32|他作箴言三千句，诗歌一千零五首。
1KGS|4|33|他讲论草木，从 黎巴嫩 的香柏树直到墙上长的牛膝草，又讲论飞禽、走兽、爬行动物和鱼类。
1KGS|4|34|地上凡曾听过他智慧的君王，都派人来；万民都有人来听 所罗门 的智慧。
1KGS|5|1|推罗 王 希兰 是 大卫 平生的好友。 希兰 听见 以色列 人膏 所罗门 接续他父亲作王，就派臣仆到他那里。
1KGS|5|2|所罗门 也派人到 希兰 那里，说：
1KGS|5|3|“你知道我父亲 大卫 因四围的战争，不能为耶和华－他上帝的名建殿，直等到耶和华使仇敌都服在他脚下。
1KGS|5|4|现在耶和华－我的上帝使我四围太平，没有仇敌，没有灾祸。
1KGS|5|5|看哪，我吩咐要为耶和华－我上帝的名建殿，是照耶和华向我父亲 大卫 说的：‘我必使你儿子接续你，坐你的王位，他必为我的名建殿。’
1KGS|5|6|现在，请吩咐人在 黎巴嫩 为我砍伐香柏木，我的仆人必帮助你的仆人。至于你仆人的工钱，我必照你所定的给你。你知道，在我们中间没有人像 西顿 人那样擅长砍伐树木。”
1KGS|5|7|希兰 听见 所罗门 的话，就很高兴，说：“今日耶和华是应当称颂的，因为他赐给 大卫 一个有智慧的儿子，治理这众多的百姓。”
1KGS|5|8|希兰 送信给 所罗门 ，说：“你派人向我所提的那事，我已听见了；论到香柏木和松木，我必照你一切的心愿去做。
1KGS|5|9|我的仆人必把这木料从 黎巴嫩 运到海里，我会把它们扎成筏子浮在海上，运到你告诉我的地方，在那里拆开，你就可以收取；你也要照我的心愿做，把食物给我的家。”
1KGS|5|10|于是 希兰 照 所罗门 的心愿，给他香柏木和松木；
1KGS|5|11|所罗门 给 希兰 二万歌珥麦子，二十歌珥 捣成的油，作他家的食物。 所罗门 每年都是这样给 希兰 。
1KGS|5|12|耶和华照着所应许的赐智慧给 所罗门 。 希兰 与 所罗门 和平相处，二人彼此立约。
1KGS|5|13|所罗门 王从全 以色列 挑取服劳役的人，征来的人有三万，
1KGS|5|14|派他们轮流每月一万人上 黎巴嫩 去；一个月在 黎巴嫩 ，两个月在家里。 亚多尼兰 管理他们。
1KGS|5|15|所罗门 有七万扛抬的，八万在山上凿石头的。
1KGS|5|16|此外， 所罗门 有三千三百个监督工作的官长，监管百姓做工。
1KGS|5|17|王下令，他们就凿出又大又贵重的石头来，用以立殿的根基。
1KGS|5|18|所罗门 的工匠和 希兰 的工匠，以及 迦巴勒 人，把石头凿好，预备了木料和石头来建殿。
1KGS|6|1|以色列 人出 埃及 地后四百八十年， 所罗门 作 以色列 王第四年西弗月，就是二月，他开工建造耶和华的殿。
1KGS|6|2|所罗门 王为耶和华所建的殿，长六十肘，宽二十肘，高三十肘。
1KGS|6|3|殿的正堂前走廊长二十肘，与殿的宽度一样，殿前宽十肘；
1KGS|6|4|他为殿做了有框嵌壁式的窗户。
1KGS|6|5|靠着殿墙，围着外殿和内殿的墙，周围建造了厢房；
1KGS|6|6|下层宽五肘，中层宽六肘，第三层宽七肘。他在殿墙的周围造坎，免得梁木插入殿墙里。
1KGS|6|7|殿是用山中凿成的石头建的，所以建殿的时候，锤子、斧子和别样铁器的响声都没有听见。
1KGS|6|8|在殿右边当中的厢房有门，可以从螺旋梯上到中层，再从中层上到第三层。
1KGS|6|9|所罗门 完成殿的建造。他用香柏木作梁木和横板，遮盖殿顶。
1KGS|6|10|靠着整个殿所造的厢房，每层高五肘，香柏木的梁板搁在殿的墙坎上。
1KGS|6|11|耶和华的话临到 所罗门 ，说：
1KGS|6|12|“论到你所建的这殿，你若遵行我的律例，谨守我的典章，遵从我的一切诫命，行在其中，我必向你应验我所应许你父亲 大卫 的话。
1KGS|6|13|我必住在 以色列 人中间，并不丢弃我的百姓 以色列 。”
1KGS|6|14|所罗门 完成殿的建造。
1KGS|6|15|他用香柏木板建造殿的内墙，从殿的地到墙顶 都贴上木板，又用松木板铺地。
1KGS|6|16|他在殿的后部建了一间内殿，长二十肘，从地到墙 用香柏木板，作为至圣所。
1KGS|6|17|殿，就在内殿的前面 ，长四十肘。
1KGS|6|18|殿里一点石头都不显露，一概用香柏木遮蔽；香柏木上刻着野瓜和绽开的花。
1KGS|6|19|他在殿的中间预备内殿，在那里安放耶和华的约柜。
1KGS|6|20|内殿 长二十肘，宽二十肘，高二十肘，都贴上纯金。他又用香柏木做坛。
1KGS|6|21|所罗门 用纯金贴殿内，又用金链子挂在内殿前，内殿也贴上金子。
1KGS|6|22|整个殿都贴上金子，直到贴满；内殿前的整个坛，也都包上金子。
1KGS|6|23|他在内殿里用橄榄木做两个基路伯，各高十肘。
1KGS|6|24|这基路伯的一个翅膀长五肘，另一个翅膀长五肘，从一个翅膀尖到另一个翅膀尖共有十肘；
1KGS|6|25|第二个基路伯也是十肘；两个基路伯的尺寸、形状都一样。
1KGS|6|26|这一个基路伯高十肘，第二个基路伯也是如此。
1KGS|6|27|他把两个基路伯安在内殿中间。基路伯的翅膀是张开的，这基路伯的一个翅膀挨着这边的墙，第二个基路伯的一个翅膀挨着那边的墙，向内的两个翅膀在殿中间彼此相接。
1KGS|6|28|二基路伯都包上金子。
1KGS|6|29|殿周围的墙上全都刻着基路伯、棕树和绽开的花，内外都是如此。
1KGS|6|30|殿的地板都贴上金子，内外都是如此。
1KGS|6|31|他用橄榄木制造内殿的入口、门楣和五边形的门柱。
1KGS|6|32|在橄榄木做的两门扇上刻着基路伯、棕树和绽开的花，都贴上金子。基路伯和棕树上也洒上金子。
1KGS|6|33|他又为外殿的入口，用橄榄木制造门柱，是四边形的。
1KGS|6|34|他用松木做两扇门。这一扇有两叶摺叠，第二扇也有两叶 摺叠。
1KGS|6|35|上面刻着基路伯、棕树和绽开的花，雕刻物都均匀地贴上金子。
1KGS|6|36|他又用三层凿成的石头、香柏木一层建造内院。
1KGS|6|37|所罗门 在位第四年西弗月，立了耶和华殿的根基。
1KGS|6|38|到十一年布勒月，就是八月，殿和一切属殿的都按着样式造成。他建殿共用了七年。
1KGS|7|1|所罗门 为自己建造宫殿，十三年方才建成整座宫殿。
1KGS|7|2|他建造 黎巴嫩林宫 ，长一百肘，宽五十肘，高三十肘，有四行香柏木柱，柱上有香柏木横梁；
1KGS|7|3|厢房以上覆盖着香柏木，在四十五根柱子之上，每行十五根。
1KGS|7|4|窗户有三排，三排的窗与窗相对。
1KGS|7|5|所有的门和门柱都有四方形的框，共有三行，彼此相对。
1KGS|7|6|他建造有柱子的厅，长五十肘，宽三十肘。在这前面有走廊，前面有柱子和顶盖 。
1KGS|7|7|他又建造一个有座位的厅，就是审判厅，他在那里审判；这厅的地板从这边到那边都铺上香柏木。
1KGS|7|8|厅后面的院内有 所罗门 自己住的宫殿，都用同样的建造方式。 所罗门 又为所娶法老的女儿建造一座宫，建造方式与这厅一样。
1KGS|7|9|建造这一切所用的石头都是贵重的，按着尺寸凿成，用锯子里外锯齐；从根基直到房檐，从外头直到大院，都是如此。
1KGS|7|10|根基是贵重的大石头，有长十肘的，有长八肘的；
1KGS|7|11|上面有香柏木和按着尺寸凿成的贵重石头。
1KGS|7|12|大院周围有凿成的石头三层、香柏木板一层，都照耶和华殿的内院和殿的走廊的样式。
1KGS|7|13|所罗门 王派人从 推罗 把 户兰 接来。
1KGS|7|14|他是 拿弗他利 支派中一个寡妇的儿子，父亲是 推罗 人，是作铜匠的。 户兰 满有智慧、聪明、技能，善作各样的铜器。他来到 所罗门 王那里，为王做一切的工。
1KGS|7|15|户兰 制造两根铜柱，一根高十八肘，第二根柱子用绳子量，周围是十二肘 ；
1KGS|7|16|他做了两个柱顶安在柱上，是用铜铸造的，一个柱顶高五肘，第二个柱顶也高五肘。
1KGS|7|17|柱子顶上有装饰的网子和编成的链子，一个柱顶有七个，第二个柱顶也有七个。
1KGS|7|18|他做了柱子 ，第一根柱子的柱顶上，周围有两行网子在柱子 上面遮盖柱顶，第二根柱顶也是这样做。
1KGS|7|19|走廊柱子顶上的柱顶高四肘，刻着百合花。
1KGS|7|20|两根柱子上面有柱顶，柱顶靠近网子的圆凸面上，有石榴的行列环绕着，共二百个，第二个柱顶也是如此。
1KGS|7|21|他把两根柱子立在殿的走廊前：右边立一根，起名叫 雅斤 ；左边立一根，起名叫 波阿斯 。
1KGS|7|22|柱顶上刻着百合花。这样，柱子的工程就完毕了。
1KGS|7|23|他又铸一个铜海，周围是圆的，直径十肘，高五肘，用绳子量周围是三十肘。
1KGS|7|24|铜海边缘下面的周围有野瓜的形状，每肘十个，共两行，绕着铜海，是造铜海的时候铸上去的。
1KGS|7|25|铜海安在十二头铜牛上：三头向北，三头向西，三头向南，三头向东。铜海安在牛上，牛尾都向内。
1KGS|7|26|铜海厚一掌，边如杯边，像百合花，容量是二千罢特。
1KGS|7|27|他用铜制造十个盆座，每座长四肘，宽四肘，高三肘。
1KGS|7|28|铜座的造法是这样：周围各有嵌边，嵌边装在框架中。
1KGS|7|29|装在框架中的嵌边上有狮子和牛，以及基路伯。框架上有小座，狮子和牛的上面和下面有锤成的花纹浮雕。
1KGS|7|30|每座有四个铜轮和铜轴，它有四个支架在盆以下，这些支架是铸成的，各边都有花纹。
1KGS|7|31|它的口在柱顶里，向上高一肘，口是圆的，做法如座一样，直径是一肘半，口上也有雕工。嵌边是方形的，不是圆的。
1KGS|7|32|四个轮子在嵌边以下，轮轴与座相连，每轮高一肘半。
1KGS|7|33|轮的样式如同车的轮子；轴、辋、辐、毂都是铸成的。
1KGS|7|34|每个座四边有四个盆形的支架，这些支架是与座从一整块铸成的。
1KGS|7|35|座顶有圆架，高半肘；座顶有支柱和嵌边，是与座从一整块铸成的。
1KGS|7|36|他在支柱和嵌边上，每个空处刻上基路伯、狮子和棕树，周围有花纹。
1KGS|7|37|他按照这样的做法造了十个盆座，它们的铸法、尺寸、样式全都相同。
1KGS|7|38|他又造十个铜盆，每盆的容量四十罢特，直径四肘。在十个座上，每座安设一盆。
1KGS|7|39|他把五个安置在殿的右边，五个安置在殿的左边，又把铜海安置在殿的右旁，在东南边。
1KGS|7|40|户兰 又造了盆、铲子和盘子。这样， 户兰 为 所罗门 王做完了耶和华殿一切的工：
1KGS|7|41|两根柱子和柱子顶上两个如碗的柱顶，以及盖着如碗柱顶的两个网子；
1KGS|7|42|四百个石榴，安在两个网子上，每网两行石榴，盖着柱子上面两个如碗的柱顶；
1KGS|7|43|十个盆座和其上的十个盆；
1KGS|7|44|铜海和其下的十二头牛；
1KGS|7|45|盆、铲子、盘子。 户兰 给 所罗门 王为耶和华殿造的这一切器皿都是用光亮的铜，
1KGS|7|46|是王在 约旦 平原、 疏割 和 撒拉但 中间的泥巴地铸成的。
1KGS|7|47|所罗门 允许这一切器皿不过秤，因为所用的铜太多，重量无法计算。
1KGS|7|48|所罗门 又为耶和华的殿造了各样的器皿：金坛和献供饼的金供桌；
1KGS|7|49|内殿前的纯金灯台，右边五个，左边五个，以及其上的花、灯盏、灯剪，都是金的；
1KGS|7|50|纯金的杯、钳子、盘子、勺子 、火盆，以及圣殿的最里面，就是至圣所的门枢和外殿的门枢，都是金的。
1KGS|7|51|所罗门 王做完了耶和华殿一切的工，就把他父亲 大卫 分别为圣的金银和器皿都带来，放在耶和华殿的库房里。
1KGS|8|1|那时， 所罗门 召集 以色列 的长老、各支派的领袖和 以色列 人的族长到 耶路撒冷 ， 所罗门 王那里，要把耶和华的约柜从 大卫城 ，就是 锡安 ，接上来。
1KGS|8|2|以他念月，就是七月，在节期时，所有的 以色列 人都聚集到 所罗门 王那里。
1KGS|8|3|以色列 众长老一来到，祭司就抬起约柜。
1KGS|8|4|祭司和 利未 人将耶和华的约柜请上来，又把会幕和会幕一切的圣器皿都带上来。
1KGS|8|5|所罗门 王和聚集到他那里的 以色列 全会众一同在约柜前献牛羊为祭，多得不可胜数，无法计算。
1KGS|8|6|祭司将耶和华的约柜请进内殿，就是至圣所，安置在两个基路伯的翅膀底下约柜的地方。
1KGS|8|7|基路伯张开翅膀在约柜上面的地方，从上面遮住约柜和抬柜的杠。
1KGS|8|8|这杠很长，从内殿前的圣所可以看见杠头，从外面却看不见。这杠直到今日还在那里。
1KGS|8|9|约柜里没有别的，只有两块石版，就是 以色列 人出 埃及 地，耶和华与他们立约的时候， 摩西 在 何烈山 放在那里的。
1KGS|8|10|祭司从圣所出来的时候，有云充满耶和华的殿，
1KGS|8|11|祭司因云彩的缘故不能站立供职，因为耶和华的荣光充满了耶和华的殿。
1KGS|8|12|那时， 所罗门 说： “耶和华曾说要住在幽暗之处 。
1KGS|8|13|我的确为你建了一座雄伟的殿宇， 作为你永远居住的地方。”
1KGS|8|14|王转过脸来为 以色列 全会众祝福， 以色列 全会众都站立。
1KGS|8|15|所罗门 说：“耶和华－ 以色列 的上帝是应当称颂的！因他亲口向我父 大卫 应许的，也亲手成就了；他曾说：
1KGS|8|16|‘自从那日我领我百姓 以色列 出 埃及 以来，我未曾在 以色列 各支派中选择一城，在那里为我的名建造殿宇，但我拣选 大卫 治理我的百姓 以色列 。’
1KGS|8|17|我父 大卫 的心意是要为耶和华－ 以色列 上帝的名建殿。
1KGS|8|18|耶和华却对我父 大卫 说：‘你有心为我的名建殿，这心意是好的；
1KGS|8|19|但你不可建殿，惟有你亲生的儿子才可为我的名建殿。’
1KGS|8|20|现在耶和华实现了他所应许的话，使我接续我父 大卫 坐 以色列 的王位，正如耶和华所说的，我也为耶和华－ 以色列 上帝的名建造了这殿。
1KGS|8|21|我也在那里为约柜预备一处。约柜那里有耶和华的约，就是他领我们列祖出 埃及 地的时候，与他们所立的约。”
1KGS|8|22|所罗门 当着 以色列 全会众，站在耶和华的坛前，向天举手，
1KGS|8|23|说：“耶和华－ 以色列 的上帝啊，天上地下没有神明可与你相比！你向那些尽心行在你面前的仆人守约施慈爱，
1KGS|8|24|这约是你向你仆人 大卫 守的，是你应许他的。你亲口应许，亲手成就，正如今日一样。
1KGS|8|25|耶和华－ 以色列 的上帝啊，你向你仆人我父 大卫 应许说：‘你的子孙若谨慎自己的行为，在我面前行事像你所行的一样，就不断有人在我面前坐 以色列 的王位。’现在求你信守这话。
1KGS|8|26|以色列 的上帝啊，现在求你成就向你仆人我父 大卫 所应许的话。
1KGS|8|27|“上帝果真住在地上吗？看哪，天和天上的天尚且不足容纳你，何况我所建的这殿呢？
1KGS|8|28|惟求耶和华－我的上帝垂顾仆人的祷告祈求，俯听仆人今日在你面前的祈祷呼求。
1KGS|8|29|愿你的眼目昼夜看顾这殿，就是你说要作为你名的居所；求你垂听祷告，你仆人向此处的祷告。
1KGS|8|30|你仆人和你百姓 以色列 向此处祈祷的时候，求你在你天上的居所垂听，垂听而赦免。
1KGS|8|31|“人若得罪邻舍，有人强迫他，要他起誓，他来到这殿，在你的坛前起誓，
1KGS|8|32|求你在天上垂听、处理，向你的仆人施行审判，定恶人有罪，照他所行的报应在他头上；定义人为义，照他的义赏赐他。
1KGS|8|33|“你的百姓 以色列 若得罪你，败在仇敌面前，却又归向你，宣认你的名，在这殿里向你祈求祷告，
1KGS|8|34|求你在天上垂听，赦免你百姓 以色列 的罪，使他们归回你赐给他们列祖的地。
1KGS|8|35|“你的百姓若得罪了你，你使天闭塞不下雨；他们若向此处祷告，宣认你的名，因你的惩罚而离开他们的罪，
1KGS|8|36|求你在天上垂听，赦免你仆人你百姓 以色列 的罪，将当行的善道教导他们，并降雨在你的地，就是你赐给你百姓为业之地。
1KGS|8|37|“这地若有饥荒、瘟疫、焚风 、霉烂、蝗虫、蚂蚱，或有仇敌围困这地的 城门，无论遭遇什么灾祸疾病，
1KGS|8|38|你的百姓 以色列 ，或众人或一人，内心知道有祸，向这殿举手，无论祈求什么，祷告什么，
1KGS|8|39|求你在天上你的居所垂听、赦免、处理。因为你知道人心，惟有你知道世人的心，求你照各人所行的一切待他们，
1KGS|8|40|使他们在你赐给我们列祖的土地上一生一世敬畏你。
1KGS|8|41|“论到不属你百姓 以色列 的外邦人，若为你的名从远方而来，
1KGS|8|42|他们因听见你的大名和大能的手，以及伸出来的膀臂，来向这殿祷告，
1KGS|8|43|求你在天上你的居所垂听，照着外邦人向你所求的一切而行，使地上万民都认识你的名，敬畏你，像你的百姓 以色列 一样，又使他们知道我所建造的是称为你名下的殿。
1KGS|8|44|“你的百姓若奉你的派遣出去，无论往何处与仇敌争战，他们若向耶和华所选择的城，以及我为你名所建造的这殿祷告，
1KGS|8|45|求你在天上垂听他们的祷告祈求，为他们伸张正义。
1KGS|8|46|“你的百姓若得罪你，因为没有人不犯罪，你向他们发怒，把他们交在仇敌面前，掳他们的人把他们带到仇敌之地，或远或近，
1KGS|8|47|他们若在被掳之地那里回心转意，在掳掠者之地悔改，向你恳求说：‘我们有罪了，我们悖逆了，我们作恶了’；
1KGS|8|48|他们若在掳他们的仇敌之地尽心尽性归向你，又向自己的地，就是你赐给他们列祖的地和你所选择的城，以及我为你名所建造的这殿祷告，
1KGS|8|49|求你在天上你的居所垂听他们的祷告祈求，为他们伸张正义，
1KGS|8|50|饶恕得罪你的子民，赦免他们向你所犯一切的过犯，使他们在掳他们的人面前蒙怜悯。
1KGS|8|51|因为他们是你的子民，你的产业，是你从 埃及 ，从铁炉中领出来的。
1KGS|8|52|愿你的眼目看顾仆人和你百姓 以色列 的祈求；他们无论何时向你呼求，愿你垂听。
1KGS|8|53|主耶和华啊，你将他们从地上万民中分别出来作你的产业，是照着你领我们列祖出 埃及 的时候，藉你仆人 摩西 所应许的。”
1KGS|8|54|所罗门 在耶和华的坛前屈膝跪着，向天举手；他在耶和华面前祷告祈求完毕的时候，就起来，
1KGS|8|55|站着，大声为 以色列 全会众祝福，说：
1KGS|8|56|“耶和华是应当称颂的！因为他照着一切所应许的赐平安给他的百姓 以色列 ，凡藉他仆人 摩西 应许赐福的话，一句都没有落空。
1KGS|8|57|愿耶和华－我们的上帝与我们同在，像与我们列祖同在一样，不撇下我们，不丢弃我们，
1KGS|8|58|使我们的心归向他，遵行他一切的道，谨守他吩咐我们列祖的诫命、律例、典章。
1KGS|8|59|愿我在耶和华面前祈求的这些话，昼夜靠近耶和华－我们的上帝，好让他每日为他仆人和他百姓 以色列 伸张正义，
1KGS|8|60|使地上的万民都知道惟独耶和华是上帝，没有别的了。
1KGS|8|61|所以你们当向耶和华－我们的上帝存纯正的心，遵行他的律例，谨守他的诫命，如同今日一样。”
1KGS|8|62|王和全 以色列 一同在耶和华面前献祭。
1KGS|8|63|所罗门 向耶和华献平安祭，二万二千头牛，十二万只羊。这样，王和全 以色列 为耶和华的殿行了奉献之礼。
1KGS|8|64|当日，王因耶和华殿前的铜坛太小，容不下燔祭、素祭和平安祭牲的脂肪，就将耶和华殿前院子的中间分别为圣，在那里献燔祭、素祭和平安祭牲的脂肪。
1KGS|8|65|那时 所罗门 守节，从 哈马口 直到 埃及 溪谷的 以色列 众人都与他同在一起，成了一个盛大的会，在耶和华－我们的上帝面前七日又七日，共十四日。
1KGS|8|66|第八日，王遣散百姓；他们都为王祝福。他们为耶和华向他仆人 大卫 和他百姓 以色列 所施的一切恩惠都心中喜乐，愉快地各回自己的帐棚去了。
1KGS|9|1|所罗门 建造耶和华的殿和王宫，以及一切所想要建造的都完毕了，
1KGS|9|2|耶和华第二次向 所罗门 显现，如先前在 基遍 向他显现一样。
1KGS|9|3|耶和华对他说：“我已听了你在我面前的祷告和祈求，将你所建的这殿分别为圣，使我的名永远立在那里；我的眼、我的心也必时常在那里。
1KGS|9|4|你若以纯正的心和正直行在我面前，效法你父 大卫 所行的，遵行我一切所吩咐你的，谨守我的律例典章，
1KGS|9|5|我就必坚固你在 以色列 国度的王位，直到永远，正如我应许你父 大卫 说：‘你的子孙必不断有人坐 以色列 的王位。’
1KGS|9|6|倘若你们和你们的子孙转去不跟从我，不守我摆在你们面前的诫命律例，去事奉别神，敬拜它们，
1KGS|9|7|我就必把 以色列 从我赐给他们的地上剪除，也必从我面前舍弃那为我名所分别为圣的殿，使 以色列 在万民中成为笑柄，被人讥诮。
1KGS|9|8|这殿虽然崇高 ，将来凡经过的人必惊讶，嗤笑，说：‘耶和华为何向这地和这殿如此行呢？’
1KGS|9|9|人必说：‘因为此地的人离弃领他们祖先出 埃及 地的耶和华－他们的上帝，去亲近别神，敬拜事奉它们，所以耶和华使这一切灾祸临到他们。’”
1KGS|9|10|所罗门 建造耶和华殿和王宫这两座殿宇，用了二十年才完成。
1KGS|9|11|推罗 王 希兰 曾照 所罗门 所要的资助他香柏木、松木和金子， 所罗门 王就把 加利利 地的二十座城给了 希兰 。
1KGS|9|12|希兰 从 推罗 出来，察看 所罗门 给他的城镇，看不顺眼，
1KGS|9|13|就说：“我兄啊，你给我的是什么城镇呢？”他就给这些城镇起名叫 迦步勒 地，直到今日。
1KGS|9|14|希兰 曾给 所罗门 一百二十他连得金子。
1KGS|9|15|所罗门 王挑取服劳役的工人，为要建造耶和华的殿、自己的宫、 米罗 、 耶路撒冷 的城墙、 夏琐 、 米吉多 和 基色 。
1KGS|9|16|先前 埃及 王法老上来攻取 基色 ，用火焚烧，杀了城内居住的 迦南 人，把城赐给他的女儿，就是 所罗门 的妻子，作为嫁妆。
1KGS|9|17|所罗门 建造 基色 、 下伯．和仑 、
1KGS|9|18|巴拉 ，和位于境内旷野的 达莫 。
1KGS|9|19|所罗门 建造一切的储货城、战车城、战马城，以及他所想要建造的，在 耶路撒冷 、 黎巴嫩 和自己治理全国中的一切建设。
1KGS|9|20|至于所有剩下的百姓，不属 以色列 人的 亚摩利 人、 赫 人、 比利洗 人、 希未 人、 耶布斯 人，
1KGS|9|21|那些 以色列 人在当地不能灭尽的人， 所罗门 征召他们剩下的后代作服劳役的奴仆，直到今日。
1KGS|9|22|惟有 以色列 人， 所罗门 不使他们作奴仆，而是作他的战士、臣仆、官长、军官、战车长、骑兵长。
1KGS|9|23|这些是 所罗门 工程的五百五十个监工，他们在百姓中监管作工的人。
1KGS|9|24|法老的女儿从 大卫城 上到 所罗门 为她建造的宫里。那时， 所罗门 才建造 米罗 。
1KGS|9|25|所罗门 每年三次在他为耶和华所筑的坛上献燔祭和平安祭，又在耶和华面前的坛上烧香。这样，他完成了建殿。
1KGS|9|26|所罗门 王在 以东 地 红海 边，靠近 以禄 的 以旬．迦别 制造船只。
1KGS|9|27|希兰 派他的仆人，就是熟悉航海的船员，与 所罗门 的仆人一同坐船航海。
1KGS|9|28|他们到了 俄斐 ，从那里得了四百二十他连得金子，运到 所罗门 王那里。
1KGS|10|1|示巴 女王听见 所罗门 因耶和华的名所得的名声，就来要用难题考问 所罗门 。
1KGS|10|2|她带着很多的随从来到 耶路撒冷 ，有骆驼驮着香料、极多金子和宝石。她来到 所罗门 那里，向他提出心中所有的问题。
1KGS|10|3|所罗门 回答了她所有的问题，没有一个问题太难，王不能向她解答的。
1KGS|10|4|示巴 女王看见 所罗门 一切的智慧，和他所建造的宫殿，
1KGS|10|5|席上的食物，坐着的群臣，侍立的仆人，他们的服装，和他的司酒长，以及他在耶和华殿里所献的燔祭 ，就诧异得神不守舍。
1KGS|10|6|她对王说：“我在本国所听到的话，论到你的事和你的智慧是真的！
1KGS|10|7|我本来不信那些话，及至我来亲眼看见了，看哪，人所告诉我的还不到一半，你的智慧和你的福分超过我所听见的传闻。
1KGS|10|8|你的人 是有福的！你这些仆人常侍立在你面前、听你智慧的话是有福的！
1KGS|10|9|耶和华－你的上帝是应当称颂的！他喜爱你，使你坐 以色列 的王位，因为他永远爱 以色列 ，所以立你作王，使你秉公行义。”
1KGS|10|10|于是， 示巴 女王把一百二十他连得金子、极多的香料和宝石送给 所罗门 王；送来的香料，从来没有像 示巴 女王送给他的那么多。
1KGS|10|11|希兰 的船只也从 俄斐 运了金子来，又从 俄斐 运了许多檀香木和宝石来。
1KGS|10|12|王用檀香木为耶和华的殿和王宫做栏杆，又为歌唱的人做琴瑟。以后再没有这样的檀香木运进来，也再没有人见过，直到如今。
1KGS|10|13|所罗门 王除了照自己的厚意馈赠 示巴 女王之外，凡她所提出的一切要求， 所罗门 王都送给她。于是女王和她臣仆转回，到本国去了。
1KGS|10|14|所罗门 每年所得的金子，重六百六十六他连得；
1KGS|10|15|另外还有来自商人 和做生意的商品，以及 阿拉伯 诸王和各地省长的。
1KGS|10|16|所罗门 王用锤出来的金子打成二百面盾牌，每面盾牌用六百舍客勒金子；
1KGS|10|17|又用锤出来的金子打成三百面小盾牌，每面小盾牌用三弥那金子。王把它们放在 黎巴嫩林宫 里。
1KGS|10|18|王又制造一个大的象牙宝座，包上纯金。
1KGS|10|19|宝座有六层台阶，座的后背是圆的，座位之处两旁有扶手，靠近扶手有两只狮子站立。
1KGS|10|20|六层台阶上有十二只狮子站立，分站左边和右边；任何国度都没有这样做的。
1KGS|10|21|所罗门 王一切的饮器都是金的， 黎巴嫩林宫 里所有的器皿都是纯金的。在 所罗门 的日子，银子算不了什么。
1KGS|10|22|王有 他施 船只与 希兰 的船只一同航海， 他施 船只每三年一次把金、银、象牙、猿猴、孔雀 运回来。
1KGS|10|23|所罗门 王的财宝与智慧胜过地上的众王。
1KGS|10|24|全地都求见 所罗门 的面，要听上帝放在他心里的智慧。
1KGS|10|25|他们各带贡物，就是银器、金器、衣服、兵器、香料、马、骡子，每年都有一定的数量。
1KGS|10|26|所罗门 聚集战车骑兵；他有一千四百辆战车，一万二千名骑兵，安置在屯车城，在 耶路撒冷 的王那里。
1KGS|10|27|王在 耶路撒冷 使银子多如石头，香柏木多如 谢非拉 的桑树。
1KGS|10|28|所罗门 的马是从 埃及 和 科威 运来的，是王的商人按着定价从 科威 买来的。
1KGS|10|29|从 埃及 进口的战车，每辆六百舍客勒银子，马每匹一百五十舍客勒； 赫 人众王和 亚兰 诸王的战车和马，也是经由他们的手出口的。
1KGS|11|1|所罗门 王在法老的女儿之外，又宠爱许多外邦女子，就是 摩押 女子、 亚扪 女子、 以东 女子、 西顿 女子、 赫 人女子。
1KGS|11|2|论到这些国的人，耶和华曾吩咐 以色列 人说：“你们不可跟他们通婚，他们也不可跟你们在一起，因为他们一定会诱惑你们的心去随从他们的神明。” 所罗门 却为了爱，紧紧跟从他们。
1KGS|11|3|所罗门 娶七百个公主，三百个妃嫔。这些妻妾诱惑他的心。
1KGS|11|4|所罗门 年老的时候，他的妻妾诱惑他的心去随从别神，不像他父亲 大卫 以纯正的心顺服耶和华－他的上帝。
1KGS|11|5|所罗门 随从 西顿 人的女神 亚斯她录 和 亚扪 人可憎的 米勒公 。
1KGS|11|6|所罗门 行耶和华眼中看为恶的事，不像他父亲 大卫 专心顺从耶和华。
1KGS|11|7|那时， 所罗门 为 摩押 可憎的 基抹 和 亚扪 人可憎的 摩洛 ，在 耶路撒冷 对面的山上建造丘坛。
1KGS|11|8|他为所有的妻妾，就是那些向自己神明烧香献祭的外邦女子，也是这样做。
1KGS|11|9|耶和华向 所罗门 发怒，因为他的心偏离了向他显现两次的耶和华－ 以色列 的上帝。
1KGS|11|10|耶和华曾吩咐他这件事，不可随从别神，他却没有遵守耶和华所吩咐的。
1KGS|11|11|所以耶和华对他说：“你既然是这样，不遵守我所吩咐你守的约和律例，我必定把国度撕裂离开你，将它赐给你的大臣。
1KGS|11|12|然而，因你父亲 大卫 的缘故，我不在你的日子行这事，而要从你儿子的手中撕裂这国。
1KGS|11|13|只是我不撕裂全国，却要因我仆人 大卫 和我所选择的 耶路撒冷 ，保留一个支派给你的儿子。”
1KGS|11|14|耶和华使 以东 人 哈达 兴起，作 所罗门 的敌人；他是 以东 王的后裔。
1KGS|11|15|大卫 在 以东 的时候， 约押 元帅上去埋葬阵亡的人，杀了 以东 所有的男丁。
1KGS|11|16|约押 和 以色列 众人在 以东 住了六个月，直到把 以东 的男丁尽都剪除。
1KGS|11|17|那时 哈达 还是幼童；他和他父亲的臣仆，以及几个 以东 人逃往 埃及 。
1KGS|11|18|他们从 米甸 起行，到了 巴兰 ，再从 巴兰 带着几个人来到 埃及 ，到 埃及 王法老那里。法老给他房屋，吩咐给他粮食，又把地赐给他。
1KGS|11|19|哈达 在法老眼前大蒙恩宠，法老就把王后 答比匿 的妹妹嫁给他。
1KGS|11|20|答比匿 的妹妹给 哈达 生了一个儿子，叫 基努拔 。 答比匿 使 基努拔 在法老的宫里断奶， 基努拔 就与法老的众子一同住在法老的宫里。
1KGS|11|21|哈达 在 埃及 听见 大卫 与他祖先同睡， 约押 元帅也死了，就对法老说：“请你让我走，我要回本国去。”
1KGS|11|22|法老对他说：“你在我这里有什么缺乏？看哪，你竟想要回你本国去！”他说：“我没有缺乏什么，只是恳求王准我回去。”
1KGS|11|23|上帝又使 以利亚大 的儿子 利逊 兴起，作 所罗门 的敌人。他曾逃避主人 琐巴 王 哈大底谢 。
1KGS|11|24|大卫 击杀 琐巴 人的时候， 利逊 召集了一群人，自己作他们的领袖。他们往 大马士革 ，住在那里，在 大马士革 建立王国。
1KGS|11|25|所罗门 活着的时候，除了 哈达 为患之外， 利逊 也作 以色列 的敌人。他憎恨 以色列 ，作了 亚兰 人的王。
1KGS|11|26|尼八 的儿子 耶罗波安 也举起手来攻击王。他是 所罗门 的臣仆， 以法莲 支派的 洗利达 人；他母亲是个寡妇，名叫 洗鲁阿 。
1KGS|11|27|他举手攻击王是因先前 所罗门 建造 米罗 ，修补他父亲 大卫城 缺口的这件事。
1KGS|11|28|耶罗波安 是个大有才能的人。 所罗门 见这青年殷勤，就派他监管 约瑟 家所有服劳役的工人。
1KGS|11|29|那时， 耶罗波安 出了 耶路撒冷 ， 示罗 人 亚希雅 先知在路上遇见他； 亚希雅 身上穿着一件新衣。田野中只有他们二人，没有其他的人。
1KGS|11|30|亚希雅 拿起穿在自己身上的新衣，把它撕成十二片，
1KGS|11|31|对 耶罗波安 说：“你可以拿十片。耶和华－ 以色列 的上帝如此说：‘看哪，我必从 所罗门 手里撕裂这国，把十个支派赐给你。
1KGS|11|32|我因我仆人 大卫 和我在 以色列 众支派中所选择的 耶路撒冷城 的缘故，仍为 所罗门 留一个支派。
1KGS|11|33|因为他们 离弃我，敬拜 西顿 人的女神 亚斯她录 、 摩押 的神明 基抹 和 亚扪 人的神明 米勒公 ，没有像他父亲 大卫 一样遵从我的道，行我眼中看为正的事，守我的律例典章。
1KGS|11|34|但我不从他手里夺走整个国家，却使他在活着的日子作君王，是因我所拣选的仆人 大卫 遵守我的诫命律例。
1KGS|11|35|我必从他儿子手里将王国夺走，赐给你十个支派，
1KGS|11|36|只留一个支派给他的儿子，使我仆人 大卫 在我所选择立我名的 耶路撒冷城 那里，在我面前常有灯光。
1KGS|11|37|我选你，使你照你心里一切所愿的作王，成为 以色列 的王。
1KGS|11|38|你若听从我一切所吩咐你的，遵行我的道，行我眼中看为正的事，谨守我的律例诫命，像我仆人 大卫 所行的，我就与你同在，为你立坚固的家，像我为 大卫 所立的一样，将 以色列 赐给你。
1KGS|11|39|我必因这事使 大卫 的后裔遭受患难，但不是永远的。’”
1KGS|11|40|所罗门 想要杀 耶罗波安 ， 耶罗波安 起身逃往 埃及 。他到了 埃及 王 示撒 那里，就住在 埃及 ，直到 所罗门 死了。
1KGS|11|41|所罗门 其余的事，凡他所做的和他的智慧，不都写在《所罗门记》上吗？
1KGS|11|42|所罗门 在 耶路撒冷 作全 以色列 的王四十年。
1KGS|11|43|所罗门 与他祖先同睡，葬在他父亲 大卫 的城里，他儿子 罗波安 接续他作王。
1KGS|12|1|罗波安 往 示剑 去，因 以色列 众人都到了 示剑 ，要立他作王。
1KGS|12|2|尼八 的儿子 耶罗波安 先前躲避 所罗门 王，逃往 埃及 ，住在那里。他还在 埃及 ，听见了这事 ，
1KGS|12|3|以色列 人派人去请他来。 耶罗波安 就和 以色列 全会众来，与 罗波安 谈话，说：
1KGS|12|4|“你父亲使我们负重轭，现在求你减轻你父亲所加给我们的苦工和重轭，我们就服事你。”
1KGS|12|5|罗波安 对他们说：“你们走吧，过三天再来见我。”百姓就走了。
1KGS|12|6|罗波安 的父亲 所罗门 在世的日子，有侍立在他面前的长者， 罗波安 王和他们商议，说：“你们出个主意，好把话带回给这百姓。”
1KGS|12|7|他们对他说：“现在王若像仆人一样服事这百姓，用好话回覆他们，他们就永远作王的仆人了。”
1KGS|12|8|王不采纳长者给他出的主意，却和那些与他一同长大、在他面前侍立的年轻人商议。
1KGS|12|9|他对他们说：“这百姓对我说：‘你父亲使我们负重轭，求你减轻一些。’你们出个什么主意，我们好把话带回给他们。”
1KGS|12|10|那些与他一同长大的年轻人对他说：“这百姓对王说：‘你父亲使我们负重轭，求你给我们减轻一些。’王要对他们如此说：‘我的小指头比我父亲的腰还粗呢！
1KGS|12|11|我父亲使你们负重轭，现在我必使你们负更重的轭！我父亲用鞭子惩罚你们，我要用蝎子惩罚你们！’”
1KGS|12|12|耶罗波安 和众百姓遵照王所说“你们第三天再来见我”的话，第三天来到 罗波安 那里。
1KGS|12|13|王严厉地回答百姓，不采纳长者给他出的主意。
1KGS|12|14|他照着年轻人所出的主意对他们说：“我父亲使你们负重轭，我必使你们负更重的轭！我父亲用鞭子惩罚你们，我却要用蝎子惩罚你们！”
1KGS|12|15|王不依从百姓，因这事件是出于耶和华，为要应验耶和华藉 示罗 人 亚希雅 对 尼八 的儿子 耶罗波安 所说的话。
1KGS|12|16|以色列 众人见王不依从他们，百姓就回话给王，说： “我们在 大卫 中有什么份呢？ 我们在 耶西 的儿子中没有产业！ 以色列 啊，回你的帐棚去吧！ 大卫 啊，现在你顾自己的家吧！” 于是， 以色列 人都回自己的帐棚去了；
1KGS|12|17|至于住 犹大 城镇的 以色列 人， 罗波安 仍作他们的王。
1KGS|12|18|罗波安 王派监管劳役的 亚多兰 去， 以色列 众人用石头打他，他就死了。 罗波安 王急忙上车，逃回 耶路撒冷 去了。
1KGS|12|19|这样， 以色列 背叛 大卫 家，直到今日。
1KGS|12|20|以色列 众人听见 耶罗波安 回来了，就派人去请他到会众那里，立他作全 以色列 的王。除了 犹大 支派，没有跟从 大卫 家的。
1KGS|12|21|罗波安 来到 耶路撒冷 ，召集了 犹大 全家和 便雅悯 支派的人共十八万，都是精选的战士，要与 以色列 家打仗，好将王国夺回，归 所罗门 的儿子 罗波安 。
1KGS|12|22|但上帝的话临到神人 示玛雅 ，说：
1KGS|12|23|“你去告诉 所罗门 的儿子 犹大 王 罗波安 ， 犹大 和 便雅悯 全家，以及其余的百姓，说：
1KGS|12|24|‘耶和华如此说：你们不可上去与你们的弟兄 以色列 人打仗。你们各自回家去吧！因为这事是出于我。’”众人就听从耶和华的话，遵照耶和华的话回去了。
1KGS|12|25|耶罗波安 在 以法莲 山区建了 示剑 ，住在其中，又从 示剑 出去，建了 毗努伊勒 。
1KGS|12|26|耶罗波安 心里说：“现在，这国恐怕仍会归 大卫 家；
1KGS|12|27|这百姓若上 耶路撒冷 去，在耶和华的殿里献祭，他们的心必归向他们的主 犹大 王 罗波安 。他们会杀了我，仍归 犹大 王 罗波安 。”
1KGS|12|28|耶罗波安 王就筹划，铸造了两个金牛犊，对众百姓说：“你们上 耶路撒冷 去实在够久了。 以色列 啊，看哪，这是领你出 埃及 地的神明。”
1KGS|12|29|他把一个安置在 伯特利 ，另一个安置在 但 。
1KGS|12|30|这事使百姓陷入罪里，因为他们甚至到 但 去拜那牛犊。
1KGS|12|31|耶罗波安 在一些丘坛建神殿，立不属 利未 人的平民百姓为祭司。
1KGS|12|32|耶罗波安 定八月十五日为节期，像在 犹大 的节期一样，自己上坛献祭。他在 伯特利 这样做，向他所铸的牛犊献祭，又把他所立丘坛的祭司安置在 伯特利 。
1KGS|12|33|他在八月十五日，就是他自己心中所定的月份，在 伯特利 上到自己所造的祭坛；他为 以色列 人定了一个节期，亲自上坛烧香。
1KGS|13|1|看哪，有一个神人遵照耶和华的话从 犹大 来到 伯特利 。 耶罗波安 正站在坛旁烧香；
1KGS|13|2|神人遵照耶和华的话向坛呼叫，说：“坛哪，坛哪！耶和华如此说：‘看哪， 大卫 家必生一个儿子，名叫 约西亚 ，他必将在你上面烧香的丘坛祭司，宰杀在你上面，人的骨头也必烧在你上面。’”
1KGS|13|3|当日，神人设个预兆，说：“这是耶和华说的预兆：‘看哪，这坛必破裂，坛上的灰必倾倒出来。’”
1KGS|13|4|耶罗波安 王听见神人向 伯特利 的坛呼叫的话，就从坛上伸手，说：“拿住他！”王向神人所伸的手却萎缩了，不能弯回。
1KGS|13|5|坛也破裂了，坛上的灰倾倒出来，正如神人遵照耶和华的话所设的预兆。
1KGS|13|6|王对神人说：“请你为我祷告，向耶和华－你的上帝恳求恩惠，使我的手复原。”于是神人向耶和华恳求，王的手就复原了，如平常一样。
1KGS|13|7|王对神人说：“请你跟我回宫，让你恢复心力，我必给你赏赐。”
1KGS|13|8|神人对王说：“你就是把你一半的王宫给我，我也不跟你进去，也不在这地方吃饭喝水，
1KGS|13|9|因为耶和华的话这样吩咐我说：‘不可吃饭喝水，也不可从你去的原路回来。’”
1KGS|13|10|于是神人从别的路回去，不从他到 伯特利 来的原路回去。
1KGS|13|11|有一个老先知住在 伯特利 ，他的儿子来，把神人当日在 伯特利 所做的一切事和他向王所说的话，都告诉了父亲。
1KGS|13|12|父亲对他们说：“神人从哪条路去了呢？”他的儿子都看到 从 犹大 来的神人所去的路。
1KGS|13|13|老先知吩咐儿子说：“你们为我备驴。”他们备好了驴，他就骑上，
1KGS|13|14|去追神人，遇见神人坐在橡树底下，就对他说：“你是不是从 犹大 来的神人？”他说：“是我。”
1KGS|13|15|老先知对他说：“请你跟我一起回家吃饭。”
1KGS|13|16|神人说：“我不能跟你回去，与你同行，也不能在这地方跟你一起吃饭喝水，
1KGS|13|17|因为有耶和华的话吩咐我说：‘你在那里不可吃饭喝水，也不可从你去的原路回来。’”
1KGS|13|18|老先知对他说：“我也是先知，和你一样。有天使遵照耶和华的话对我说：‘你去带他一同回你的家，给他吃饭喝水。’”老先知在欺骗他。
1KGS|13|19|于是神人跟老先知回去，在他家里吃饭喝水。
1KGS|13|20|他们坐席的时候，耶和华的话临到那带神人回来的先知，
1KGS|13|21|他就对从 犹大 来的神人宣告说：“耶和华如此说：‘你既违背耶和华的指示，不遵守耶和华－你上帝的命令，
1KGS|13|22|反倒回来，在耶和华禁止你吃饭喝水的地方吃了饭喝了水，因此你的尸体必不得葬在你祖先的坟墓里。’”
1KGS|13|23|神人吃喝完了，老先知为他带回来的先知备驴。
1KGS|13|24|神人就去了，在路上有只狮子遇见他，把他咬死。他的尸体倒在路上，驴站在尸体旁边，狮子也站在尸体旁边。
1KGS|13|25|看哪，有人经过，看见尸体倒在路上，狮子站在尸体旁边，就来到老先知所住的城里述说这事。
1KGS|13|26|那带神人回来的先知听见了，就说：“这是那违背了耶和华指示的神人，所以耶和华把他交给狮子；狮子撕裂他，咬死他，正如耶和华对他说的话。”
1KGS|13|27|老先知吩咐他儿子说：“你们为我备驴。”他们就备了驴。
1KGS|13|28|他去了，发现神人的尸体倒在路上，驴和狮子站在尸体旁边，狮子却没有吃尸体，也没有撕裂驴。
1KGS|13|29|老先知把神人的尸体抬起，驮在驴上，带回自己的城里，要为他哀哭，为他安葬。
1KGS|13|30|老先知把尸体葬在自己的坟里，为他哀哭，说：“哀哉！我的弟兄啊！”
1KGS|13|31|安葬之后，老先知对他儿子说：“我死了，你们要把我葬在神人所葬的坟里，使我的尸骨在他的尸骨旁边，
1KGS|13|32|因为他遵照耶和华的话，指着 伯特利 的坛和 撒玛利亚 各城丘坛神殿所宣告的话必定应验。”
1KGS|13|33|这事以后， 耶罗波安 仍不离开他的恶道，立平民百姓为丘坛的祭司；凡愿意的，他都分别为圣，立为丘坛的祭司。
1KGS|13|34|这事使 耶罗波安 的家陷入罪里，甚至他的家被剪除，从地面上消灭了。
1KGS|14|1|那时， 耶罗波安 的儿子 亚比雅 病了。
1KGS|14|2|耶罗波安 对他的妻子说：“你起来改装，使人认不出你是 耶罗波安 的妻子。你往 示罗 去，看哪，那里有先知 亚希雅 ，他曾告诉我说，你必作这百姓的王。
1KGS|14|3|现在你手里要带十个饼、几个薄饼和一瓶蜜到他那里去，他必告诉你，孩子会怎样。”
1KGS|14|4|耶罗波安 的妻子就照样做，起身往 示罗 去，到了 亚希雅 的家。 亚希雅 因年纪老迈，两眼发直，不能看见。
1KGS|14|5|耶和华对 亚希雅 说：“看哪， 耶罗波安 的妻子来问你她儿子的事，因她儿子病了，你当如此如此告诉她。她进来的时候会扮成别的妇人。”
1KGS|14|6|她刚进门， 亚希雅 听见她的脚步声，就说：“ 耶罗波安 的妻子，进来吧！你为何扮成别的妇人呢？我奉差遣将凶信告诉你。
1KGS|14|7|你回去告诉 耶罗波安 说：‘耶和华－ 以色列 的上帝如此说：我从百姓中提拔了你，立你作我百姓 以色列 的君王，
1KGS|14|8|将 大卫 家的国撕裂，赐给你，你却不效法我仆人 大卫 ，遵守我的诫命，全心顺从我，行我眼中看为正的事。
1KGS|14|9|你反倒行恶，比在你之前所有的人更严重；你离开了我，为自己立了别神，铸了偶像，惹我发怒，将我丢在背后。
1KGS|14|10|因此，看哪，我必使灾祸临到 耶罗波安 的家，把属 耶罗波安 的男丁，无论是奴役的、自由的，都从 以色列 中剪除。我必除灭 耶罗波安 的家，如同人扫除粪土，直到消灭。
1KGS|14|11|凡属 耶罗波安 的人，死在城中的必被狗吃，死在田野的必被空中的鸟吃。这是耶和华说的。’
1KGS|14|12|你起身回家去吧！你的脚一进城，孩子就死了。
1KGS|14|13|以色列 众人必为他哀哭，为他安葬。凡属 耶罗波安 的人，只有他可以葬入坟墓，因为在 耶罗波安 的家中，只有他向耶和华－ 以色列 的上帝表现出好的行为。
1KGS|14|14|耶和华必另立一王治理 以色列 ，这一天，他必剪除 耶罗波安 的家；什么时候呢？现在就是了。
1KGS|14|15|耶和华必击打 以色列 ，使他们摇动，像水中的芦苇一样，又将他们从耶和华赐给他们列祖的美地上拔出来，分散在 大河 那边，因为他们造了 亚舍拉 ，惹耶和华发怒。
1KGS|14|16|因 耶罗波安 所犯的罪，又因他使 以色列 陷入罪里，耶和华必将 以色列 交出来。”
1KGS|14|17|耶罗波安 的妻子起身回去，到了 得撒 ，刚到门槛，孩子就死了。
1KGS|14|18|以色列 众人为他安葬，为他哀哭，正如耶和华藉他仆人 亚希雅 先知所说的话。
1KGS|14|19|耶罗波安 其余的事，他怎样打仗，怎样作王，看哪，都写在《以色列诸王记》上。
1KGS|14|20|耶罗波安 作王二十二年，就与他祖先同睡，他儿子 拿答 接续他作王。
1KGS|14|21|所罗门 的儿子 罗波安 作 犹大 王。他登基的时候年四十一岁，在 耶路撒冷 ，就是耶和华从 以色列 众支派中所选择立他名的城，作王十七年。 罗波安 的母亲名叫 拿玛 ，是 亚扪 人。
1KGS|14|22|犹大 人行耶和华眼中看为恶的事，以所犯的罪惹动他的妒忌，比他们的祖先所犯的一切更严重。
1KGS|14|23|因为他们在各高冈上，各青翠树下筑丘坛，立柱像和 亚舍拉 。
1KGS|14|24|国中也有男的庙妓。他们效法耶和华在 以色列 人面前所赶出的外邦人，行一切可憎恶的事。
1KGS|14|25|罗波安 王第五年， 埃及 王 示撒 上来攻打 耶路撒冷 ，
1KGS|14|26|夺了耶和华殿和王宫里的宝物，尽都带走，又夺走 所罗门 制造的一切金盾牌。
1KGS|14|27|罗波安 王制造铜盾牌代替那些金盾牌，交给看守王宫宫门的护卫长看管。
1KGS|14|28|每逢王进耶和华的殿，护卫兵就举起这些盾牌；随后仍将盾牌送回护卫室。
1KGS|14|29|罗波安 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
1KGS|14|30|罗波安 与 耶罗波安 时常交战。
1KGS|14|31|罗波安 与他祖先同睡，与他祖先同葬在 大卫城 。他母亲名叫 拿玛 ，是 亚扪 人，他儿子 亚比央 接续他作王。
1KGS|15|1|尼八 的儿子 耶罗波安 王十八年， 亚比央 登基作 犹大 王，
1KGS|15|2|在 耶路撒冷 作王三年。他母亲名叫 玛迦 ，是 押沙龙 的女儿。
1KGS|15|3|亚比央 行他父亲从前所犯一切的罪，他的心不像他曾祖父 大卫 以纯正的心顺服耶和华－他的上帝。
1KGS|15|4|然而耶和华－他的上帝因 大卫 的缘故，仍使大卫在 耶路撒冷 有灯光，立他儿子接续他作王，又坚立 耶路撒冷 。
1KGS|15|5|因为 大卫 除了 赫 人 乌利亚 那件事，都行耶和华眼中看为正的事，一生没有违背耶和华一切所吩咐的。
1KGS|15|6|罗波安 在世的日子常与 耶罗波安 交战。
1KGS|15|7|亚比央 其余的事，凡他所做的，不都写在《犹大列王记》上吗？ 亚比央 常与 耶罗波安 交战。
1KGS|15|8|亚比央 与他祖先同睡，葬在 大卫城 ，他儿子 亚撒 接续他作王。
1KGS|15|9|以色列 王 耶罗波安 第二十年， 亚撒 登基作 犹大 王，
1KGS|15|10|在 耶路撒冷 作王四十一年。他祖母名叫 玛迦 ，是 押沙龙 的女儿。
1KGS|15|11|亚撒 效法他的高祖父 大卫 行耶和华眼中看为正的事，
1KGS|15|12|从国中除去男的庙妓，又除掉他祖先所造的一切偶像。
1KGS|15|13|他甚至废了他祖母 玛迦 太后的位，因 玛迦 造了可憎的 亚舍拉 。 亚撒 砍下她的偶像，在 汲沦溪 边烧了，
1KGS|15|14|只是丘坛还没有废去。 亚撒 一生向耶和华存纯正的心。
1KGS|15|15|亚撒 将他父亲所分别为圣与自己所分别为圣的金银和器皿都奉到耶和华的殿里。
1KGS|15|16|亚撒 和 以色列 王 巴沙 在世的日子常常交战。
1KGS|15|17|以色列 王 巴沙 上来攻击 犹大 ，修筑 拉玛 ，不许人从 犹大 王 亚撒 那里出入。
1KGS|15|18|于是 亚撒 把耶和华殿和王宫府库里所剩下的金银都交在他臣仆手中，派他们到住在 大马士革 的 亚兰 王，就是 希旬 的孙子， 他伯利门 的儿子 便．哈达 那里去，说：
1KGS|15|19|“你父曾与我父立约，我与你也要这样立约。看哪，我把金银送给你作礼物，请你废掉你与 以色列 王 巴沙 所立的约，使他从我这里撤退。”
1KGS|15|20|便．哈达 听从了 亚撒 王，就派遣他的军官去攻打 以色列 的城镇，攻下了 以云 、 但 、 亚伯．伯．玛迦 、全 基尼烈 、 拿弗他利 全地。
1KGS|15|21|巴沙 听见了，就停工不修筑 拉玛 ，仍住在 得撒 。
1KGS|15|22|于是 亚撒 王向 犹大 众人宣布，不准任何人推辞，吩咐他们运走 巴沙 修筑 拉玛 所用的石头和木料。 亚撒 王用它们来修筑 便雅悯 的 迦巴 和 米斯巴 。
1KGS|15|23|亚撒 其余的事，他英勇的事迹，凡他所做的，以及他所建筑的城镇，不都写在《犹大列王记》上吗？只是 亚撒 年老的时候患有脚疾。
1KGS|15|24|亚撒 与他祖先同睡，与他祖先同葬在 大卫城 ，他儿子 约沙法 接续他作王。
1KGS|15|25|犹大 王 亚撒 第二年， 耶罗波安 的儿子 拿答 登基作 以色列 王二年，
1KGS|15|26|拿答 行耶和华眼中看为恶的事，行他父亲所行的道，犯他父亲使 以色列 陷入罪里的那罪。
1KGS|15|27|以萨迦 人 亚希雅 的儿子 巴沙 背叛 拿答 ，在 非利士 人的 基比顿 杀了他，那时 拿答 和 以色列 众人正围困 基比顿 。
1KGS|15|28|犹大 王 亚撒 第三年， 巴沙 杀了 拿答 ，篡了他的位。
1KGS|15|29|巴沙 一作王就杀了 耶罗波安 全家， 耶罗波安 家凡有气息的，一个也没有留下，都杀灭了，正如耶和华藉他仆人 示罗 人 亚希雅 所说的话。
1KGS|15|30|这是因为 耶罗波安 所犯的罪，他使 以色列 陷入罪里，激怒了耶和华－ 以色列 的上帝。
1KGS|15|31|拿答 其余的事，凡他所做的，不都写在《以色列诸王记》上吗？
1KGS|15|32|亚撒 和 以色列 王 巴沙 在世的日子常常交战。
1KGS|15|33|犹大 王 亚撒 第三年， 亚希雅 的儿子 巴沙 在 得撒 登基，作全 以色列 的王二十四年。
1KGS|15|34|他行耶和华眼中看为恶的事，行 耶罗波安 所行的道，犯他使 以色列 陷入罪里的那罪。
1KGS|16|1|耶和华的话临到 哈拿尼 的儿子 耶户 ，责备 巴沙 说：
1KGS|16|2|“我既从尘埃中提拔你，立你作我百姓 以色列 的君王，你竟行 耶罗波安 所行的道，使我的百姓 以色列 陷入罪里，以他们的罪惹我发怒，
1KGS|16|3|看哪，我必除尽 巴沙 和他的家，使你的家像 尼八 的儿子 耶罗波安 的家一样。
1KGS|16|4|凡属 巴沙 的人，死在城中的必被狗吃，死在田野的必被空中的鸟吃。”
1KGS|16|5|巴沙 其余的事，凡他所做的和他英勇的事迹，不都写在《以色列诸王记》上吗？
1KGS|16|6|巴沙 与他祖先同睡，葬在 得撒 ，他儿子 以拉 接续他作王。
1KGS|16|7|耶和华的话临到 哈拿尼 的儿子 耶户 先知，责备 巴沙 和他的家，因他行耶和华眼中看为恶的一切事，以他手所做的惹耶和华发怒，像 耶罗波安 的家一样，又因他杀了 耶罗波安 全家。
1KGS|16|8|犹大 王 亚撒 第二十六年， 巴沙 的儿子 以拉 在 得撒 登基，作 以色列 王二年。
1KGS|16|9|他的大臣 心利 ，就是管理他一半战车的军官背叛他。当他在 得撒 ，在王宫的管家 亚杂 家里喝醉的时候，
1KGS|16|10|心利 进去击杀他，把他杀死，篡了他的位。这是 犹大 王 亚撒 第二十七年的事。
1KGS|16|11|心利 一坐上王位就杀了 巴沙 全家，连他的亲属和朋友，一个男丁也没有留下。
1KGS|16|12|心利 灭绝 巴沙 全家，正如耶和华藉 耶户 先知责备 巴沙 的话。
1KGS|16|13|这是因为 巴沙 和他儿子 以拉 的一切罪，就是他们使 以色列 陷入罪里的那罪，以虚无的神明 惹耶和华－ 以色列 的上帝发怒。
1KGS|16|14|以拉 其余的事，凡他所做的，不都写在《以色列诸王记》上吗？
1KGS|16|15|犹大 王 亚撒 第二十七年， 心利 在 得撒 作王七日。那时军兵正安营围攻 非利士 人的 基比顿 。
1KGS|16|16|军兵在营中听说 心利 已经背叛，杀了王， 以色列 众人当日就在营中立 暗利 元帅作 以色列 王。
1KGS|16|17|暗利 率领 以色列 众人，从 基比顿 上去，围困 得撒 。
1KGS|16|18|心利 见城被攻陷，就进了王宫的堡垒，放火焚烧宫殿，自焚而死。
1KGS|16|19|这是因为他犯罪，行耶和华眼中看为恶的事，行 耶罗波安 所行的道，犯他使 以色列 陷入罪里的那罪。
1KGS|16|20|心利 其余的事和他背叛的事，不都写在《以色列诸王记》上吗？
1KGS|16|21|那时， 以色列 百姓分为两半：一半随从 基纳 的儿子 提比尼 ，要拥立他作王；另一半随从 暗利 。
1KGS|16|22|但随从 暗利 的百姓胜过随从 基纳 儿子 提比尼 的百姓。 提比尼 死了， 暗利 就作了王。
1KGS|16|23|犹大 王 亚撒 第三十一年， 暗利 登基作 以色列 王十二年；他在 得撒 作王六年。
1KGS|16|24|暗利 用二他连得银子向 撒玛 买了 撒玛利亚山 ，在山上建城，按着山的原主 撒玛 的名，给所建的城起名叫 撒玛利亚 。
1KGS|16|25|暗利 行耶和华眼中看为恶的事，比他以前所有的王作恶更严重。
1KGS|16|26|因为他行了 尼八 的儿子 耶罗波安 所行的道，犯他使 以色列 陷入罪里的那罪，以虚无的神明惹耶和华－ 以色列 的上帝发怒。
1KGS|16|27|暗利 其余的事，他所做的和所显出的英勇事迹，不都写在《以色列诸王记》上吗？
1KGS|16|28|暗利 与他祖先同睡，葬在 撒玛利亚 ，他儿子 亚哈 接续他作王。
1KGS|16|29|犹大 王 亚撒 第三十八年， 暗利 的儿子 亚哈 登基作 以色列 王。 暗利 的儿子 亚哈 在 撒玛利亚 作 以色列 王二十二年。
1KGS|16|30|暗利 的儿子 亚哈 行耶和华眼中看为恶的事，比他以前所有的王更严重。
1KGS|16|31|他犯了 尼八 的儿子 耶罗波安 所犯的罪，还当作是小事，又娶了 西顿 王 谒巴力 的女儿 耶洗别 为妻，去事奉 巴力 ，敬拜它，
1KGS|16|32|又在 撒玛利亚 建 巴力庙 ，在庙里为 巴力 筑坛。
1KGS|16|33|亚哈 又造 亚舍拉 ，他所做的惹耶和华－ 以色列 的上帝发怒，比他以前所有的 以色列 王更严重。
1KGS|16|34|亚哈 的日子， 伯特利 人 希伊勒 重修 耶利哥 。立根基的时候，他丧了长子 亚比兰 ；安门的时候，他丧了幼子 西割 ，正如耶和华藉 嫩 的儿子 约书亚 所说的话。
1KGS|17|1|住在 基列 的 提斯比 人 以利亚 对 亚哈 说：“我指着所事奉永生的耶和华－ 以色列 的上帝起誓，这几年我若不祷告，必不降露水，也不下雨。”
1KGS|17|2|耶和华的话临到 以利亚 ，说：
1KGS|17|3|“你离开这里往东去，躲在 约旦河 东边的 基立溪 旁。
1KGS|17|4|你要喝那溪里的水，我已吩咐乌鸦在那里供养你。”
1KGS|17|5|于是 以利亚 去了，他遵照耶和华的话做，去住在 约旦河 东的 基立溪 旁。
1KGS|17|6|乌鸦早上给他叼饼和肉来，晚上也有饼和肉，他又喝溪里的水。
1KGS|17|7|过了些日子溪水干了，因为雨没有下在地上。
1KGS|17|8|耶和华的话临到他，说：
1KGS|17|9|“你起身到 西顿 的 撒勒法 去，住在那里，看哪，我已吩咐那里的一个寡妇供养你。”
1KGS|17|10|以利亚 就起身往 撒勒法 去。他到了城门，看哪，有一个寡妇在那里捡柴。 以利亚 呼唤她说：“请你用器皿取点水来给我喝。”
1KGS|17|11|她去取水的时候， 以利亚 又呼唤她说：“请你手里也拿点饼来给我。”
1KGS|17|12|她说：“我指着永生的耶和华－你的上帝起誓，我没有饼，坛内只有一把面，瓶里只有一点油。看哪，我去找两根柴，带回家为我和我儿子做饼。我们吃了，就等死吧！”
1KGS|17|13|以利亚 对她说：“不要怕！你去照你所说的做吧！只要先为我做一个小饼，拿来给我，然后为你和你的儿子做饼；
1KGS|17|14|因为耶和华－ 以色列 的上帝如此说：‘坛内的面必不用尽，瓶里的油必不短缺，直到耶和华使雨降在地上的日子。’”
1KGS|17|15|妇人就照 以利亚 的话去做。她和 以利亚 ，以及她家中的人，吃了许多日子。
1KGS|17|16|坛内的面果然没有用尽，瓶里的油也不短缺，正如耶和华藉 以利亚 所说的话。
1KGS|17|17|这事以后，那妇人，就是那家的女主人，她的儿子病了，病得很重，甚至没有气息。
1KGS|17|18|妇人对 以利亚 说：“神人哪，我跟你有什么关系，你竟到我这里来，使上帝记起我的罪，以致我的儿子死了呢？”
1KGS|17|19|以利亚 对她说：“把你儿子交给我。” 以利亚 就从妇人怀中接过孩子来，抱到他所住的顶楼，放在自己的床上。
1KGS|17|20|他求告耶和华说：“耶和华－我的上帝啊，我寄居在这寡妇的家里，你却降祸于她，使她的儿子死了吗？”
1KGS|17|21|以利亚 三次伏在孩子的身上，求告耶和华说：“耶和华－我的上帝啊，求你使这孩子的生命归回给他吧！”
1KGS|17|22|耶和华听了 以利亚 的呼求，孩子的生命归回给他，他就活了。
1KGS|17|23|以利亚 把孩子从楼上抱下来，进了房间交给他母亲，说：“看，你的儿子活了！”
1KGS|17|24|妇人对 以利亚 说：“现在我知道你是神人，耶和华藉你口所说的话是真的。”
1KGS|18|1|过了许多日子，到了第三年，耶和华的话临到 以利亚 ，说：“你去，让 亚哈 看见你，我要降雨在地面上。”
1KGS|18|2|以利亚 就去，要让 亚哈 见到他。那时， 撒玛利亚 的饥荒非常严重。
1KGS|18|3|亚哈 召来他的管家 俄巴底 。 俄巴底 非常敬畏耶和华。
1KGS|18|4|耶洗别 杀耶和华先知的时候， 俄巴底 把一百个先知藏了，每五十人藏在一个洞里，拿饼和水供养他们。
1KGS|18|5|亚哈 对 俄巴底 说：“我们要走遍这地，到一切水泉旁和一切溪边，或者能找到青草，可以救活马和骡子，免得丧失一些牲畜。”
1KGS|18|6|于是二人分地巡查， 亚哈 独自走一路， 俄巴底 独自走另一路。
1KGS|18|7|俄巴底 在路上时，看哪， 以利亚 遇见他。 俄巴底 认出他来，就脸伏于地，说：“你是我主 以利亚 吗？”
1KGS|18|8|以利亚 对他说：“我是。你去，告诉你主人说：‘看哪， 以利亚 在这里。’”
1KGS|18|9|俄巴底 说：“仆人犯了什么罪，你竟要把我交在 亚哈 手里，使他杀我呢？
1KGS|18|10|我指着永生的耶和华－你的上帝起誓，无论哪一邦哪一国，我主都派人去找你。若他们说：‘不在这里’，他就叫那邦那国的人起誓说，他们实在找不到你。
1KGS|18|11|现在你说：‘你去告诉你主人说，看哪， 以利亚 在这里’；
1KGS|18|12|恐怕我一离开你，耶和华的灵就把你提到我所不知道的地方去。这样，我去告诉 亚哈 ，他若找不到你，就必杀我。仆人是自幼敬畏耶和华的。
1KGS|18|13|耶洗别 杀耶和华先知的时候，我把耶和华的一百个先知藏了，每五十人藏在一个洞里，拿饼和水供养他们，难道没有人把我做的这事告诉我主吗？
1KGS|18|14|现在你说：‘你去告诉你主人说，看哪， 以利亚 在这里’，他一定会杀我。”
1KGS|18|15|以利亚 说：“我指着所事奉永生的万军之耶和华起誓，我今日要让 亚哈 见到我。”
1KGS|18|16|于是 俄巴底 去迎见 亚哈 ，告诉他这事。 亚哈 就去见 以利亚 。
1KGS|18|17|亚哈 见了 以利亚 ，就说：“真的是你吗？你这使 以色列 遭殃的人！”
1KGS|18|18|以利亚 说：“使 以色列 遭殃的不是我，而是你和你的父家，因为你们离弃耶和华的诫命 ，去随从 巴力 。
1KGS|18|19|现在你要派人去召集 以色列 众人，以及 耶洗别 所供养的四百五十个 巴力 的先知和四百个 亚舍拉 的先知，叫他们都上 迦密山 到我这里来。”
1KGS|18|20|亚哈 就派人到 以色列 众人那里，召集先知上 迦密山 。
1KGS|18|21|以利亚 近前来对众百姓说：“你们心持二意要到几时呢？如果耶和华是上帝，就当顺从耶和华；如果是 巴力 ，就当顺从 巴力 。”百姓一言不答。
1KGS|18|22|以利亚 对百姓说：“作耶和华先知的只剩下我一个； 巴力 的先知却有四百五十人。
1KGS|18|23|请给我们两头牛犊， 巴力 的先知可以为自己挑选一头牛犊，切成小块，放在柴上，不要点火；我也预备一头牛犊放在柴上，也不点火。
1KGS|18|24|你们求告你们神明的名，我也求告耶和华的名。那应允祷告降火的就是上帝。”众百姓回答说：“好主意。”
1KGS|18|25|以利亚 对 巴力 的先知说：“因为你们人多，先挑选一头牛犊，预备好了，求告你们神明的名，却不要点火。”
1KGS|18|26|他们把所给他们的牛犊预备好了，从早晨到中午，求告 巴力 的名说：“ 巴力 啊，求你应允我们！”却没有声音，也没有回应。他们就在所筑的坛四围蹦跳。
1KGS|18|27|到了正午， 以利亚 嘲笑他们，说：“大声求告吧！因为它是神明，它或许在默想，或许正忙着 ，或许在路上，或许在睡觉，它该醒过来了。”
1KGS|18|28|他们大声求告，按着他们的仪式，用刀枪刺割自己，直到浑身流血。
1KGS|18|29|中午过去了，他们狂呼乱叫，直到献晚祭的时候，却没有声音，没有回应的，也没有理睬的。
1KGS|18|30|以利亚 对众百姓说：“你们到我这里来。”众百姓就到他那里，他把那已经毁坏了的耶和华的坛修好。
1KGS|18|31|以利亚 按照 雅各 子孙支派的数目，取了十二块石头；耶和华的话曾临到 雅各 ，说：“你的名要叫 以色列 。”
1KGS|18|32|以利亚 用这些石头为耶和华的名筑一座坛，在坛的四围挖沟，可容纳二细亚谷种。
1KGS|18|33|他又在坛上摆好了柴，把牛犊切成小块放在柴上，说：“你们用四个桶盛满水，倒在燔祭和柴上。”
1KGS|18|34|他又说：“倒第二次。”他们就倒第二次。他又说：“倒第三次。”他们就倒第三次。
1KGS|18|35|水流到坛的四围，沟里也满了水。
1KGS|18|36|到了献晚祭的时候，先知 以利亚 近前来，说：“耶和华－ 亚伯拉罕 、 以撒 、 以色列 的上帝啊，求你今日使人知道你是 以色列 的上帝，我是你的仆人，我遵照你的话做这一切事。
1KGS|18|37|求你应允我，耶和华啊，应允我，使这百姓知道你－耶和华是上帝，是你叫他们回心转意的。”
1KGS|18|38|于是，耶和华降下火来，烧尽燔祭、木柴、石头、尘土，又烧干了沟里的水。
1KGS|18|39|众百姓看见了，就脸伏于地，说：“耶和华是上帝！耶和华是上帝！”
1KGS|18|40|以利亚 对他们说：“拿住 巴力 的先知，不让任何人逃走！”众人就拿住他们。 以利亚 带他们到 基顺河 边，在那里杀了他们。
1KGS|18|41|以利亚 对 亚哈 说：“你现在可以上去吃喝，因为有暴雨的响声了。”
1KGS|18|42|亚哈 就上去吃喝。 以利亚 上了 迦密山 顶，屈身在地，把脸伏在两膝之中。
1KGS|18|43|他对仆人说：“你上去，向海观看。”仆人就上去观看，说：“没有什么。” 以利亚 说：“你再去。”如此七次。
1KGS|18|44|第七次，仆人说：“看哪，有一小片云从海里上来，好像人的手掌那么大。” 以利亚 说：“你上去告诉 亚哈 ，当套车下去，免得被雨阻挡。”
1KGS|18|45|霎时间，天因风云黑暗，降下大雨。 亚哈 就坐上车，往 耶斯列 去了。
1KGS|18|46|耶和华的手按在 以利亚 身上，他就束上腰，奔在 亚哈 前头，一路到 耶斯列 。
1KGS|19|1|亚哈 把 以利亚 一切所做的和他用刀杀众先知的事都告诉 耶洗别 。
1KGS|19|2|耶洗别 就派使者到 以利亚 那里，说：“明日约这时候，我若不使你的性命像那些人的性命一样，愿神明重重惩罚我。”
1KGS|19|3|以利亚 害怕 ，就起来逃命，到了 犹大 的 别是巴 ，把仆人留在那里。
1KGS|19|4|他自己在旷野走了一日的路程，来到一棵罗腾 树下，就坐在那里求死，说：“耶和华啊，现在够了！求你取我的性命吧，因为我不比我的祖先好。”
1KGS|19|5|他躺在罗腾树下睡着了。看哪，有一个天使拍他，对他说：“起来吃吧！”
1KGS|19|6|他观看，看哪，头旁有烧热的石头烤的饼和一壶水，他就吃了喝了，又再躺下。
1KGS|19|7|耶和华的使者回来，第二次拍他，说：“起来吃吧！因为你要走的路很远。”
1KGS|19|8|他就起来吃了喝了，仗着这饮食的力走了四十昼夜，到了上帝的山，就是 何烈山 。
1KGS|19|9|他在那里进了一个洞，在洞中过夜。看哪，耶和华的话临到他，说：“ 以利亚 ，你在这里做什么？”
1KGS|19|10|他说：“我为耶和华－万军之上帝大发热心，因为 以色列 人背弃了你的约，毁坏了你的坛，用刀杀了你的先知，只剩下我一人，他们还要追杀我。”
1KGS|19|11|耶和华说：“你出来站在山上，在耶和华面前。”看哪，耶和华从那里经过。在耶和华面前有烈风大作，山崩石裂，耶和华却不在风中；风后有地震，耶和华也不在其中；
1KGS|19|12|地震后有火，耶和华也不在火中；火以后，有轻微细小的声音。
1KGS|19|13|以利亚 听见，就用外衣蒙脸，出来站在洞口。听啊，有声音向他说：“ 以利亚 ，你在这里做什么？”
1KGS|19|14|他说：“我为耶和华－万军之上帝大发热心，因为 以色列 人背弃了你的约，毁坏了你的坛，用刀杀了你的先知，只剩下我一人，他们还要追杀我。”
1KGS|19|15|耶和华对他说：“去吧，从原路回去，往 大马士革 的旷野去。到了那里，你要膏 哈薛 作 亚兰 王，
1KGS|19|16|又膏 宁示 的孙子 耶户 作 以色列 王，并膏 亚伯．米何拉 人 沙法 的儿子 以利沙 作先知接续你。
1KGS|19|17|将来逃过 哈薛 之刀的，必被 耶户 所杀；逃过 耶户 之刀的，必被 以利沙 所杀。
1KGS|19|18|但我在 以色列 中留下七千人，是未曾向 巴力 屈膝，未曾亲吻 巴力 的。”
1KGS|19|19|于是， 以利亚 离开那里走了，遇见 沙法 的儿子 以利沙 ；他正在耕田，在他前头有十二对牛，自己赶着第十二对。 以利亚 经过他，把自己的外衣搭在他身上。
1KGS|19|20|以利沙 就离开牛，跑到 以利亚 那里，说：“请你让我先与父母吻别，然后我就跟随你。” 以利亚 对他说：“因我对你所做的事，你去吧，然后回来。 ”
1KGS|19|21|以利沙 离开他回去，宰了一对牛，用套牛的器具煮肉给百姓吃，随后就起身跟随 以利亚 ，服事他。
1KGS|20|1|亚兰 王 便．哈达 召集他的全军，率领三十二个王，带着马和战车，上来围困 撒玛利亚 ，要攻打它。
1KGS|20|2|他派使者进城到 以色列 王 亚哈 那里，对他说：“ 便．哈达 如此说：
1KGS|20|3|‘你的金银都要归我，你妻妾儿女中最美的也要归我。’”
1KGS|20|4|以色列 王回答说：“我主我王啊，就照着你的话，我和我所有的都归你。”
1KGS|20|5|使者又来说：“ 便．哈达 如此说：‘我已派人到你那里，要你把你的金银、妻妾、儿女都归我。’
1KGS|20|6|但明日约在这时候，我还要派臣仆到你那里，搜查你的家和你仆人的家，你眼中一切所喜爱的都由他们的手拿走。”
1KGS|20|7|以色列 王召了国内所有的长老来，说：“你们要知道，看哪，这人是来找麻烦的！他派人到我这里来，要我的妻妾、儿女和金银，我并没有拒绝他。”
1KGS|20|8|所有的长老和众百姓对王说：“不要听从他，也不要答应他。”
1KGS|20|9|以色列 王对 便．哈达 的使者说：“你们告诉我主我王说：‘王头一次派人向仆人所要的一切，仆人都依从，但这事我不能依从。’”使者就去回覆 便．哈达 。
1KGS|20|10|便．哈达 又派人到 亚哈 那里，说：“ 撒玛利亚 的尘土若足够跟从我的军兵每人手拿一把，愿神明重重惩罚我！”
1KGS|20|11|以色列 王回答说：“你们告诉他说，‘刚束上腰带的，不要像已卸下的那样夸口。’”
1KGS|20|12|便．哈达 和诸王正在帐幕里喝酒，听见这话，就对他臣仆说：“摆阵吧！”他们就摆阵攻城。
1KGS|20|13|看哪，一个先知靠近 以色列 王 亚哈 ，说：“耶和华如此说：‘这一大群人你看见了吗？看哪，今日我必把他们交在你手里，你就知道我是耶和华。’”
1KGS|20|14|亚哈 说：“藉着谁呢？”他说：“耶和华如此说：‘藉着跟从省长的年轻人。’” 亚哈 说：“谁要开战呢？”他说：“你！”
1KGS|20|15|于是 亚哈 数点跟从省长的年轻人，共二百三十二名，然后又数点 以色列 的众军兵，共七千名。
1KGS|20|16|中午，他们出了城； 便．哈达 和帮助他的三十二个王正在帐幕里畅饮。
1KGS|20|17|跟从省长的年轻人先出城。 便．哈达 派人去，他们回报说：“有人从 撒玛利亚 出来了。”
1KGS|20|18|他说：“他们若为求和出来，要活捉他们，若为打仗出来，也要活捉他们。”
1KGS|20|19|跟从省长的年轻人，和跟随他们的军兵，都出了城，
1KGS|20|20|各人遇见敌人就击杀。 亚兰 人逃跑， 以色列 人追赶他们； 亚兰 王 便．哈达 骑着马和骑兵一同逃跑。
1KGS|20|21|以色列 王出城攻击 马和战车，大大击杀 亚兰 人。
1KGS|20|22|那先知靠近 以色列 王，对他说：“去吧，你当自强，看清楚，也要知道你所要做的事，因为再过一年， 亚兰 王会上来攻击你。”
1KGS|20|23|亚兰 王的臣仆对他说：“他们的神是山神，所以他们胜过我们。但在平原与他们打仗，我们一定胜过他们。
1KGS|20|24|王当做这样的事，把诸王革去，派军官代替他们，
1KGS|20|25|又照着王丧失军兵的数目，再招募一支军队，马补马，车补车。然后在平原与他们打仗，我们一定胜过他们。”王就听臣仆的话，照样去做。
1KGS|20|26|过了一年， 便．哈达 果然召集 亚兰 人上 亚弗 去，要与 以色列 人打仗。
1KGS|20|27|以色列 人也召集军兵，预备食物，去迎战 亚兰 人。 以色列 人对着他们安营，好像两小群的山羊； 亚兰 人却布满了地面。
1KGS|20|28|有神人靠近，对 以色列 王说：“耶和华如此说：‘ 亚兰 人既说我－耶和华是山神，不是平原之神，我必将这一大群人全都交在你手中，你们就知道我是耶和华。’”
1KGS|20|29|以色列 人与 亚兰 人相对安营七日，到第七日两军开战。那一日 以色列 人杀了 亚兰 的十万步兵，
1KGS|20|30|其余的都逃向 亚弗 ，到了城里，城墙倒塌，压死了剩下的二万七千人。 便．哈达 也逃入城内，藏在严密的内室里。
1KGS|20|31|他的臣仆对他说：“看哪，我们听说 以色列 家的王都是仁慈的王；让我们腰束麻布，头套绳索，出去到 以色列 王那里，也许他会存留王的性命。”
1KGS|20|32|于是他们腰束麻布，头套绳索，来到 以色列 王那里，说：“王的仆人 便．哈达 说：‘求王饶我一命。’” 亚哈 说：“他还活着吗？他是我的兄弟。”
1KGS|20|33|这些人正在探测吉凶，就立即抓住他的话说：“ 便．哈达 是王的兄弟！”王说：“你们去请他来。” 便．哈达 出来到王那里，王就请他上车。
1KGS|20|34|便．哈达 对王说：“我父从你父那里所夺的城镇，我必归还给你。你可以在 大马士革 为你自己设立街市，像我父在 撒玛利亚 所设立的一样。” 亚哈 说：“我照此立约，放你回去。”王就与他立约，放了他。
1KGS|20|35|有一个人是先知的门徒，遵照耶和华的话对他同伴说：“你打我吧！”那人不肯打他。
1KGS|20|36|他就对那人说：“你既不听从耶和华的话，看哪，你一离开我，必有狮子咬死你。”那人一离开他，果然遇见狮子，把他咬死了。
1KGS|20|37|先知的门徒又遇见一个人，对他说：“你打我吧！”那人就打他，把他打伤。
1KGS|20|38|那先知就去了，用头巾蒙眼，改了装，在路旁等候王。
1KGS|20|39|王从那里经过，他向王呼叫说：“仆人出战的时候，看哪，有人转过来，带了一个人到我这里来，说：‘你要看守这人，若他真的失踪了，你的性命必代替他的性命，否则，你就要交出一他连得银子来。’
1KGS|20|40|仆人正在到处忙碌的时候，那人就不见了。” 以色列 王对他说：“你自己决定了，就必照样判你。”
1KGS|20|41|他急忙除掉蒙眼的头巾， 以色列 王就认出他是一个先知。
1KGS|20|42|他对王说：“耶和华如此说：‘因你把我决定要消灭的人从你手中放走，所以你的命必代替他的命，你的百姓必代替他的百姓。’”
1KGS|20|43|于是 以色列 王生气，忧闷地回 撒玛利亚 ，到自己的宫去了。
1KGS|21|1|这些事以后，又有一事。 耶斯列 人 拿伯 在 耶斯列 有一个葡萄园，靠近 撒玛利亚 ， 亚哈 王的宫。
1KGS|21|2|亚哈 对 拿伯 说：“把你的葡萄园给我作菜园，因为它靠近我的宫，我就把更好的葡萄园换给你。你若要银子，我就按着价钱给你。”
1KGS|21|3|拿伯 对 亚哈 说：“耶和华不准我把我祖先留下的产业给你。”
1KGS|21|4|亚哈 因 耶斯列 人 拿伯 说“我不把我祖先留下的产业给你”，就生气，忧闷地回宫，躺在床上，脸转向内，也不吃饭。
1KGS|21|5|耶洗别 王后来对他说：“你为什么心里这样生气，不吃饭呢？”
1KGS|21|6|他对王后说：“我向 耶斯列 人 拿伯 说：‘把你的葡萄园按价钱卖给我，或是你愿意，我可以把别的葡萄园换给你。’他却说：‘我不把我的葡萄园给你。’”
1KGS|21|7|耶洗别 王后对王说：“你现在是不是治理 以色列 国呢？只管起来，心里畅畅快快地吃饭，我会把 耶斯列 人 拿伯 的葡萄园给你。”
1KGS|21|8|于是王后以 亚哈 的名义写信，盖上王的印，把信送给那些与 拿伯 同城居住的长老和贵族。
1KGS|21|9|她在信上写着说：“你们当宣告禁食，叫 拿伯 坐在百姓的高位上，
1KGS|21|10|又叫两个无赖坐在 拿伯 对面，作证告他说：‘你诅咒了上帝和王。’然后把他拉出去用石头打死。”
1KGS|21|11|那些与 拿伯 同城居住的长老和贵族，照 耶洗别 送给他们的信去做。正如她送的信上所写，
1KGS|21|12|他们宣告禁食，叫 拿伯 坐在百姓的高位上。
1KGS|21|13|有两个无赖来，坐在 拿伯 对面。无赖当着百姓作证告他说：“ 拿伯 诅咒上帝和王了！”众人就把他拉到城外，用石头打他，他就死了。
1KGS|21|14|于是他们派人到 耶洗别 那里，说：“ 拿伯 被石头打死了。”
1KGS|21|15|耶洗别 听见 拿伯 被石头打死，就对 亚哈 说：“你起来，去取得 耶斯列 人 拿伯 不肯出价卖给你的葡萄园吧！因为 拿伯 不在了，他已经死了。”
1KGS|21|16|亚哈 听见 拿伯 死了，就起来，下去要取得 耶斯列 人 拿伯 的葡萄园。
1KGS|21|17|耶和华的话临到 提斯比 人 以利亚 ，说：
1KGS|21|18|“你起来，去见在 撒玛利亚 的 以色列 王 亚哈 。看哪，他下去要取得 拿伯 的葡萄园，他正在那园里。
1KGS|21|19|你要对他说：‘耶和华如此说：你杀了人，还要取得他的产业吗？’又要对他说：‘耶和华如此说：狗在何处舔 拿伯 的血，狗也必在何处舔你的血。’”
1KGS|21|20|亚哈 对 以利亚 说：“我的仇敌啊，你找到我了吗？”他说：“我找到你了。因为你出卖自己，行了耶和华眼中看为恶的事。
1KGS|21|21|耶和华说：‘看哪，我必使灾祸临到你，把你除灭。 以色列 中凡属 亚哈 的男丁，无论是奴役的、自由的，我都要剪除。
1KGS|21|22|我必使你的家像 尼八 的儿子 耶罗波安 的家，又像 亚希雅 的儿子 巴沙 的家，因为你惹我发怒，又使 以色列 陷入罪里。’
1KGS|21|23|论到 耶洗别 ，耶和华说：‘狗必在 耶斯列 的城郭 吃 耶洗别 。
1KGS|21|24|凡属 亚哈 的人，死在城中的必被狗吃，死在田野的必被空中的鸟吃。’”
1KGS|21|25|（只是从来没有像 亚哈 的，因他受 耶洗别 王后的唆使，出卖自己，行了耶和华眼中看为恶的事。
1KGS|21|26|他行了最可憎的事，随从偶像，正如耶和华在 以色列 人面前赶出的 亚摩利 人所行的一切。）
1KGS|21|27|亚哈 听见这些话，就撕裂衣服，禁食，贴身穿着麻布，也睡在麻布上，沮丧地走来走去。
1KGS|21|28|耶和华的话临到 提斯比 人 以利亚 ，说：
1KGS|21|29|“ 亚哈 在我面前这样谦卑，你看见了吗？因为他在我面前谦卑，所以在他的日子，我不降这祸；到他儿子的时候，我必降这祸于他的家。”
1KGS|22|1|亚兰 和 以色列 之间连续三年没有战争。
1KGS|22|2|到了第三年， 犹大 王 约沙法 下去见 以色列 王。
1KGS|22|3|以色列 王对臣仆说：“你们不知道 基列 的 拉末 是属我们的吗？我们岂可不采取行动，把它从 亚兰 王手里夺回来呢？”
1KGS|22|4|亚哈 问 约沙法 说：“你肯同我去攻打 基列 的 拉末 吗？” 约沙法 对 以色列 王说：“你我不分彼此，我的军队就是你的军队，我的马就是你的马。”
1KGS|22|5|约沙法 对 以色列 王说：“请你先求问耶和华的话。”
1KGS|22|6|于是 以色列 王召集先知，约有四百人，问他们说：“我可以上去攻打 基列 的 拉末 吗？还是不要上去呢？”他们说：“可以上去，因为主必将那城交在王的手里。”
1KGS|22|7|约沙法 说：“这里还有没有耶和华的先知，我们好求问他呢？”
1KGS|22|8|以色列 王对 约沙法 说：“还有一个人，是 音拉 的儿子 米该雅 ，我们可以托他求问耶和华。只是我真的很恨他，因为他对我说预言，从不说吉言，总是说凶信。” 约沙法 说：“请王不要这么说。”
1KGS|22|9|以色列 王召了一个官员来，说：“你快去，把 音拉 的儿子 米该雅 召来。”
1KGS|22|10|以色列 王和 犹大 王 约沙法 在 撒玛利亚 城门前的禾场，各穿朝服，坐在宝座上，所有的先知都在他们面前说预言。
1KGS|22|11|基拿拿 的儿子 西底家 造了铁角，说：“耶和华如此说：‘你要用这些角抵触 亚兰 人，直到将他们灭尽。’”
1KGS|22|12|所有的先知也都这样预言说：“可以上 基列 的 拉末 去，必然得胜，因为耶和华必将那城交在王的手中。”
1KGS|22|13|那去召 米该雅 的使者对他说：“看哪，众先知都异口同声向王说吉言，你也跟他们说一样的话，说吉言吧！”
1KGS|22|14|米该雅 说：“我指着永生的耶和华起誓，耶和华向我说什么，我就说什么。”
1KGS|22|15|米该雅 来到王那里，王问他：“ 米该雅 ，我们可以上去攻打 基列 的 拉末 吗？还是不要上去呢？”他对王说：“你可以上去，必然得胜，耶和华必将那城交在王的手中。”
1KGS|22|16|王对他说：“我要你发誓多少次，你才会奉耶和华的名向我说实话呢？”
1KGS|22|17|米该雅 说：“我看见 以色列 众人散布在山上，如同没有牧人的羊群一般。耶和华说：‘这些人没有主人，他们可以平安地各自回家去。’”
1KGS|22|18|以色列 王对 约沙法 说：“我岂没有告诉你，这人对我说预言，从不说吉言，只说凶信吗？”
1KGS|22|19|米该雅 说：“因此你要听耶和华的话！我看见耶和华坐在宝座上，天上的万军侍立在他左右。
1KGS|22|20|耶和华说：‘谁去引诱 亚哈 上 基列 的 拉末 去阵亡呢？’这个这样说，那个那样说。
1KGS|22|21|随后有一个灵出来，站在耶和华面前，说：‘我去引诱他。’
1KGS|22|22|耶和华问他：‘用什么方法呢？’他说：‘我要出去，在他众先知的口中成为谎言的灵。’耶和华说：‘这样，你去引诱他，必能成功。你出去，照样做吧！’
1KGS|22|23|现在，看哪，耶和华使谎言的灵入了你所有的这些先知的口，并且耶和华已经宣告要降祸于你。”
1KGS|22|24|基拿拿 的儿子 西底家 前来，打 米该雅 一巴掌，说：“耶和华的灵从哪里离开我向你说话呢？”
1KGS|22|25|米该雅 说：“看哪，你进入严密的内室躲藏的那日，就必看见。”
1KGS|22|26|以色列 王说：“把 米该雅 带走，交回给 亚们 市长和 约阿施 王子。
1KGS|22|27|你们要说：‘王如此说，把这个人关在监狱里，使他受苦，吃不饱喝不足，直等到我平安回来。’”
1KGS|22|28|米该雅 说：“你若真的能平安回来，那就是耶和华没有藉我说这话了。”他又说：“众百姓啊，你们都要听！”
1KGS|22|29|以色列 王和 犹大 王 约沙法 上 基列 的 拉末 去。
1KGS|22|30|以色列 王对 约沙法 说：“我要改装上阵，你可以仍穿王袍。” 以色列 王就改装上阵去了。
1KGS|22|31|亚兰 王吩咐他的三十二个战车长说：“你们不要与他们的大将或小兵交战，只要单单攻击 以色列 王。”
1KGS|22|32|那些战车长看见 约沙法 就说：“这一定是 以色列 王！”他们转过去与他交战， 约沙法 就呼喊起来。
1KGS|22|33|战车长见他不是 以色列 王，就转身不追他了。
1KGS|22|34|有一人开弓，并不知情，箭恰巧射入 以色列 王铠甲的缝里。王对驾车的说：“我受重伤了，你掉过车来，载我离开战场！”
1KGS|22|35|那日，战况越来越猛，有人扶着王站在战车上，面对 亚兰 人。到了傍晚，王就死了，血从伤处流入车底。
1KGS|22|36|约在日落的时候，有喊声传遍军中，说：“大家各归本城，各归本地吧！”
1KGS|22|37|王死了，人把他送到 撒玛利亚 ，葬在 撒玛利亚 。
1KGS|22|38|他们在 撒玛利亚 的水池旁洗他的车，有狗来舔他的血，有妓女在那里洗澡，正如耶和华所说的话。
1KGS|22|39|亚哈 其余的事，凡他所做的、他所修造的象牙宫和所建筑的一切城镇，不都写在《以色列诸王记》上吗？
1KGS|22|40|亚哈 与他祖先同睡，他儿子 亚哈谢 接续他作王。
1KGS|22|41|以色列 王 亚哈 第四年， 亚撒 的儿子 约沙法 登基作 犹大 王。
1KGS|22|42|约沙法 登基的时候年三十五岁，在 耶路撒冷 作王二十五年。他母亲名叫 阿苏巴 ，是 示利希 的女儿。
1KGS|22|43|约沙法 效法他父亲 亚撒 所行的道，不偏离左右，行耶和华眼中看为正的事。只是丘坛还没有废去，百姓仍在那里献祭烧香。
1KGS|22|44|约沙法 与 以色列 王和平相处。
1KGS|22|45|约沙法 其余的事和他所行的英勇事迹，以及他的战役，不都写在《犹大列王记》上吗？
1KGS|22|46|约沙法 把他父亲 亚撒 的日子所剩下男的庙妓都从国中除去了。
1KGS|22|47|那时 以东 没有立王，由总督治理。
1KGS|22|48|约沙法 造了 他施 船只，要往 俄斐 去，把金子运来，却没有启航，因为船在 以旬．迦别 毁坏了。
1KGS|22|49|亚哈 的儿子 亚哈谢 对 约沙法 说：“让我的仆人和你的仆人坐船同去吧！” 约沙法 却不肯。
1KGS|22|50|约沙法 与他祖先同睡，与他祖先同葬在 大卫城 ，他儿子 约兰 接续他作王。
1KGS|22|51|犹大 王 约沙法 第十七年， 亚哈 的儿子 亚哈谢 在 撒玛利亚 登基作 以色列 王；他作 以色列 王二年。
1KGS|22|52|他行耶和华眼中看为恶的事，行他父母的道，又行 尼八 的儿子 耶罗波安 的道，使 以色列 陷入罪里。
1KGS|22|53|他事奉 巴力 ，敬拜它，惹耶和华－ 以色列 的上帝发怒，正如他父亲一切所行的。
2KGS|1|1|亚哈 死后， 摩押 背叛 以色列 。
2KGS|1|2|亚哈谢 在 撒玛利亚 ，一日从楼上的栏杆跌下来，就病了。于是他派使者，对他们说：“你们去问 以革伦 的神明 巴力．西卜 ，我这病是否能痊愈。”
2KGS|1|3|但耶和华的使者对 提斯比 人 以利亚 说：“你起来，上去迎见 撒玛利亚 王的使者，对他们说：‘你们去问 以革伦 的神明 巴力．西卜 ，是因为 以色列 中没有上帝吗？’
2KGS|1|4|所以耶和华如此说：‘你必不能下你所上的床，因为你一定会死！’” 以利亚 就去了。
2KGS|1|5|使者回到王那里，王对他们说：“你们为什么回来了呢？”
2KGS|1|6|他们对王说：“有一个人上来迎见我们，对我们说：‘去，回到差你们来的王那里，对他说：耶和华如此说，你派人去问 以革伦 的神明 巴力．西卜 ，是因为 以色列 中没有上帝吗？所以你必不能下所上的床，你一定会死。’”
2KGS|1|7|王对他们说：“上来迎见你们，告诉你们这些话的人是什么样子呢？”
2KGS|1|8|他们对王说：“这人身穿毛衣 ，腰束皮带。”王说：“他一定是 提斯比 人 以利亚 。”
2KGS|1|9|于是，王派了一个五十夫长，带领五十人到 以利亚 那里。他上来，看哪， 以利亚 正坐在山顶上。五十夫长对他说：“神人哪，王吩咐你下来！”
2KGS|1|10|以利亚 回答五十夫长说：“我若是神人，愿火从天上降下来，吞灭你和你的五十个人！”于是有火从天上降下来，吞灭五十夫长和他的五十个人。
2KGS|1|11|王又派另一个五十夫长，带领五十人到 以利亚 那里。五十夫长对他说：“神人哪，王这样吩咐，快快下来！”
2KGS|1|12|以利亚 回答他们说：“我若是神人，愿火从天上降下来，吞灭你和你的五十个人！”于是上帝的火 从天上降下来，吞灭五十夫长和他的五十个人。
2KGS|1|13|王第三次又派一个五十夫长，带领五十人去。第三个五十夫长上去，双膝跪在 以利亚 面前，哀求他说：“神人哪，愿我的性命和你这五十个仆人的性命在你眼中看为宝贵！
2KGS|1|14|看哪，已经有火从天上降下来，吞灭前两次来的五十夫长和他们的五十个人，现在愿我的性命在你眼中看为宝贵！”
2KGS|1|15|耶和华的使者对 以利亚 说：“你跟他下去，不要怕他！” 以利亚 就起来，跟他下到王那里去。
2KGS|1|16|他对王说：“耶和华如此说：‘你派人去问 以革伦 的神明 巴力．西卜 ，是因为 以色列 中没有上帝可以让你求问他的话吗？所以你必不能下所上的床，你一定会死！’”
2KGS|1|17|亚哈谢 死了，正如耶和华藉 以利亚 所说的话。 犹大 王 约沙法 的儿子 约兰 第二年， 亚哈谢 的兄弟 约兰 接续他作王，因 亚哈谢 没有儿子。
2KGS|1|18|亚哈谢 其余所做的事，不都写在《以色列诸王记》上吗？
2KGS|2|1|耶和华要用旋风接 以利亚 升天的时候， 以利亚 与 以利沙 从 吉甲 往前行。
2KGS|2|2|以利亚 对 以利沙 说：“耶和华差遣我往 伯特利 去，你可以留在这里。” 以利沙 说：“我指着永生的耶和华，又指着你的性命起誓，我必不离开你。”于是二人下到 伯特利 。
2KGS|2|3|在 伯特利 的先知的门徒出来，到 以利沙 那里，对他说：“耶和华今日要接你的师父离开你 ，你知不知道？”他说：“我知道，你们不要作声。”
2KGS|2|4|以利亚 对 以利沙 说：“耶和华差遣我往 耶利哥 去，你可以留在这里。” 以利沙 说：“我指着永生的耶和华，又指着你的性命起誓，我必不离开你。”于是二人到了 耶利哥 。
2KGS|2|5|在 耶利哥 的先知的门徒来靠近 以利沙 ，对他说：“耶和华今日要接你的师父离开你，你知不知道？”他说：“我知道，你们不要作声。”
2KGS|2|6|以利亚 对 以利沙 说：“耶和华差遣我往 约旦河 去，你可以留在这里。” 以利沙 说：“我指着永生的耶和华，又指着你的性命起誓，我必不离开你。”于是二人一同往前行。
2KGS|2|7|有五十个先知的门徒同去，远远地站在他们对面；他们二人在 约旦河 边站住。
2KGS|2|8|以利亚 卷起自己的外衣，用来打水，水就左右分开，二人走干地过去。
2KGS|2|9|过去之后， 以利亚 对 以利沙 说：“我未被接去离开你以前，你要我为你做什么，只管求。” 以利沙 说：“愿感动你的灵双倍感动我。”
2KGS|2|10|以利亚 说：“你求的是一件难事。我被接去离开你的时候，你若看见我，就必得着；若不然，就得不着了。”
2KGS|2|11|他们边走边说话的时候，看哪，有火马和火焰车出现，把二人隔开， 以利亚 就乘旋风升天去了。
2KGS|2|12|以利沙 看见，就呼叫说：“我父啊！我父啊！ 以色列 的战车骑兵啊！” 以利沙 不再看见他的时候，就把自己的衣服撕为两片。
2KGS|2|13|他拾起 以利亚 身上掉下来的外衣，回去站在 约旦河 边。
2KGS|2|14|他用 以利亚 身上掉下来的外衣打水，说：“耶和华－ 以利亚 的上帝在哪里呢？”打水之后，水也左右分开， 以利沙 就过去了。
2KGS|2|15|在 耶利哥 的先知的门徒从对面看见他，说：“感动 以利亚 的灵临到 以利沙 身上了。”他们就来迎接他，俯伏于地，向他下拜，
2KGS|2|16|对他说：“看哪，仆人这里有五十个壮士，请你让他们去寻找你师父，或者耶和华的灵将他提起来，投在某山某谷。” 以利沙 说：“你们不必派人去。”
2KGS|2|17|他们再三催促，直到他不好意思，就说：“你们派人去吧！”他们就派了五十个人去，寻找了三天，也没有找着他。
2KGS|2|18|以利沙 仍然留在 耶利哥 ，他们回到他那里，他对他们说：“我不是告诉你们不必去吗？”
2KGS|2|19|耶利哥城 的人对 以利沙 说：“看哪，这城的地势美好，正如我主所看见的，只是水质恶劣，地也没有生产。”
2KGS|2|20|以利沙 说：“你们拿一个新的瓶子来，里面装盐。”他们就拿给他。
2KGS|2|21|他出去到了水源，把盐倒在那里，说：“耶和华如此说：‘我治好了这水，从那里不会再有死亡和不生产的事了。’”
2KGS|2|22|于是那水治好了，直到今日，正如 以利沙 所说的话。
2KGS|2|23|以利沙 从那里上 伯特利 去。正上路的时候，有些孩童从城里出来，讥笑他，对他说：“秃头的，上去吧！秃头的，上去吧！”
2KGS|2|24|他转过身来瞪着他们，奉耶和华的名诅咒他们。于是有两只母熊从林中出来，撕裂他们当中的四十二个孩童。
2KGS|2|25|以利沙 从 伯特利 上 迦密山 ，又从那里回到 撒玛利亚 。
2KGS|3|1|犹大 王 约沙法 第十八年， 亚哈 的儿子 约兰 在 撒玛利亚 登基，作 以色列 王十二年。
2KGS|3|2|他行耶和华眼中看为恶的事，但不致像他父母所行的，因为他除掉他父所造 巴力 的柱像。
2KGS|3|3|然而，他依恋 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的那罪，总不离开。
2KGS|3|4|摩押 王 米沙 牧养许多羊，曾向 以色列 王进贡十万羔羊和十万公绵羊的毛。
2KGS|3|5|亚哈 死后， 摩押 王背叛 以色列 王。
2KGS|3|6|那时 约兰 王出 撒玛利亚 ，数点 以色列 众人。
2KGS|3|7|他向前行，派人到 犹大 王 约沙法 那里，说：“ 摩押 王背叛我，你肯同我去攻打 摩押 吗？” 约沙法 说：“我肯上去，你我不分彼此，我的军队就是你的军队，我的马就是你的马。”
2KGS|3|8|然后 约沙法 说：“我们从哪条路上去呢？” 约兰 说：“从 以东 旷野的路上去。”
2KGS|3|9|于是， 以色列 王和 犹大 王，以及 以东 王，都一同去。他们绕行了七日的路程，军队和所带的牲畜都没有水喝。
2KGS|3|10|以色列 王说：“哀哉！耶和华召集我们这三王，是要交在 摩押 人的手里。”
2KGS|3|11|约沙法 说：“这里不是有耶和华的先知吗？我们可以托他求问耶和华。” 以色列 王的一个大臣回答说：“这里有 沙法 的儿子 以利沙 ，就是从前服事 以利亚 的 。”
2KGS|3|12|约沙法 说：“他必有耶和华的话。”于是 以色列 王、 约沙法 和 以东 王都下去见他。
2KGS|3|13|以利沙 对 以色列 王说：“我跟你有什么关系呢？去问你父亲的先知和你母亲的先知吧！” 以色列 王对他说：“不，因为耶和华召集我们这三王，是要交在 摩押 人的手里。”
2KGS|3|14|以利沙 说：“我指着所事奉永生的万军之耶和华起誓，我若不看 犹大 王 约沙法 的情面，必不理你，不睬你。
2KGS|3|15|现在你们给我找一个弹琴的人来。”弹琴的人弹奏的时候，耶和华的手就按在 以利沙 身上。
2KGS|3|16|他就说：“耶和华如此说：‘你们要在这谷中到处挖沟。’
2KGS|3|17|因为耶和华如此说：‘你们虽不见风，也不见雨，这谷却必满了水，使你们和你们的牛羊牲畜都有水喝。’
2KGS|3|18|在耶和华眼中这还算是小事，他也必将 摩押 人交在你们手中。
2KGS|3|19|你们必攻破一切堡垒和美好的城镇，砍伐各种好树，塞住一切水泉，用石头毁坏一切良田。”
2KGS|3|20|到了早晨，约在献祭的时候，看哪，有水从 以东 而来，遍地就满了水。
2KGS|3|21|摩押 众人听见这三王上来要与他们打仗，凡能束上腰带的，无论老少，都被召集站在边界上。
2KGS|3|22|摩押 人清早起来，日光照在水上，他们看见对面水红如血，
2KGS|3|23|就说：“这是血啊！必是三王互相击杀，全都灭亡了。 摩押 人哪，我们现在去抢夺财物吧！”
2KGS|3|24|摩押 人到了 以色列 营， 以色列 人起来攻打他们，他们就在 以色列 人面前逃跑。 以色列 人追杀 摩押 人，直杀入 摩押 境内 。
2KGS|3|25|他们拆毁 摩押 的城镇，各人抛石头填满一切良田，塞住一切水泉，砍伐各种好树，只剩下 吉珥．哈列设 的石墙，但甩石的兵仍然包围攻打那城。
2KGS|3|26|摩押 王见战事激烈，对他不利，就率领七百个拿刀的兵，想突围逃到 以东 王那里，却没有成功。
2KGS|3|27|于是他在城墙上，把那应当接续他作王的长子献为燔祭。 有极大的愤怒临到 以色列 ，于是三王离开 摩押 王，各自回本地去了。
2KGS|4|1|有个先知门徒的妻子哀求 以利沙 说：“你的仆人，我丈夫死了，他敬畏耶和华是你所知道的。现在有债主来，要带走我的两个孩子给他作奴隶。”
2KGS|4|2|以利沙 对她说：“我可以为你做什么呢？告诉我，你家里有什么？”她说：“婢女家中除了一瓶油之外，什么也没有。”
2KGS|4|3|以利沙 说：“你到外面去向所有的邻舍借器皿，要空的器皿，不要少借。
2KGS|4|4|然后你回家，关上门，你和你儿子在里面把油倒在所有的器皿里，倒满了就放在一边。”
2KGS|4|5|于是妇人离开 以利沙 去了。她关上门，把自己和儿子关在家里。他们把器皿拿给她，她就倒油。
2KGS|4|6|器皿都满了，她对儿子说：“再给我拿器皿来。”儿子对她说：“没有器皿了。”油就止住了。
2KGS|4|7|妇人去告诉神人，神人说：“你去卖了油还债，你和你两个儿子可以靠着所剩的过活。”
2KGS|4|8|一日， 以利沙 经过 书念 ，在那里有一个富有的妇人强留他吃饭。此后， 以利沙 每次经过就转到那里去吃饭。
2KGS|4|9|妇人对丈夫说：“看哪，我知道那常从我们这里经过的是神圣的神人。
2KGS|4|10|我们可以为他盖一间有墙的小阁楼，里面安放床榻、桌子、椅子、灯台。每当他来到我们这里，就可以住在那里。”
2KGS|4|11|一日， 以利沙 来到那里，转进那阁楼，躺卧在那里。
2KGS|4|12|以利沙 吩咐仆人 基哈西 说：“你叫这 书念 妇人来。”他把妇人叫了来，妇人就站在 以利沙 面前。
2KGS|4|13|以利沙 吩咐仆人说：“你对她说：‘看哪，你为我们费了许多心思，我可以为你做什么呢？我可以为你向王或元帅求什么呢？’”她说：“我已住在自己百姓之中。”
2KGS|4|14|以利沙 说：“究竟可以为她做什么呢？” 基哈西 说：“她真的没有儿子，她丈夫也老了。”
2KGS|4|15|以利沙 说：“叫她回来。”于是他叫了她来，她就站在门口。
2KGS|4|16|以利沙 说：“明年这时候 ，你必抱一个儿子。”她说：“神人，我主啊，不要这样欺哄婢女。”
2KGS|4|17|妇人果然怀孕，到了明年那时候，生了一个儿子，正如 以利沙 向她所说的。
2KGS|4|18|孩子长大，一日出去到他父亲和收割的人那里。
2KGS|4|19|他对父亲说：“我的头啊，我的头啊！”他父亲对仆人说：“把他抱到他母亲那里。”
2KGS|4|20|仆人抱去，交给他母亲。孩子坐在母亲的膝上，到中午就死了。
2KGS|4|21|他母亲上去，把他放在神人的床上，关了门出来，
2KGS|4|22|呼叫她丈夫说：“你叫一个仆人给我牵一匹驴来，我要赶去见神人，然后回来。”
2KGS|4|23|丈夫说：“今日不是初一，也不是安息日，你为何要到他那里去呢？”妇人说：“平安无事。”
2KGS|4|24|于是她备上驴，对仆人说：“走，赶紧走，除非我吩咐你，不要为了我而慢下来。”
2KGS|4|25|妇人往 迦密山 去，到了神人那里。 神人远远看见她，对仆人 基哈西 说：“看哪， 书念 的妇人来了！
2KGS|4|26|现在你跑去迎接她，对她说，你平安吗？你丈夫平安吗？孩子平安吗？”她说：“平安。”
2KGS|4|27|妇人上了山，到神人那里，就抱住神人的脚。 基哈西 前来要推开她，神人说：“由她吧！因为她心里愁苦。但耶和华向我隐瞒这事，没有告诉我。”
2KGS|4|28|妇人说：“我何尝向我主求过儿子呢？我岂不是说过，不要欺哄我吗？”
2KGS|4|29|以利沙 吩咐 基哈西 说：“你束上腰，手拿我的杖前去。若遇见人，不要向他问安，人若向你问安，也不要回答。要把我的杖放在孩子脸上。”
2KGS|4|30|孩子的母亲说：“我指着永生的耶和华，又指着你的性命起誓，我必不离开你。”于是 以利沙 起身，随着她去了。
2KGS|4|31|基哈西 在他们以先去了，把杖放在孩子脸上，却没有声音，也没有动静。 基哈西 回去，迎见 以利沙 ，告诉他说：“孩子还没有醒过来。”
2KGS|4|32|以利沙 进了屋子，看哪，孩子死了，放在自己的床上。
2KGS|4|33|他进去，关上门，只有他们两个人，他就向耶和华祈祷。
2KGS|4|34|他上去伏在孩子身上，口对口，眼对眼，手对手。他伏在孩子身上，孩子的身体就渐渐暖和了。
2KGS|4|35|然后他下来，在屋里来回走了一趟，又上去伏在孩子身上。孩子打了七个喷嚏，眼睛就睁开了。
2KGS|4|36|以利沙 叫 基哈西 说：“你叫这 书念 妇人来。”于是他叫了她来。妇人来到 以利沙 那里， 以利沙 说：“把你儿子抱起来。”
2KGS|4|37|妇人就进来，在 以利沙 脚前俯伏于地，向他下拜，然后抱起她儿子出去了。
2KGS|4|38|以利沙 回到 吉甲 ，那地正有饥荒。先知的门徒坐在他面前，他吩咐仆人说：“你把大锅放在火上，给先知的门徒熬汤。”
2KGS|4|39|有一个人去到田野摘菜，发现一棵野瓜藤，就摘了满满一兜的野瓜回来，切了放进熬汤的锅中，并不知道那是什么。
2KGS|4|40|他们把汤倒出来给大家吃。他们吃汤里东西的时候，喊叫说：“神人哪，锅子里的东西会死人！”所以他们不能吃了。
2KGS|4|41|以利沙 说：“拿点面来。”他把面撒在锅中，说：“倒出来，给大家吃吧！”锅中就没有毒了。
2KGS|4|42|有一个人从 巴力．沙利沙 来，带着初熟果子的食物、二十个大麦做的饼和新麦穗，装在袋子里送给神人。神人说：“把这些给大家吃。”
2KGS|4|43|仆人说：“这些岂可摆在一百人面前呢？” 以利沙 说：“你只管给大家吃吧！因为耶和华如此说，他们必吃了，还有剩下的。”
2KGS|4|44|仆人就摆在他们面前，他们吃了，还有剩下，正如耶和华所说的。
2KGS|5|1|亚兰 王的元帅 乃缦 在他主人面前是一个伟大的人，得王的喜悦，因为耶和华曾藉他使 亚兰 人得胜。他虽然是大能的勇士，却染上了痲疯 。
2KGS|5|2|亚兰 人成群出征的时候，从 以色列 地掳了一个小女孩，她就服事 乃缦 的妻子。
2KGS|5|3|她对女主人说：“我希望主人去见 撒玛利亚 的先知，他必能治好主人的痲疯。”
2KGS|5|4|乃缦 去告诉他主人说，从 以色列 地来的女孩如此如此说。
2KGS|5|5|亚兰 王说：“你可以去，我也会送信给 以色列 王。”于是 乃缦 手里带十他连得银子、六千舍客勒金子和十套衣裳去了。
2KGS|5|6|他带着这信给 以色列 王，说：“现在你接到这信，看哪，我派臣仆 乃缦 到你这里来，你要治好他的痲疯。”
2KGS|5|7|以色列 王读了信就撕裂衣服，说：“我岂是上帝，能使人死使人活呢？这人竟派人来，叫我治好一个人的痲疯。你们要知道，看，这人是找机会来跟我吵架的。”
2KGS|5|8|神人 以利沙 听见 以色列 王撕裂衣服，就派人到王那里，说：“你为什么撕裂衣服呢？让那人到我这里来，他会知道 以色列 中有先知。”
2KGS|5|9|于是 乃缦 带着车马到了 以利沙 的家，站在门前。
2KGS|5|10|以利沙 派一个使者，对 乃缦 说：“去，在 约旦河 中沐浴七次，你的肉就必复原，你会得洁净。”
2KGS|5|11|乃缦 却发怒走了。他说：“看哪，我以为他必定会出来，到我这里，站着求告耶和华－他上帝的名，在患处上摇手，治好这痲疯。
2KGS|5|12|大马士革 的 亚玛拿河 和 法珥法河 岂不比 以色列 的一切水更好吗？我难道不可以在那里沐浴而得洁净吗？”于是他生气，转身走了。
2KGS|5|13|他的仆人近前来，对他说：“我父啊，先知若吩咐你做一件大事，你岂不做吗？何况是吩咐你去沐浴，得洁净呢？”
2KGS|5|14|于是 乃缦 下去，照着神人的话，在 约旦河 里浸了七次。他的肉复原，好像小孩的肉，他就洁净了。
2KGS|5|15|乃缦 带着所有跟随他的人，回到神人那里，站在他面前，说：“看哪，我知道，除了 以色列 ，全地没有上帝。现在请你收下仆人的礼物。”
2KGS|5|16|以利沙 说：“我指着所事奉永生的耶和华起誓，我必不接受。” 乃缦 再三请他收下，他却不肯。
2KGS|5|17|乃缦 说：“你若不肯，请把两匹骡子能驮的土赐给仆人，仆人必不再把燔祭或祭物献给别神，只献给耶和华。
2KGS|5|18|惟有一件事，愿耶和华饶恕你仆人：我主人进 临门 庙在那里叩拜的时候，他总是扶着我的手，所以我也在 临门 庙叩拜。我在 临门 庙叩拜的这事，愿耶和华饶恕你仆人。”
2KGS|5|19|以利沙 对他说：“你平安地回去吧！” 乃缦 离开他去了。走了一小段路，
2KGS|5|20|神人 以利沙 的仆人 基哈西 说：“看哪，我主人不愿从这 亚兰 人 乃缦 手里接受他带来的礼物，我指着永生的耶和华起誓，我必跑去追上他，向他拿些东西。”
2KGS|5|21|于是 基哈西 去追 乃缦 。 乃缦 看见有人追来，就下车迎着他，说：“都平安吗？”
2KGS|5|22|他说：“都平安！我主人派我来说：‘看哪，现在有两个年轻人，是先知的门徒，从 以法莲 山区来到我这里，请你给他们一他连得银子，两套衣裳。’”
2KGS|5|23|乃缦 说：“好啊，请收下二他连得。”他再三请求，就把二他连得银子装在两个袋子里，连同两套衣裳交给两个仆人；他们就在 基哈西 前头抬着走。
2KGS|5|24|到了山冈， 基哈西 从他们手中接过来，放在屋里，打发这些人走了。
2KGS|5|25|基哈西 进去，站在主人面前。 以利沙 对他说：“ 基哈西 ，你从哪里来？”他说：“仆人哪里也没去。”
2KGS|5|26|以利沙 对他说：“那人下车转过来迎着你的时候，我的心岂没有去呢？这岂是接受银子，接受衣裳、橄榄园、葡萄园、牛羊、仆婢的时候呢？
2KGS|5|27|因此， 乃缦 的痲疯必紧随你和你的后裔，直到永远。” 基哈西 从 以利沙 面前出去，就长了痲疯，像雪一样。
2KGS|6|1|先知的门徒对 以利沙 说：“看哪，我们在你面前居住的地方，那里对我们太窄小了。
2KGS|6|2|让我们往 约旦河 去，各人从那里取一根木料，在那里为自己建造居住的地方。”他说：“你们去吧！”
2KGS|6|3|有一人说：“请你与仆人同去。”他说：“我可以去。”
2KGS|6|4|于是 以利沙 与他们同去。到了 约旦河 ，他们砍伐树木。
2KGS|6|5|有一人砍树的时候，斧子的头掉在水里，他就喊着说：“不好了！我主啊，斧子是借来的。”
2KGS|6|6|神人说：“掉在哪里了？”他把那地方指给 以利沙 看。 以利沙 砍了一块木头，抛在水里，就使斧子的头浮上来了。
2KGS|6|7|以利沙 说：“拿起来吧！”那人就伸手拿起来了。
2KGS|6|8|亚兰 王与 以色列 作战，他和臣仆商议说：“我要在某处某处安营 。”
2KGS|6|9|神人派人到 以色列 王那里，说：“你要小心，不要从某处经过，因为 亚兰 人下到那里去了。”
2KGS|6|10|以色列 王派人到神人告诉他的地方去。神人警告他，他就在那里有所防备，不止一两次。
2KGS|6|11|亚兰 王因这事心里气愤，召了臣仆来，对他们说：“我们当中有谁帮助 以色列 王，你们不告诉我吗？”
2KGS|6|12|有一个臣仆说：“不，我主，我王！只有 以色列 中的先知 以利沙 ，把王在卧房所说的话告诉 以色列 王。”
2KGS|6|13|王说：“你们去查看他在哪里，我好派人去捉拿他。”有人告诉王说：“看哪，他在 多坍 。”
2KGS|6|14|王就派遣车马和大军往那里去，夜间他们到了，围困那城。
2KGS|6|15|神人的仆人清早起来出去，看哪，车马军兵围困了城。仆人对神人说：“不好了！我主啊，我们该怎么办呢？”
2KGS|6|16|神人说：“不要惧怕！因与我们同在的比与他们同在的更多。”
2KGS|6|17|以利沙 祷告说：“耶和华啊，求你开他的眼目，使他能看见。”耶和华开了这年轻人的眼目，他就看见了，看哪，满山有火马和火焰车围绕 以利沙 。
2KGS|6|18|亚兰 人下到 以利沙 那里， 以利沙 向耶和华祷告说：“求你击打这国，使他们眼目失明。”耶和华就照 以利沙 的话，击打他们，使他们眼目失明。
2KGS|6|19|以利沙 对他们说：“这不是那条路，也不是那座城。你们跟我走，我必领你们到你们要寻找的人那里。”于是他领他们到了 撒玛利亚 。
2KGS|6|20|他们进了 撒玛利亚 ， 以利沙 说：“耶和华啊，求你开这些人的眼目，使他们能看见。”耶和华开了他们的眼目，他们就看见了，看哪，是在 撒玛利亚城 中。
2KGS|6|21|以色列 王看见他们，就对 以利沙 说：“我父啊，我真的可以击杀他们吗？”
2KGS|6|22|他说：“不可击杀！这些人岂是你用刀用弓掳来给你击杀的呢？当在他们面前摆设饮食给他们吃喝，让他们回到他们主人那里。”
2KGS|6|23|王为他们预备了盛大的宴席。他们吃喝完了，王就送他们回到他们主人那里。此后， 亚兰 的军队不再侵犯 以色列 地了。
2KGS|6|24|此后， 亚兰 王 便．哈达 召集他的全军，上来围困 撒玛利亚 。
2KGS|6|25|看哪，被围困的时候， 撒玛利亚 有大饥荒，甚至一个驴头值八十舍客勒，四分之一卡布 的鸽子粪值五舍客勒。
2KGS|6|26|一日， 以色列 王在城墙上经过，有一个妇人向他呼叫说：“我主，我王啊！求你帮助。”
2KGS|6|27|王说：“耶和华不帮助你，我从哪里帮助你呢？是从禾场，或从压酒池吗？”
2KGS|6|28|王对妇人说：“你有什么事？”她说：“这妇人对我说：‘把你的儿子交出来，我们今日可以吃他，明日可以吃我的儿子。’
2KGS|6|29|我们就煮了我的儿子吃了。次日我对她说：‘要把你的儿子交出来，我们可以吃。’她却把她的儿子藏起来。”
2KGS|6|30|王听见妇人的话，就撕裂衣服；那时，王在城墙上经过，百姓看见了，看哪，王贴身穿着麻布。
2KGS|6|31|王说：“我今日若容许 沙法 的儿子 以利沙 的头还留在他身上，愿上帝重重惩罚我！”
2KGS|6|32|那时， 以利沙 正坐在家中，有长老与他同坐。王派一个人先去，使者还没有到， 以利沙 对长老说：“你们看，这凶手之子派人来斩我的头。你们注意，当使者来到，你们就关上门，把他关在门外。在他后头不就是他主人的脚步声吗？”
2KGS|6|33|正与他们说话的时候，看哪，使者 下到他那里，说：“看哪，这灾祸是从耶和华来的，我何必再仰望耶和华呢？”
2KGS|7|1|以利沙 说：“你们要听耶和华的话，耶和华如此说：明日约这时候，在 撒玛利亚 城门口，一细亚细面只卖一舍客勒，二细亚大麦也卖一舍客勒。”
2KGS|7|2|有一个搀扶王的军官回答神人说：“看哪，即使耶和华打开天上的窗户，也不可能有这事。” 以利沙 说：“看哪，你必亲眼看见，在那里却吃不到什么。”
2KGS|7|3|在城门口有四个长痲疯的人，他们彼此说：“我们为何坐在这里等死呢？
2KGS|7|4|我们若说要进城去，城里有饥荒，我们必死在那里。若我们在这里坐着不动，也必死。现在，来吧，我们去向 亚兰 人的军队投降。若他们饶我们的命，我们就活着；若杀我们，我们就死吧！”
2KGS|7|5|黄昏的时候，他们起来往 亚兰 人的军营去；到了营边，看哪，没有一人在那里。
2KGS|7|6|因为主使 亚兰 人的军队听见战车战马的声音，大军的声音，他们就彼此说：“看哪，这必是 以色列 王雇用 赫 人诸王和 埃及 诸王来攻击我们。”
2KGS|7|7|所以，在黄昏的时候他们起来逃跑，撇下帐棚、马、驴，把军营留在原处，只顾逃命。
2KGS|7|8|那些长痲疯的人到了营边，进了一座帐棚，吃了喝了，从当中拿走金银和衣服，收藏起来。他们又回来，进了另一座帐棚，从当中拿走财物去收藏。
2KGS|7|9|那时，他们彼此说：“我们所做的不对了！这一天是有好消息的日子，我们竟不作声！若等到天亮，我们就有罪了。现在，来，我们去向王室报信吧！”
2KGS|7|10|他们就去叫守城门的人，告诉他们说：“我们到了 亚兰 人的军营，看哪，没有一人在那里，也无人声，只有拴着的马和驴，帐棚都留在原处。”
2KGS|7|11|守城门的人就呼叫，他们向城内的王室报信。
2KGS|7|12|王夜间起来，对臣仆说：“我告诉你们 亚兰 人向我们做的事。他们知道我们饥饿，所以离营，埋伏在田野，说：‘ 以色列 人出城的时候，我们活捉他们，我们就可以进到城里去。’”
2KGS|7|13|王的一个臣仆回答说：“不如叫人从城里剩下的马中取五匹，看哪，这些马像 以色列 大众一样 ，快要灭亡了；我们派人去窥探吧！”
2KGS|7|14|于是他们取了两辆车和马，王派人去跟踪 亚兰 人的军队，说：“你们去窥探吧。”
2KGS|7|15|他们去跟踪 亚兰 人，直到 约旦河 。看哪，整条路上都是 亚兰 人匆忙逃跑时所丢弃的衣服和器具，使者就回来向王报告。
2KGS|7|16|百姓就出去，掳掠 亚兰 人的军营。于是一细亚细面只卖一舍客勒，二细亚大麦也卖一舍客勒，正如耶和华所说的。
2KGS|7|17|王派搀扶他的那军官在城门指挥，百姓在城门把他踩死了，正如神人在王下到他那里的时候所说的。
2KGS|7|18|神人曾对王说：“明日约这时候，在 撒玛利亚 城门口，二细亚大麦只卖一舍客勒，一细亚细面也卖一舍客勒。”
2KGS|7|19|那军官回答神人说：“看哪，即使耶和华打开天上的窗户，也不可能有这事。”神人说：“看哪，你必亲眼看见，在那里却吃不到什么。”
2KGS|7|20|这话果然应验在他身上，因为百姓在城门把他踩死了。
2KGS|8|1|以利沙 曾对他救活的孩子的母亲说：“你和你的全家要起身，往你可住的地方去住，因为耶和华已令饥荒降在这地七年。”
2KGS|8|2|妇人就起身，照神人的话去做，带着全家往 非利士 人的地去，寄居了七年。
2KGS|8|3|过了七年，那妇人从 非利士 人的地回来，就出去为自己的房屋田地哀求王。
2KGS|8|4|那时王正与神人的仆人 基哈西 谈话，说：“你把 以利沙 所做的一切大事告诉我。”
2KGS|8|5|基哈西 告诉王 以利沙 如何使死人复活，看哪， 以利沙 所救活的孩子的母亲正为自己的房屋田地来哀求王。 基哈西 说：“我主我王，这就是那妇人，这是她的儿子，就是 以利沙 所救活的。”
2KGS|8|6|王问那妇人，她就把事情告诉王。于是王为她派一个官员，说：“凡属这妇人的都还给她，自从她离开本地直到今日，她田地的出产也都还给她。”
2KGS|8|7|以利沙 来到 大马士革 ， 亚兰 王 便．哈达 正患病。有人告诉王说：“神人来到这里了。”
2KGS|8|8|王就吩咐 哈薛 说：“你带着礼物去见神人，托他求问耶和华，我这病能不能好？”
2KGS|8|9|于是 哈薛 用四十匹骆驼，驮着 大马士革 的各样美物为礼物，去迎见 以利沙 。 哈薛 到了那里，站在他面前，说：“你儿子 亚兰 王 便．哈达 派我到你这里，问说：‘我这病会不会好？’”
2KGS|8|10|以利沙 对 哈薛 说：“你回去告诉他说：‘你一定会好。’但耶和华指示我，他必定会死。”
2KGS|8|11|神人定睛看着 哈薛 ，直到他感到羞愧。神人就哭了。
2KGS|8|12|哈薛 说：“我主为什么哭？”他说：“因为我知道你必虐待 以色列 人，用火焚烧他们的堡垒，用刀杀死他们的壮丁，摔死他们的婴孩，剖开他们的孕妇。”
2KGS|8|13|哈薛 说：“仆人算什么，不过是一条狗，怎么能行这大事呢？” 以利沙 说：“耶和华指示我，你必作 亚兰 王。”
2KGS|8|14|哈薛 离开 以利沙 ，回到他主人那里。主人对他说：“ 以利沙 对你说了什么？”他说：“他告诉我你必能好。”
2KGS|8|15|次日， 哈薛 拿被子浸在水中，蒙住王的脸，王就死了。于是 哈薛 篡了他的位。
2KGS|8|16|亚哈 的儿子 以色列 王 约兰 第五年－ 约沙法 曾作 犹大 王 － 犹大 王 约沙法 的儿子 约兰 登基作了 犹大 王。
2KGS|8|17|约兰 登基的时候年三十二岁，在 耶路撒冷 作王八年。
2KGS|8|18|他行 以色列 诸王的道，正如 亚哈 家所行的，因他娶了 亚哈 的女儿为妻，行耶和华眼中看为恶的事。
2KGS|8|19|耶和华却因他仆人 大卫 的缘故，不肯灭绝 犹大 ，要照他所应许的，永远赐灯光给 大卫 和他的子孙。
2KGS|8|20|约兰 在位期间， 以东 背叛，自己立王治理他们，脱离 犹大 的权势。
2KGS|8|21|约兰 率领他所有的战车过到 撒益 去。他夜间起来，攻打围困他的 以东 人和战车长； 犹大 军兵逃跑，各回自己的帐棚去了；
2KGS|8|22|这样， 以东 背叛，脱离 犹大 的管辖，直到今日。那时 立拿 也背叛了。
2KGS|8|23|约兰 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
2KGS|8|24|约兰 与他祖先同睡，与他祖先同葬在 大卫城 ，他儿子 亚哈谢 接续他作王。
2KGS|8|25|亚哈 的儿子 以色列 王 约兰 第十二年， 犹大 王 约兰 的儿子 亚哈谢 登基。
2KGS|8|26|他登基的时候年二十二岁，在 耶路撒冷 作王一年。他母亲名叫 亚她利雅 ，是 以色列 王 暗利 的孙女。
2KGS|8|27|亚哈谢 行 亚哈 家的道，行耶和华眼中看为恶的事，与 亚哈 家一样，因为他是 亚哈 家的女婿。
2KGS|8|28|他与 亚哈 的儿子 约兰 同往 基列 的 拉末 去，与 亚兰 王 哈薛 交战。 亚兰 人打伤了 约兰 ，
2KGS|8|29|约兰 王回到 耶斯列 ，医治在 拉末 与 亚兰 王 哈薛 打仗时，被 亚兰 人击打所受的伤。 约兰 的儿子 犹大 王 亚哈谢 因为 亚哈 的儿子 约兰 病了，就下到 耶斯列 看望他。
2KGS|9|1|以利沙 先知叫了一个先知的门徒来，吩咐他：“你束上腰，手拿这瓶膏油往 基列 的 拉末 去。
2KGS|9|2|你到了那里，要在那里寻找 宁示 的孙子， 约沙法 的儿子 耶户 。你去，使他从弟兄中起来，带他进最里面的内室，
2KGS|9|3|把瓶里的膏油倒在他头上，说：‘耶和华如此说：我膏你作 以色列 王。’然后你就开门逃跑，不要等候。”
2KGS|9|4|于是那青年，那年轻的先知往 基列 的 拉末 去了。
2KGS|9|5|他到了那里，看哪，众军官都坐着，就说：“长官，我有话对你说。” 耶户 说：“你要对我们哪一个说呢？”他说：“长官，我要对你说。”
2KGS|9|6|耶户 就起来，进了内室，那青年把膏油倒在他头上，对他说：“耶和华－ 以色列 的上帝如此说：‘我膏你作耶和华百姓 以色列 的王。
2KGS|9|7|你要击杀你主人 亚哈 的全家，我好在 耶洗别 身上，为我仆人众先知和耶和华所有仆人的血伸冤。
2KGS|9|8|亚哈 全家都必灭亡，凡属 亚哈 的男丁，无论是奴役的、自由的，我必从 以色列 中剪除。
2KGS|9|9|我必使 亚哈 的家像 尼八 儿子 耶罗波安 的家，又像 亚希雅 儿子 巴沙 的家。
2KGS|9|10|至于 耶洗别 ，狗必在 耶斯列 田里吃她，无人埋葬。’”于是那青年就开门逃跑了。
2KGS|9|11|耶户 出来，回到他主人的臣仆那里，有一人问他说：“平安吗？这疯狂的人为什么到你这里来呢？”他对他们说：“你们认得那人，也知道他在胡说。”
2KGS|9|12|他们说：“说谎！告诉我们吧。”他说：“他如此如此对我说：‘耶和华如此说：我膏你作 以色列 的王。’”
2KGS|9|13|他们各人就急忙把自己的衣服铺在台阶的上层，在 耶户 的下面；他们吹角，说：“ 耶户 作王了！”
2KGS|9|14|这样， 宁示 的孙子， 约沙法 的儿子 耶户 背叛了 约兰 。先前 约兰 和 以色列 众人因为 亚兰 王 哈薛 的缘故，把守 基列 的 拉末 。
2KGS|9|15|后来 约兰 王回到 耶斯列 ，医治他与 亚兰 王 哈薛 打仗时，被 亚兰 人击打所受的伤。 耶户 说：“若你们有这样的意思，就不要让人溜出城，到 耶斯列 去报信。”
2KGS|9|16|于是 耶户 驾战车往 耶斯列 去，因为 约兰 卧病在那里。 犹大 王 亚哈谢 已经下去看望他。
2KGS|9|17|有一个守望的人站在 耶斯列 的城楼上，看见 耶户 带着一队人来，就说：“我看见一队人。” 约兰 说：“派一个骑兵去迎接他们，问说：‘平安吗？’”
2KGS|9|18|骑兵就去迎接 耶户 ，说：“王如此说：‘平安吗？’”耶户说：“平安不平安跟你有什么关系呢？转身跟在我后面吧！”守望的人说：“使者到了他们那里，却不回来。”
2KGS|9|19|王又派第二个骑兵去。这人到了他们那里，说：“王如此说：‘平安吗？’” 耶户 说：“平安不平安跟你有什么关系呢？转身跟在我后面吧！”
2KGS|9|20|守望的人又说：“他到了他们那里，也不回来。车驾得很凶猛，好像 宁示 的孙子 耶户 在驾车。”
2KGS|9|21|约兰 吩咐说：“套车！”人就给他套车。 以色列 王 约兰 和 犹大 王 亚哈谢 各坐自己的车出去迎接 耶户 ，在 耶斯列 人 拿伯 的田那里遇见他。
2KGS|9|22|约兰 见 耶户 就说：“ 耶户 ，平安吗？” 耶户 说：“你母亲 耶洗别 的淫行邪术这样多，怎么能平安呢？”
2KGS|9|23|约兰 用手转过车来逃跑，对 亚哈谢 说：“ 亚哈谢 啊，反了！”
2KGS|9|24|耶户 全力拉弓，射中 约兰 两臂中间，箭从心窝穿出， 约兰 就仆倒在车上。
2KGS|9|25|耶户 对他的军官 毕甲 说：“把他抛在 耶斯列 人 拿伯 的田里。你当记得，你我一同驾车跟随他父亲 亚哈 的时候，耶和华对 亚哈 说了预言，
2KGS|9|26|耶和华说：‘我昨日看见 拿伯 的血和他众子的血，我发誓我必在这块田上报应你。’这是耶和华说的。现在你要照着耶和华的话，把他抛在这田里。”
2KGS|9|27|犹大 王 亚哈谢 看见了，就沿着 伯．哈干 的路逃跑。 耶户 追赶他，说：“把这人也击杀在车上，在靠近 以伯莲 的 姑珥 坡上 。”他逃到 米吉多 ，就死在那里。
2KGS|9|28|他的臣仆用车把他的尸体运回 耶路撒冷 ，与他祖先同葬在 大卫城 ，他自己的坟墓里。
2KGS|9|29|亚哈 的儿子 约兰 第十一年， 亚哈谢 登基作了 犹大 王。
2KGS|9|30|耶户 到了 耶斯列 。 耶洗别 听见了，就画眼影、梳头，从窗户往外观看。
2KGS|9|31|耶户 进了城门， 耶洗别 说：“杀主人的 心利 啊，平安吗？”
2KGS|9|32|耶户 向窗户抬头，说：“有谁顺从我？谁？”有两三个太监向外看他。
2KGS|9|33|耶户 说：“把她抛下来！”他们就把她抛下来。她的血溅在墙上和马上， 耶户 践踏在她身上。
2KGS|9|34|耶户 进去，吃了喝了，说：“你们去处理这被诅咒的妇人，埋了她，因为她是王的女儿。”
2KGS|9|35|他们去了，要埋葬她，却只找到她的头骨和脚，以及手掌。
2KGS|9|36|他们回来报告 耶户 ， 耶户 说：“这正应验耶和华藉他仆人 提斯比 人 以利亚 所说的话，说：‘在 耶斯列 田里，狗必吃 耶洗别 的肉，
2KGS|9|37|耶洗别 的尸体必在 耶斯列 田里的地面上如同粪土，甚至没有人可说：这是 耶洗别 。’”
2KGS|10|1|亚哈 有七十个儿子在 撒玛利亚 。 耶户 写信送到 撒玛利亚 ，给 耶斯列 的领袖和长老 ，以及教养 亚哈 众儿子的人，说：
2KGS|10|2|“你们主人的众儿子既然在你们那里，你们又有战车、马匹、兵器、坚固城，现在你们接了这信，
2KGS|10|3|可以在你们主人的众儿子中选一个贤能正直的，使他坐他父亲的王位，你们也可以为你们主人的家作战。”
2KGS|10|4|他们却非常惧怕，说：“看哪，两个王在他面前尚且站立不住，我们怎能站立得住呢？”
2KGS|10|5|王宫总管、市长和长老，并教养众儿子的人，派人到 耶户 那里，说：“我们是你的仆人，凡你所吩咐的，我们都必遵行。我们不立谁作王，你看怎样好就怎样做吧。”
2KGS|10|6|耶户 写第二封信给他们，说：“你们若归顺我，听从我的话，明日这时候，要带着你们主人众儿子的首级，来到 耶斯列 我这里。”那时王的儿子七十人都住在城中教养他们的那些尊贵人家里。
2KGS|10|7|信一到他们那里，他们就把王的七十个儿子杀了，将首级装在筐里，送到 耶斯列 ， 耶户 那里。
2KGS|10|8|有使者来告诉 耶户 说：“他们把王众儿子的首级送来了。” 耶户 说：“把首级分成两堆，放在城门口，直到早晨。”
2KGS|10|9|次日早晨， 耶户 出来，站着对众百姓说：“你们都是公义的！看哪，我背叛了我的主人，把他杀了，但这所有的人又是谁杀的呢？
2KGS|10|10|由此可知，耶和华指着 亚哈 家所说的话一句也没有落空，因为耶和华实现了他藉他仆人 以利亚 所说的话。”
2KGS|10|11|凡 亚哈 家在 耶斯列 所剩下的，他的大臣、密友、祭司， 耶户 全都杀了，没有留下一个幸存者。
2KGS|10|12|耶户 起身往 撒玛利亚 去。路途中，在牧人聚集的 伯．艾克特 ，
2KGS|10|13|耶户 遇见 犹大 王 亚哈谢 的兄弟，说：“你们是谁？”他们说：“我们是 亚哈谢 的兄弟，现在下去要向王和太后的众儿子问安。”
2KGS|10|14|耶户 说：“活捉他们！”人就活捉了他们，把他们杀在 伯．艾克特 的坑边，共四十二人，一个也没有留下。
2KGS|10|15|耶户 从那里往前行，遇见 利甲 的儿子 约拿达 来迎接他， 耶户 向他问安，对他说：“你的心 ，像我的心待你的心那样正直吗？” 约拿达 说：“是。” 耶户 说：“若是这样，请你伸出手来。”他伸出手， 耶户 就拉他上车。
2KGS|10|16|耶户 说：“你和我同去，看我为耶和华怎样热心。”于是他们请他坐在车上。
2KGS|10|17|到了 撒玛利亚 ， 耶户 把 亚哈 家在 撒玛利亚 剩下的人全都杀了，直到灭尽，正如耶和华对 以利亚 所说的话。
2KGS|10|18|耶户 召集众百姓，对他们说：“ 亚哈 事奉 巴力 还不够热心， 耶户 更要热心。
2KGS|10|19|现在你们召集 巴力 的众先知和所有拜 巴力 的人，以及 巴力 的众祭司，都到我这里来，一个也不可缺少，因为我要给 巴力 献大祭；凡不来的必不得活。” 耶户 行诡诈，为要消灭拜 巴力 的人。
2KGS|10|20|耶户 说：“要为 巴力 召集严肃会！”于是他们宣告了。
2KGS|10|21|耶户 派人走遍 以色列 ；凡拜 巴力 的人都来齐了，没有留下一个不来的。他们进了 巴力 庙， 巴力 庙中前后都挤满了人。
2KGS|10|22|耶户 对掌管服装的人说：“拿出袍子来，给所有拜 巴力 的人穿。”他就拿出礼服来给了他们。
2KGS|10|23|耶户 和 利甲 的儿子 约拿达 进了 巴力 庙，对拜 巴力 的人说：“你们要搜查察看，不可以有耶和华的仆人在你们这里，只可以有拜 巴力 的人。”
2KGS|10|24|他们进去，献上祭物和燔祭． 耶户 先安排八十人在庙外，说：“我把这些人交在你们手中，谁放走其中一人，谁就要以命偿命！”
2KGS|10|25|耶户 献完了燔祭，就对护卫兵和众军官说：“进去杀他们，不要让一人逃脱！”护卫兵和军官用刀杀了他们，将尸体抛出去，然后进入 巴力 庙的堡垒，
2KGS|10|26|将 巴力 庙中的柱像都 拿出来焚烧。
2KGS|10|27|他们毁坏 巴力 的柱像，拆毁了 巴力 庙当厕所，直到今日。
2KGS|10|28|这样， 耶户 在 以色列 中消灭了 巴力 。
2KGS|10|29|只是 耶户 不离开 尼八 的儿子 耶罗波安 使 以色列 人陷入罪里的那罪，就是拜 伯特利 和 但 的金牛犊。
2KGS|10|30|耶和华对 耶户 说：“因你办好我眼中看为正的事，照我的心意待 亚哈 家，你的子孙必接续你坐 以色列 的王位，直到第四代。”
2KGS|10|31|只是 耶户 不尽心遵守耶和华－ 以色列 上帝的律法，不离开 耶罗波安 使 以色列 人陷入罪里的那罪。
2KGS|10|32|在那些日子，耶和华开始削弱 以色列 。 哈薛 在 以色列 各边界攻击他们，
2KGS|10|33|就是 约旦河 东 基列 全地，从靠近 亚嫩谷 边的 亚罗珥 起，包括 基列 和 巴珊 ，就是 迦得 人、 吕便 人、 玛拿西 人的地。
2KGS|10|34|耶户 其余的事，凡他所做的和他英勇的事迹，不都写在《以色列诸王记》上吗？
2KGS|10|35|耶户 与他祖先同睡，葬在 撒玛利亚 ，他儿子 约哈斯 接续他作王。
2KGS|10|36|耶户 在 撒玛利亚 作 以色列 王二十八年。
2KGS|11|1|亚哈谢 的母亲 亚她利雅 见她儿子死了，就起来剿灭王室所有的后裔。
2KGS|11|2|但 约兰 王的女儿， 亚哈谢 的妹妹 约示巴 ，将 亚哈谢 的儿子 约阿施 从被杀的王子中偷出来，把他和他的奶妈藏在卧房里，躲避了 亚她利雅 ，没有被杀。
2KGS|11|3|亚她利雅 治理这地的时候， 约阿施 和他的奶妈在耶和华的殿里藏了六年。
2KGS|11|4|第七年， 耶何耶大 派人叫 迦利 人和护卫兵的众百夫长来，领他们进耶和华的殿，与他们立约，使他们在耶和华殿里起誓，又把王的儿子指给他们看，
2KGS|11|5|吩咐他们说：“你们要这样做：你们当中在安息日值班的，三分之一要把守王宫，
2KGS|11|6|三分之一要在 苏珥门 ，三分之一要在护卫兵院的后门；你们要这样轮流把守王宫。
2KGS|11|7|你们安息日所有不值班的两队人员要在耶和华的殿里护卫王；
2KGS|11|8|各人手拿兵器，四围保护王。凡擅自闯入你们行列的，要被处死。王出入的时候，你们当跟随他。”
2KGS|11|9|众百夫长就照着 耶何耶大 祭司一切所吩咐的去做，各带自己的人，无论安息日值班或不值班的，都到 耶何耶大 祭司那里。
2KGS|11|10|祭司就把耶和华殿里所藏 大卫 王的枪和盾牌交给百夫长。
2KGS|11|11|护卫兵手中各拿兵器，在祭坛和殿那里，从殿南到殿北，站在王的四围。
2KGS|11|12|耶何耶大 领 约阿施 出来，给他戴上冠冕，把律法书交给他，膏他作王；众人都鼓掌说：“愿王万岁！”
2KGS|11|13|亚她利雅 听见护卫兵和百姓的声音，就进耶和华的殿，到百姓那里。
2KGS|11|14|她观看，看哪，王照仪式站在柱旁，百夫长和号手在王旁边，国中的众百姓欢乐吹号。 亚她利雅 就撕裂衣服，喊着说：“反了！反了！”
2KGS|11|15|耶何耶大 祭司吩咐管军兵的百夫长，对他们说：“把她从行列之间赶出去，凡跟随她的必用刀杀死！”因为祭司说：“不可在耶和华殿里杀她。”
2KGS|11|16|他们就下手拿住她；她进入通往王宫的 马门 ，就在那里被杀。
2KGS|11|17|耶何耶大 使王和百姓与耶和华立约，作耶和华的子民，又使王与百姓立约。
2KGS|11|18|于是国中的众百姓都到 巴力 庙去，拆毁了庙，彻底打碎祭坛和偶像，又在坛前把 巴力 的祭司 玛坦 杀了。 耶何耶大 祭司派官员看守耶和华的殿，
2KGS|11|19|又率领百夫长， 迦利 人和护卫兵，以及国中的众百姓，请王从耶和华的殿下来，由护卫兵的门进入王宫，他就坐上王位。
2KGS|11|20|国中的众百姓都欢乐，合城也都平静。他们已将 亚她利雅 在王宫那里用刀杀了。
2KGS|11|21|约阿施 登基的时候年方七岁。
2KGS|12|1|耶户 第七年， 约阿施 登基，在 耶路撒冷 作王四十年。他母亲名叫 西比亚 ，是 别是巴 人。
2KGS|12|2|约阿施 在 耶何耶大 祭司教导他的一切日子，行耶和华眼中看为正的事。
2KGS|12|3|只是丘坛还没有废去，百姓仍在丘坛献祭烧香。
2KGS|12|4|约阿施 对众祭司说：“凡献到耶和华殿分别为圣的银子，无论是人的赎价，各人生命的赎价， 或自愿献给耶和华殿的银子，
2KGS|12|5|祭司可以各自从认识的人收取，用来修理殿的破坏之处，就是在那里发现的一切破坏之处。”
2KGS|12|6|然而，到了 约阿施 王第二十三年，祭司仍未修理殿的破坏之处。
2KGS|12|7|所以 约阿施 王召了 耶何耶大 祭司和众祭司来，对他们说：“你们怎么不修理殿的破坏之处呢？现在，不要再从认识的人收银子了，但要为了殿的破坏之处，把银子交出来。”
2KGS|12|8|众祭司答应不再收百姓的银子，也不再修理殿的破坏之处。
2KGS|12|9|耶何耶大 祭司取了一个柜子，在柜盖上钻了一个洞，放在祭坛旁，在进耶和华殿的右边；守门的祭司将献到耶和华殿的一切银子投在柜里。
2KGS|12|10|他们见柜里的银子多了，就叫王的书记和大祭司上来，将耶和华殿里所得的银子数点了，包起来。
2KGS|12|11|他们把秤好了的银子交在管理耶和华殿督工的手里，督工就支付给木匠和建造耶和华殿的工人，
2KGS|12|12|瓦匠和石匠，又买木料和凿成的石头，用来修理耶和华殿的破坏之处，以及其他修理殿的各项费用。
2KGS|12|13|但这些献到耶和华殿的银子，并没有用来造耶和华殿里的银杯、钳子、盘子、号筒和其他的金银器皿。
2KGS|12|14|他们把这银子交给工人，用来整修耶和华的殿。
2KGS|12|15|他们不用跟这些经手接受银子去支付工人的人算账，因为这些人办事诚实。
2KGS|12|16|赎愆祭和赎罪祭的银子没有献到耶和华的殿里，都归给祭司。
2KGS|12|17|那时， 亚兰 王 哈薛 上来攻打 迦特 ，攻取了它。 哈薛 就定意上来攻打 耶路撒冷 。
2KGS|12|18|犹大 王 约阿施 将他祖先 犹大 王 约沙法 、 约兰 、 亚哈谢 所分别为圣的物和自己所分别为圣的物，以及耶和华殿与王宫府库里所有的金子都送给 亚兰 王 哈薛 ； 哈薛 就不上 耶路撒冷 来了。
2KGS|12|19|约阿施 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
2KGS|12|20|约阿施 的臣仆起来背叛，在下到 悉拉 路上的 米罗 宫那里把他杀了。
2KGS|12|21|杀他的臣仆就是 示米押 的儿子 约撒拔 和 朔默 的儿子 约萨拔 。他与祖先同葬在 大卫城 ，他儿子 亚玛谢 接续他作王。
2KGS|13|1|亚哈谢 的儿子 犹大 王 约阿施 第二十三年， 耶户 的儿子 约哈斯 在 撒玛利亚 登基作 以色列 王十七年。
2KGS|13|2|约哈斯 行耶和华眼中看为恶的事，效法 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的那罪，总不离开。
2KGS|13|3|于是，耶和华的怒气向 以色列 发作，将他们屡次交在 亚兰 王 哈薛 和他儿子 便．哈达 的手里。
2KGS|13|4|约哈斯 恳求耶和华，耶和华就应允他，因为耶和华看见 以色列 所受的欺压，因 亚兰 王欺压他们。
2KGS|13|5|耶和华赐给 以色列 一位拯救者，使他们脱离 亚兰 人的手，于是 以色列 人仍旧安居在自己的帐棚里。
2KGS|13|6|然而他们不离开 耶罗波安 家使 以色列 陷入罪里的那罪，仍行在罪中，并且在 撒玛利亚 留下 亚舍拉 。
2KGS|13|7|亚兰 王灭绝 约哈斯 的军队，践踏他们如禾场上的尘沙，只给 约哈斯 留下五十骑兵，十辆战车，一万步兵。
2KGS|13|8|约哈斯 其余的事，凡他所做的和他英勇的事迹，不都写在《以色列诸王记》上吗？
2KGS|13|9|约哈斯 与他祖先同睡，葬在 撒玛利亚 ，他儿子 约阿施 接续他作王。
2KGS|13|10|犹大 王 约阿施 第三十七年， 约哈斯 的儿子 约阿施 在 撒玛利亚 登基作 以色列 王十六年。
2KGS|13|11|他行耶和华眼中看为恶的事，不离开 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的一切罪，仍行在罪中。
2KGS|13|12|约阿施 其余的事，凡他所做的和他与 犹大 王 亚玛谢 交战的英勇事迹，不都写在《以色列诸王记》上吗？
2KGS|13|13|约阿施 与他祖先同睡， 耶罗波安 坐上他的王位。 约阿施 与 以色列 诸王一同葬在 撒玛利亚 。
2KGS|13|14|以利沙 得了致命的病， 以色列 王 约阿施 下来看他，伏在他脸上哭泣，说：“我父啊！我父啊！ 以色列 的战车和骑兵啊！”
2KGS|13|15|以利沙 对他说：“把弓箭拿来。”王就拿了弓箭来。
2KGS|13|16|以利沙 对 以色列 王说：“你用手开弓。”王就用手开弓。 以利沙 按手在王的手上，
2KGS|13|17|说：“打开朝东的窗户。”他就打开。 以利沙 说：“射箭！”他就射箭。 以利沙 说：“这是耶和华得胜的箭，是战胜 亚兰 人的箭，因为你必在 亚弗 攻打 亚兰 人，直到灭尽他们。”
2KGS|13|18|以利沙 又说：“拿几枝箭来。”他就拿了来。 以利沙 对 以色列 王说：“打地吧！”他打了三次，就停止了。
2KGS|13|19|神人向他发怒，说：“你应当击打五六次，就能攻打 亚兰 人直到灭尽；现在你只能打败 亚兰 人三次。”
2KGS|13|20|以利沙 死了，人把他埋葬了。新的一年， 摩押 人成群结队入侵境内。
2KGS|13|21|有人正在埋葬死人，看哪，他们看见一群人来，就把死人抛在 以利沙 的坟墓里，逃跑了。死人一碰到 以利沙 的骸骨，就活过来，用脚站了起来。
2KGS|13|22|约哈斯 在位年间， 亚兰 王 哈薛 屡次欺压 以色列 。
2KGS|13|23|耶和华却因与 亚伯拉罕 、 以撒 、 雅各 所立的约，仍施恩给 以色列 人，怜悯他们，眷顾他们，不肯灭尽他们，直到现在 仍不赶逐他们离开自己面前。
2KGS|13|24|亚兰 王 哈薛 死了，他儿子 便．哈达 接续他作王。
2KGS|13|25|从前 哈薛 和 约阿施 的父亲 约哈斯 交战，攻取了些城镇，现在 约哈斯 的儿子 约阿施 三次打败 哈薛 的儿子 便．哈达 ，从他手中收回了 以色列 的城镇。
2KGS|14|1|约哈斯 的儿子 以色列 王 约阿施 第二年， 犹大 王 约阿施 的儿子 亚玛谢 登基。
2KGS|14|2|他登基的时候年二十五岁，在 耶路撒冷 作王二十九年。他母亲名叫 约耶但 ，是 耶路撒冷 人。
2KGS|14|3|亚玛谢 行耶和华眼中看为正的事，但不如他祖先 大卫 。他效法他父亲 约阿施 一切所行的。
2KGS|14|4|只是丘坛还没有废去，百姓仍在丘坛献祭烧香。
2KGS|14|5|王国在他手里巩固的时候，他就把杀他父王的臣仆杀了，
2KGS|14|6|却没有处死杀王凶手的儿子，正如 摩西 律法书上耶和华所吩咐的说：“不可因子杀父，也不可因父杀子，各人要为自己的罪而死。”
2KGS|14|7|亚玛谢 在 盐谷 杀了一万 以东 人，又在战役中攻取了 西拉 ，称它为 约帖 ，直到今日。
2KGS|14|8|那时， 亚玛谢 派使者到 耶户 的孙子， 约哈斯 的儿子 以色列 王 约阿施 那里，说：“来，让我们面对面较量吧！”
2KGS|14|9|以色列 王 约阿施 派人去见 犹大 王 亚玛谢 ，说：“ 黎巴嫩 的蒺藜派人去见 黎巴嫩 的香柏树，说：‘将你的女儿嫁给我的儿子。’但有一只野兽经过 黎巴嫩 ，把蒺藜践踏了。
2KGS|14|10|你果然打败了 以东 ，就心高气傲。你以此为荣，就待在自己家里算了吧，为何要惹祸，使自己和 犹大 一同败亡呢？”
2KGS|14|11|亚玛谢 却不肯听从。于是 以色列 王 约阿施 上来，在 犹大 的 伯．示麦 与 犹大 王 亚玛谢 面对面较量。
2KGS|14|12|犹大 败在 以色列 面前，他们逃跑，各人逃回自己的帐棚去了。
2KGS|14|13|以色列 王 约阿施 在 伯．示麦 擒住 亚哈谢 的孙子， 约阿施 的儿子 犹大 王 亚玛谢 ，就来到 耶路撒冷 ，拆毁 耶路撒冷 的城墙，从 以法莲门 直到 角门 共四百肘。
2KGS|14|14|他又拿了耶和华殿里与王宫府库里所有的金银和器皿，并带着人质，回 撒玛利亚 去了。
2KGS|14|15|约阿施 其余所做的事和他英勇的事迹，以及他与 犹大 王 亚玛谢 交战的事，不都写在《以色列诸王记》上吗？
2KGS|14|16|约阿施 与他祖先同睡，与 以色列 诸王一同葬在 撒玛利亚 ，他儿子 耶罗波安 接续他作王。
2KGS|14|17|约哈斯 的儿子 以色列 王 约阿施 死后， 犹大 王 约阿施 的儿子 亚玛谢 又活了十五年。
2KGS|14|18|亚玛谢 其余的事，不都写在《犹大列王记》上吗？
2KGS|14|19|耶路撒冷 有人背叛 亚玛谢 ， 亚玛谢 逃往 拉吉 ；他们却派人追到 拉吉 ，在那里杀了他。
2KGS|14|20|有人用马将他驮回，葬在 耶路撒冷 ，与他祖先一同葬在 大卫城 。
2KGS|14|21|犹大 众百姓立 亚撒利雅 接续他父亲 亚玛谢 作王，那时他年十六岁。
2KGS|14|22|亚玛谢 王与他祖先同睡之后， 亚撒利雅 收复 以拉他 回归 犹大 ，又重新整修。
2KGS|14|23|约阿施 的儿子 犹大 王 亚玛谢 第十五年， 以色列 王 约阿施 的儿子 耶罗波安 在 撒玛利亚 登基，作王四十一年。
2KGS|14|24|他行耶和华眼中看为恶的事，不离开 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的一切罪。
2KGS|14|25|他收回 以色列 边界之地，从 哈马口 直到 亚拉巴海 ，正如耶和华－ 以色列 的上帝藉他仆人 迦特．希弗 人 亚米太 的儿子 约拿 先知所说的。
2KGS|14|26|因耶和华看见 以色列 非常艰苦的困境；没有奴役的，没有自由的，也没有人来帮助 以色列 。
2KGS|14|27|耶和华并没有说要将 以色列 的名从天下涂抹，却要藉 约阿施 的儿子 耶罗波安 拯救他们。
2KGS|14|28|耶罗波安 其余的事，凡他所做的和他英勇的事迹，他怎样作战，怎样收复 大马士革 和先前属 犹大 的 哈马 回归 以色列 ，不都写在《以色列诸王记》上吗？
2KGS|14|29|耶罗波安 与他祖先 以色列 诸王同睡，他儿子 撒迦利雅 接续他作王。
2KGS|15|1|以色列 王 耶罗波安 第二十七年， 犹大 王 亚玛谢 的儿子 亚撒利雅 登基。
2KGS|15|2|他登基的时候年十六岁，在 耶路撒冷 作王五十二年。他母亲名叫 耶可利雅 ，是 耶路撒冷 人。
2KGS|15|3|亚撒利雅 行耶和华眼中看为正的事，效法他父亲 亚玛谢 一切所行的。
2KGS|15|4|只是丘坛还没有废去，百姓仍在丘坛献祭烧香。
2KGS|15|5|耶和华降灾于王，使他长了痲疯，直到死的那日。他住在隔离的行宫里，他儿子 约坦 管理王的家，治理这地的百姓。
2KGS|15|6|亚撒利雅 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
2KGS|15|7|亚撒利雅 与他祖先同睡，与他祖先同葬在 大卫城 ，他儿子 约坦 接续他作王。
2KGS|15|8|犹大 王 亚撒利雅 第三十八年， 耶罗波安 的儿子 撒迦利雅 登基，在 撒玛利亚 作 以色列 王六个月。
2KGS|15|9|他行耶和华眼中看为恶的事，效法他祖先所行的，不离开 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的那罪。
2KGS|15|10|雅比 的儿子 沙龙 背叛他，在百姓面前 击杀他，篡了他的位。
2KGS|15|11|撒迦利雅 其余的事，看哪，都写在《以色列诸王记》上。
2KGS|15|12|这就是耶和华应许 耶户 的话：“你的子孙必坐 以色列 的王位，直到第四代。”这事果然发生了。
2KGS|15|13|犹大 王 乌西雅 第三十九年， 雅比 的儿子 沙龙 登基，在 撒玛利亚 作王一个月。
2KGS|15|14|迦底 的儿子 米拿现 从 得撒 上 撒玛利亚 ，杀了 雅比 的儿子 沙龙 ，篡了他的位。
2KGS|15|15|沙龙 其余的事和他阴谋背叛的事，看哪，都写在《以色列诸王记》上。
2KGS|15|16|那时， 米拿现 从 得撒 起击杀 提斐萨 和城中所有的人，以及它周围的地区，因为他们没有给他开城门。他击杀他们，剖开其中所有的孕妇。
2KGS|15|17|犹大 王 亚撒利雅 第三十九年， 迦底 的儿子 米拿现 登基，在 撒玛利亚 作 以色列 王十年。
2KGS|15|18|他行耶和华眼中看为恶的事，终生不离开 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的那罪。
2KGS|15|19|亚述 王 普勒 来攻击这地， 米拿现 给他一千他连得银子，为了请 普勒 帮助他巩固他所掌握的国度。
2KGS|15|20|米拿现 向 以色列 所有的富豪索取银子，要他们各出五十舍客勒，交给 亚述 王。于是 亚述 王回去了，不在境内停留。
2KGS|15|21|米拿现 其余的事，凡他所做的，不都写在《以色列诸王记》上吗？
2KGS|15|22|米拿现 与他祖先同睡，他儿子 比加辖 接续他作王。
2KGS|15|23|犹大 王 亚撒利雅 第五十年， 米拿现 的儿子 比加辖 登基，在 撒玛利亚 作 以色列 王二年。
2KGS|15|24|他行耶和华眼中看为恶的事，不离开 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的那罪。
2KGS|15|25|比加辖 的将军， 利玛利 的儿子 比加 背叛他，在 撒玛利亚 王宫的堡垒杀了他。 亚珥歌伯 和 亚利耶 并 基列 的五十人帮助 比加 ； 比加 击杀他，篡了他的位。
2KGS|15|26|比加辖 其余的事，凡他所做的，看哪，都写在《以色列诸王记》上。
2KGS|15|27|犹大 王 亚撒利雅 第五十二年， 利玛利 的儿子 比加 登基，在 撒玛利亚 作 以色列 王二十年。
2KGS|15|28|他行耶和华眼中看为恶的事，不离开 尼八 的儿子 耶罗波安 使 以色列 陷入罪里的那罪。
2KGS|15|29|在 以色列 王 比加 的日子， 亚述 王 提革拉．毗列色 来夺取 以云 、 亚伯．伯．玛迦 、 亚挪 、 基低斯 、 夏琐 、 基列 、 加利利 和 拿弗他利 全地，把这些地方的居民都掳到 亚述 去了。
2KGS|15|30|乌西雅 的儿子 约坦 第二十年， 以拉 的儿子 何细亚 背叛 利玛利 的儿子 比加 ，击杀他，篡了他的位。
2KGS|15|31|比加 其余的事，凡他所做的，看哪，都写在《以色列诸王记》上。
2KGS|15|32|利玛利 的儿子 以色列 王 比加 第二年， 犹大 王 乌西雅 的儿子 约坦 登基。
2KGS|15|33|他登基的时候年二十五岁，在 耶路撒冷 作王十六年。他母亲名叫 耶路沙 ，是 撒督 的女儿。
2KGS|15|34|约坦 行耶和华眼中看为正的事，效法他父亲 乌西雅 一切所行的。
2KGS|15|35|只是丘坛还没有废去，百姓仍在丘坛献祭烧香。 约坦 建了耶和华殿的 上门 。
2KGS|15|36|约坦 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
2KGS|15|37|在那些日子，耶和华开始差 亚兰 王 利汛 和 利玛利 的儿子 比加 去攻击 犹大 。
2KGS|15|38|约坦 与他祖先同睡，与他祖先同葬在 大卫城 ，他儿子 亚哈斯 接续他作王。
2KGS|16|1|利玛利 的儿子 比加 第十七年， 犹大 王 约坦 的儿子 亚哈斯 登基。
2KGS|16|2|他登基的时候年二十岁，在 耶路撒冷 作王十六年。他不像他祖先 大卫 行耶和华－他上帝眼中看为正的事，
2KGS|16|3|却行 以色列 诸王的道，又照着耶和华从 以色列 人面前赶出的外邦人所行可憎的事，使他的儿子经火，
2KGS|16|4|并在丘坛上、山冈上、各青翠树下献祭烧香。
2KGS|16|5|那时， 亚兰 王 利汛 和 利玛利 的儿子 以色列 王 比加 上来攻打 耶路撒冷 ，围困 亚哈斯 ，却不能打胜。
2KGS|16|6|当时 亚兰 王 利汛 收复 以拉他 回归 亚兰 ，把 犹大 人从 以拉他 赶出去。 以东 人来到 以拉他 ，住在那里，直到今日。
2KGS|16|7|亚哈斯 派使者到 亚述 王 提革拉．毗列色 那里，说：“我是你的仆人，你的儿子。现在 亚兰 王和 以色列 王攻击我，求你上来，救我脱离他们的手。”
2KGS|16|8|亚哈斯 将耶和华殿里和王宫府库里所有的金银都送给 亚述 王为礼物。
2KGS|16|9|亚述 王答应了他，上去攻打 大马士革 ，攻下了城，杀了 利汛 ，把居民掳到 吉珥 。
2KGS|16|10|亚哈斯 王到 大马士革 迎接 亚述 王 提革拉．毗列色 ，在 大马士革 看见一座坛。 亚哈斯 王把坛的规模和样式，以及作法的细节，送到 乌利亚 祭司那里。
2KGS|16|11|乌利亚 祭司照着 亚哈斯 王从 大马士革 所送来的一切，在 亚哈斯 王还未从 大马士革 回来之前，筑了一座坛。
2KGS|16|12|王从 大马士革 回来，看见坛，走近坛前，在坛上献祭。
2KGS|16|13|他烧燔祭和素祭，献浇酒祭，将平安祭牲的血洒在坛上。
2KGS|16|14|他移动耶和华面前的铜坛，从殿的前面，新坛和耶和华殿的中间，搬到新坛的北边。
2KGS|16|15|亚哈斯 王吩咐 乌利亚 祭司说：“早晨的燔祭、晚上的素祭，王的燔祭、素祭，国内众百姓的燔祭、素祭、浇酒祭都要烧在大坛上。燔祭牲和其他祭牲的血全都要洒在这坛上。至于铜坛，我要作求问之用。”
2KGS|16|16|乌利亚 祭司就照着 亚哈斯 王所吩咐的一切做了。
2KGS|16|17|亚哈斯 王把盆座四面的嵌边拆下来，把盆从座上挪下来，又将铜海从驮铜海的铜牛上搬下来，放在石板铺的地上。
2KGS|16|18|他为了 亚述 王的缘故，在耶和华的殿里移动 殿里为安息日所盖的遮棚 和王从外面进来的入口。
2KGS|16|19|亚哈斯 其余所做的事，不都写在《犹大列王记》上吗？
2KGS|16|20|亚哈斯 与他祖先同睡， 与他祖先同葬在 大卫城 ，他儿子 希西家 接续他作王。
2KGS|17|1|犹大 王 亚哈斯 第十二年， 以拉 的儿子 何细亚 在 撒玛利亚 登基作 以色列 王九年。
2KGS|17|2|他行耶和华眼中看为恶的事，只是不像在他以前的 以色列 诸王。
2KGS|17|3|亚述 王 撒缦以色 上来攻击 何细亚 ， 何细亚 就服事他，向他进贡。
2KGS|17|4|何细亚 背叛，派使者到 埃及 王 梭 那里 ，不照往年所行的向 亚述 王进贡。 亚述 王知道了，就逮捕他，把他囚在监里。
2KGS|17|5|亚述 王上来攻击 以色列 全地，上到 撒玛利亚 ，围困这城三年。
2KGS|17|6|何细亚 第九年， 亚述 王攻取了 撒玛利亚 ，把 以色列 人掳到 亚述 ，安置在 哈腊 与 歌散 的 哈博河 边，以及 玛代 人的城镇。
2KGS|17|7|这是因为 以色列 人得罪了那领他们出 埃及 地、脱离 埃及 王法老之手的耶和华－他们的上帝，去敬畏别神，
2KGS|17|8|随从耶和华在 以色列 人面前所赶出外邦人的风俗和 以色列 诸王所立的规条。
2KGS|17|9|以色列 人暗中行不正的事，违背耶和华－他们的上帝，在他们所有的城镇，从了望楼直到坚固城，建筑丘坛；
2KGS|17|10|在各高冈上、各青翠树下立柱像和 亚舍拉 ；
2KGS|17|11|在各丘坛上烧香，效法耶和华在他们面前赶出的外邦人所行的，又行恶事，惹耶和华发怒。
2KGS|17|12|他们事奉偶像，耶和华对他们说：“你们不可做这事。”
2KGS|17|13|耶和华藉众先知、先见劝戒 以色列 和 犹大 说：“当离开你们的恶行，谨守我的诫命律例，遵行我吩咐你们祖先、藉我仆人众先知所传给你们的一切律法。”
2KGS|17|14|他们却不听从，竟硬着颈项，像他们祖先一样，不信服耶和华－他们的上帝。
2KGS|17|15|他们厌弃他的律例，和他与他们列祖所立的约，以及他劝戒他们的话，去随从虚无的神明 ，自己成为虚妄，效法周围的列国，就是耶和华嘱咐他们不可效法的。
2KGS|17|16|他们离弃耶和华－他们上帝的一切诫命，为自己铸造了两个牛犊的像，立了 亚舍拉 ，敬拜天上的万象，事奉 巴力 ，
2KGS|17|17|使他们的儿女经火，占卜，行法术，出卖自己，行耶和华眼中看为恶的事，惹他发怒。
2KGS|17|18|所以耶和华向 以色列 大大发怒，从自己面前赶出他们，只剩下 犹大 一个支派。
2KGS|17|19|但是， 犹大 也不遵守耶和华－他们上帝的诫命，效法 以色列 所立的规条。
2KGS|17|20|耶和华就厌弃 以色列 所有的后裔，使他们受苦，把他们交在抢夺他们的人手中，直到他把他们从自己面前赶出去。
2KGS|17|21|当他使 以色列 从 大卫 家分离出来的时候，他们立 尼八 的儿子 耶罗波安 作王。 耶罗波安 引诱 以色列 不随从耶和华，陷入大罪中。
2KGS|17|22|以色列 人行 耶罗波安 所犯的一切罪，总不离开，
2KGS|17|23|以致耶和华把他们从自己面前赶出去，正如他藉他仆人众先知所说的。这样， 以色列 人从自己的土地被掳到 亚述 ，直到今日。
2KGS|17|24|亚述 王从 巴比伦 、 古他 、 亚瓦 、 哈马 和 西法瓦音 迁移人来，安置在 撒玛利亚 的城镇，代替 以色列 人；他们就占据了 撒玛利亚 ，住在城中。
2KGS|17|25|他们开始住在那里的时候，不敬畏耶和华，所以耶和华叫狮子进入他们中间，咬死了一些人。
2KGS|17|26|有人对 亚述 王说：“你所迁移安置在 撒玛利亚 城镇的各国的人，他们不知道那地之上帝的规矩，所以他叫狮子进入他们中间。看哪，狮子咬死了他们，因为他们不知道那地之上帝的规矩。”
2KGS|17|27|亚述 王吩咐说：“当派一个从那里掳来的祭司回去，叫他住在那里，将那地之上帝的规矩指导他们。”
2KGS|17|28|于是有一个从 撒玛利亚 掳去的祭司回来，住在 伯特利 ，教导他们怎样敬畏耶和华。
2KGS|17|29|然而，各国的人在所住的城里为自己制造神像，安置在 撒玛利亚 人所建有丘坛的庙中。
2KGS|17|30|巴比伦 人造 疏割．比讷 像； 古他 人造 匿甲 像； 哈马 人造 亚示玛 像；
2KGS|17|31|亚瓦 人造 匿哈 和 他珥他 像； 西法瓦音 人用火焚烧儿女，献给 西法瓦音 的神明 亚得米勒 和 亚拿米勒 。
2KGS|17|32|他们惧怕耶和华，却从他们中间立丘坛的祭司，在丘坛的庙中为他们献祭。
2KGS|17|33|他们惧怕耶和华，但又事奉自己的神明，从何邦迁来，就随从那里的风俗，
2KGS|17|34|直到如今仍照先前的风俗去行。 他们不敬畏耶和华，不遵守耶和华吩咐 雅各 后裔的律例、典章、律法、诫命； 雅各 就是从前耶和华起名叫 以色列 的。
2KGS|17|35|耶和华曾与他们立约，吩咐他们说：“不可敬畏别神，不可跪拜事奉它们，也不可向它们献祭。
2KGS|17|36|惟有那用大能和伸出来的膀臂领你们出 埃及 地的耶和华，你们当敬畏他，向他跪拜，向他献祭。
2KGS|17|37|他给你们写的律例、典章、律法、诫命，你们应当永远谨守遵行。你们不可敬畏别神。
2KGS|17|38|你们不可忘记我与你们所立的约，也不可敬畏别神。
2KGS|17|39|只要敬畏耶和华－你们的上帝，他必救你们脱离一切仇敌的手。”
2KGS|17|40|他们却不听从，仍照先前的风俗去行。
2KGS|17|41|这样，这些国家又惧怕耶和华，又事奉他们的偶像。他们子子孙孙也都照样行，效法他们的祖宗，直到今日。
2KGS|18|1|以拉 的儿子 以色列 王 何细亚 第三年， 犹大 王 亚哈斯 的儿子 希西家 登基。
2KGS|18|2|他登基的时候年二十五岁，在 耶路撒冷 作王二十九年。他母亲名叫 亚比 ，是 撒迦利雅 的女儿。
2KGS|18|3|希西家 行耶和华眼中看为正的事，效法他祖先 大卫 一切所行的。
2KGS|18|4|他废去丘坛，毁坏柱像，砍下 亚舍拉 ，打碎 摩西 所造的铜蛇，因为到那时 以色列 人仍向铜蛇烧香。人叫铜蛇为 尼忽士但 。
2KGS|18|5|希西家 倚靠耶和华－ 以色列 的上帝，在他之前和在他之后的 犹大 列王中没有一个像他一样的。
2KGS|18|6|因为他紧紧跟随耶和华，谨守耶和华所吩咐 摩西 的诫命，总不离开。
2KGS|18|7|耶和华与他同在，他无论往何处去尽都亨通。他背叛 亚述 王，不服事他。
2KGS|18|8|希西家 攻击 非利士 人，直到 迦萨 ，以及所属的领土，从了望楼到坚固城。
2KGS|18|9|希西家 王第四年，也就是 以拉 的儿子 以色列 王 何细亚 第七年， 亚述 王 撒缦以色 上来围困 撒玛利亚 。
2KGS|18|10|过了三年，他们攻取了城。 希西家 第六年， 以色列 王 何细亚 第九年， 撒玛利亚 被攻取了。
2KGS|18|11|亚述 王把 以色列 人掳到 亚述 ，安置在 哈腊 与 歌散 的 哈博河 边，以及 玛代 人的城镇。
2KGS|18|12|这是因为他们不听从耶和华－他们的上帝的话，违背了他的约；他们既不听从，也不遵行耶和华仆人 摩西 一切所吩咐的。
2KGS|18|13|希西家 王十四年， 亚述 王 西拿基立 上来攻击 犹大 的一切坚固的城，将城攻取。
2KGS|18|14|犹大 王 希西家 派人到 拉吉 ， 亚述 王那里，说：“我错了，求你撤退离开我；凡你罚我的，我必承当。”于是 亚述 王罚 犹大 王 希西家 三百他连得银子，三十他连得金子。
2KGS|18|15|希西家 把耶和华殿里和王宫府库里所有的银子都给了他。
2KGS|18|16|那时， 犹大 王 希西家 将耶和华殿门上的金子和他自己包在柱子上的金子都刮下来，给了 亚述 王。
2KGS|18|17|亚述 王从 拉吉 差遣元帅 、太监长 和将军 率领大军前往 耶路撒冷 ，到 希西家 王那里去。他们上来，到 耶路撒冷 。他们上来之后，站在 上池 的水沟旁，在往漂布地的大路上。
2KGS|18|18|他们呼叫王， 希勒家 的儿子 以利亚敬 宫廷总管， 舍伯那 书记和 亚萨 的儿子 约亚 史官就出来见他们。
2KGS|18|19|将军对他们说：“你们去告诉 希西家 ，大王 亚述 王如此说：‘你倚靠什么，让你如此自信满满？
2KGS|18|20|你说，你有打仗的计谋和能力，我看不过是空话。你到底倚靠谁，竟敢背叛我呢？
2KGS|18|21|现在，看哪，你自己所倚靠的 埃及 是那断裂的苇杖，人若倚靠这杖，它就刺进他的手，穿透它。 埃及 王法老向所有倚靠他的人都是这样。
2KGS|18|22|你们若对我说：我们倚靠耶和华－我们的上帝， 希西家 岂不是将上帝的丘坛和祭坛废去，并且吩咐 犹大 和 耶路撒冷 的人说：你们当在 耶路撒冷 这坛前敬拜吗？
2KGS|18|23|现在你与我主 亚述 王打赌，我给你两千匹马，看你能否派得出骑士来骑它们。
2KGS|18|24|若不然，怎能使我主臣仆中最小的一个军官转脸而逃呢？你难道要倚靠 埃及 的战车和骑兵吗？
2KGS|18|25|现在我上来攻击毁灭这地方，岂不是出于耶和华吗？耶和华吩咐我说，你上去攻击这地，毁灭它吧！’”
2KGS|18|26|希勒家 的儿子 以利亚敬 ， 舍伯那 和 约亚 对将军说：“求你用 亚兰 话对仆人说，因为我们听得懂；不要用 犹大 话对我们说，免得传到城墙上百姓的耳中。”
2KGS|18|27|将军对他们说：“我主差遣我来，岂是单对你和你的主人说这些话吗？不也是对这些坐在城墙上、要与你们一同吃自己粪、喝自己尿的人说的吗？”
2KGS|18|28|于是 亚述 将军站着，用 犹大 话大声喊着说：“你们当听大王 亚述 王的话，
2KGS|18|29|王如此说：‘你们不要被 希西家 欺哄了，因他不能救你们脱离我的手。
2KGS|18|30|不要听凭 希西家 说服你们倚靠耶和华，他说，耶和华必要拯救我们，这城必不交在 亚述 王的手中。’
2KGS|18|31|你们不要听 希西家 的话！因 亚述 王如此说：‘你们要与我讲和，出来投降我，各人就可以吃自己葡萄树和无花果树的果子，喝自己井里的水，
2KGS|18|32|等我来领你们到一个地方，与你们本地一样，就是有五谷和新酒之地，有粮食和葡萄园之地，有橄榄树和蜂蜜之地，好使你们存活，不至于死。不要听 希西家 的话，因为他误导你们说：耶和华必拯救我们。
2KGS|18|33|列国的神明有哪一个曾救它本国脱离 亚述 王的手呢？
2KGS|18|34|哈马 、 亚珥拔 的神明在哪里呢？ 西法瓦音 、 希拿 、 以瓦 的神明在哪里呢？ 它们曾救 撒玛利亚 脱离我的手吗？
2KGS|18|35|这些国的神明有谁曾救自己的国脱离我的手呢？难道耶和华能救 耶路撒冷 脱离我的手吗？’”
2KGS|18|36|百姓静默不言，一句不答，因为 希西家 王曾吩咐说：“不要回答他。”
2KGS|18|37|当下， 希勒家 的儿子 以利亚敬 宫廷总管、 舍伯那 书记和 亚萨 的儿子 约亚 史官，都撕裂衣服，来到 希西家 那里，将 亚述 将军的话告诉他。
2KGS|19|1|希西家 王听见了，就撕裂衣服，披上麻布，进了耶和华的殿。
2KGS|19|2|他差遣 以利亚敬 宫廷总管和 舍伯那 书记，并祭司中年长的，都披上麻布，到 亚摩斯 的儿子 以赛亚 先知那里去。
2KGS|19|3|他们对他说：“ 希西家 如此说：‘今日是急难、惩罚、凌辱的日子，就如婴孩快要出生，却没有力气生产。
2KGS|19|4|或许耶和华－你的上帝听见 亚述 将军一切的话，就是他主人 亚述 王差他来辱骂永生上帝的话，耶和华－你的上帝就斥责所听见的这些话。求你为幸存的余民扬声祷告。’”
2KGS|19|5|希西家 王的臣仆来到 以赛亚 那里的时候，
2KGS|19|6|以赛亚 对他们说：“要对你们的主人这样说，耶和华如此说：‘你听见 亚述 王的仆人亵渎我的话，不要惧怕。
2KGS|19|7|看哪，我必惊动他的心 ，他要听见风声就归回本地，在那里我必使他倒在刀下。’”
2KGS|19|8|亚述 将军听见 亚述 王已拔营离开 拉吉 ，就启程返回，正遇见 亚述 王去攻打 立拿 。
2KGS|19|9|亚述 王听见有人谈论 古实 王 特哈加 说：“看哪，他出来要与你争战。”于是 亚述 王又差使者去见 希西家 ，说：
2KGS|19|10|“你们要对 犹大 王 希西家 如此说：‘不要听你所倚靠的上帝欺哄你说： 耶路撒冷 必不交在 亚述 王的手中。
2KGS|19|11|看哪，你总听说 亚述 诸王向列国所行的是尽行灭绝，难道你能幸免吗？
2KGS|19|12|我祖先所毁灭的，就是 歌散 、 哈兰 、 利色 和 提．拉撒 的 伊甸 人；这些国的神明何曾拯救他们呢？
2KGS|19|13|哈马 的王， 亚珥拔 的王， 西法瓦音城 的王， 希拿 和 以瓦 的王，都在哪里呢？’”
2KGS|19|14|希西家 从使者手里接过书信，读完了，就上耶和华的殿，在耶和华面前展开书信。
2KGS|19|15|希西家 向耶和华祷告说：“坐在基路伯之上耶和华－ 以色列 的上帝啊，你，惟有你是地上万国的上帝，你创造了天和地。
2KGS|19|16|耶和华啊，求你侧耳而听；耶和华啊，求你睁眼而看，听 西拿基立 差遣使者辱骂永生上帝的话。
2KGS|19|17|耶和华啊， 亚述 诸王果然使列国和列国之地变为荒芜，
2KGS|19|18|将列国的神像扔在火里，因为它们不是上帝，是人手所造的，是木头、石头，所以被灭绝了。
2KGS|19|19|耶和华－我们的上帝啊，现在求你救我们脱离 亚述 王的手，使地上万国都知道惟独你－耶和华是上帝！”
2KGS|19|20|亚摩斯 的儿子 以赛亚 差人去见 希西家 ，说：“耶和华－ 以色列 的上帝如此说：你因 亚述 王 西拿基立 的事向我祈求，我已听见了。
2KGS|19|21|耶和华论他这样说： ‘少女 锡安 藐视你，嘲笑你； 耶路撒冷 向你摇头。
2KGS|19|22|‘你辱骂谁，亵渎谁， 扬起声来，高举眼目攻击谁呢？ 你攻击的是 以色列 的圣者。
2KGS|19|23|你藉你的使者辱骂主说： 我率领许多战车登上高山， 到 黎巴嫩 的顶端； 我要砍伐其中高大的香柏树 和上好的松树； 我必进到极遥远的住所， 进入最茂盛的森林里。
2KGS|19|24|我已经在外邦挖井喝水； 我必用脚掌踏干 埃及 一切的河流。
2KGS|19|25|‘你岂没有听见 我早先所定、古时所立、现今实现的事吗？ 就是让你去毁坏坚固的城镇，使它们变为废墟；
2KGS|19|26|城里的居民力量微小， 他们惊惶羞愧； 像野草，像青菜， 如房顶上的草， 又如未长成而枯干的禾稼。
2KGS|19|27|‘你坐下，你出去，你进来， 你向我发烈怒，我都知道。
2KGS|19|28|因你向我发烈怒， 你的狂傲上达我耳中， 我要用钩子钩住你的鼻子， 将嚼环放在你口里， 使你从原路转回去。’
2KGS|19|29|“这是给你的预兆：你们今年要吃野生的，明年也要吃自长的；后年，你们就要耕种收割，栽葡萄园，吃其中的果子。
2KGS|19|30|犹大 家所逃脱剩余的，仍要往下扎根，向上结果。
2KGS|19|31|必有剩余的民从 耶路撒冷 而出，有逃脱的人从 锡安山 而来。万军之耶和华的热心必成就这事。
2KGS|19|32|“所以耶和华论 亚述 王如此说：他必不得来到这城，也不在这里射箭，不得拿盾牌到城前，也不建土堆攻城。
2KGS|19|33|他从哪条路来，必从那条路回去，必不得来到这城。这是耶和华说的。
2KGS|19|34|因我为自己的缘故，又为我仆人 大卫 的缘故，必保护拯救这城。”
2KGS|19|35|当夜，耶和华的使者出去，在 亚述 营中杀了十八万五千人。清早有人起来，看哪，都是死尸。
2KGS|19|36|亚述 王 西拿基立 就拔营回去，住在 尼尼微 。
2KGS|19|37|一日，他在他的神明 尼斯洛 庙里叩拜，他儿子 亚得米勒 和 沙利色 用刀杀了他，然后逃到 亚拉腊 地；他儿子 以撒．哈顿 接续他作王。
2KGS|20|1|那些日子， 希西家 病得要死， 亚摩斯 的儿子 以赛亚 先知来见他，对他说：“耶和华如此说：‘你当留遗嘱给你的家，因为你必死，不能活了。’”
2KGS|20|2|希西家 转脸朝墙，向耶和华祷告说：
2KGS|20|3|“耶和华啊，求你记念我在你面前怎样存完全的心，按诚实行事，又做你眼中看为善的事。” 希西家 就痛哭。
2KGS|20|4|以赛亚 出来，还没有离开中院，耶和华的话就临到他，说：
2KGS|20|5|“你回去告诉我百姓的君王 希西家 说：耶和华－你祖先 大卫 的上帝如此说：‘我听见了你的祷告，看见了你的眼泪。看哪，我必医治你；到第三日，你必上到耶和华的殿。
2KGS|20|6|我必加添你十五年的寿数，并且我要救你和这城脱离 亚述 王的手。我为自己和我仆人 大卫 的缘故，必保护这城。’”
2KGS|20|7|以赛亚 说：“取一块无花果饼来。”人就取了来，贴在疮上，王就痊愈了。
2KGS|20|8|希西家 对 以赛亚 说：“耶和华必医治我，到第三日我能上耶和华的殿，有什么预兆呢？”
2KGS|20|9|以赛亚 说：“耶和华必成就他所说的这话。这是耶和华给你的预兆：你要日影向前进十度呢？或是要往后退十度呢？”
2KGS|20|10|希西家 说：“日影向前进十度容易；不，让日影往后退十度吧。”
2KGS|20|11|以赛亚 先知求告耶和华，耶和华就使 亚哈斯 日晷上照下来的日影，往后退了十度。
2KGS|20|12|那时， 巴拉但 的儿子， 巴比伦 王 米罗达．巴拉但 听见 希西家 生病了，就送书信和礼物给他。
2KGS|20|13|希西家 听使者的话 ，就将自己一切宝库里的金子、银子、香料、贵重的膏油和他军械库里的兵器，以及他所有的财宝，都给他们看；在他家中和全国之内， 希西家 没有一样东西不给他们看的。
2KGS|20|14|于是 以赛亚 先知到 希西家 王那里去，对他说：“这些人说了些什么？他们从哪里来见你？” 希西家 说：“他们从远方的 巴比伦 来。”
2KGS|20|15|以赛亚 说：“他们在你家里看见了什么？” 希西家 说：“凡我家中所有的，他们都看见了；我财宝中没有一样东西不给他们看的。”
2KGS|20|16|以赛亚 对 希西家 说：“你要听耶和华的话：
2KGS|20|17|耶和华说：‘看哪，日子将到，凡你家里所有的，并你祖先积蓄到如今的一切，都要被掳到 巴比伦 去，不留下一样；
2KGS|20|18|从你本身所生的孩子，其中必有被掳到 巴比伦 王宫当太监的。’”
2KGS|20|19|希西家 对 以赛亚 说：“你所说耶和华的话甚好。”因为他想：“在我有生之年岂不是有太平和安稳吗？”
2KGS|20|20|希西家 其余的事和他一切英勇的事迹，他怎样造池、挖沟、引水入城，不都写在《犹大列王记》上吗？
2KGS|20|21|希西家 与他祖先同睡，他儿子 玛拿西 接续他作王。
2KGS|21|1|玛拿西 登基的时候年十二岁，在 耶路撒冷 作王五十五年。他母亲名叫 协西巴 。
2KGS|21|2|玛拿西 行耶和华眼中看为恶的事，效法耶和华在 以色列 人面前赶出的列国那些可憎的事。
2KGS|21|3|他重新建筑他父亲 希西家 所毁坏的丘坛，又为 巴力 筑坛，造 亚舍拉 ，效法 以色列 王 亚哈 所行的，敬拜天上的万象，事奉它们。
2KGS|21|4|他在耶和华殿中筑坛，耶和华曾指着这殿说：“我必立我的名在 耶路撒冷 。”
2KGS|21|5|他在耶和华殿的两个院子为天上的万象筑坛，
2KGS|21|6|并使他的儿子经火，又观星象，行法术，求问招魂的和行巫术的，多行耶和华眼中看为恶的事，惹他发怒。
2KGS|21|7|他又把自己所造的 亚舍拉 雕像立在殿内，耶和华曾对 大卫 和他儿子 所罗门 说：“我在 以色列 众支派中所选择的 耶路撒冷 和这殿，必立我的名，直到永远。
2KGS|21|8|只要 以色列 人谨守遵行我一切所吩咐的和我仆人 摩西 所吩咐的一切律法，我就不再使他们的脚挪移，离开我所赐给他们列祖之土地。”
2KGS|21|9|他们却不听从，并且 玛拿西 引诱他们行恶，比耶和华在 以色列 人面前所灭的列国更严重。
2KGS|21|10|耶和华藉他仆人众先知说：
2KGS|21|11|“因 犹大 王 玛拿西 行这些可憎的恶事，比先前 亚摩利 人所行的一切更坏，使 犹大 人拜偶像，陷入罪里，
2KGS|21|12|所以耶和华－ 以色列 的上帝如此说：看哪，我必降祸于 耶路撒冷 和 犹大 ，凡听见的人都必双耳齐鸣。
2KGS|21|13|我必用量 撒玛利亚 的准绳和 亚哈 家的铅垂线拉在 耶路撒冷 之上；我必擦拭 耶路撒冷 ，如人擦盘子，把盘子翻过来。
2KGS|21|14|我必撇弃我产业中的余民，把他们交在仇敌手中，使他们成为所有仇敌的掳物和掠物，
2KGS|21|15|因为自从他们的祖先出 埃及 的那日直到今日，他们常行我眼中看为恶的事，惹我发怒。”
2KGS|21|16|玛拿西 行耶和华眼中看为恶的事，使 犹大 陷入罪里，又流许多无辜人的血，直到这血充满了 耶路撒冷 ，从这边到那边。
2KGS|21|17|玛拿西 其余的事，凡他所做的和他所犯的罪，不都写在《犹大列王记》上吗？
2KGS|21|18|玛拿西 与他祖先同睡，葬在自己王宫的园子， 乌撒 园里，他儿子 亚们 接续他作王。
2KGS|21|19|亚们 登基的时候年二十二岁，在 耶路撒冷 作王二年。他母亲名叫 米舒利密 ，是 约提巴 人 哈鲁斯 的女儿。
2KGS|21|20|亚们 行耶和华眼中看为恶的事，效法他父亲 玛拿西 所行的。
2KGS|21|21|他行他父亲一切所行的道，事奉他父亲所事奉的偶像，敬拜它们，
2KGS|21|22|离弃耶和华－他列祖的上帝，不遵行耶和华的道。
2KGS|21|23|亚们 的臣仆背叛他，在宫里杀了王。
2KGS|21|24|但这地的百姓杀了所有背叛 亚们 王的人；这地的百姓立他儿子 约西亚 接续他作王。
2KGS|21|25|亚们 其余所做的事，不都写在《犹大列王记》上吗？
2KGS|21|26|亚们 葬在 乌撒 园内自己的坟墓里，他儿子 约西亚 接续他作王。
2KGS|22|1|约西亚 登基的时候年八岁，在 耶路撒冷 作王三十一年。他母亲名叫 耶底大 ，是 波斯加 人 亚大雅 的女儿。
2KGS|22|2|约西亚 行耶和华眼中看为正的事，行他祖先 大卫 一切所行的道，不偏左右。
2KGS|22|3|约西亚 王十八年，王派 米书兰 的孙子， 亚萨利雅 的儿子 沙番 书记上耶和华殿去，说：
2KGS|22|4|“你上到 希勒家 大祭司那里，请他把奉献到耶和华殿的银子，就是门口的守卫从百姓中收来的银子，结算清楚，
2KGS|22|5|交在管理耶和华殿督工的手里，由他们支付给在耶和华殿里做工的人，好修理殿的破坏之处，
2KGS|22|6|就是木匠、工人和瓦匠，又买木料和凿成的石头，来整修殿宇。
2KGS|22|7|但他们不用跟这些经手接受银子的人算帐，因为这些人办事诚实。”
2KGS|22|8|希勒家 大祭司对 沙番 书记说：“我在耶和华殿里发现了律法书。” 希勒家 把书递给 沙番 ， 沙番 就读了。
2KGS|22|9|沙番 书记到王那里，把这事回覆王说：“你的仆人已把殿里所发现的银子倒出来，交在管理耶和华殿督工的手里了。”
2KGS|22|10|沙番 书记又向王报告说：“ 希勒家 祭司递给我一卷书。” 沙番 就在王面前朗读那书。
2KGS|22|11|王听见律法书上的话，就撕裂衣服。
2KGS|22|12|王吩咐 希勒家 祭司与 沙番 的儿子 亚希甘 、 米该亚 的儿子 亚革波 、 沙番 书记和王的臣仆 亚撒雅 ，说：
2KGS|22|13|“你们去，以所发现这书上的话，为我、为百姓、为全 犹大 求问耶和华；因为我们祖先没有听从这书上的话，没有遵照一切所写有关我们的 去行，耶和华就向我们大发烈怒。”
2KGS|22|14|于是， 希勒家 祭司和 亚希甘 、 亚革波 、 沙番 、 亚撒雅 都去见 户勒大 女先知，她是掌管礼服的 沙龙 的妻子； 沙龙 是 哈珥哈斯 的孙子， 特瓦 的儿子。 户勒大 住在 耶路撒冷 第二区。他们向她请教。
2KGS|22|15|她对他们说：“耶和华－ 以色列 的上帝如此说：‘你们可以回覆那派你们来见我的人说，
2KGS|22|16|耶和华如此说：看哪，我必照着 犹大 王所读那书上的一切话，降祸于这地方和其上的居民。
2KGS|22|17|因为他们离弃我，向别神烧香，用他们手所做的一切惹我发怒，所以我的愤怒必向这地方发作，总不止息。’
2KGS|22|18|然而，派你们来求问耶和华的 犹大 王，你们要这样回覆他：‘耶和华－ 以色列 的上帝如此说：至于你所听见的话，
2KGS|22|19|就是听见我指着这地方和其上的居民说，要使这地方变为荒芜、百姓受诅咒的话，你的心就软化，在耶和华面前谦卑下来，撕裂衣服，向我哭泣，因此我应允你。这是耶和华说的。
2KGS|22|20|因此，看哪，我必使你归到你祖先那里，平安地进入坟墓；我要降于这地方的一切灾祸，你不会亲眼看见。’”他们就去把这话回覆王。
2KGS|23|1|王派人召集 犹大 和 耶路撒冷 的众长老来。
2KGS|23|2|王和 犹大 众人、 耶路撒冷 的居民、祭司、先知，以及所有的百姓，无论大小，都一同上到耶和华的殿去；王把耶和华殿里所发现的约书上一切的话读给他们听。
2KGS|23|3|王站在柱子旁边，在耶和华面前立约，要尽心尽性跟从耶和华，遵守他的诫命、法度、律例，实行这书上所写这约的话。全体百姓都愿遵守所立的约。
2KGS|23|4|王吩咐 希勒家 大祭司和副祭司，以及把守殿门的，把那些为 巴力 和 亚舍拉 ，以及天上万象所造的器皿，都从耶和华殿里搬出来，在 耶路撒冷 外 汲沦 的田间烧了，把灰拿到 伯特利 去。
2KGS|23|5|从前 犹大 列王所立拜偶像的祭司，在 犹大 城镇的丘坛和 耶路撒冷 周围烧香，现在王都废去，他们是向 巴力 和日、月、行星，以及天上万象烧香的人。
2KGS|23|6|他把 亚舍拉 从耶和华殿里搬到 耶路撒冷 外的 汲沦溪 ，在 汲沦溪 边焚烧，打碎成灰，把灰撒在平民的坟上。
2KGS|23|7|他又拆毁耶和华殿里男的庙妓的屋子，就是妇女在那里为 亚舍拉 编织衣服的屋子。
2KGS|23|8|他从 犹大 的城镇将众祭司带来，从 迦巴 直到 别是巴 ，玷污祭司烧香的丘坛。他又拆毁城门旁的丘坛，这丘坛是在 约书亚 市长的城门前，在人进城门的左边。
2KGS|23|9|只是丘坛的祭司不登 耶路撒冷 耶和华的坛，仅在他们弟兄中间吃无酵饼。
2KGS|23|10|他又玷污 欣嫩子谷 的 陀斐特 ，不许人在那里使儿女经火献给 摩洛 。
2KGS|23|11|他把在耶和华殿门旁、靠近 拿单．米勒 官员走廊的屋子， 犹大 列王献给太阳的马废去，且用火焚烧献给太阳的战车。
2KGS|23|12|犹大 列王在 亚哈斯 楼房顶上所筑的坛和 玛拿西 在耶和华殿两院中所筑的坛，王都拆毁，从那里移走 ，把灰倒在 汲沦溪 中。
2KGS|23|13|从前 以色列 王 所罗门 在 耶路撒冷 东边、 邪僻山 南边为 西顿 人可憎的 亚斯她录 、 摩押 人可憎的 基抹 、 亚扪 人可憎的 米勒公 所筑的丘坛，王都玷污了，
2KGS|23|14|又打碎柱像，砍下 亚舍拉 ，用人的骨头填满那地方。
2KGS|23|15|此外，在 伯特利 丘坛的坛，就是 尼八 的儿子 耶罗波安 所筑、使 以色列 人陷入罪里的，他也把这坛和丘坛都拆毁了，又焚烧丘坛 ，打碎成灰，并焚烧了 亚舍拉 。
2KGS|23|16|约西亚 转头，看见山上的坟墓，就派人取出坟墓里的骸骨，烧在坛上，玷污了坛，正如从前 耶罗波安 在节期中站在坛旁时，耶和华藉神人所宣告的话。 约西亚 转头看见了宣告这些话的神人的坟墓。
2KGS|23|17|他说：“我看见的这碑是什么呢？”那城里的人对他说：“这是神人的坟墓，他从 犹大 来，宣告了王向 伯特利 的坛所做的这些事。”
2KGS|23|18|约西亚 说：“让他安息吧！不要挪移他的骸骨。”他们就保存了他的骸骨和从 撒玛利亚 来的那先知的骸骨。
2KGS|23|19|从前 以色列 诸王在 撒玛利亚 的城镇所建一切惹动怒气的丘坛的庙， 约西亚 也都废去了，正如他在 伯特利 所做的。
2KGS|23|20|他又把在那里所有丘坛的祭司都杀在坛上，并在坛上烧人的骨头。于是他回 耶路撒冷 去了。
2KGS|23|21|王吩咐众百姓说：“你们当照这约书上所写的，向耶和华－你们的上帝守逾越节。”
2KGS|23|22|自从士师治理 以色列 ，到 以色列 诸王、 犹大 列王在位的一切日子，从来没有守过这样的逾越节，
2KGS|23|23|只有在 约西亚 王十八年，才在 耶路撒冷 向耶和华守这逾越节。
2KGS|23|24|此外，在 犹大 地和 耶路撒冷 所见那些招魂的、行巫术的，家中的神像和偶像，以及一切可憎之物， 约西亚 尽都除掉，实行了 希勒家 祭司在耶和华殿里所发现的律法书上所写的话。
2KGS|23|25|在 约西亚 以前，没有王像他尽心、尽性、尽力地归向耶和华，遵行 摩西 的一切律法；在他以后，也没有兴起一个王像他。
2KGS|23|26|然而，耶和华向 犹大 所发猛烈的怒气仍不止息，因为 玛拿西 种种的恶事激怒了他。
2KGS|23|27|耶和华说：“我也必将 犹大 从我面前赶出，如同赶出 以色列 一样。我必撇弃我从前所选择的这城 耶路撒冷 和我所说我的名必留在那里的殿。”
2KGS|23|28|约西亚 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
2KGS|23|29|约西亚 的日子， 埃及 王法老 尼哥 上到 幼发拉底河 ，到 亚述 王那里； 约西亚 王去迎击他。 埃及 王在 米吉多 看见 约西亚 ，就杀了他。
2KGS|23|30|他的臣仆用车把他的尸体从 米吉多 送到 耶路撒冷 ，葬在他自己的坟墓里。这地的百姓选 约西亚 的儿子 约哈斯 ，膏立他，接续他父亲作王。
2KGS|23|31|约哈斯 登基的时候年二十三岁，在 耶路撒冷 作王三个月。他母亲名叫 哈慕她 ，是 立拿 人 耶利米 的女儿。
2KGS|23|32|约哈斯 行耶和华眼中看为恶的事，效法他祖先一切所行的。
2KGS|23|33|法老 尼哥 把 约哈斯 监禁在 哈马 地的 利比拉 ，不许他在 耶路撒冷 作王 ，又罚这地一百他连得银子，一他连得金子。
2KGS|23|34|法老 尼哥 立 约西亚 的儿子 以利亚敬 接续他父亲 约西亚 作王，给他改名叫 约雅敬 ，却把 约哈斯 带到 埃及 ，他就死在那里。
2KGS|23|35|约雅敬 进贡金银给法老，照着法老的指示在这地征收银子，向这地的百姓按各人的能力索取金银，要送给法老 尼哥 。
2KGS|23|36|约雅敬 登基的时候年二十五岁，在 耶路撒冷 作王十一年。他母亲名叫 西布大 ，是 鲁玛 人 毗大雅 的女儿。
2KGS|23|37|约雅敬 行耶和华眼中看为恶的事，效法他祖先一切所行的。
2KGS|24|1|约雅敬 的日子， 巴比伦 王 尼布甲尼撒 上来； 约雅敬 服事他三年，以后又背叛他。
2KGS|24|2|耶和华派 迦勒底 、 亚兰 、 摩押 和 亚扪 人的军队来攻击 约雅敬 ；耶和华派他们来攻击 犹大 ，要毁灭它，正如耶和华藉他仆人众先知所说的话。
2KGS|24|3|这事临到 犹大 ，诚然是出于耶和华的命令 ，要把 犹大 从自己面前赶出去，是因 玛拿西 所犯的一切罪，
2KGS|24|4|又因他流无辜人的血，使无辜人的血充满 耶路撒冷 ；耶和华不愿赦免。
2KGS|24|5|约雅敬 其余的事，凡他所做的，不都写在《犹大列王记》上吗？
2KGS|24|6|约雅敬 与他祖先同睡，他儿子 约雅斤 接续他作王。
2KGS|24|7|埃及 王不再从他的国出征，因为 巴比伦 王把 埃及 王所管之地，从 埃及 溪谷直到 幼发拉底河 都夺去了。
2KGS|24|8|约雅斤 登基的时候年十八岁，在 耶路撒冷 作王三个月。他母亲名叫 尼护施她 ，是 耶路撒冷 人 以利拿单 的女儿。
2KGS|24|9|约雅斤 行耶和华眼中看为恶的事，效法他父亲一切所行的。
2KGS|24|10|那时， 巴比伦 王 尼布甲尼撒 的军兵上到 耶路撒冷 ，城被围困。
2KGS|24|11|当他的军兵围困城的时候， 巴比伦 王 尼布甲尼撒 亲自来到 耶路撒冷 。
2KGS|24|12|犹大 王 约雅斤 和他母亲、臣仆、王子、官员一同出来，向 巴比伦 王投降。 巴比伦 王俘掳了他，那时是 巴比伦 王第八年。
2KGS|24|13|巴比伦 王把耶和华殿里和王宫里一切的宝物从那里拿走，又把 以色列 王 所罗门 所造耶和华殿里一切的金器都毁坏了，正如耶和华所说的。
2KGS|24|14|他把全 耶路撒冷 众领袖和所有大能的勇士，共一万人，连同所有的木匠和铁匠都掳了去，只留下这地最贫穷的百姓。
2KGS|24|15|他把 约雅斤 和他的母亲、后妃、官员，以及这地的贵族，都从 耶路撒冷 掳到 巴比伦 去了，
2KGS|24|16|又把所有的勇士七千人，木匠和铁匠一千人，全是能上阵的勇士，都掳到 巴比伦 去了。
2KGS|24|17|巴比伦 王立 约雅斤 的叔父 玛探雅 取代他作王，给 玛探雅 改名叫 西底家 。
2KGS|24|18|西底家 登基的时候年二十一岁，在 耶路撒冷 作王十一年。他母亲名叫 哈慕她 ，是 立拿 人 耶利米 的女儿。
2KGS|24|19|西底家 行耶和华眼中看为恶的事，正如 约雅敬 一切所行的。
2KGS|24|20|因此，耶和华向 耶路撒冷 和 犹大 发怒，以致把他们从自己面前赶出去。 西底家 背叛 巴比伦 王。
2KGS|25|1|西底家 作王第九年十月初十， 巴比伦 王 尼布甲尼撒 率领全军前来攻击 耶路撒冷 ，对城安营，四围筑堡垒攻城。
2KGS|25|2|城被围困，直到 西底家 王十一年。
2KGS|25|3|四月初九，城里的饥荒非常严重，当地的百姓都没有粮食。
2KGS|25|4|城被攻破，士兵全都在夜间从靠近王的花园、两城墙中间的门逃跑。 迦勒底 人正在四围攻城，王就往 亚拉巴 逃去。
2KGS|25|5|迦勒底 的军队追赶王，在 耶利哥 的平原追上他；他的全军都离开他溃散了。
2KGS|25|6|迦勒底 人就拿住王，带他到 利比拉 的 巴比伦 王那里；他们就判他的罪。
2KGS|25|7|他们在 西底家 眼前杀了他的儿女，挖了 西底家 的眼睛，用铜链锁着他，带到 巴比伦 去。
2KGS|25|8|巴比伦 王 尼布甲尼撒 十九年五月初七， 巴比伦 王的臣仆 尼布撒拉旦 护卫长进入 耶路撒冷 ，
2KGS|25|9|他焚烧了耶和华的殿、王宫和 耶路撒冷 一切的房屋；用火焚烧所有大户人家的房屋。
2KGS|25|10|跟从护卫长的 迦勒底 全军拆毁了 耶路撒冷 四围的城墙。
2KGS|25|11|那时 尼布撒拉旦 护卫长将城里剩下的百姓和那些投降 巴比伦 王的人，以及其余的众人，都掳去了。
2KGS|25|12|但护卫长留下一些当地最穷的人，叫他们修整葡萄园，耕种田地。
2KGS|25|13|耶和华殿的铜柱并殿内的盆座和铜海， 迦勒底 人都打碎了，把那些铜运到 巴比伦 去。
2KGS|25|14|他们又带走锅、铲子、钳子、勺子和供奉用的一切铜器；
2KGS|25|15|火盆和碗，无论金的银的，护卫长都带走了；
2KGS|25|16|还有 所罗门 为耶和华殿所造的两根柱子、一个铜海和盆座，这一切器皿的铜多得无法可秤。
2KGS|25|17|这一根柱子高十八肘，柱上有铜顶，铜顶高三肘；铜顶的周围有网子和石榴，也都是铜的。第二根柱子与此相同，也有网子。
2KGS|25|18|护卫长拿住 西莱雅 大祭司、 西番亚 副祭司和门口的三个守卫，
2KGS|25|19|又从城中拿住一个管理士兵的官 ，并在城里所找到王面前的五个亲信，和召募当地百姓之将军的书记官，以及在城中找到的六十个当地百姓。
2KGS|25|20|尼布撒拉旦 护卫长把这些人带到 利比拉 的 巴比伦 王那里。
2KGS|25|21|巴比伦 王击杀他们，在 哈马 地的 利比拉 把他们处死。这样， 犹大 人就被掳去离开本地。
2KGS|25|22|至于 犹大 地剩下的百姓，就是 巴比伦 王 尼布甲尼撒 所留下的， 巴比伦 王立了 沙番 的孙子， 亚希甘 的儿子 基大利 作他们的省长。
2KGS|25|23|所有的军官和属他们的人听见 巴比伦 王立了 基大利 作省长， 尼探雅 的儿子 以实玛利 、 加利亚 的儿子 约哈难 、 尼陀法 人 单户蔑 的儿子 西莱雅 、 玛迦 人的儿子 雅撒尼亚 ，和属他们的人，都来到 米斯巴 的 基大利 那里。
2KGS|25|24|基大利 向他们和属他们的人起誓说：“你们不必惧怕 迦勒底 臣仆，只管住在这地，服事 巴比伦 王，就可以得福。”
2KGS|25|25|七月中，王室后裔 以利沙玛 的孙子， 尼探雅 的儿子 以实玛利 带着十个人来，击杀了 基大利 和同他在 米斯巴 的 犹大 人与 迦勒底 人，把他们杀死。
2KGS|25|26|于是众人，无论大小，连同军官，因为惧怕 迦勒底 人，都起身逃到 埃及 去了。
2KGS|25|27|巴比伦 王 以未．米罗达 作王的元年，就是 犹大 王 约雅斤 被掳后三十七年，十二月二十七日，他使 犹大 王 约雅斤 抬起头来，提他出监，
2KGS|25|28|对他说好话，使他的位高过与他一同被掳在 巴比伦 众王的位；
2KGS|25|29|又给他脱了囚服，使他终身常在 巴比伦 王面前吃饭。
2KGS|25|30|王赐给他日常需用的食物，每日一份，终身都是这样。
1CHR|1|1|亚当 ， 塞特 ， 以挪士 ，
1CHR|1|2|该南 ， 玛勒列 ， 雅列 ，
1CHR|1|3|以诺 ， 玛土撒拉 ， 拉麦 ，
1CHR|1|4|挪亚 ， 闪 ， 含 ， 雅弗 。
1CHR|1|5|雅弗 的儿子是 歌篾 、 玛各 、 玛代 、 雅完 、 土巴 、 米设 和 提拉 。
1CHR|1|6|歌篾 的儿子是 亚实基拿 、 低法 和 陀迦玛 。
1CHR|1|7|雅完 的儿子是 以利沙 、 他施 、 基提 和 罗单 人 。
1CHR|1|8|含 的儿子是 古实 、 麦西 、 弗 和 迦南 。
1CHR|1|9|古实 的儿子是 西巴 、 哈腓拉 、 撒弗他 、 拉玛 和 撒弗提迦 。 拉玛 的儿子是 示巴 和 底但 。
1CHR|1|10|古实 又生 宁录 ，他是地上第一个勇士。
1CHR|1|11|麦西 生 路低 人、 亚拿米 人、 利哈比 人、 拿弗土希 人、
1CHR|1|12|帕斯鲁细 人、 迦斯路希 人和 迦斐托 人； 非利士 人是从 迦斐托 人 出来的。
1CHR|1|13|迦南 生了长子 西顿 ，又生 赫
1CHR|1|14|和 耶布斯 人、 亚摩利 人、 革迦撒 人、
1CHR|1|15|希未 人、 亚基 人、 西尼 人、
1CHR|1|16|亚瓦底 人、 洗玛利 人和 哈马 人。
1CHR|1|17|闪 的儿子是 以拦 、 亚述 、 亚法撒 、 路德 、 亚兰 、 乌斯 、 户勒 、 基帖 和 米设 。
1CHR|1|18|亚法撒 生 沙拉 ； 沙拉 生 希伯 。
1CHR|1|19|希伯 生了两个儿子：一个名叫 法勒 ，因为那时人分地居住； 法勒 的兄弟名叫 约坍 。
1CHR|1|20|约坍 生 亚摩答 、 沙列 、 哈萨玛非 、 耶拉 、
1CHR|1|21|哈多兰 、 乌萨 、 德拉 、
1CHR|1|22|以巴录 、 亚比玛利 、 示巴 、
1CHR|1|23|阿斐 、 哈腓拉 和 约巴 。这些都是 约坍 的儿子。
1CHR|1|24|闪 ， 亚法撒 ， 沙拉 ，
1CHR|1|25|希伯 ， 法勒 ， 拉吴 ，
1CHR|1|26|西鹿 ， 拿鹤 ， 他拉 ，
1CHR|1|27|亚伯兰 ， 亚伯兰 就是 亚伯拉罕 。
1CHR|1|28|亚伯拉罕 的儿子是 以撒 和 以实玛利 。
1CHR|1|29|以实玛利 的后代如下： 以实玛利 的长子是 尼拜约 ，又有 基达 、 亚德别 、 米比衫 、
1CHR|1|30|米施玛 、 度玛 、 玛撒 、 哈大 、 提玛 、
1CHR|1|31|伊突 、 拿非施 和 基底玛 。这些都是 以实玛利 的儿子。
1CHR|1|32|亚伯拉罕 的妾 基土拉 所生的儿子，就是 心兰 、 约珊 、 米但 、 米甸 、 伊施巴 和 书亚 。 约珊 的儿子是 示巴 和 底但 。
1CHR|1|33|米甸 的儿子是 以法 、 以弗 、 哈诺 、 亚比大 和 以勒大 。这些都是 基土拉 的子孙。
1CHR|1|34|亚伯拉罕 生 以撒 ； 以撒 的儿子是 以扫 和 以色列 。
1CHR|1|35|以扫 的儿子是 以利法 、 流珥 、 耶乌施 、 雅兰 和 可拉 。
1CHR|1|36|以利法 的儿子是 提幔 、 阿抹 、 洗玻 、 迦坦 、 基纳斯 、 亭纳 和 亚玛力 。
1CHR|1|37|流珥 的儿子是 拿哈 、 谢拉 、 沙玛 和 米撒 。
1CHR|1|38|西珥 的儿子是 罗坍 、 朔巴 、 祭便 、 亚拿 、 底顺 、 以察 和 底珊 。
1CHR|1|39|罗坍 的儿子是 何利 和 荷幔 ； 罗坍 的妹妹是 亭纳 。
1CHR|1|40|朔巴 的儿子是 亚勒文 、 玛拿辖 、 以巴录 、 示非 和 阿南 。 祭便 的儿子是 爱亚 和 亚拿 。
1CHR|1|41|亚拿 的儿子是 底顺 。 底顺 的儿子是 哈默兰 、 伊是班 、 益兰 和 基兰 。
1CHR|1|42|以察 的儿子是 辟罕 、 撒番 ，和 亚干 。 底珊 的儿子是 乌斯 和 亚兰 。
1CHR|1|43|以色列 人未有君王治理之前，这些是在 以东 地作王的。有 比珥 的儿子 比拉 ，他的城名叫 亭哈巴 。
1CHR|1|44|比拉 死了， 波斯拉 人 谢拉 的儿子 约巴 接续他作王。
1CHR|1|45|约巴 死了， 提幔 人之地的 户珊 接续他作王。
1CHR|1|46|户珊 死了， 比达 的儿子 哈达 接续他作王， 哈达 曾在 摩押 地击败 米甸 人，他的城名叫 亚未得 。
1CHR|1|47|哈达 死了， 玛士利加 人 桑拉 接续他作王。
1CHR|1|48|桑拉 死了， 大河 边的 利河伯 人 扫罗 接续他作王。
1CHR|1|49|扫罗 死了， 亚革波 的儿子 巴勒．哈南 接续他作王。
1CHR|1|50|巴勒．哈南 死了， 哈达 接续他作王，他的城名叫 巴伊 。他的妻子名叫 米希她别 ，是 米．萨合 的孙女， 玛特列 的女儿。
1CHR|1|51|哈达 死了。 以东 的族长有： 亭纳 族长、 亚勒瓦 族长、 耶帖 族长、
1CHR|1|52|阿何利巴玛 族长、 以拉 族长、 比嫩 族长、
1CHR|1|53|基纳斯 族长、 提幔 族长、 米比萨 族长、
1CHR|1|54|玛基叠 族长、 以兰 族长。这些都是 以东 的族长。
1CHR|2|1|以色列 的儿子是 吕便 、 西缅 、 利未 、 犹大 、 以萨迦 、 西布伦 、
1CHR|2|2|但 、 约瑟 、 便雅悯 、 拿弗他利 、 迦得 和 亚设 。
1CHR|2|3|犹大 的儿子是 珥 、 俄南 和 示拉 ，这三人是 迦南 女子 拔．书亚 所生的。 犹大 的长子 珥 在耶和华眼中看为恶，耶和华就杀死了他。
1CHR|2|4|犹大 的媳妇 她玛 为 犹大 生了 法勒斯 和 谢拉 。 犹大 共有五个儿子。
1CHR|2|5|法勒斯 的儿子是 希斯仑 和 哈母勒 。
1CHR|2|6|谢拉 的儿子是 心利 、 以探 、 希幔 、 甲各 和 大拉 ，共五人。
1CHR|2|7|迦米 的儿子是 亚迦 ，他在当灭的物上犯了罪，连累了 以色列 人。
1CHR|2|8|以探 的儿子是 亚撒利雅 。
1CHR|2|9|希斯仑 所生的儿子是 耶拉篾 、 兰 和 基路拜 。
1CHR|2|10|兰 生 亚米拿达 ； 亚米拿达 生 拿顺 ， 拿顺 是 犹大 人的领袖。
1CHR|2|11|拿顺 生 撒门 ； 撒门 生 波阿斯 ；
1CHR|2|12|波阿斯 生 俄备得 ； 俄备得 生 耶西 ；
1CHR|2|13|耶西 生长子 以利押 ，次子 亚比拿达 ，三子 示米亚 ，
1CHR|2|14|四子 拿坦业 ，五子 拉代 ，
1CHR|2|15|六子 阿鲜 ，七子 大卫 。
1CHR|2|16|他们的姊妹是 洗鲁雅 和 亚比该 。 洗鲁雅 的儿子是 亚比筛 、 约押 和 亚撒黑 ，共三人。
1CHR|2|17|亚比该 生 亚玛撒 ； 亚玛撒 的父亲是 以实玛利 人 益帖 。
1CHR|2|18|希斯仑 的儿子 迦勒 娶 阿苏巴 和 耶略 为妻， 阿苏巴 的儿子是 耶设 、 朔罢 和 押墩 。
1CHR|2|19|阿苏巴 死了， 迦勒 又娶 以法她 ，生了 户珥 。
1CHR|2|20|户珥 生 乌利 ； 乌利 生 比撒列 。
1CHR|2|21|后来， 希斯仑 六十岁时娶了 基列 的父亲 玛吉 的女儿，与她同房； 玛吉 的女儿为他生了 西割 ；
1CHR|2|22|西割 生 睚珥 。 睚珥 在 基列 地有二十三座城。
1CHR|2|23|后来 基述 和 亚兰 夺了 哈倭特．睚珥 ，以及 基纳 和所属的乡镇 ，共六十个。这些城镇的人全都是 基列 的父亲 玛吉 的子孙。
1CHR|2|24|希斯仑 在 迦勒．以法他 死后，他的妻子 亚比雅 为他生了 提哥亚 的父亲 亚施户 。
1CHR|2|25|希斯仑 的长子 耶拉篾 的儿子有长子 兰 、 布拿 、 阿连 、 阿鲜 和 亚希雅 。
1CHR|2|26|耶拉篾 又娶一妻名叫 亚她拉 ，是 阿南 的母亲。
1CHR|2|27|耶拉篾 的长子 兰 的儿子有 玛斯 、 雅悯 和 以结 。
1CHR|2|28|阿南 的儿子是 沙买 和 雅大 。 沙买 的儿子是 拿答 和 亚比述 。
1CHR|2|29|亚比述 的妻子名叫 亚比孩 ，为他生了 亚办 和 摩利 。
1CHR|2|30|拿答 的儿子是 西列 和 亚遍 ； 西列 死了，没有儿子。
1CHR|2|31|亚遍 的儿子是 以示 ； 以示 的儿子是 示珊 ； 示珊 的儿子是 亚来 。
1CHR|2|32|沙买 的兄弟 雅大 的儿子是 益帖 和 约拿单 ； 益帖 死了，没有儿子。
1CHR|2|33|约拿单 的儿子是 比勒 和 撒萨 。这些都是 耶拉篾 的子孙。
1CHR|2|34|示珊 没有儿子，只有女儿。 示珊 有一个仆人名叫 耶哈 ，是 埃及 人。
1CHR|2|35|示珊 把女儿嫁给仆人 耶哈 ，她为他生了 亚太 。
1CHR|2|36|亚太 生 拿单 ； 拿单 生 撒拔 ；
1CHR|2|37|撒拔 生 以弗拉 ； 以弗拉 生 俄备得 ；
1CHR|2|38|俄备得 生 耶户 ； 耶户 生 亚撒利雅 ；
1CHR|2|39|亚撒利雅 生 希利斯 ； 希利斯 生 以利亚萨 ；
1CHR|2|40|以利亚萨 生 西斯买 ； 西斯买 生 沙龙 ；
1CHR|2|41|沙龙 生 耶加米雅 ； 耶加米雅 生 以利沙玛 。
1CHR|2|42|耶拉篾 的兄弟 迦勒 的众儿子：长子是 米沙 ， 米沙 是 西弗 的父亲，还有 希伯伦 的父亲 玛利沙 的众儿子。
1CHR|2|43|希伯伦 的儿子是 可拉 、 他普亚 、 利肯 和 示玛 。
1CHR|2|44|示玛 生 拉含 ，是 约干 之祖。 利肯 生 沙买 。
1CHR|2|45|沙买 的儿子是 玛云 ； 玛云 是 伯．夙 的父亲。
1CHR|2|46|迦勒 的妾 以法 生 哈兰 、 摩撒 和 迦谢 ； 哈兰 生 迦卸 。
1CHR|2|47|雅代 的儿子是 利健 、 约坦 、 基珊 、 毗力 、 以法 和 沙亚弗 。
1CHR|2|48|迦勒 的妾 玛迦 生 示别 和 特哈拿 ，
1CHR|2|49|又生 麦玛拿 的父亲 沙亚弗 ，又生 抹比拿 和 基比亚 的父亲 示法 。 迦勒 的女儿是 押撒 。
1CHR|2|50|这些都是 迦勒 的子孙。 以法她 的长子 户珥 的子孙： 基列．耶琳 之祖 朔巴 ，
1CHR|2|51|伯利恒 之祖 萨玛 ， 伯．迦得 之祖 哈勒 。
1CHR|2|52|基列．耶琳 之祖 朔巴 的子孙是 哈罗以 和一半的 米努哈 人 。
1CHR|2|53|基列．耶琳 的宗族有 以帖 人、 布特 人、 舒玛 人、 密来 人，又从这些宗族生出 琐拉 人和 以实陶 人。
1CHR|2|54|萨玛 的子孙有 伯利恒 人、 尼陀法 人、 亚他绿．伯．约押 人、一半的 玛拿哈 人、 琐利 人。
1CHR|2|55|住 雅比斯 的文士的宗族有 特拉 人、 示米押 人和 苏甲 人。这些都是 利甲 家之祖 哈末 所生的 基尼 人。
1CHR|3|1|大卫 在 希伯仑 所生的儿子如下：长子 暗嫩 是 耶斯列 人 亚希暖 生的。次子 但以利 是 迦密 人 亚比该 生的。
1CHR|3|2|三子 押沙龙 是 基述 王 达买 的女儿 玛迦 生的。四子 亚多尼雅 是 哈及 生的。
1CHR|3|3|五子 示法提雅 是 亚比她 生的。六子 以特念 是 大卫 的妻子 以格拉 生的。
1CHR|3|4|这六人都是 大卫 在 希伯仑 生的。 大卫 在 希伯仑 作王七年六个月，在 耶路撒冷 作王三十三年。
1CHR|3|5|大卫 在 耶路撒冷 所生的儿子是 示米亚 、 朔罢 、 拿单 和 所罗门 。这四人是 亚米利 的女儿 拔．书亚 生的。
1CHR|3|6|还有 益辖 、 以利沙玛 、 以利法列 、
1CHR|3|7|挪迦 、 尼斐 、 雅非亚 、
1CHR|3|8|以利沙玛 、 以利雅大 、 以利法列 ，共九人。
1CHR|3|9|这些全都是 大卫 的儿子，妃嫔的儿子不在其内； 她玛 是他们的妹妹。
1CHR|3|10|所罗门 的后裔如下： 罗波安 ，他的儿子 亚比雅 ，他的儿子 亚撒 ，他的儿子 约沙法 ，
1CHR|3|11|他的儿子 约兰 ，他的儿子 亚哈谢 ，他的儿子 约阿施 ，
1CHR|3|12|他的儿子 亚玛谢 ，他的儿子 亚撒利雅 ，他的儿子 约坦 ；
1CHR|3|13|他的儿子 亚哈斯 ，他的儿子 希西家 ，他的儿子 玛拿西 ，
1CHR|3|14|他的儿子 亚们 ，他的儿子 约西亚 ，
1CHR|3|15|他的长子 约哈难 ，次子 约雅敬 ，三子 西底家 ，四子 沙龙 。
1CHR|3|16|约雅敬 的后裔：他的儿子 耶哥尼雅 ，他的儿子 西底家 。
1CHR|3|17|被掳的 耶哥尼雅 的后裔如下：他的儿子 撒拉铁 、
1CHR|3|18|玛基兰 、 毗大雅 、 示拿萨 、 耶加米 、 何沙玛 和 尼大比雅 。
1CHR|3|19|毗大雅 的儿子是 所罗巴伯 和 示每 。 所罗巴伯 的儿子是 米书兰 和 哈拿尼雅 ， 示罗密 是他们的妹妹；
1CHR|3|20|还有 哈舒巴 、 阿黑 、 比利家 、 哈撒底 、 于沙．希悉 ，共五人。
1CHR|3|21|哈拿尼雅 的儿子是 毗拉提 和 耶筛亚 。还有 利法雅 的众儿子， 亚珥难 的众儿子， 俄巴底亚 的众儿子， 示迦尼 的众儿子。
1CHR|3|22|示迦尼 的后裔： 示玛雅 ， 示玛雅 的儿子 哈突 、 以甲 、 巴利亚 、 尼利雅 、 沙法 ，共六人。
1CHR|3|23|尼利雅 的儿子是 以利约乃 、 希西家 、 亚斯利干 ，共三人。
1CHR|3|24|以利约乃 的儿子是 何大雅 、 以利亚实 、 毗莱雅 、 阿谷 、 约哈难 、 第莱雅 、 阿拿尼 ，共七人。
1CHR|4|1|犹大 的儿子是 法勒斯 、 希斯仑 、 迦米 、 户珥 和 朔巴 。
1CHR|4|2|朔巴 的儿子 利亚雅 生 雅哈 ； 雅哈 生 亚户买 和 拉哈 。这些是 琐拉 人的宗族。
1CHR|4|3|以坦 之祖 是 耶斯列 、 伊施玛 和 伊得巴 ；他们的妹妹名叫 哈悉勒玻尼 。
1CHR|4|4|基多 之祖是 毗努伊勒 。 户沙 之祖是 以谢珥 。这些都是 伯利恒 之祖， 以法她 的长子 户珥 的后裔。
1CHR|4|5|提哥亚 的父亲 亚施户 有两个妻子， 希拉 和 拿拉 。
1CHR|4|6|拿拉 为 亚施户 生 亚户撒 、 希弗 、 提米尼 和 哈辖斯他利 。这些都是 拿拉 的儿子。
1CHR|4|7|希拉 生的是 洗列 、 琐辖 和 伊提南 。
1CHR|4|8|哥斯 生 亚诺 、 琐比巴 和 哈仑 的儿子 亚哈黑 的宗族。
1CHR|4|9|雅比斯 比他众兄弟更尊贵，他母亲给他起名叫 雅比斯 ，意思说：“我生他甚是痛苦。”
1CHR|4|10|雅比斯 求告 以色列 的上帝说：“甚愿你赐福与我，扩张我的疆界，你的手常与我同在，保佑我不遭患难，不受艰苦。”上帝就应允他所求的。
1CHR|4|11|书哈 的兄弟 基绿 生 米黑 ， 米黑 是 伊施屯 的父亲。
1CHR|4|12|伊施屯 生 伯拉巴 、 巴西亚 和 珥．拿辖 之祖 提欣拿 。这些都是 利迦 人。
1CHR|4|13|基纳斯 的儿子是 俄陀聂 和 西莱雅 。 俄陀聂 的儿子是 哈塔 。
1CHR|4|14|悯挪太 生 俄弗拉 ； 西莱雅 生 革．夏纳欣 之祖 约押 。他们都是工匠。
1CHR|4|15|耶孚尼 的儿子 迦勒 的后裔： 以路 、 以拉 和 拿安 。 以拉 的儿子是 基纳斯 。
1CHR|4|16|耶哈利勒 的儿子是 西弗 、 西法 、 提利 和 亚撒列 。
1CHR|4|17|以斯拉 的儿子是 益帖 、 米列 、 以弗 和 雅伦 。 米列 所娶法老的女儿 比提雅 的后裔如下：她怀了 米利暗 、 沙买 ，和 以实提摩 之祖 益巴 。 米列 的 犹大 妻子生 基多 之祖 雅列 ， 梭哥 之祖 希伯 ，和 撒挪亚 之祖 耶古铁 。
1CHR|4|18|
1CHR|4|19|拿含 的妹妹， 荷第雅 的妻子所生的是 达利亚 ， 迦米 人 基伊拉 和 玛迦 人 以实提摩 的祖先。
1CHR|4|20|示门 的儿子是 暗嫩 、 林拿 、 便．哈南 和 提伦 。 以示 的儿子是 梭黑 和 便．梭黑 。
1CHR|4|21|犹大 的儿子 示拉 的后裔： 利迦 之祖 珥 ， 玛利沙 之祖 拉大 ，和住在 伯．亚实比 织细麻布的各宗族。
1CHR|4|22|还有 约敬 、 哥西巴 人、 约阿施 ，和那在 摩押 娶妻，回到 利恒 的 萨拉 。这都是古时的记载。
1CHR|4|23|这些人都是陶匠，是 尼他应 和 基底拉 的居民。他们住在王那里，为王做工。
1CHR|4|24|西缅 的后裔如下： 尼母利 、 雅悯 、 雅立 、 谢拉 和 扫罗 ；
1CHR|4|25|他的儿子 沙龙 ，他的儿子 米比衫 ，他的儿子 米施玛 ；
1CHR|4|26|米施玛 的后裔：他的儿子 哈母利 ，他的儿子 撒刻 ，他的儿子 示每 。
1CHR|4|27|示每 有十六个儿子和六个女儿，但他兄弟的儿女不多，他们各家族也不如 犹大 族那样人丁兴旺。
1CHR|4|28|西缅 人住在 别是巴 、 摩拉大 、 哈萨．书亚 、
1CHR|4|29|辟拉 、 以森 、 陀腊 、
1CHR|4|30|彼土利 、 何珥玛 、 洗革拉 、
1CHR|4|31|伯．玛加博 、 哈萨．苏撒 、 伯．比利 和 沙拉音 ，这些城镇直到 大卫 作王的时候都是属 西缅 人的；
1CHR|4|32|还有所属的村庄 以坦 、 亚因 、 临门 、 陀健 、 亚珊 ，共五个城镇；
1CHR|4|33|连同环绕这些城镇的一切乡村，直到 巴力 。这是他们的住处，他们都有家谱。
1CHR|4|34|还有 米所巴 、 雅米勒 、 亚玛谢 的儿子 约沙 、
1CHR|4|35|约珥 ，和 亚薛 的曾孙， 西莱雅 的孙子， 约示比 的儿子 耶户 。
1CHR|4|36|还有 以利约乃 、 雅哥巴 、 约朔海 、 亚帅雅 、 亚底业 、 耶西篾 、 比拿雅 、
1CHR|4|37|细撒 ； 细撒 是 示非 的儿子， 示非 是 亚龙 的儿子， 亚龙 是 耶大雅 的儿子， 耶大雅 是 申利 的儿子， 申利 是 示玛雅 的儿子。
1CHR|4|38|以上所记的人名都是作族长的，他们父系的家属大量增加。
1CHR|4|39|他们往平原东边 基多口 去，寻找牧放羊群的草场，
1CHR|4|40|找到了肥沃优美的草场，又宽阔又平静安宁之地；从前住那里的是 含 族的人。
1CHR|4|41|以上纪录上有名的人，在 犹大 王 希西家 的日子，来攻击 含 族人的帐棚和那里所有的 米乌尼 人，把他们灭尽，就住在他们的地方，直到今日，因为那里有草场可以牧放羊群。
1CHR|4|42|这些 西缅 人中有五百人上 西珥山 ，率领他们的是 以示 的儿子 毗拉提 、 尼利雅 、 利法雅 和 乌薛 。
1CHR|4|43|他们杀了 亚玛力 剩下的残存之民，就住在那里，直到今日。
1CHR|5|1|以色列 的长子 吕便 的后裔。 吕便 玷污了父亲的床，他长子的名分就归了 以色列 的儿子 约瑟 的后裔；因此，家谱就不按出生顺序登录。
1CHR|5|2|虽然 犹大 比他兄弟强盛，君王也从他而出，然而长子的名分却归 约瑟 。
1CHR|5|3|以色列 长子 吕便 的后裔如下： 哈诺 、 法路 、 希斯伦 和 迦米 。
1CHR|5|4|约珥 的后裔：他的儿子 示玛雅 ，他的儿子 歌革 ，他的儿子 示每 ，
1CHR|5|5|他的儿子 米迦 ，他的儿子 利亚雅 ，他的儿子 巴力 ，
1CHR|5|6|他的儿子 备拉 ；这 备拉 作 吕便 支派的领袖，被 亚述 王 提革拉．毗列色 掳去。
1CHR|5|7|他的弟兄照着宗族，按着家谱作族长的是 耶利 、 撒迦利雅 、
1CHR|5|8|比拉 ； 比拉 是 亚撒 的儿子， 亚撒 是 示玛 的儿子， 示玛 是 约珥 的儿子； 约珥 住在 亚罗珥 ，直到 尼波 和 巴力．免 。
1CHR|5|9|他也住在东边，直到 幼发拉底河 这边的旷野边界，因为他们在 基列 地牲畜增多。
1CHR|5|10|扫罗 年间，他们与 夏甲 人争战， 夏甲 人倒在他们手下，他们就在 基列 东边的全地，住在 夏甲 人的帐棚里。
1CHR|5|11|迦得 的后裔在 吕便 对面，住在 巴珊 地，延伸到 撒迦 ：
1CHR|5|12|有作族长的 约珥 ，有作副族长的 沙番 ，还有 雅乃 和住在 巴珊 的 沙法 。
1CHR|5|13|按着家族，他们的弟兄是 米迦勒 、 米书兰 、 示巴 、 约赖 、 雅干 、 细亚 和 希伯 ，共七人。
1CHR|5|14|这些都是 亚比孩 的儿子； 亚比孩 是 户利 的儿子， 户利 是 耶罗亚 的儿子， 耶罗亚 是 基列 的儿子， 基列 是 米迦勒 的儿子， 米迦勒 是 耶示筛 的儿子， 耶示筛 是 耶哈多 的儿子， 耶哈多 是 布斯 的儿子；
1CHR|5|15|古尼 的孙子， 押比叠 的儿子 亚希 是他们的族长。
1CHR|5|16|他们住在 基列 、 巴珊 和所属的乡镇，以及 沙仑 一切的郊野，直到四围的交界。
1CHR|5|17|这些人在 犹大 王 约坦 和 以色列 王 耶罗波安 年间，都载入家谱。
1CHR|5|18|吕便 人、 迦得 人和 玛拿西 半支派的人，能拿盾牌和刀剑、拉弓、出征善战的勇士共有四万四千七百六十名。
1CHR|5|19|他们与 夏甲 人、 伊突 人、 拿非施 人、 挪答 人打仗。
1CHR|5|20|他们在打仗的时候得了上帝的帮助， 夏甲 人和所有跟随 夏甲 人的人都交在他们手中；因为他们在阵上呼求上帝，倚赖他，他就应允他们。
1CHR|5|21|他们掳掠了 夏甲 人的牲畜，有五万匹骆驼，二十五万只羊，二千匹驴，又有十万人；
1CHR|5|22|被杀仆倒的很多，因为这战争是出乎上帝。他们就住在 夏甲 人的地上，直到被掳的时候。
1CHR|5|23|玛拿西 半支派的人住在那地，从 巴珊 延到 巴力．黑门 、 示尼珥 和 黑门山 ，他们人数增多 。
1CHR|5|24|他们的族长如下： 以弗 、 以示 、 以利业 、 亚斯列 、 耶利米 、 何达威雅 和 雅叠 ；他们都是大能的勇士，有名的人，是作族长的。
1CHR|5|25|但他们得罪了他们列祖的上帝，随从当地百姓的神明而行淫，这百姓就是上帝在他们面前所除灭的。
1CHR|5|26|因此， 以色列 的上帝激发 亚述 王 普勒 ，就是 亚述 王 提革拉．毗列色 的心，他掳掠了 吕便 人、 迦得 人、 玛拿西 半支派的人，把他们带到 哈腊 、 哈博 、 哈拉 与 歌散河 边，直到今日。
1CHR|6|1|利未 的后裔： 革顺 、 哥辖 和 米拉利 。
1CHR|6|2|哥辖 的儿子是 暗兰 、 以斯哈 、 希伯伦 和 乌薛 。
1CHR|6|3|暗兰 的儿女是 亚伦 、 摩西 和 米利暗 。 亚伦 的儿子是 拿答 、 亚比户 、 以利亚撒 和 以他玛 。
1CHR|6|4|以利亚撒 生 非尼哈 ； 非尼哈 生 亚比书 ；
1CHR|6|5|亚比书 生 布基 ； 布基 生 乌西 ；
1CHR|6|6|乌西 生 西拉希雅 ； 西拉希雅 生 米拉约 ；
1CHR|6|7|米拉约 生 亚玛利雅 ； 亚玛利雅 生 亚希突 ；
1CHR|6|8|亚希突 生 撒督 ； 撒督 生 亚希玛斯 ；
1CHR|6|9|亚希玛斯 生 亚撒利雅 ； 亚撒利雅 生 约哈难 ；
1CHR|6|10|约哈难 生 亚撒利雅 ， 亚撒利雅 在 所罗门 建造的 耶路撒冷 殿中担任祭司的职分；
1CHR|6|11|亚撒利雅 生 亚玛利雅 ； 亚玛利雅 生 亚希突 ；
1CHR|6|12|亚希突 生 撒督 ； 撒督 生 沙龙 ；
1CHR|6|13|沙龙 生 希勒家 ； 希勒家 生 亚撒利雅 ；
1CHR|6|14|亚撒利雅 生 西莱雅 ； 西莱雅 生 约萨答 。
1CHR|6|15|当耶和华藉 尼布甲尼撒 的手掳掠 犹大 和 耶路撒冷 的时候， 约萨答 也被掳去。
1CHR|6|16|利未 的后裔： 革顺 、 哥辖 和 米拉利 。
1CHR|6|17|革顺 的儿子名叫 立尼 和 示每 。
1CHR|6|18|哥辖 的儿子是 暗兰 、 以斯哈 、 希伯伦 和 乌薛 。
1CHR|6|19|米拉利 的儿子是 抹利 和 母示 。这是按着父系所分 利未 人的宗族。
1CHR|6|20|属 革顺 的：他的儿子 立尼 ，他的儿子 雅哈 ，他的儿子 薪玛 ，
1CHR|6|21|他的儿子 约亚 ，他的儿子 易多 ，他的儿子 谢拉 ，他的儿子 耶特赖 。
1CHR|6|22|哥辖 的后裔：他的儿子 亚米拿达 ，他的儿子 可拉 ，他的儿子 亚惜 ，
1CHR|6|23|他的儿子 以利加拿 ，他的儿子 以比雅撒 ，他的儿子 亚惜 ，
1CHR|6|24|他的儿子 他哈 ，他的儿子 乌列 ，他的儿子 乌西雅 ，他的儿子 少罗 。
1CHR|6|25|以利加拿 的儿子是 亚玛赛 、 亚希摩 、
1CHR|6|26|以利加拿 。 以利加拿 的后裔：他的儿子 琐菲 ，他的儿子 拿哈 ，
1CHR|6|27|他的儿子 以利押 ，他的儿子 耶罗罕 ，他的儿子 以利加拿 ，他的儿子 撒母耳 。
1CHR|6|28|撒母耳 的儿子是长子 约珥 和次子 亚比亚 。
1CHR|6|29|米拉利 的后裔： 抹利 ，他的儿子 立尼 ，他的儿子 示每 ，他的儿子 乌撒 ，
1CHR|6|30|他的儿子 示米亚 ，他的儿子 哈基雅 ，他的儿子 亚帅雅 。
1CHR|6|31|这些是约柜安设之后， 大卫 派在耶和华殿中管理歌唱事奉的人。
1CHR|6|32|他们在会幕前负责歌唱的事奉，及至 所罗门 在 耶路撒冷 建造了耶和华的殿，他们就按着班次供职。
1CHR|6|33|供职的人和他们的子孙如下： 哥辖 的子孙中有歌唱的 希幔 ； 希幔 是 约珥 的儿子， 约珥 是 撒母耳 的儿子，
1CHR|6|34|撒母耳 是 以利加拿 的儿子， 以利加拿 是 耶罗罕 的儿子， 耶罗罕 是 以利业 的儿子， 以利业 是 陀亚 的儿子，
1CHR|6|35|陀亚 是 苏弗 的儿子， 苏弗 是 以利加拿 的儿子， 以利加拿 是 玛哈 的儿子， 玛哈 是 亚玛赛 的儿子，
1CHR|6|36|亚玛赛 是 以利加拿 的儿子， 以利加拿 是 约珥 的儿子， 约珥 是 亚撒利雅 的儿子， 亚撒利雅 是 西番雅 的儿子，
1CHR|6|37|西番雅 是 他哈 的儿子， 他哈 是 亚惜 的儿子， 亚惜 是 以比雅撒 的儿子， 以比雅撒 是 可拉 的儿子，
1CHR|6|38|可拉 是 以斯哈 的儿子， 以斯哈 是 哥辖 的儿子， 哥辖 是 利未 的儿子， 利未 是 以色列 的儿子。
1CHR|6|39|希幔 的弟兄 亚萨 在 希幔 的右边供职； 亚萨 是 比利家 的儿子， 比利家 是 示米亚 的儿子，
1CHR|6|40|示米亚 是 米迦勒 的儿子， 米迦勒 是 巴西雅 的儿子， 巴西雅 是 玛基雅 的儿子，
1CHR|6|41|玛基雅 是 伊特尼 的儿子， 伊特尼 是 谢拉 的儿子， 谢拉 是 亚大雅 的儿子，
1CHR|6|42|亚大雅 是 以探 的儿子， 以探 是 薪玛 的儿子， 薪玛 是 示每 的儿子，
1CHR|6|43|示每 是 雅哈 的儿子， 雅哈 是 革顺 的儿子， 革顺 是 利未 的儿子。
1CHR|6|44|他们的弟兄 米拉利 的子孙，在他们左边供职的有 以探 ； 以探 是 基示 的儿子， 基示 是 亚伯底 的儿子， 亚伯底 是 玛鹿 的儿子，
1CHR|6|45|玛鹿 是 哈沙比雅 的儿子， 哈沙比雅 是 亚玛谢 的儿子， 亚玛谢 是 希勒家 的儿子，
1CHR|6|46|希勒家 是 暗西 的儿子， 暗西 是 巴尼 的儿子， 巴尼 是 沙麦 的儿子，
1CHR|6|47|沙麦 是 末力 的儿子， 末力 是 母示 的儿子， 母示 是 米拉利 的儿子， 米拉利 是 利未 的儿子。
1CHR|6|48|他们的弟兄 利未 人也被派办理上帝殿中帐幕的一切事务。
1CHR|6|49|亚伦 和他的子孙在燔祭坛和香坛上献祭烧香，办理至圣所一切的事，为 以色列 赎罪，正如上帝仆人 摩西 所吩咐的一切。
1CHR|6|50|亚伦 的后裔如下：他的儿子 以利亚撒 ，他的儿子 非尼哈 ，他的儿子 亚比书 ，
1CHR|6|51|他的儿子 布基 ，他的儿子 乌西 ，他的儿子 西拉希雅 ，
1CHR|6|52|他的儿子 米拉约 ，他的儿子 亚玛利雅 ，他的儿子 亚希突 ，
1CHR|6|53|他的儿子 撒督 ，他的儿子 亚希玛斯 。
1CHR|6|54|他们的住处按着境内的营寨如下： 亚伦 的子孙 哥辖 族先抽签得地，
1CHR|6|55|得了 犹大 地的 希伯仑 和四围的郊野；
1CHR|6|56|只是这城的田地和所属的村庄都为 耶孚尼 的儿子 迦勒 所得。
1CHR|6|57|亚伦 的子孙所得逃城如下： 希伯仑 、 立拿 与其郊野、 雅提珥 、 以实提莫 与其郊野、
1CHR|6|58|希仑 与其郊野、 底璧 与其郊野、
1CHR|6|59|亚珊 与其郊野、 伯．示麦 与其郊野。
1CHR|6|60|他们也从 便雅悯 支派中得了 迦巴 与其郊野、 阿勒篾 与其郊野、 亚拿突 与其郊野。他们宗族所得的城共十三座。
1CHR|6|61|哥辖 族其余的人抽签，按支派的宗族，从半个支派，就是 玛拿西 半支派中得了十座城。
1CHR|6|62|革顺 族按着宗族，从 以萨迦 支派、 亚设 支派、 拿弗他利 支派、 巴珊 内的 玛拿西 支派中，得了十三座城。
1CHR|6|63|米拉利 族按着宗族抽签，从 吕便 支派、 迦得 支派、 西布伦 支派中，得了十二座城。
1CHR|6|64|以色列 人把这些城与其郊野给了 利未 人。
1CHR|6|65|以色列 人用抽签的方式，从 犹大 人、 西缅 人、 便雅悯 人三支派中，把以上提到名字的城给了他们。
1CHR|6|66|哥辖 子孙中有几个宗族从 以法莲 支派中也得了城镇作为他们的区域。
1CHR|6|67|他们在 以法莲 山区所得的逃城： 示剑 与其郊野、 基色 与其郊野、
1CHR|6|68|约缅 与其郊野、 伯．和仑 与其郊野、
1CHR|6|69|亚雅仑 与其郊野、 迦特．临门 与其郊野。
1CHR|6|70|哥辖 其余的子孙从 玛拿西 半支派中得了 亚乃 与其郊野、 比连 与其郊野。
1CHR|6|71|革顺 子孙从 玛拿西 半支派中得了 巴珊 的 哥兰 与其郊野、 亚斯她录 与其郊野；
1CHR|6|72|从 以萨迦 支派中得了 基低斯 与其郊野、 大比拉 与其郊野、
1CHR|6|73|拉末 与其郊野、 亚年 与其郊野；
1CHR|6|74|从 亚设 支派中得了 玛沙 与其郊野、 押顿 与其郊野、
1CHR|6|75|户割 与其郊野、 利合 与其郊野；
1CHR|6|76|从 拿弗他利 支派中得了 加利利 的 基低斯 与其郊野、 哈们 与其郊野、 基列亭 与其郊野。
1CHR|6|77|米拉利 其余的子孙从 西布伦 支派中得了 临摩挪 与其郊野、 他泊 与其郊野；
1CHR|6|78|又在 耶利哥 的 约旦河 东，从 吕便 支派中得了旷野的 比悉 与其郊野、 雅杂 与其郊野，
1CHR|6|79|基底莫 与其郊野、 米法押 与其郊野；
1CHR|6|80|又从 迦得 支派中得了 基列 的 拉末 与其郊野、 玛哈念 与其郊野、
1CHR|6|81|希实本 与其郊野、 雅谢 与其郊野。
1CHR|7|1|以萨迦 的后裔： 陀拉 、 普瓦 、 雅述 和 伸仑 ，共四人。
1CHR|7|2|陀拉 的后裔： 乌西 、 利法雅 、 耶勒 、 雅买 、 易伯散 和 示母利 ，都是 陀拉 的族长，在他们世代中是大能的勇士。到 大卫 年间，他们的人数共有二万二千六百名。
1CHR|7|3|乌西 的后裔： 伊斯拉希 ， 伊斯拉希 的儿子 米迦勒 、 俄巴底亚 、 约珥 和 伊示雅 ，共五人，全都是族长。
1CHR|7|4|他们所率领的，按着家谱，照着父家，可作战的军队共有三万六千人，因为他们的妻子和儿子众多。
1CHR|7|5|他们的弟兄在 以萨迦 各族中的大能勇士，登记在家谱中的全部共有八万七千人。
1CHR|7|6|便雅悯 ： 比拉 、 比结 和 耶叠 ，共三人。
1CHR|7|7|比拉 的儿子： 以斯本 、 乌西 、 乌薛 、 耶利末 和 以利 ，共五人，都是族长，是大能的勇士。登记在家谱中的人共有二万二千零三十四人。
1CHR|7|8|比结 的儿子： 细米拉 、 约阿施 、 以利以谢 、 以利约乃 、 暗利 、 耶列末 、 亚比雅 、 亚拿突 和 亚拉篾 ；这些全都是 比结 的儿子。
1CHR|7|9|登记在家谱中，按家谱的族长，大能的勇士，共有二万零二百人。
1CHR|7|10|耶叠 的后裔： 比勒罕 ， 比勒罕 的儿子 耶乌施 、 便雅悯 、 以笏 、 基拿拿 、 细坦 、 他施 和 亚希沙哈 。
1CHR|7|11|这些全都是 耶叠 的后裔，都是族长，是大能的勇士，能上阵打仗的共有一万七千二百人。
1CHR|7|12|还有 以珥 的儿子 书品 和 户品 ，以及 亚黑 的儿子 户伸 。
1CHR|7|13|拿弗他利 的后裔： 雅薛 、 沽尼 、 耶色 和 沙龙 ，都是 辟拉 的子孙。
1CHR|7|14|玛拿西 的儿子 亚斯烈 是他的妾 亚兰 女子所生的；她又生了 玛吉 ，是 基列 的父亲。
1CHR|7|15|玛吉 为 户品 和 书品 各娶了一妻，他的姊妹名叫 玛迦 。第二个名叫 西罗非哈 ； 西罗非哈 只有女儿。
1CHR|7|16|玛吉 的妻子 玛迦 生了一个儿子， 玛迦 给他起名叫 毗利施 。 毗利施 的弟弟名叫 示利施 ； 示利施 的儿子是 乌兰 和 利金 。
1CHR|7|17|乌兰 的儿子是 比但 。这些都是 基列 的子孙； 基列 是 玛吉 的儿子， 玛吉 是 玛拿西 的儿子。
1CHR|7|18|基列 的妹妹 哈摩利吉 生了 伊施荷 、 亚比以谢 和 玛拉 。
1CHR|7|19|示米大 的儿子是 亚现 、 示剑 、 利克希 和 阿尼安 。
1CHR|7|20|以法莲 的后裔： 书提拉 ，他的儿子 比列 ，他的儿子 他哈 ，他的儿子 以拉大 ，他的儿子 他哈 ，
1CHR|7|21|他的儿子 撒拔 ，他的儿子 书提拉 。 以法莲 又生 以谢 和 以列 ；这二人因为下去夺取 迦特 人的牲畜，被本地的 迦特 人杀了。
1CHR|7|22|他们的父亲 以法莲 为他们悲哀了多日，他的兄弟都来安慰他。
1CHR|7|23|以法莲 与妻子同房，妻子怀孕生了一子， 以法莲 因为家里遭祸，就给这儿子起名叫 比利亚 。
1CHR|7|24|他的女儿名叫 舍伊拉 ， 舍伊拉 建筑了 上伯．和仑 、 下伯．和仑 和 乌羡．舍伊拉 。
1CHR|7|25|他的儿子 利法 和 利悉 ，他的儿子 他拉 ，他的儿子 他罕 ，
1CHR|7|26|他的儿子 拉但 ，他的儿子 亚米忽 ，他的儿子 以利沙玛 ，
1CHR|7|27|他的儿子 嫩 ，他的儿子 约书亚 。
1CHR|7|28|以法莲 人的地业和住处是 伯特利 和所属的乡镇，东边 拿兰 ，西边 基色 和所属的乡镇， 示剑 和所属的乡镇，直到 艾雅 和所属的乡镇；
1CHR|7|29|还有靠近 玛拿西 人的边界， 伯．善 和所属的乡镇， 他纳 和所属的乡镇， 米吉多 和所属的乡镇， 多珥 和所属的乡镇。 以色列 儿子 约瑟 的子孙住在这些地方。
1CHR|7|30|亚设 的后裔： 音拿 、 亦施瓦 、 亦施韦 和 比利亚 ，还有他们的妹妹 西拉 。
1CHR|7|31|比利亚 的儿子是 希别 和 玛结 ； 玛结 是 比撒威 的父亲。
1CHR|7|32|希别 生 雅弗勒 、 朔默 、 何坦 和他们的妹妹 书雅 。
1CHR|7|33|雅弗勒 的儿子是 巴萨 、 宾哈 和 亚施法 ；这些都是 雅弗勒 的儿子。
1CHR|7|34|朔默 的儿子是 亚希 、 罗迦 、 耶户巴 和 亚兰 。
1CHR|7|35|朔默 的兄弟 希连 的儿子是 琐法 、 音那 、 示利斯 和 亚抹 。
1CHR|7|36|琐法 的儿子是 书亚 、 哈尼弗 、 书阿勒 、 比利 、 音拉 、
1CHR|7|37|比悉 、 河得 、 珊玛 、 施沙 、 益兰 和 比拉 。
1CHR|7|38|益帖 的儿子是 耶孚尼 、 毗斯巴 和 亚拉 。
1CHR|7|39|乌拉 的儿子是 亚拉 、 汉尼业 和 利写 。
1CHR|7|40|这些全都是 亚设 的子孙，都是族长，是精壮大能的勇士，也是领袖中的领袖。登记在家谱中，能上阵打仗的共有二万六千人。
1CHR|8|1|便雅悯 生长子 比拉 ，次子 亚实别 ，三子 亚哈拉 ，
1CHR|8|2|四子 挪哈 ，五子 拉法 。
1CHR|8|3|比拉 的儿子是 亚大 、 基拉 、 亚比忽 、
1CHR|8|4|亚比书 、 乃幔 、 亚何亚 、
1CHR|8|5|基拉 、 示孚汛 和 户兰 。
1CHR|8|6|以忽 的后裔如下，他们是 迦巴 居民的族长，曾被掳到 玛拿辖 ：
1CHR|8|7|乃幔 、 亚希亚 、 基拉 ；他掳了他们，又生了 乌撒 和 亚希忽 。
1CHR|8|8|沙哈连 休了两个妻子 户伸 和 巴拉 之后，在 摩押 地生了儿子。
1CHR|8|9|他与妻子 贺得 生了 约巴 、 洗比雅 、 米沙 、 玛拉干 、
1CHR|8|10|耶乌斯 、 沙迦 和 米玛 ；这些是他的儿子，都是族长。
1CHR|8|11|户伸 为他生了 亚比突 和 以利巴力 。
1CHR|8|12|以利巴力 的儿子是 希伯 、 米珊 和 沙麦 ； 沙麦 建立 阿挪 、 罗德 和所属的乡镇。
1CHR|8|13|比利亚 和 示玛 是 亚雅仑 居民的族长，他们驱逐了 迦特 的居民。
1CHR|8|14|亚希约 、 沙煞 、 耶列末 、
1CHR|8|15|西巴第雅 、 亚拉得 、 亚得 、
1CHR|8|16|米迦勒 、 伊施巴 和 约哈 都是 比利亚 的儿子。
1CHR|8|17|西巴第雅 、 米书兰 、 希西基 、 希伯 、
1CHR|8|18|伊施米莱 、 伊斯利亚 和 约巴 都是 以利巴力 的儿子。
1CHR|8|19|雅金 、 细基利 、 撒底 、
1CHR|8|20|以利乃 、 洗勒太 、 以利业 、
1CHR|8|21|亚大雅 、 比拉雅 和 申拉 都是 示每 的儿子。
1CHR|8|22|伊施班 、 希伯 、 以利业 、
1CHR|8|23|亚伯顿 、 细基利 、 哈难 、
1CHR|8|24|哈拿尼雅 、 以拦 、 安陀提雅 、
1CHR|8|25|伊弗底雅 、 毗努伊勒 都是 沙煞 的儿子。
1CHR|8|26|珊示莱 、 示哈利 、 亚他利雅 、
1CHR|8|27|雅利西 、 以利亚 和 细基利 都是 耶罗罕 的儿子。
1CHR|8|28|这些人按照他们的家谱都是族长，是领袖，都住在 耶路撒冷 。
1CHR|8|29|在 基遍 住的有 基遍 的父亲 耶利 ，他的妻子名叫 玛迦 ；
1CHR|8|30|他的长子是 亚伯顿 ，还有 苏珥 、 基士 、 巴力 、 拿答 、
1CHR|8|31|基多 、 亚希约 和 撒迦 。
1CHR|8|32|米基罗 生 示米暗 。这些人在他们弟兄的对面，和他们的弟兄同住在 耶路撒冷 。
1CHR|8|33|尼珥 生 基士 ； 基士 生 扫罗 ； 扫罗 生 约拿单 、 麦基．舒亚 、 亚比拿达 和 伊施巴力 。
1CHR|8|34|约拿单 的儿子是 米力．巴力 ； 米力．巴力 生 米迦 。
1CHR|8|35|米迦 的儿子是 毗敦 、 米勒 、 他利亚 和 亚哈斯 ；
1CHR|8|36|亚哈斯 生 耶何阿达 ； 耶何阿达 生 亚拉篾 、 亚斯玛威 和 心利 ； 心利 生 摩撒 ；
1CHR|8|37|摩撒 生 比尼亚 ； 比尼亚 的儿子是 拉法 ， 拉法 的儿子是 以利亚萨 ， 以利亚萨 的儿子是 亚悉 。
1CHR|8|38|亚悉 有六个儿子，他们的名字是 亚斯利干 、 波基路 、 以实玛利 、 示亚利雅 、 俄巴底雅 和 哈难 ；这些全都是 亚悉 的儿子。
1CHR|8|39|亚悉 兄弟 以设 的儿子：长子是 乌兰 ，次子是 耶乌施 ，三子是 以利法列 。
1CHR|8|40|乌兰 的儿子都是大能的勇士，是弓箭手，他们有许多的子孙，共一百五十名，都是 便雅悯 人。
1CHR|9|1|以色列 众人按家谱登记，看哪，都写在《以色列诸王记》上。 犹大 人因背叛被掳到 巴比伦 。
1CHR|9|2|从 巴比伦 先回来，住在自己地业城镇中的有 以色列 人、祭司、 利未 人和殿役。
1CHR|9|3|住在 耶路撒冷 的有 犹大 人、 便雅悯 人、 以法莲 人和 玛拿西 人：
1CHR|9|4|犹大 儿子 法勒斯 的子孙中有 乌太 ， 乌太 是 亚米忽 的儿子， 亚米忽 是 暗利 的儿子， 暗利 是 音利 的儿子， 音利 是 巴尼 的儿子；
1CHR|9|5|示罗 人中有长子 亚帅雅 和他的众儿子；
1CHR|9|6|谢拉 的子孙中有 耶乌利 和他的弟兄，共六百九十人；
1CHR|9|7|便雅悯 人中有 哈西努亚 的曾孙， 何达威雅 的孙子， 米书兰 的儿子 撒路 ；
1CHR|9|8|又有 耶罗罕 的儿子 伊比内雅 ； 米基立 的孙子， 乌西 的儿子 以拉 ； 伊比尼雅 的曾孙， 流珥 的孙子， 示法提雅 的儿子 米书兰 ；
1CHR|9|9|和他们的弟兄，按着家谱登记，共有九百五十六名；这些人都是族长。
1CHR|9|10|祭司中有 耶大雅 、 耶何雅立 、 雅斤 ，
1CHR|9|11|还有管理上帝殿的 亚撒利雅 ， 亚撒利雅 是 希勒家 的儿子， 希勒家 是 米书兰 的儿子， 米书兰 是 撒督 的儿子， 撒督 是 米拉约 的儿子， 米拉约 是 亚希突 的儿子。
1CHR|9|12|还有 玛基雅 的曾孙， 巴施户珥 的孙子， 耶罗罕 的儿子 亚大雅 ；又有 玛赛 ， 玛赛 是 亚第业 的儿子， 亚第业 是 雅希细拉 的儿子， 雅希细拉 是 米书兰 的儿子， 米书兰 是 米实利密 的儿子， 米实利密 是 音麦 的儿子。
1CHR|9|13|他们和他们的弟兄都是族长，共有一千七百六十人，都善于做上帝殿的事工。
1CHR|9|14|利未 人 米拉利 的子孙中有 哈沙比雅 的曾孙， 押利甘 的孙子， 哈述 的儿子 示玛雅 ；
1CHR|9|15|有 拔巴甲 、 黑勒施 、 加拉 和 亚萨 的曾孙， 细基利 的孙子， 米迦 的儿子 玛探雅 ；
1CHR|9|16|又有 耶杜顿 的曾孙， 加拉 的孙子， 示玛雅 的儿子 俄巴底 ，还有 以利加拿 的孙子， 亚撒 的儿子 比利家 。他们都住在 尼陀法 人的村庄。
1CHR|9|17|守卫是 沙龙 、 亚谷 、 达们 、 亚希幔 和他们的弟兄； 沙龙 是领袖。
1CHR|9|18|从前这些人看守朝东的王门，如今是 利未 人营中的守卫。
1CHR|9|19|可拉 的曾孙， 以比雅撒 的孙子， 可利 的儿子 沙龙 ，和他父家的弟兄 可拉 人管理事务，看守会幕的门。他们的祖宗曾管理耶和华的军营，把守营的入口。
1CHR|9|20|从前 以利亚撒 的儿子 非尼哈 管理他们，耶和华也与他同在。
1CHR|9|21|米施利米雅 的儿子 撒迦利雅 是看守会幕门口的。
1CHR|9|22|被选作门口守卫的总共有二百一十二名。他们在自己的村庄，按着家谱登记，是 大卫 和 撒母耳 先见所派担当这受托之职任的。
1CHR|9|23|他们和他们的子孙看守耶和华殿的门，就是会幕的门口。
1CHR|9|24|在东西南北，四方 都有守卫。
1CHR|9|25|他们的弟兄住在村庄，每七日来与他们换班。
1CHR|9|26|这些守卫的四个领袖都是 利未 人，各有受托的职任，看守上帝殿的房间和宝库。
1CHR|9|27|他们住在上帝殿的四围，受托看守圣殿，负责每日早晨开门。
1CHR|9|28|利未 人中有人管理所使用的器皿，拿出拿入都按数目点算。
1CHR|9|29|又有人管理器具和圣所一切的器皿，以及细面、酒、油、乳香和香料。
1CHR|9|30|祭司的子孙中有人用香料做膏油。
1CHR|9|31|利未 人 玛他提雅 是 可拉 族 沙龙 的长子，他受托做烤饼。
1CHR|9|32|他们弟兄 哥辖 子孙中，有人负责每安息日排列供饼。
1CHR|9|33|歌唱的有 利未 人的族长，住在殿的房间，昼夜供职，不做别样的工。
1CHR|9|34|以上都是 利未 人的族长，按各世系作领袖，他们都住在 耶路撒冷 。
1CHR|9|35|在 基遍 住的有 基遍 的父亲 耶利 ，他的妻子名叫 玛迦 ；
1CHR|9|36|他的长子是 亚伯顿 ，还有 苏珥 、 基士 、 巴力 、 尼珥 、 拿答 、
1CHR|9|37|基多 、 亚希约 、 撒迦利雅 和 米基罗 。
1CHR|9|38|米基罗 生 示米暗 。这些人在他们弟兄的对面，和他们的弟兄同住在 耶路撒冷 。
1CHR|9|39|尼珥 生 基士 ； 基士 生 扫罗 ； 扫罗 生 约拿单 、 麦基．舒亚 、 亚比拿达 和 伊施巴力 。
1CHR|9|40|约拿单 的儿子是 米力．巴力 ； 米力．巴力 生 米迦 。
1CHR|9|41|米迦 的儿子是 毗敦 、 米勒 、 他利亚 和 亚哈斯 。
1CHR|9|42|亚哈斯 生 雅拉 ； 雅拉 生 亚拉篾 、 亚斯玛威 和 心利 ； 心利 生 摩撒 ；
1CHR|9|43|摩撒 生 比尼亚 ； 比尼亚 的儿子是 利法雅 ， 利法雅 的儿子是 以利亚萨 ， 以利亚萨 的儿子是 亚悉 。
1CHR|9|44|亚悉 有六个儿子，他们的名字是 亚斯利干 、 波基路 、 以实玛利 、 示亚利雅 、 俄巴底雅 和 哈难 ；这些都是 亚悉 的儿子。
1CHR|10|1|非利士 人攻打 以色列 。 以色列 人在 非利士 人面前逃跑，很多人 在 基利波山 被杀仆倒。
1CHR|10|2|非利士 人紧追 扫罗 和他的儿子，杀了 扫罗 的儿子 约拿单 、 亚比拿达 、 麦基．舒亚 。
1CHR|10|3|攻击 扫罗 的战事激烈， 扫罗 被弓箭手射中，被他们射伤。
1CHR|10|4|扫罗 吩咐拿他兵器的人说：“你拔出刀来，把我刺死，免得那些未受割礼的人来凌辱我。”但拿兵器的人非常惧怕，不肯刺他。于是 扫罗 拿起刀来，伏在刀上。
1CHR|10|5|拿兵器的人见 扫罗 已死，也伏在刀上死了。
1CHR|10|6|这样， 扫罗 和他三个儿子，以及他的全家都一起阵亡了。
1CHR|10|7|住平原的 以色列 众人见 以色列 军兵 逃跑， 扫罗 和他儿子都死了，就弃城逃跑。 非利士 人前来，占据了他们的城。
1CHR|10|8|次日， 非利士 人来剥那些被杀之人的衣服，看见 扫罗 和他儿子仆倒在 基利波山 。
1CHR|10|9|他们剥了他的军装，拿着他的首级和盔甲，派人到 非利士 人之地的四境，报信给他们的偶像和百姓。
1CHR|10|10|他们将 扫罗 的盔甲放在他们神明的庙里，把他的首级钉在 大衮 庙中。
1CHR|10|11|基列 的 雅比 居民听见 非利士 人向 扫罗 所行的一切事，
1CHR|10|12|他们中间所有的勇士就起身，把 扫罗 和他儿子的尸身送到 雅比 ，把他们的尸骨葬在 雅比 的橡树下，禁食七日。
1CHR|10|13|这样， 扫罗 为了他的不忠死了；因为他干犯耶和华，没有遵守耶和华的话，又因他求问招魂的妇人，
1CHR|10|14|不求问耶和华，所以耶和华使他被杀，把王国给了 耶西 的儿子 大卫 。
1CHR|11|1|以色列 众人聚集到 希伯仑 见 大卫 ，说：“看哪，我们是你的骨肉。
1CHR|11|2|从前 扫罗 作王的时候，率领 以色列 人出入的是你；耶和华－你的上帝也曾对你说：‘你必牧养我的百姓 以色列 ，你必作我百姓 以色列 的君王。’”
1CHR|11|3|于是 以色列 的众长老都来到 希伯仑 见王。 大卫 在 希伯仑 ，在耶和华面前与他们立约，他们就膏 大卫 作 以色列 的王，正如耶和华藉 撒母耳 所说的话。
1CHR|11|4|大卫 和 以色列 众人到了 耶路撒冷 ，就是 耶布斯 ；那时 耶布斯 人住在那里。
1CHR|11|5|耶布斯 人对 大卫 说：“你必不能进到这里。”然而 大卫 攻取了 锡安 的堡垒，就是 大卫 的城。
1CHR|11|6|大卫 说：“谁先攻打 耶布斯 人，必作领袖，作元帅。” 洗鲁雅 的儿子 约押 先上去，就作了领袖。
1CHR|11|7|大卫 住在堡垒里，所以那堡垒叫作 大卫城 。
1CHR|11|8|大卫 又从 米罗 起，四围建筑城墙，其余的由 约押 修建。
1CHR|11|9|大卫 日见强大，万军之耶和华与他同在。
1CHR|11|10|以下是跟随 大卫 勇士的领袖；他们奋勇帮助他得到国度，并照着耶和华吩咐 以色列 的话，与 以色列 众人一同立他作王。
1CHR|11|11|大卫 勇士的名单如下： 哈革摩尼 的儿子 雅朔班 ，他是军官的统领 ，曾一次举枪杀了三百人。
1CHR|11|12|其次是 亚何亚 人 朵多 的儿子 以利亚撒 ，他是三个勇士里的一个。
1CHR|11|13|他从前与 大卫 在 巴斯．大悯 ， 非利士 人聚集要打仗。那里有一块长满大麦的田。百姓在 非利士 人面前逃跑，
1CHR|11|14|他们 却站在那块田的中间，防守那田，击败了 非利士 人。耶和华大获全胜。
1CHR|11|15|三十个领袖中的三个人下到磐石那里，进了 亚杜兰洞 见 大卫 ； 非利士 的军队在 利乏音谷 安营。
1CHR|11|16|那时 大卫 在山寨， 非利士 人的驻军在 伯利恒 。
1CHR|11|17|大卫 渴想着说：“但愿有人从 伯利恒 城门旁的井里打水来给我喝！”
1CHR|11|18|这三个勇士就闯过 非利士 人的军营，从 伯利恒 城门旁的井里打水，拿来给 大卫 喝。 大卫 却不肯喝，将水浇在耶和华面前，
1CHR|11|19|说：“我的上帝啊，我绝不做这事！这些人冒死去打水，这水是他们用生命换来的，我怎能喝他们的血呢？” 大卫 不肯喝这水。这是三个勇士所做的事。
1CHR|11|20|约押 的兄弟 亚比筛 是这三个 勇士的领袖；他曾举枪杀了三百人，就在三个勇士中得了名。
1CHR|11|21|他在这三个勇士里比其他两个更有名望，所以作他们的领袖，只是不及前三个勇士。
1CHR|11|22|耶何耶大 的儿子 比拿雅 是来自 甲薛 的勇士，曾行了大事。他杀了 摩押 人 亚利伊勒 的两个儿子，又在下雪的时候下到坑里去，杀了一只狮子。
1CHR|11|23|他又杀了一个身高五肘的 埃及 人； 埃及 人手里拿着枪，枪杆粗如织布机的轴。 比拿雅 只拿着棍子下到他那里去，从 埃及 人手里夺过枪来，用那枪杀死了他。
1CHR|11|24|这些是 耶何耶大 的儿子 比拿雅 所做的事，就在三个勇士里得了名。
1CHR|11|25|看哪，他比那三十个勇士更有名望，只是不及前三个勇士。 大卫 立他作护卫长。
1CHR|11|26|军中的勇士有 约押 的兄弟 亚撒黑 ， 伯利恒 人 朵多 的儿子 伊勒哈难 ，
1CHR|11|27|哈律 人 沙玛 ， 比伦 人 希利斯 ，
1CHR|11|28|提哥亚 人 益吉 的儿子 以拉 ， 亚拿突 人 亚比以谢 ，
1CHR|11|29|户沙 人 西比该 ， 亚何亚 人 以来 ，
1CHR|11|30|尼陀法 人 玛哈莱 ， 尼陀法 人 巴拿 的儿子 希立 ，
1CHR|11|31|便雅悯 族 基比亚 人 利拜 的儿子 以太 ， 比拉顿 人 比拿雅 ，
1CHR|11|32|迦实溪 人 户莱 ， 亚拉巴 人 亚比 ，
1CHR|11|33|巴路米 人 押斯玛弗 ， 沙本 人 以利雅哈巴 ，
1CHR|11|34|基孙 人 哈深 的众儿子， 哈拉 人 沙基 的儿子 约拿单 ，
1CHR|11|35|哈拉 人 沙甲 的儿子 亚希暗 ， 吾珥 的儿子 以利法勒 ，
1CHR|11|36|米基拉 人 希弗 ， 比伦 人 亚希雅 ，
1CHR|11|37|迦密 人 希斯罗 ， 伊斯拜 的儿子 拿莱 ，
1CHR|11|38|拿单 的兄弟 约珥 ， 哈基利 的儿子 弥伯哈 ，
1CHR|11|39|亚扪 人 洗勒 ， 比录 人 拿哈莱 ，他是给 洗鲁雅 的儿子 约押 拿兵器的，
1CHR|11|40|以帖 人 以拉 ， 以帖 人 迦立 ，
1CHR|11|41|赫 人 乌利亚 ， 亚莱 的儿子 撒拔 ，
1CHR|11|42|吕便 人 示撒 的儿子 亚第拿 ，是 吕便 支派中的一个领袖，率领三十人，
1CHR|11|43|玛迦 的儿子 哈难 ， 弥特尼 人 约沙法 ，
1CHR|11|44|亚施他拉 人 乌西亚 ， 亚罗珥 人 何坦 的儿子 沙玛 和 耶利 ，
1CHR|11|45|提洗 人 申利 的儿子 耶叠 和他的兄弟 约哈 ，
1CHR|11|46|玛哈未 人 以利业 ， 伊利拿安 的儿子 耶利拜 和 约沙未雅 ， 摩押 人 伊特玛 、
1CHR|11|47|以利业 、 俄备得 ，以及 米琐八 人 雅西业 。
1CHR|12|1|以下是 大卫 因 基士 的儿子 扫罗 的缘故被放逐到 洗革拉 的时候，到他那里帮助他打仗的勇士；
1CHR|12|2|他们是弓箭手，能左右甩石，开弓射箭，都是 便雅悯 人 扫罗 同族的弟兄：
1CHR|12|3|为首的是 亚希以谢 ，其次是 约阿施 ，都是 基比亚 人 示玛 的儿子。还有 亚斯玛威 的儿子 耶薛 和 毗力 ， 比拉迦 ， 亚拿突 人 耶户 ，
1CHR|12|4|基遍 人 以实买雅 ，他在三十人中是勇士，管理这三十人，又有 耶利米 ， 雅哈悉 ， 约哈难 ， 基底拉 人 约撒拔 ，
1CHR|12|5|伊利乌赛 ， 耶利末 ， 比亚利雅 ， 示玛利雅 ， 哈律弗 人 示法提雅 ，
1CHR|12|6|可拉 人 以利加拿 、 耶西亚 、 亚萨列 、 约以谢 、 雅朔班 ，
1CHR|12|7|基多 人 耶罗罕 的儿子 犹拉 和 西巴第雅 。
1CHR|12|8|迦得 人中有人到旷野的山寨投奔 大卫 ，都是大能的勇士，能拿盾牌和枪的战士。他们的面貌好像狮子，敏捷如山上的鹿。
1CHR|12|9|第一 以薛 ，第二 俄巴底雅 ，第三 以利押 ，
1CHR|12|10|第四 弥施玛拿 ，第五 耶利米 ，
1CHR|12|11|第六 亚太 ，第七 以利业 ，
1CHR|12|12|第八 约哈难 ，第九 以利萨巴 ，
1CHR|12|13|第十 耶利米 ，第十一 末巴奈 。
1CHR|12|14|这些都是 迦得 人中的军官，小的能抵一百人，大的能抵一千人 。
1CHR|12|15|正月， 约旦河 水涨过两岸的时候，他们过河，使所有住河谷的人东奔西逃。
1CHR|12|16|便雅悯 人和 犹大 人中有人来到山寨 大卫 那里。
1CHR|12|17|大卫 出去迎接他们，回答他们说：“你们若和平地来帮助我，我的心就与你们契合；但你们若把我这双手无辜的人卖给敌人，愿我们列祖的上帝察看责罚。”
1CHR|12|18|那时军官 的领袖 亚玛撒 受灵的感动说： “ 大卫 啊，我们归向你！ 耶西 的儿子啊，我们帮助你！ 愿你平平安安， 愿帮助你的也都平安！ 因为你的上帝帮助你。” 大卫 就收留他们，派他们作军官。
1CHR|12|19|大卫 从前与 非利士 人同去，要与 扫罗 争战，有些 玛拿西 人来投奔 大卫 。其实他们并没有帮助 非利士 人，因为 非利士 人的领袖商议，打发他回去，说：“恐怕 大卫 拿我们的首级去向他的主人 扫罗 投诚。”
1CHR|12|20|大卫 往 洗革拉 去的时候，有 玛拿西 人的千夫长 押拿 、 约撒拔 、 耶叠 、 米迦勒 、 约撒拔 、 以利户 、 洗勒太 都来投奔他。
1CHR|12|21|他们帮助 大卫 攻击敌军；因为他们都是大能的勇士，又作军官。
1CHR|12|22|那时天天有人来帮助 大卫 ，以致成了强大的军队，如上帝的军队一样。
1CHR|12|23|以下是来到 希伯仑 见 大卫 ，要照耶和华的话把 扫罗 的国位归给 大卫 的武装士兵的数目：
1CHR|12|24|犹大 人，拿盾牌和枪的武装战士有六千八百人。
1CHR|12|25|西缅 人中，能上阵的大能勇士有七千一百人。
1CHR|12|26|利未 人中，有四千六百人。
1CHR|12|27|耶何耶大 是 亚伦 家的领袖，跟从他的有三千七百人。
1CHR|12|28|还有大能的青年勇士 撒督 ，同他本族的二十二个军官。
1CHR|12|29|便雅悯 人中， 扫罗 同族的弟兄也有三千人；直到现在他们大部分仍然效忠 扫罗 家。
1CHR|12|30|以法莲 人中，在本族中著名的大能勇士有二万零八百人。
1CHR|12|31|玛拿西 半支派，册上有名来拥立 大卫 作王的，有一万八千人。
1CHR|12|32|以萨迦 人中，通达时务，知道 以色列 所当行，同族弟兄也都听从他们命令的族长有二百人。
1CHR|12|33|西布伦 中，能上阵用各样作战的兵器、不生二心帮助打仗的有五万人。
1CHR|12|34|拿弗他利 中，有一千个军官；跟从他们、拿盾牌和枪的有三万七千人。
1CHR|12|35|但 人中，能摆阵的有二万八千六百人。
1CHR|12|36|亚设 中，能上阵打仗的有四万人。
1CHR|12|37|约旦河 东的 吕便 人、 迦得 人、 玛拿西 半支派，拿各样兵器打仗的有十二万人。
1CHR|12|38|以上都是能列队上阵的战士，他们都全心来到 希伯仑 ，要拥立 大卫 作全 以色列 的王。 以色列 其余的人也都一心要拥立 大卫 作王。
1CHR|12|39|他们在那里三日，与 大卫 一同吃喝，因为他们同族的弟兄已经为他们预备好了。
1CHR|12|40|他们附近的人，以及 以萨迦 、 西布伦 、 拿弗他利 人，都将食物，许多面饼、无花果饼、干葡萄、酒、油，用驴、骆驼、骡子、牛驮来，又带了许多的牛和羊来，因为在 以色列 中充满了欢乐。
1CHR|13|1|大卫 与千夫长、百夫长，以及所有的领袖商议。
1CHR|13|2|大卫 对 以色列 全会众说：“你们若以为好，见这事是出于耶和华－我们的上帝，我们就派人到远近各处去见仍留在 以色列 各地我们的弟兄，以及住在有郊野之城的祭司和 利未 人，使他们都到我们这里来聚集。
1CHR|13|3|我们要把上帝的约柜接到这里来；因为在 扫罗 年间，我们没有去寻求约柜 。”
1CHR|13|4|全会众都说可以这么做，因这事在众百姓眼中都看为好。
1CHR|13|5|于是， 大卫 把 以色列 众人从 埃及 的 西曷河 直到 哈马口 都召集了来，要从 基列．耶琳 将上帝的约柜接来。
1CHR|13|6|大卫 率领 以色列 众人上到 巴拉 ，就是属 犹大 的 基列．耶琳 ，要将耶和华上帝的约柜从那里接上来，他坐在二基路伯之上，这约柜是以他的名来命名的。
1CHR|13|7|他们将上帝的约柜从 亚比拿达 的家里抬出来，放在新车上，由 乌撒 和 亚希约 赶车。
1CHR|13|8|大卫 和 以色列 众人在上帝面前随着诗歌、琴、瑟、鼓、钹、号，极力跳舞。
1CHR|13|9|到了 基顿 的禾场，因为牛失前蹄 ， 乌撒 就伸手扶住约柜。
1CHR|13|10|耶和华的怒气向 乌撒 发作，因他伸手扶住约柜而击杀他，他就死在那里，在上帝面前。
1CHR|13|11|大卫 因耶和华突然冲出撞死 乌撒 就生气，称那地方为 毗列斯．乌撒 ，直到今日。
1CHR|13|12|那日， 大卫 惧怕上帝，说：“我怎能将上帝的约柜接到我这里来呢？”
1CHR|13|13|于是 大卫 不将约柜接进 大卫城 他自己的地方，却转送到 迦特 人 俄别．以东 的家中。
1CHR|13|14|上帝的约柜停在 俄别．以东 家中三个月，耶和华赐福给 俄别．以东 的家和他一切所有的。
1CHR|14|1|推罗 王 希兰 派使者把香柏木运到 大卫 那里，又派石匠和木匠给 大卫 建造宫殿。
1CHR|14|2|大卫 知道耶和华坚立他作 以色列 王，又为自己百姓 以色列 的缘故，使他的国兴盛。
1CHR|14|3|大卫 在 耶路撒冷 又立后妃，又生儿女。
1CHR|14|4|在 耶路撒冷 所生的孩子名字是 沙母亚 、 朔罢 、 拿单 、 所罗门 、
1CHR|14|5|益辖 、 以利书亚 、 以法列 、
1CHR|14|6|挪迦 、 尼斐 、 雅非亚 、
1CHR|14|7|以利沙玛 、 比利雅大 、 以利法列 。
1CHR|14|8|非利士 人听见 大卫 受膏作全 以色列 的王， 非利士 众人就上来寻索 大卫 。 大卫 听见了，就出去迎敌。
1CHR|14|9|非利士 人来了，侵犯 利乏音谷 。
1CHR|14|10|大卫 求问上帝说：“我可以上去攻打 非利士 人吗？你将他们交在我手里吗？”耶和华对他说：“你可以上去，我必将他们交在你手里。”
1CHR|14|11|非利士 人上到 巴力．毗拉心 ， 大卫 在那里击败他们。 大卫 说：“上帝藉我的手冲破敌人，如水冲破一样。”因此那地方称为 巴力．毗拉心 。
1CHR|14|12|非利士 人把神像抛弃在那里， 大卫 吩咐人用火焚烧了。
1CHR|14|13|非利士 人又侵犯 利乏音谷 。
1CHR|14|14|大卫 再求问上帝。上帝对他说：“不要从他们后头追上去，要绕道离开他们，从桑树林对面攻打他们。
1CHR|14|15|你听见桑树梢上有脚步的声音，那时你就要出战，因为上帝已经出去，在你前头攻打 非利士 人的军队了。”
1CHR|14|16|大卫 就遵照上帝所吩咐的去做，攻打 非利士 人的军队，从 基遍 直到 基色 。
1CHR|14|17|于是 大卫 的名传扬到万邦，耶和华使万国都惧怕他。
1CHR|15|1|大卫 在 大卫城 为自己建造宫殿，又为上帝的约柜预备地方，支搭帐幕。
1CHR|15|2|那时 大卫 说：“除了 利未 人之外，无人可抬上帝的约柜，因为耶和华拣选他们抬上帝的约柜，永远事奉他。”
1CHR|15|3|大卫 召集 以色列 众人到 耶路撒冷 ，要将耶和华的约柜接到他所预备的地方。
1CHR|15|4|大卫 又召集 亚伦 的子孙和 利未 人：
1CHR|15|5|哥辖 子孙中有领袖 乌列 和他的弟兄一百二十人，
1CHR|15|6|米拉利 子孙中有领袖 亚帅雅 和他的弟兄二百二十人，
1CHR|15|7|革顺 子孙中有领袖 约珥 和他的弟兄一百三十人，
1CHR|15|8|以利撒反 子孙中有领袖 示玛雅 和他的弟兄二百人，
1CHR|15|9|希伯伦 子孙中有领袖 以利业 和他的弟兄八十人，
1CHR|15|10|乌薛 子孙中有领袖 亚米拿达 和他的弟兄一百一十二人。
1CHR|15|11|大卫 召来 撒督 和 亚比亚他 二位祭司，以及 利未 人 乌列 、 亚帅雅 、 约珥 、 示玛雅 、 以利业 、 亚米拿达 ，
1CHR|15|12|对他们说：“你们是 利未 人的族长，你们和你们的弟兄应当使自己分别为圣，好将耶和华－ 以色列 上帝的约柜接到我所预备的地方。
1CHR|15|13|因为你们上一次没有抬这约柜，并且我们没有按规矩求问耶和华－我们的上帝，所以他冲出来攻击我们。”
1CHR|15|14|于是祭司和 利未 人使自己分别为圣，将耶和华－ 以色列 上帝的约柜接上来。
1CHR|15|15|利未 子孙用杠，把上帝的约柜抬在肩上，正如 摩西 按照耶和华的话所吩咐的。
1CHR|15|16|大卫 吩咐 利未 人的领袖派他们歌唱的弟兄用琴瑟和钹的乐器奏乐，欢欢喜喜地大声歌颂。
1CHR|15|17|于是 利未 人派 约珥 的儿子 希幔 和他弟兄中 比利家 的儿子 亚萨 ，以及他们同族弟兄 米拉利 子孙里 古沙雅 的儿子 以探 。
1CHR|15|18|其次还有跟随他们的弟兄 撒迦利雅 、 便．雅薛 、 示米拉末 、 耶歇 、 乌尼 、 以利押 、 比拿雅 、 玛西雅 、 玛他提雅 、 以利斐利户 、 弥克尼雅 ，以及门口的守卫 俄别．以东 和 耶利 。
1CHR|15|19|歌唱的 希幔 、 亚萨 和 以探 ，敲铜钹，声音响亮；
1CHR|15|20|撒迦利雅 、 雅薛 、 示米拉末 、 耶歇 、 乌尼 、 以利押 、 玛西雅 、 比拿雅 鼓瑟，调用女音；
1CHR|15|21|玛他提雅 、 以利斐利户 、 弥克尼雅 、 俄别．以东 、 耶利 、 亚撒西雅 用琴指挥，调用第八。
1CHR|15|22|基拿尼雅 是 利未 人圣咏团的领袖，又教导人唱歌，因为他精通此事。
1CHR|15|23|比利家 和 以利加拿 是约柜的守卫。
1CHR|15|24|示巴尼 、 约沙法 、 拿坦业 、 亚玛赛 、 撒迦利雅 、 比拿亚 、 以利以谢 众祭司在上帝的约柜前吹号。 俄别．以东 和 耶希亚 也是约柜的守卫。
1CHR|15|25|于是， 大卫 和 以色列 的长老，以及千夫长都去，欢欢喜喜地将耶和华的约柜从 俄别．以东 家中接上来。
1CHR|15|26|上帝赐恩给抬耶和华约柜的 利未 人，他们就献上七头公牛，七只公羊。
1CHR|15|27|大卫 和所有抬约柜的 利未 人，以及圣咏团的领袖 基拿尼雅 和歌唱的人，都穿着细麻布外袍； 大卫 另外穿着细麻布以弗得。
1CHR|15|28|这样， 以色列 众人欢呼、吹角、吹号、敲钹、鼓瑟、弹琴，声音响亮，将耶和华的约柜接上来。
1CHR|15|29|耶和华的约柜进 大卫城 的时候， 扫罗 的女儿 米甲 从窗户里往外观看，见 大卫 王踊跃跳舞，心里就轻视他。
1CHR|16|1|众人将上帝的约柜请进去，安放在 大卫 为它搭的帐幕中，就在上帝面前献燔祭和平安祭。
1CHR|16|2|大卫 献完了燔祭和平安祭，就奉耶和华的名祝福百姓，
1CHR|16|3|并且分给每一个 以色列 人，无论男女，每人一个饼，一个枣子饼 ，一个葡萄饼。
1CHR|16|4|大卫 派几个 利未 人在耶和华的约柜前事奉，颂扬，称谢，赞美耶和华－ 以色列 的上帝：
1CHR|16|5|为首的是 亚萨 ，其次是 撒迦利雅 、 耶利 、 示米拉末 、 耶歇 、 玛他提雅 、 以利押 、 比拿雅 、 俄别．以东 、 耶利 ；他们鼓瑟弹琴， 亚萨 敲钹，声音响亮；
1CHR|16|6|比拿雅 和 雅哈悉 二位祭司常在上帝的约柜前吹号。
1CHR|16|7|那日， 大卫 初次指派 亚萨 和他的弟兄称谢耶和华。
1CHR|16|8|你们要称谢耶和华，求告他的名， 在万民中传扬他的作为！
1CHR|16|9|要向他唱诗，向他歌颂， 述说他一切奇妙的作为！
1CHR|16|10|要夸耀他的圣名！ 愿寻求耶和华的人心中欢喜！
1CHR|16|11|要寻求耶和华与他的能力， 时常寻求他的面。
1CHR|16|12|他仆人 以色列 的后裔， 他所拣选 雅各 的子孙哪， 要记念他奇妙的作为和他的奇事， 并他口中的判语。
1CHR|16|13|
1CHR|16|14|他是耶和华－我们的上帝， 全地都有他的判断。
1CHR|16|15|要记念他的约，直到永远； 记念他吩咐的话，直到千代，
1CHR|16|16|就是他与 亚伯拉罕 所立的约， 向 以撒 所起的誓。
1CHR|16|17|他将这约向 雅各 定为律例， 向 以色列 定为永远的约，
1CHR|16|18|说：“我必将 迦南 地赐给你， 作你们应得的产业。”
1CHR|16|19|当时，你们人丁有限， 数目稀少，在那地寄居。
1CHR|16|20|他们从这邦游到那邦， 从这国去到另一民族。
1CHR|16|21|他不容人欺负他们， 为他们的缘故责备君王：
1CHR|16|22|“不可伤害我的受膏者， 也不可恶待我的先知。”
1CHR|16|23|全地都要向耶和华歌唱！ 天天传扬他的救恩！
1CHR|16|24|在列国中述说他的荣耀！ 在万民中述说他的奇事！
1CHR|16|25|因耶和华本为大，当受极大的赞美； 他在万神之上，当受敬畏。
1CHR|16|26|因万民的神明都属虚无； 惟独耶和华创造诸天。
1CHR|16|27|有尊荣和威严在他面前， 有能力和喜乐在他自己的地方。
1CHR|16|28|民中的万族啊，要将荣耀、能力归给耶和华， 都归给耶和华！
1CHR|16|29|要将耶和华的名所当得的荣耀归给他， 拿供物来献在他面前； 当敬拜神圣荣耀的耶和华 。
1CHR|16|30|全地都要在他面前战抖！ 世界坚定，不得动摇。
1CHR|16|31|愿天欢喜，愿地快乐！ 愿人在列国中说： “耶和华作王了！”
1CHR|16|32|愿海和其中所充满的澎湃！ 愿田和其中所有的都欢乐！
1CHR|16|33|那时，林中的树木都要在耶和华面前欢呼， 因为他来要审判全地。
1CHR|16|34|你们要称谢耶和华，因他本为善， 他的慈爱永远长存！
1CHR|16|35|你们要说： “拯救我们的上帝啊，求你拯救我们， 聚集我们，救我们脱离列国， 我们好颂扬你的圣名， 以赞美你为夸胜。
1CHR|16|36|耶和华－ 以色列 的上帝是应当称颂的， 从亘古直到永远。” 全体百姓都说：“阿们！”并且赞美耶和华。
1CHR|16|37|大卫 把 亚萨 和他的弟兄留在耶和华的约柜那里，经常在约柜前事奉，天天尽本分供职，
1CHR|16|38|又有 俄别．以东 和他的弟兄六十八人； 耶杜顿 的儿子 俄别．以东 ，以及 何萨 作门口的守卫。
1CHR|16|39|还有 撒督 祭司和他弟兄众祭司在 基遍 的丘坛、耶和华的帐幕前，
1CHR|16|40|在燔祭坛上，每日早晚，照着写在耶和华律法书上所吩咐 以色列 的，经常献燔祭给耶和华。
1CHR|16|41|与他们一同的还有 希幔 、 耶杜顿 ，和其余被选、名字录在册上的，为要称谢耶和华，因他的慈爱永远长存。
1CHR|16|42|希幔 、 耶杜顿 同他们吹号、敲钹，声音响亮，并用其他乐器配合，歌颂上帝。 耶杜顿 的子孙作门口的守卫。
1CHR|16|43|于是众百姓各自回家， 大卫 也回去为家人祝福。
1CHR|17|1|大卫 住在自己宫中，对 拿单 先知说：“看哪，我住在香柏木的宫中，耶和华的约柜却在幔子里。”
1CHR|17|2|拿单 对 大卫 说：“你可以完全照你的心意去做，因为上帝与你同在。”
1CHR|17|3|当夜上帝的话临到 拿单 ，说：
1CHR|17|4|“你去对我仆人 大卫 说：‘耶和华如此说：你不可建造殿宇给我居住。
1CHR|17|5|自从我领 以色列 人上来，直到今日，我未曾住过殿宇；我从这会幕到那会幕，从这帐幕到那帐幕 。
1CHR|17|6|凡我同 以色列 人所走的地方，我何曾向 以色列 的一个士师，就是我吩咐牧养我百姓的，说过这话：你们为何不给我建造香柏木的殿宇呢？’
1CHR|17|7|现在，你要对我仆人 大卫 这样说：‘万军之耶和华如此说：我从羊圈中将你召来，叫你不再牧放羊群，立你作我百姓 以色列 的君王。
1CHR|17|8|你无论往哪里去，我都与你同在，剪除你所有的仇敌。我必使你得大名，好像世上伟人的名一样。
1CHR|17|9|我必为我百姓 以色列 选定一个地方，栽植他们，使他们住自己的地方，不再受搅扰；凶恶之子也不再像从前那样扰乱他们，
1CHR|17|10|并不像我命令士师治理我百姓 以色列 的日子。我必制伏你所有的仇敌，并且我应许你 ，耶和华必为你建立家室。
1CHR|17|11|当你寿数满足归你祖先的时候，我必使你的后裔，你自己的儿子接续你；我也必坚定他的国。
1CHR|17|12|他必为我建造殿宇，我必坚定他的王位，直到永远。
1CHR|17|13|我要作他的父，他要作我的子；我必不使我的慈爱离开他，像离开在你以前的那位一样。
1CHR|17|14|我要永远坚立他在我的家和我的国里；他的王位也必坚定，直到永远。’”
1CHR|17|15|拿单 就按这一切话，照这一切异象告诉 大卫 。
1CHR|17|16|于是 大卫 王进去，坐在耶和华面前，说：“耶和华上帝啊，我是谁，我的家算什么，你竟带领我到这地步呢？
1CHR|17|17|上帝啊，这在你眼中还看为小，你又说到你仆人的家将来的情况。耶和华上帝啊，你看顾我好像看顾尊贵的人。
1CHR|17|18|你加于仆人的尊荣， 大卫 还有什么可以对你说呢？你是知道你仆人的。
1CHR|17|19|耶和华啊，因你仆人的缘故，也照着你的心意，你行这一切大事，为了显明这一切伟大的事。
1CHR|17|20|耶和华啊，照我们耳中一切所听见的，没有可比你的，除你以外再没有上帝。
1CHR|17|21|世上有何国能比你的百姓 以色列 呢？上帝亲自去救赎世上的一国 ，作自己的子民，又行大而可畏的事，显出你的大名，在你从 埃及 赎出来的子民面前驱逐了列国。
1CHR|17|22|你使你的百姓 以色列 作你的子民，直到永远；你－耶和华也作他们的上帝。
1CHR|17|23|现在，耶和华啊，你所应许仆人和仆人家的话，求你坚定，直到永远；求你照你所说的而行。
1CHR|17|24|愿你的名永远坚立，被尊为大，人要说：‘万军之耶和华－ 以色列 的上帝，是 以色列 的上帝。’这样，你仆人 大卫 的家必在你面前坚立。
1CHR|17|25|我的上帝啊，因你启示你的仆人，要为他建立家室，所以仆人大胆在你面前祈祷。
1CHR|17|26|现在，耶和华啊，惟有你是上帝！你应许将这福气赐给仆人。
1CHR|17|27|现在，你喜悦赐福给仆人的家，可以永存在你面前。耶和华啊，因你已经赐福，还要赐福到永远。”
1CHR|18|1|此后， 大卫 攻打 非利士 人，制伏了他们，从 非利士 人手中夺取了 迦特 和所属的乡镇。
1CHR|18|2|他又攻打 摩押 ， 摩押 人就臣服 大卫 ，向他进贡。
1CHR|18|3|琐巴 王 哈大底谢 往 幼发拉底河 去，要巩固自己的国权。 大卫 攻打他，直到 哈马 ，
1CHR|18|4|夺了他的战车一千，俘掳了骑兵七千人，步兵二万人。 大卫 把所有战马的蹄筋砍断，只留下一百辆战车。
1CHR|18|5|大马士革 的 亚兰 人来帮助 琐巴 王 哈大底谢 ， 大卫 杀了 亚兰 人二万二千。
1CHR|18|6|于是 大卫 在 大马士革 的 亚兰 地设立军营 ， 亚兰 人就臣服 大卫 ，向他进贡。 大卫 无论往哪里去，耶和华都使他得胜。
1CHR|18|7|大卫 夺了 哈大底谢 臣仆拥有的金盾牌，带到 耶路撒冷 。
1CHR|18|8|大卫 又从 哈大底谢 的 提巴 和 均 二城夺取了许多的铜；后来 所罗门 用这些铜制造铜海、铜柱和铜器。
1CHR|18|9|哈马 王 陀乌 听见 大卫 击败 琐巴 王 哈大底谢 的全军，
1CHR|18|10|就派他儿子 哈多兰 到 大卫 王那里，向他请安，为他祝福，因他与 哈大底谢 争战，并且击败了他；原来 哈大底谢 与 陀乌 常常争战。 哈多兰 带了金银铜的各样器皿来。
1CHR|18|11|大卫 王把这些器皿，以及从各国夺来的金银，就是从 以东 、 摩押 、 亚扪 人、 非利士 人、 亚玛力 所夺来的，都分别为圣献给耶和华。
1CHR|18|12|洗鲁雅 的儿子 亚比筛 在 盐谷 击杀了一万八千 以东 人。
1CHR|18|13|大卫 在 以东 设立军营， 以东 人就都臣服他。 大卫 无论往哪里去，耶和华都使他得胜。
1CHR|18|14|大卫 作全 以色列 的王，又向众百姓秉公行义。
1CHR|18|15|洗鲁雅 的儿子 约押 作元帅； 亚希律 的儿子 约沙法 作史官；
1CHR|18|16|亚希突 的儿子 撒督 和 亚比亚他 的儿子 亚希米勒 作祭司； 沙威沙 作书记；
1CHR|18|17|耶何耶大 的儿子 比拿雅 管辖 基利提 人和 比利提 人。 大卫 的众儿子都在王的左右作领袖。
1CHR|19|1|此后， 亚扪 人的王 拿辖 死了，他儿子接续他作王。
1CHR|19|2|大卫 说：“ 哈嫩 的父亲 拿辖 怎样向我施恩，我也要怎样向 哈嫩 施恩。”于是 大卫 派使者为他的父亲安慰他。 大卫 的臣仆到了 亚扪 人的境内来见 哈嫩 ，要安慰他。
1CHR|19|3|但 亚扪 人的领袖对 哈嫩 说：“ 大卫 派人来安慰你，你看他是要尊敬你父亲吗？他的臣仆来见你，不是为了要窥探侦察，而倾覆这地吗？”
1CHR|19|4|哈嫩 就抓住 大卫 的臣仆，剃去他们的胡须，又割断他们下半截的衣服，露出臀部，然后放了他们。
1CHR|19|5|他们走了，有人把臣仆所遭遇的事告诉 大卫 ，他就派人去迎接他们，因为这些人觉得很羞耻。王说：“可以住在 耶利哥 ，等到胡须长出来再回来。”
1CHR|19|6|亚扪 人看到 大卫 憎恶他们， 哈嫩 和 亚扪 人就派人拿一千他连得银子，从 美索不达米亚 、 亚兰．玛迦 、 琐巴 雇用战车和骑兵。
1CHR|19|7|他们雇了三万二千辆战车，以及 玛迦 王和他的军兵；这些部队来安营在 米底巴 前。 亚扪 人也从他们的城里出来，聚集预备作战。
1CHR|19|8|大卫 听见了，就派 约押 和所有勇猛的军队出去。
1CHR|19|9|亚扪 人出来，在城门前摆阵，前来的诸王另在郊野摆阵。
1CHR|19|10|约押 看见战阵对着他前后摆列，就把从 以色列 所有精兵中挑选出来的，摆阵迎战 亚兰 人。
1CHR|19|11|他把其余的兵交在他兄弟 亚比筛 手里，他们就摆阵迎战 亚扪 人。
1CHR|19|12|约押 说：“ 亚兰 人若强过我，你就来帮助我； 亚扪 人若强过你，我就去帮助你。
1CHR|19|13|你要刚强，我们要为自己的百姓，为我们上帝的城镇奋勇。愿耶和华照他所看为好的去做！”
1CHR|19|14|于是， 约押 和跟随他的士兵前进攻打 亚兰 人； 亚兰 人在他面前逃跑。
1CHR|19|15|亚扪 人见 亚兰 人逃跑，他们也在 约押 的兄弟 亚比筛 面前逃跑进城。 约押 就回 耶路撒冷 去了。
1CHR|19|16|亚兰 人见自己被 以色列 打败，就派使者把 大河 那边的 亚兰 人调来，由 哈大底谢 的将军 朔法 在他们前面率领。
1CHR|19|17|有人告诉 大卫 ，他就聚集 以色列 众人过 约旦河 ，来到 亚兰 人那里，迎着他们摆阵。 大卫 摆阵攻击 亚兰 人， 亚兰 人就与他打仗。
1CHR|19|18|亚兰 人在 以色列 人面前逃跑。 大卫 杀了 亚兰 七千辆战车的士兵，四万步兵，又杀死 亚兰 的将军 朔法 。
1CHR|19|19|哈大底谢 的臣仆见自己被 以色列 打败，就与 大卫 讲和，臣服他。于是 亚兰 人不愿再帮助 亚扪 人了。
1CHR|20|1|到了年初，诸王出征的时候， 约押 率领军兵蹂躏 亚扪 人的地，前来围攻 拉巴 ； 大卫 仍住在 耶路撒冷 。 约押 攻打 拉巴 ，把它毁坏。
1CHR|20|2|大卫 夺了 米勒公 所戴的冠冕，其上的金子重一他连得，又嵌着宝石。这冠冕就戴在 大卫 头上。 大卫 又从城里夺了许多财物，
1CHR|20|3|把城里的百姓拉出来，放在锯下，或铁耙下，或斧 的下面； 大卫 待 亚扪 各城的居民都是如此。于是， 大卫 和全军都回 耶路撒冷 去了。
1CHR|20|4|后来， 以色列 人在 基色 与 非利士 人打仗。 户沙 人 西比该 杀了巨人族的后裔 细派 ， 非利士 人就被制伏了。
1CHR|20|5|他们又与 非利士 人打仗。 睚珥 的儿子 伊勒哈难 杀了 迦特 人 歌利亚 的兄弟 拉哈米 ；这人的枪杆粗如织布机的轴。
1CHR|20|6|又有一次，他们在 迦特 打仗。那里有一个身材高大的人，手指脚趾都是六根，共有二十四根；他也是巨人族的后裔。
1CHR|20|7|他向 以色列 骂阵， 大卫 的哥哥 示米亚 的儿子 约拿单 就杀了他。
1CHR|20|8|这些人是 迦特 巨人族的后裔，都仆倒在 大卫 和他仆人的手下。
1CHR|21|1|撒但起来攻击 以色列 ，激起 大卫 数点以色列人。
1CHR|21|2|大卫 对 约押 和百姓的领袖说：“去，数点 以色列 人，从 别是巴 直到 但 ，回来告诉我，我好知道他们的数目。”
1CHR|21|3|约押 说：“愿耶和华使他的百姓比现在加增百倍。我主我王啊，他们不都是我主的仆人吗？我主为何吩咐行这事，为何使 以色列 陷入罪里呢？”
1CHR|21|4|但王坚持他对 约押 的命令。 约押 就出去，来回走遍 以色列 ，然后回到 耶路撒冷 。
1CHR|21|5|约押 向 大卫 报告百姓的总数：全 以色列 拿刀的有一百一十万人； 犹大 拿刀的有四十七万人。
1CHR|21|6|惟有 利未 人和 便雅悯 人没有算在其中，因为 约押 厌恶王的这命令。
1CHR|21|7|这件事在上帝眼中看为恶，上帝就降灾给 以色列 。
1CHR|21|8|大卫 对上帝说：“我做这事大大有罪了。现在求你除掉仆人的罪孽，因为我所做的非常愚昧。”
1CHR|21|9|耶和华吩咐 迦得 ， 大卫 的先见，说：
1CHR|21|10|“你去告诉 大卫 说：‘耶和华如此说：我列出三样灾祸给你，随你选择一样，我好降与你。’”
1CHR|21|11|于是， 迦得 来到 大卫 那里，对他说：“耶和华如此说：‘你可以随意选择：
1CHR|21|12|三年的饥荒，或败在敌人面前，被敌人的刀追杀三个月，或在国中三日有耶和华的刀，就是瘟疫，让耶和华的使者在 以色列 全境施行毁灭呢？’现在你要想一想，我怎样去回覆那差我来的。”
1CHR|21|13|大卫 对 迦得 说：“我很为难。我宁愿落在耶和华的手里，因为他有丰盛的怜悯；我不愿落在人的手里。”
1CHR|21|14|于是，耶和华降瘟疫给 以色列 ， 以色列 中死了七万人。
1CHR|21|15|上帝派遣使者去毁灭 耶路撒冷 ，刚要毁灭的时候，耶和华看见就改变心意，不降这灾了。他吩咐那灭城的天使说：“够了，住手吧！”耶和华的使者正站在 耶布斯 人 阿珥楠 的禾场那里。
1CHR|21|16|大卫 举目，看见耶和华的使者站在天和地之间，手里有拔出来的刀，伸在 耶路撒冷 以上。 大卫 和长老都披上麻布，脸伏于地。
1CHR|21|17|大卫 向上帝说：“吩咐数点百姓的不是我吗？是我犯了罪，行了大恶，但这群羊做了什么呢？耶和华－我的上帝啊，愿你的手攻击我和我的父家，不要降瘟疫给你的百姓。”
1CHR|21|18|耶和华的使者吩咐 迦得 去告诉 大卫 ，叫他上去，在 耶布斯 人 阿珥楠 的禾场上为耶和华立一座坛。
1CHR|21|19|大卫 就照着 迦得 奉耶和华名所说的话上去。
1CHR|21|20|阿珥楠 回头看见天使，跟他在一起的四个儿子都藏起来了， 阿珥楠 继续打麦子。
1CHR|21|21|大卫 到了 阿珥楠 那里， 阿珥楠 观看，看见 大卫 ，就从禾场上出去，脸伏于地，向他下拜。
1CHR|21|22|大卫 对 阿珥楠 说：“你把这禾场的地方给我，照着十足的价钱卖给我，我好在其上为耶和华筑一座坛，使瘟疫在百姓中停止。”
1CHR|21|23|阿珥楠 对 大卫 说：“请用这禾场吧，愿我主我王照你眼中看为好的去做。看，我提供牛作燔祭，打粮的器具作柴，麦子作素祭，这一切我全都提供。”
1CHR|21|24|大卫 王对 阿珥楠 说：“不，我一定要按十足的价钱买；因我不能用你的东西献给耶和华，也不能用白得之物献为燔祭。”
1CHR|21|25|于是 大卫 为那个地方付了六百舍客勒重的金子给 阿珥楠 。
1CHR|21|26|大卫 在那里为耶和华筑了一座坛，献燔祭和平安祭，求告耶和华。耶和华就应允他，使火从天降在燔祭坛上。
1CHR|21|27|耶和华吩咐使者，他就收刀入鞘。
1CHR|21|28|那时， 大卫 见耶和华在 耶布斯 人 阿珥楠 的禾场上应允了他，就在那里献祭。
1CHR|21|29|摩西 在旷野所造之耶和华的帐幕和燔祭坛，当时都在 基遍 的丘坛，
1CHR|21|30|只是 大卫 不能前去求问上帝，因为他惧怕耶和华使者的刀。
1CHR|22|1|大卫 说：“这是耶和华上帝的殿，这是 以色列 献燔祭的坛。”
1CHR|22|2|大卫 吩咐人召集住 以色列 地的寄居者，又派石匠凿石头，要建造上帝的殿。
1CHR|22|3|大卫 预备许多铁，要做门上的钉子和钩子，又预备许多铜，多得无法可秤；
1CHR|22|4|还有无数的香柏木，因为 西顿 人和 推罗 人给 大卫 运了许多香柏木来。
1CHR|22|5|大卫 说：“我儿子 所罗门 还年幼脆弱，要为耶和华建造的殿宇必须高大辉煌，使名声荣耀传遍万国，所以我要为殿预备。”于是， 大卫 在未死之前预备了许多材料。
1CHR|22|6|大卫 召了他儿子 所罗门 来，吩咐他为耶和华－ 以色列 的上帝建造殿宇。
1CHR|22|7|大卫 对 所罗门 说：“我儿啊，我心里本想为耶和华－我上帝的名建造殿宇，
1CHR|22|8|可是耶和华的话临到我说：‘你流了许多的血，打了多次大仗；你不可为我的名建造殿宇，因为你在我面前使许多血流在地上。
1CHR|22|9|看哪，你要生一个儿子，他必成为安宁的人；我必使他得享安宁，不被四围仇敌扰乱。他的名字要叫 所罗门 ，在他的日子，我必使 以色列 平安康泰。
1CHR|22|10|他必为我的名建造殿宇。他要作我的子，我要作他的父。我必坚定他国度的王位，使他治理 以色列 ，直到永远。’
1CHR|22|11|我儿啊，现今愿耶和华与你同在，使你亨通，建造耶和华－你上帝的殿，正如他指着你所说的。
1CHR|22|12|但愿耶和华赐你聪明智慧，好按着他吩咐你的去治理 以色列 ，遵行耶和华－你上帝的律法。
1CHR|22|13|那时候，你若谨守遵行耶和华藉 摩西 吩咐 以色列 的律例典章，就得亨通。你当刚强壮胆，不要惧怕，也不要惊惶。
1CHR|22|14|看哪，我辛苦地为耶和华的殿预备了十万他连得金子，一百万他连得银子，铜和铁多得无法可秤；我也预备了木头、石头，你还可以增添。
1CHR|22|15|你有许多工匠，就是石匠、木匠，和一切能做各样工的巧匠，
1CHR|22|16|以及无数的金银铜铁。你当起来做工，愿耶和华与你同在。”
1CHR|22|17|大卫 又吩咐 以色列 的众官长帮助他儿子 所罗门 ：
1CHR|22|18|“耶和华－你们的上帝不是与你们同在吗？他不是使你们四围都平安吗？因他已将这地的居民交在我手中，这地已在耶和华与他百姓面前制伏了。
1CHR|22|19|现在你们应当立定心意，寻求耶和华－你们的上帝。你们当起来建造耶和华上帝的圣所，好将耶和华的约柜和上帝神圣的器皿都搬进为耶和华的名建造的殿里。”
1CHR|23|1|大卫 年纪老迈，日子满足，就立他儿子 所罗门 作 以色列 的王。
1CHR|23|2|大卫 召集 以色列 的众领袖、祭司和 利未 人。
1CHR|23|3|利未 人三十岁以上的都被数点，他们男丁的数目共有三万八千；
1CHR|23|4|其中有二万四千人管理耶和华殿的事务，有六千人作官长和审判官，
1CHR|23|5|有四千人作门口的守卫，又有四千人颂赞耶和华，用 大卫 造的乐器来颂赞。
1CHR|23|6|大卫 把 利未 人 革顺 、 哥辖 、 米拉利 的子孙分了班次。
1CHR|23|7|属 革顺 的有 拉但 和 示每 。
1CHR|23|8|拉但 的长子是 耶歇 ，还有 西坦 和 约珥 ，共三人。
1CHR|23|9|示每 的儿子是 示罗密 、 哈薛 、 哈兰 三人。这是 拉但 族的族长。
1CHR|23|10|示每 的儿子是 雅哈 、 细拿 、 耶乌施 、 比利亚 ，这四人是 示每 的儿子。
1CHR|23|11|雅哈 是长子， 细撒 是次子。但 耶乌施 和 比利亚 的子孙不多，所以算为一族。
1CHR|23|12|哥辖 的儿子是 暗兰 、 以斯哈 、 希伯伦 、 乌薛 ，共四人。
1CHR|23|13|暗兰 的儿子是 亚伦 和 摩西 。 亚伦 被分别出来，把至圣之物分别为圣，使他和他的子孙在耶和华面前烧香、事奉他，奉他的名祝福，直到永远。
1CHR|23|14|至于神人 摩西 ，他的子孙记名在 利未 支派下。
1CHR|23|15|摩西 的儿子是 革舜 和 以利以谢 。
1CHR|23|16|革舜 的儿子，长子是 细布业 ；
1CHR|23|17|以利以谢 的儿子，长子是 利哈比雅 。 以利以谢 没有别的儿子，但 利哈比雅 的子孙很多。
1CHR|23|18|以斯哈 的儿子，长子是 示罗密 。
1CHR|23|19|希伯伦 的儿子，长子是 耶利雅 ，次子是 亚玛利亚 ，三子是 雅哈悉 ，四子是 耶加面 。
1CHR|23|20|乌薛 的儿子，长子是 米迦 ，次子是 耶西雅 。
1CHR|23|21|米拉利 的儿子是 抹利 和 母示 。 抹利 的儿子是 以利亚撒 和 基士 。
1CHR|23|22|以利亚撒 死了，没有儿子，只有女儿，他们本族 基士 的几个儿子娶了她们为妻。
1CHR|23|23|母示 的儿子是 末力 、 以得 、 耶列末 ，共三人。
1CHR|23|24|以上是 利未 子孙作族长的，按着父系、照着男丁的数目，二十岁以上登记的，都办理耶和华殿的事务。
1CHR|23|25|大卫 说：“耶和华－ 以色列 的上帝已经使他的百姓得享安宁，他永远住在 耶路撒冷 。
1CHR|23|26|因此， 利未 人不必再抬帐幕和其中所使用的一切器皿了。”
1CHR|23|27|照着 大卫 临终的话， 利未 人二十岁以上的都被数点。
1CHR|23|28|他们的职务是作 亚伦 子孙的帮手，在耶和华的殿事奉，照管院子和屋子，洁净一切圣物，办理上帝殿的事务。
1CHR|23|29|他们负责预备供饼、素祭的细面和无酵薄饼，或用盘烤，或用油调和的祭物，确认其数量和大小。
1CHR|23|30|每日早晚、安息日、初一，以及节期，按数照例，经常献燔祭给耶和华的时候，他们站立称谢赞美耶和华。
1CHR|23|31|
1CHR|23|32|他们照管会幕和圣所，服事他们的弟兄 亚伦 的子孙，办理耶和华殿的事务。
1CHR|24|1|亚伦 子孙的班次如下： 亚伦 的儿子是 拿答 、 亚比户 、 以利亚撒 、 以他玛 。
1CHR|24|2|拿答 和 亚比户 死在他们父亲之先，没有留下儿子；因此， 以利亚撒 和 以他玛 担任祭司的职分。
1CHR|24|3|大卫 和 以利亚撒 的子孙 撒督 ，以及 以他玛 的子孙 亚希米勒 ，把他们按照任务分成班次，
1CHR|24|4|发现 以利亚撒 子孙中作领袖的，比 以他玛 子孙中作领袖的更多，就分班如下： 以利亚撒 的子孙中有十六个族长， 以他玛 的子孙中有八个族长。
1CHR|24|5|他们抽签分配，彼此一样。在圣所和上帝面前作领袖的有 以利亚撒 的子孙，也有 以他玛 的子孙。
1CHR|24|6|作书记的 利未 人 拿坦业 的儿子 示玛雅 在王和领袖，与 撒督 祭司、 亚比亚他 的儿子 亚希米勒 ，以及祭司和 利未 人的族长面前记录他们的名字；在 以利亚撒 的子孙中取一族，在 以他玛 的子孙中也取一族。
1CHR|24|7|抽签的时候，第一签抽到的是 耶何雅立 ，第二是 耶大雅 ，
1CHR|24|8|第三是 哈琳 ，第四是 梭琳 ，
1CHR|24|9|第五是 玛基雅 ，第六是 米雅民 ，
1CHR|24|10|第七是 哈歌斯 ，第八是 亚比雅 ，
1CHR|24|11|第九是 耶书亚 ，第十是 示迦尼 ，
1CHR|24|12|第十一是 以利亚实 ，第十二是 雅金 ，
1CHR|24|13|第十三是 胡巴 ，第十四是 耶是比押 ，
1CHR|24|14|第十五是 璧迦 ，第十六是 音麦 ，
1CHR|24|15|第十七是 希悉 ，第十八是 哈辟悉 ，
1CHR|24|16|第十九是 毗他希雅 ，第二十是 以西结 ，
1CHR|24|17|第二十一是 雅斤 ，第二十二是 迦末 ，
1CHR|24|18|第二十三是 第来雅 ，第二十四是 玛西亚 。
1CHR|24|19|这就是他们事奉的班次，要照耶和华－ 以色列 的上帝藉他们祖宗 亚伦 所吩咐的条例，进入耶和华的殿办理事务。
1CHR|24|20|利未 其余的子孙如下： 暗兰 的子孙中有 书巴业 ； 书巴业 的子孙中有 耶希底亚 。
1CHR|24|21|属 利哈比雅 ， 利哈比雅 的儿子中有长子 伊示雅 。
1CHR|24|22|属 以斯哈 人的有 示罗摩 ； 示罗摩 的子孙中有 雅哈 。
1CHR|24|23|希伯伦 的儿子中有长子 耶利雅 ，次子 亚玛利亚 ，三子 雅哈悉 ，四子 耶加面 。
1CHR|24|24|乌薛 的子孙中有 米迦 ； 米迦 的子孙中有 沙密 。
1CHR|24|25|米迦 的兄弟是 伊示雅 ； 伊示雅 的子孙中有 撒迦利雅 。
1CHR|24|26|米拉利 的儿子是 抹利 和 母示 ； 雅西雅 的子孙中有 比挪 ；
1CHR|24|27|米拉利 的子孙中有属 雅西雅 的 比挪 、 朔含 、 撒刻 、 伊比利 。
1CHR|24|28|属 抹利 的有 以利亚撒 ； 以利亚撒 没有儿子。
1CHR|24|29|属 基士 ， 基士 的子孙中有 耶拉篾 。
1CHR|24|30|母示 的儿子是 末力 、 以得 、 耶利末 。按着宗族，这些都是 利未 的子孙。
1CHR|24|31|他们在 大卫 王和 撒督 ，以及 亚希米勒 与祭司和 利未 人的族长面前也抽签，正如他们弟兄 亚伦 的子孙一样。各族的族长与最年轻的兄弟都一样。
1CHR|25|1|大卫 和事奉团队的众领袖分派 亚萨 、 希幔 ，以及 耶杜顿 的子孙唱歌 ，以弹琴、鼓瑟、敲钹伴奏。他们供职的人数如下：
1CHR|25|2|亚萨 的儿子 撒刻 、 约瑟 、 尼探雅 、 亚萨利拉 ， 亚萨 的儿子都在 亚萨 的指导下，遵王的指示唱歌。
1CHR|25|3|属 耶杜顿 ， 耶杜顿 的儿子 基大利 、 西利 、 耶筛亚 、 示每 、 哈沙比雅 、 玛他提雅 共六人，都在他们父亲 耶杜顿 的指导下唱歌，以弹琴伴奏，称谢，颂赞耶和华。
1CHR|25|4|属 希幔 ， 希幔 的儿子是 布基雅 、 玛探雅 、 乌薛 、 细布业 、 耶利末 、 哈拿尼雅 、 哈拿尼 、 以利亚他 、 基大利提 、 罗幔提．以谢 、 约施比加沙 、 玛罗提 、 何提 、 玛哈秀 。
1CHR|25|5|这些都是 希幔 的儿子； 希幔 奉上帝之命作王的先见，吹角颂赞。上帝赐给 希幔 十四个儿子，三个女儿，
1CHR|25|6|他们都在父亲的指导下，在耶和华的殿唱歌，以敲钹、弹琴、鼓瑟伴奏，遵从王的指示，在上帝的殿里事奉。 亚萨 、 耶杜顿 、 希幔 ，
1CHR|25|7|他们和他们的弟兄学习颂赞耶和华，精通者的数目共有二百八十八人。
1CHR|25|8|这些人无论大小，为师的、为徒的，都一同抽签分了班次。
1CHR|25|9|抽签的时候，第一签抽到的是 亚萨 的儿子 约瑟 。第二是 基大利 ；他和他兄弟，以及儿子共十二人。
1CHR|25|10|第三是 撒刻 ，他儿子和他兄弟共十二人。
1CHR|25|11|第四是 伊洗利 ，他儿子和他兄弟共十二人。
1CHR|25|12|第五是 尼探雅 ，他儿子和他兄弟共十二人。
1CHR|25|13|第六是 布基雅 ，他儿子和他兄弟共十二人。
1CHR|25|14|第七是 耶萨利拉 ，他儿子和他兄弟共十二人。
1CHR|25|15|第八是 耶筛亚 ，他儿子和他兄弟共十二人。
1CHR|25|16|第九是 玛探雅 ，他儿子和他兄弟共十二人。
1CHR|25|17|第十是 示每 ，他儿子和他兄弟共十二人。
1CHR|25|18|第十一是 亚萨烈 ，他儿子和他兄弟共十二人。
1CHR|25|19|第十二是 哈沙比雅 ，他儿子和他兄弟共十二人。
1CHR|25|20|第十三是 书巴业 ，他儿子和他兄弟共十二人。
1CHR|25|21|第十四是 玛他提雅 ，他儿子和他兄弟共十二人。
1CHR|25|22|第十五是 耶列末 ，他儿子和他兄弟共十二人。
1CHR|25|23|第十六是 哈拿尼雅 ，他儿子和他兄弟共十二人。
1CHR|25|24|第十七是 约施比加沙 ，他儿子和他兄弟共十二人。
1CHR|25|25|第十八是 哈拿尼 ，他儿子和他兄弟共十二人。
1CHR|25|26|第十九是 玛罗提 ，他儿子和他兄弟共十二人。
1CHR|25|27|第二十是 以利亚他 ，他儿子和他兄弟共十二人。
1CHR|25|28|第二十一是 何提 ，他儿子和他兄弟共十二人。
1CHR|25|29|第二十二是 基大利提 ，他儿子和他兄弟共十二人。
1CHR|25|30|第二十三是 玛哈秀 ，他儿子和他兄弟共十二人。
1CHR|25|31|第二十四是 罗幔提．以谢 ，他儿子和他兄弟共十二人。
1CHR|26|1|门口守卫的班次如下： 可拉 族 以比雅撒 的子孙中，有 可利 的儿子 米施利米雅 。
1CHR|26|2|米施利米雅 的长子是 撒迦利亚 ，次子是 耶叠 ，三子是 西巴第雅 ，四子是 耶提聂 ，
1CHR|26|3|五子是 以拦 ，六子是 约哈难 ，七子是 以利约乃 。
1CHR|26|4|俄别．以东 的长子是 示玛雅 ，次子是 约萨拔 ，三子是 约亚 ，四子是 沙甲 ，五子是 拿坦业 ，
1CHR|26|5|六子是 亚米利 ，七子是 以萨迦 ，八子是 毗乌利太 ，因为上帝赐福给 俄别．以东 。
1CHR|26|6|他的儿子 示玛雅 生了几个儿子，都是大能的勇士，管理父亲的家。
1CHR|26|7|示玛雅 的儿子是 俄得尼 、 利法益 、 俄备得 、 以利萨巴 。 以利萨巴 的兄弟 以利户 和 西玛迦 是能人。
1CHR|26|8|这些都是 俄别．以东 的子孙，他们和他们的儿子，以及兄弟，都是善于办事的能人。属 俄别．以东 的共六十二人。
1CHR|26|9|米施利米雅 的儿子和兄弟都是能人，共十八人。
1CHR|26|10|米拉利 子孙中的 何萨 有几个儿子：为首的是 申利 ；他原不是长子，是他父亲立他为首的，
1CHR|26|11|次子是 希勒家 ，三子是 底巴利雅 ，四子是 撒迦利亚 。 何萨 的儿子和兄弟共十三人。
1CHR|26|12|这些是门口守卫的班次，各随他们的班长，与他们的兄弟一同在耶和华殿里按班供职。
1CHR|26|13|他们无论大小，都按着父系抽签，分守各门。
1CHR|26|14|抽到东门的是 示利米雅 ；他的儿子 撒迦利亚 是精明的谋士，抽到北门。
1CHR|26|15|俄别．以东 守南门，他的儿子守仓库。
1CHR|26|16|书聘 与 何萨 守西门，在靠近 沙利基 门、通往上去的街道上，守卫与守卫相对。
1CHR|26|17|东门有六个 利未 人 ，北门每日有四人，南门每日有四人，库房有两人轮流替换。
1CHR|26|18|至于走廊，在西面街道上有四人，在走廊上有两人。
1CHR|26|19|以上是 可拉 子孙和 米拉利 子孙门口守卫的班次。
1CHR|26|20|利未 人中有 亚希雅 管理上帝殿的库房和圣物的库房。
1CHR|26|21|拉但 子孙中， 革顺 族属 拉但 、作族长的是 革顺 族属 拉但 的 耶希伊利 。
1CHR|26|22|耶希伊利 的儿子 西坦 和他兄弟 约珥 管理耶和华殿的库房。
1CHR|26|23|暗兰 人、 以斯哈 人、 希伯伦 人、 乌薛 人也有职务。
1CHR|26|24|摩西 的孙子， 革舜 的儿子 细布业 管理库房。
1CHR|26|25|还有他的弟兄： 以利以谢 ， 以利以谢 的儿子 利哈比雅 ， 利哈比雅 的儿子 耶筛亚 ， 耶筛亚 的儿子 约兰 ， 约兰 的儿子 细基利 ， 细基利 的儿子 示罗密 。
1CHR|26|26|这 示罗密 和他的兄弟管理一切库房的圣物，就是 大卫 王和众族长、千夫长、百夫长，以及军官所分别为圣之物。
1CHR|26|27|他们把打仗时夺取的一些财物分别为圣，用来修造耶和华的殿。
1CHR|26|28|凡 撒母耳 先见、 基士 的儿子 扫罗 、 尼珥 的儿子 押尼珥 、 洗鲁雅 的儿子 约押 分别为圣的，一切分别为圣之物都归 示罗密 和他的兄弟掌管。
1CHR|26|29|以斯哈 人有 基拿尼雅 和他众儿子作官长和审判官，管理 以色列 对外的事务。
1CHR|26|30|希伯伦 人有 哈沙比雅 和他弟兄一千七百人，都是能人，在 约旦河 西监督 以色列 人，办理耶和华的一切工作和王的事务。
1CHR|26|31|希伯伦 人中有 耶利雅 作族长。 大卫 作王第四十年在各族各家从事寻访，在 基列 的 雅谢 ，从这族中发现大能的勇士。
1CHR|26|32|耶利雅 的弟兄有二千七百人，都是能人，又是族长； 大卫 王派他们在 吕便 人、 迦得 人、 玛拿西 半支派中管理上帝和王的一切事务。
1CHR|27|1|以色列 人的族长、千夫长、百夫长和官长都分配班次，每班二万四千人，整年按月轮流出入，按班次服事王。
1CHR|27|2|正月第一班的班长是 撒巴第业 的儿子 雅朔班 ；他班内有二万四千人。
1CHR|27|3|他是 法勒斯 的后裔，统管正月军队所有的官长。
1CHR|27|4|二月的班长是 亚何亚 人 朵代 ，他的班有总长 密基罗 ；他班内有二万四千人。
1CHR|27|5|三月第三班的班长是 耶何耶大 祭司长的儿子 比拿雅 ；他班内有二万四千人。
1CHR|27|6|这 比拿雅 是那三十人中的勇士，管理那三十人；他班内又有他儿子 暗米萨拔 。
1CHR|27|7|四月第四班的班长是 约押 的兄弟 亚撒黑 。接续他的是他儿子 西巴第雅 ；他班内有二万四千人。
1CHR|27|8|五月第五班的班长是 伊斯拉 人 珊合 ；他班内有二万四千人。
1CHR|27|9|六月第六班的班长是 提哥亚 人 益吉 的儿子 以拉 ；他班内有二万四千人。
1CHR|27|10|七月第七班的班长是 以法莲 族 比伦 人 希利斯 ；他班内有二万四千人。
1CHR|27|11|八月第八班的班长是 谢拉 族 户沙 人 西比该 ；他班内有二万四千人。
1CHR|27|12|九月第九班的班长是 便雅悯 族 亚拿突 人 亚比以谢 ；他班内有二万四千人。
1CHR|27|13|十月第十班的班长是 谢拉 族 尼陀法 人 玛哈莱 ；他班内有二万四千人。
1CHR|27|14|十一月第十一班的班长是 以法莲 族 比拉顿 人 比拿雅 ；他班内有二万四千人。
1CHR|27|15|十二月第十二班的班长是 俄陀聂 族 尼陀法 人 黑玳 ；他班内有二万四千人。
1CHR|27|16|管理 以色列 众支派的如下：管 吕便 人的是 细基利 的儿子 以利以谢 ；管 西缅 人的是 玛迦 的儿子 示法提雅 ；
1CHR|27|17|管 利未 的是 基摩利 的儿子 哈沙比雅 ；管 亚伦 子孙的是 撒督 ；
1CHR|27|18|管 犹大 的是 大卫 的一个哥哥 以利户 ；管 以萨迦 的是 米迦勒 的儿子 暗利 ；
1CHR|27|19|管 西布伦 的是 俄巴第雅 的儿子 伊施玛雅 ；管 拿弗他利 的是 亚斯列 的儿子 耶利摩 ；
1CHR|27|20|管 以法莲 的是 阿撒细雅 的儿子 何细亚 ；管 玛拿西 半支派的是 毗大雅 的儿子 约珥 ；
1CHR|27|21|管 基列 地 玛拿西 半支派的是 撒迦利亚 的儿子 易多 ；管 便雅悯 的是 押尼珥 的儿子 雅西业 ；
1CHR|27|22|管 但 的是 耶罗罕 的儿子 亚萨列 。以上是 以色列 众支派的领袖。
1CHR|27|23|以色列 人二十岁以下的， 大卫 没有记其数目；因耶和华曾应许，必加增 以色列 人如天上的星那样多。
1CHR|27|24|洗鲁雅 的儿子 约押 开始数点，却还没有数完。为了这事，烈怒临到 以色列 ，数点的数目也没有写在《大卫王记》上。
1CHR|27|25|管理王的库房的是 亚叠 的儿子 押斯马威 。管理田野、城镇、村庄、堡垒之仓库的是 乌西雅 的儿子 约拿单 。
1CHR|27|26|管理耕田种地的是 基绿 的儿子 以斯利 。
1CHR|27|27|管理葡萄园的是 拉玛 人 示每 。管理葡萄园酒窖的是 实弗米 人 撒巴底 。
1CHR|27|28|管理 谢非拉 橄榄树和桑树的是 基第利 人 巴勒．哈南 。管理油库的是 约阿施 。
1CHR|27|29|管理 沙仑 牧放牛群的是 沙仑 人 施提莱 。管理山谷牧养牛群的是 亚第莱 的儿子 沙法 。
1CHR|27|30|管理骆驼群的是 以实玛利 人 阿比勒 。管理驴群的是 米仑 人 耶希底亚 。管理羊群的是 夏甲 人 雅悉 。
1CHR|27|31|这些都是为 大卫 王管理产业的领袖。
1CHR|27|32|大卫 的叔父 约拿单 作谋士；这人有智慧，又作书记。 哈摩尼 的儿子 耶歇 陪伴王的众儿子。
1CHR|27|33|亚希多弗 作王的谋士。 亚基 人 户筛 作王的顾问。
1CHR|27|34|亚希多弗 之后，有 比拿雅 的儿子 耶何耶大 ，以及 亚比亚他 接续他。 约押 作王的元帅。
1CHR|28|1|大卫 召集 以色列 所有的领袖，各支派的领袖、轮班服事王的官长、千夫长、百夫长、掌管王和王子一切产业牲畜的、宫廷官员、勇士，和所有大能的勇士，都到 耶路撒冷 来。
1CHR|28|2|大卫 王站起来，说：“我的弟兄，我的百姓啊，请听我说！我心里本想建造殿宇，安放耶和华的约柜，作为我们上帝的脚凳，并且我已经预备了建造的材料。
1CHR|28|3|只是上帝对我说：‘你不可为我的名建造殿宇，因你是战士，流了人的血。’
1CHR|28|4|然而，耶和华－ 以色列 的上帝在我父的全家拣选我作 以色列 的王，直到永远。因他拣选 犹大 为领袖，在 犹大 家中拣选我父家，在我父的众儿子里喜悦我，立我作全 以色列 的王。
1CHR|28|5|耶和华赐我许多儿子，在我儿子中拣选我儿子 所罗门 坐耶和华国度的王位，治理 以色列 。
1CHR|28|6|耶和华对我说：‘你儿子 所罗门 必建造我的殿和院宇，因为我拣选他作我的子，我也必作他的父。
1CHR|28|7|他若恒久遵行我的诫命典章如今日一样，我就必坚定他的国，直到永远。’
1CHR|28|8|现今在 以色列 众人眼前，在耶和华的会中，在我们上帝的垂听下，你们务要遵行并寻求耶和华－你们上帝的一切诫命，如此你们就可以承受这美地，并留给你们的子孙，永远为业。
1CHR|28|9|“我儿 所罗门 哪，你当认识耶和华－你父的上帝，全心乐意地事奉他，因为耶和华鉴察众人的心，知道一切心思意念。你若寻求他，他必使你寻见；你若离弃他，他必永远丢弃你。
1CHR|28|10|现在你当谨慎，因耶和华拣选你建造殿宇作为圣所。你当刚强去做。”
1CHR|28|11|大卫 指示他儿子 所罗门 有关殿的走廊、屋子、库房、楼房、内殿和柜盖 之处的样式，
1CHR|28|12|被灵感动所得的一切样式：耶和华殿的院子、周围一切的房屋、上帝殿的库房和圣物库房；
1CHR|28|13|祭司和 利未 人的班次，耶和华殿里各样事奉的工作，耶和华殿里一切事奉用的器皿，
1CHR|28|14|以及各样事奉所用金器的重量，和各样事奉所用银器的重量，
1CHR|28|15|金灯台和金灯的重量，按每一个灯台和灯的重量；银灯台和银灯的重量，按每一个灯台和灯的重量，都按照每一个灯台的用途；
1CHR|28|16|每张供饼桌子的金子重量，和银桌子的银子重量，
1CHR|28|17|纯金的肉叉子、盘子，和壶的重量，金碗，按每个金碗的重量，和银碗，按每个银碗的重量，
1CHR|28|18|纯金香坛的重量，金基路伯座车的样式，基路伯张开翅膀，遮盖耶和华的约柜。
1CHR|28|19|大卫 说：“这一切，所有工作的样式，是耶和华用手写的文件使我明白的。”
1CHR|28|20|大卫 又对他儿子 所罗门 说：“你当刚强壮胆去做！不要惧怕，也不要惊惶，因为耶和华上帝，我的上帝与你同在。他必不撇下你，也不丢弃你，直到耶和华殿的工作都完毕。
1CHR|28|21|看哪，有祭司和 利未 人的班次，为要办理上帝殿各样的事务，又有擅长做各样事务的人，乐意在各样工作上帮助你，并且领袖和众百姓也都听从你的一切命令。”
1CHR|29|1|大卫 王对全会众说：“我儿子 所罗门 是上帝特选的，还年幼脆弱，但这工程浩大，因这殿不是为人，而是为耶和华上帝建造的。
1CHR|29|2|我为我上帝的殿已经尽力，预备金子做金器，银子做银器，铜做铜器，铁做铁器，木做木器，还有红玛瑙、可镶嵌的宝石、彩石、各样的宝石和许多大理石。
1CHR|29|3|此外，因我爱慕我上帝的殿，在预备建造圣殿的一切材料之外，又将我自己积蓄的金银献给我上帝的殿，
1CHR|29|4|就是三千他连得 俄斐 金子、七千他连得纯银，用来贴殿的墙；
1CHR|29|5|金子做金器，银子做银器，并藉工匠的手做一切的工。今日有谁愿意将自己献给耶和华呢？”
1CHR|29|6|于是，众族长和 以色列 各支派的领袖、千夫长、百夫长，以及监管王工作的官长，都乐意奉献。
1CHR|29|7|他们为上帝殿的工程献上五千他连得又一万达利克 金子，一万他连得银子，一万八千他连得铜，十万他连得铁。
1CHR|29|8|凡有宝石的都送入耶和华殿的库房，由 革顺 人 耶歇 的手管理。
1CHR|29|9|因这些人全心乐意献给耶和华，百姓就欢喜， 大卫 王也大大欢喜。
1CHR|29|10|大卫 在全会众眼前称颂耶和华； 大卫 说：“耶和华－ 以色列 的上帝，我们的父，你是应当称颂的，直到永永远远！
1CHR|29|11|耶和华啊，尊大、能力、荣耀、胜利、威严都是你的；天上地下的一切都是你的；耶和华啊，国度是你的，并且你为至高，为万有之首。
1CHR|29|12|丰富尊荣都从你而来，你也治理万物。在你手里有大能大力，你的手使人尊大强盛。
1CHR|29|13|我们的上帝啊，现在我们称谢你，赞美你荣耀之名！
1CHR|29|14|“我算什么，我的百姓算什么，竟然能够如此乐意奉献？因为万物都从你而来，我们把从你的手得来的献给你。
1CHR|29|15|我们在你面前是客旅，是寄居的，与我们的列祖一样。我们在世的日子如影子，没有盼望。
1CHR|29|16|耶和华－我们的上帝啊，我们预备这许多材料，要为你的圣名建造殿宇，都是从你的手而来，都是属你的。
1CHR|29|17|我的上帝啊，我知道你察验人心，喜悦正直；我以正直的心乐意献上这一切。现在我欢喜见你的百姓在此乐意奉献给你。
1CHR|29|18|耶和华－我们列祖 亚伯拉罕 、 以撒 、 以色列 的上帝啊，求你使你的百姓心中常存这样的心思意念，坚定他们的心归向你，
1CHR|29|19|又求你赐我儿子 所罗门 全心遵守你的命令、法度、律例，成就这一切的事，用我所预备的建造殿宇。”
1CHR|29|20|大卫 对全会众说：“你们应当称颂耶和华－你们的上帝。”于是全会众称颂耶和华－他们列祖的上帝，低头向耶和华和王下拜。
1CHR|29|21|次日，他们向耶和华献平安祭和燔祭，献一千头公牛，一千只公绵羊，一千只羔羊，以及同献的浇酒祭，并为 以色列 众人献许多的祭。
1CHR|29|22|那日，他们在耶和华面前吃喝，大大欢乐。 他们再次立 大卫 的儿子 所罗门 作王，膏他归耶和华作君王，又膏 撒督 作祭司。
1CHR|29|23|于是 所罗门 坐在耶和华所赐的王位上，接续他父亲 大卫 作王；他万事亨通，全 以色列 都听从他。
1CHR|29|24|众领袖和勇士，以及 大卫 王的众儿子，都顺服 所罗门 王。
1CHR|29|25|耶和华使 所罗门 在 以色列 众人眼前非常尊大，赐他君王的威严，胜过他以前任何一位 以色列 王。
1CHR|29|26|耶西 的儿子 大卫 作全 以色列 的王。
1CHR|29|27|他作 以色列 王的时期共四十年：在 希伯仑 作王七年，在 耶路撒冷 作王三十三年。
1CHR|29|28|他死的时候年纪老迈，日子满足，享尽荣华富贵。他的儿子 所罗门 接续他作王。
1CHR|29|29|大卫 王自始至终的事迹，看哪，都写在 撒母耳 先见的书上、 拿单 先知的书上和 迦得 先见的书上，
1CHR|29|30|包括他治国的一切和他英勇的事迹，以及他和 以色列 与世上列国所经历的事。
2CHR|1|1|大卫 的儿子 所罗门 巩固他的国度；耶和华－他的上帝与他同在，使他极其尊大。
2CHR|1|2|所罗门 吩咐全 以色列 ，就是千夫长、百夫长、审判官、全 以色列 的众领袖和族长前来。
2CHR|1|3|所罗门 率领全会众往 基遍 的丘坛去，因那里有上帝的会幕，就是耶和华的仆人 摩西 在旷野所造的。
2CHR|1|4|只是上帝的约柜， 大卫 已经从 基列．耶琳 接到他所预备的地方，因他曾在 耶路撒冷 为约柜支搭了帐幕，
2CHR|1|5|把 户珥 的孙子， 乌利 的儿子 比撒列 所造的铜坛摆在 基遍 耶和华的会幕前。 所罗门 和会众求告耶和华。
2CHR|1|6|所罗门 上到耶和华面前会幕的铜坛那里，在坛上献一千祭牲为燔祭。
2CHR|1|7|当夜，上帝向 所罗门 显现，对他说：“你愿我赐你什么，你可以求。”
2CHR|1|8|所罗门 对上帝说：“你曾向我父亲 大卫 大施慈爱，使我接续他作王。
2CHR|1|9|耶和华上帝啊，现在求你实现向我父亲 大卫 所应许的话；因你立我作这百姓的王，他们如同地上的尘沙那样多。
2CHR|1|10|现在，求你赐我智慧聪明，好在这百姓面前出入；不然，谁能判断你这么多的百姓呢？”
2CHR|1|11|上帝对 所罗门 说：“你有这心意，不求资财、丰富、尊荣，也不求灭绝恨你之人的性命，又不求长寿；我既立你作我百姓的王，你只求智慧聪明，好审判我的百姓，
2CHR|1|12|我必赐你智慧聪明，也必赐你资财、丰富、尊荣，在你以前的列王未曾有过，在你以后也不会再有。”
2CHR|1|13|于是， 所罗门 从 基遍 丘坛会幕前回到 耶路撒冷 ，治理 以色列 。
2CHR|1|14|所罗门 聚集战车骑兵；他有一千四百辆战车，一万二千名骑兵，安置在屯车城，在 耶路撒冷 的王那里。
2CHR|1|15|王在 耶路撒冷 使金银多如石头，香柏木多如 谢非拉 的桑树。
2CHR|1|16|所罗门 的马是从 埃及 和 科威 运来的，是王的商人按着定价从 科威 买来的。
2CHR|1|17|他们从 埃及 进口战车，每辆六百舍客勒银子，马每匹一百五十舍客勒； 赫 人众王和 亚兰 诸王的战车和马，也是经由他们的手出口的。
2CHR|2|1|所罗门 吩咐要为耶和华的名建造殿宇，又为自己的王国建造宫殿。
2CHR|2|2|所罗门 征召七万名扛抬的，八万个在山上凿石头的人，三千六百个监工。
2CHR|2|3|所罗门 派人去见 推罗 王 希兰 ，说：“你曾运香柏木给我父亲 大卫 建造宫殿居住，请你也这样待我。
2CHR|2|4|看哪，我要为耶和华－我上帝的名建造殿宇，分别为圣献给他，在他面前烧芬芳的香，经常献供饼，每早晚、安息日、初一，以及耶和华－我们上帝所定的节期献燔祭。这是 以色列 人永远的定例。
2CHR|2|5|我所要建造的殿宇宏大，因为我们的上帝至大，超乎众神。
2CHR|2|6|天和天上的天，尚且不足他居住，谁能为他建造殿宇呢？我是谁，能为他建造殿宇吗？不过在他面前烧香而已！
2CHR|2|7|现在请你派一个巧匠来，就是善用金、银、铜、铁，和紫色、朱红色、蓝色线做工，并精于雕刻之工的巧匠，与跟我一起在 犹大 和 耶路撒冷 、我父亲 大卫 所预备的巧匠一同做工；
2CHR|2|8|又请你从 黎巴嫩 运香柏木、松木、檀香木到我这里来，因我知道你的仆人擅长砍伐 黎巴嫩 的树木。看哪，我的仆人必帮助你的仆人，
2CHR|2|9|好为我预备许多的木料，因我要建造的殿宇高大出奇。
2CHR|2|10|看哪，我必给你仆人，就是砍伐树木的伐木工，二万歌珥压碎的小麦 ，二万歌珥大麦，二万罢特酒，二万罢特油。”
2CHR|2|11|推罗 王 希兰 写信回答 所罗门 说：“耶和华因为爱他的百姓，所以立你作他们的王。”
2CHR|2|12|又说：“创造天和地的耶和华－ 以色列 的上帝是应当称颂的！他赐给 大卫 王一个有智慧的儿子，使他有见识，有聪明，可以为耶和华建造殿宇，又为自己的王国建造宫殿。
2CHR|2|13|“现在我派一个精巧聪明的人去，他是我的师父 户兰 ，
2CHR|2|14|是 但 支派一个妇人的儿子，父亲是 推罗 人。他善用金、银、铜、铁、石、木，和紫色、蓝色、细麻和朱红色线制造各物，并精于雕刻，又能设计各样交给他做的图案。我派这人与你的巧匠和你父亲－我主 大卫 的巧匠一同做工。
2CHR|2|15|我主所说的小麦、大麦、酒、油，请运来给众仆人。
2CHR|2|16|我们必照你所需用的，从 黎巴嫩 砍伐树木，扎成筏子，浮海运到 约帕 ；你可以从那里运到 耶路撒冷 。”
2CHR|2|17|所罗门 仿照他父亲 大卫 数点所有在 以色列 地寄居的外邦人，共有十五万三千六百名。
2CHR|2|18|他叫其中的七万人作扛抬，八万人在山上凿石头，三千六百人监督百姓工作。
2CHR|3|1|所罗门 在 耶路撒冷 开工建造耶和华的殿，就在耶和华向他父亲 大卫 显现的 摩利亚山 上， 耶布斯 人 阿珥楠 的禾场， 大卫 指定的地方。
2CHR|3|2|所罗门 作王第四年二月初二 开工建造。
2CHR|3|3|所罗门 所建筑的上帝殿的根基是这样：长六十肘，宽二十肘，都按着古时的尺寸。
2CHR|3|4|前面的 走廊长二十肘，与殿的宽度一样，高一百二十肘；里面贴上纯金。
2CHR|3|5|大殿的墙都用松木板遮蔽，又贴上纯金，上面刻着棕树和链子。
2CHR|3|6|他用宝石装饰这殿，使殿华美；金子都是 巴瓦音 的金子。
2CHR|3|7|他用金子贴殿和殿的栋梁、门槛、墙壁、门扇；墙上刻着基路伯。
2CHR|3|8|他建造至圣所，长二十肘，与殿的宽度一样，宽二十肘，都贴上纯金，共用了六百他连得金子。
2CHR|3|9|金的钉子重五十舍客勒。楼房都贴上金子。
2CHR|3|10|他又在至圣所用雕刻的手艺造两个基路伯，包上金子。
2CHR|3|11|两个基路伯的翅膀共长二十肘。这基路伯的一个翅膀长五肘，挨着殿这边的墙；另一个翅膀也长五肘，与那基路伯翅膀相接。
2CHR|3|12|那基路伯的一个翅膀长五肘，挨着殿那边的墙；另一个翅膀也长五肘，与这基路伯的翅膀相接。
2CHR|3|13|这两个基路伯张开翅膀，共长二十肘，用脚站立，脸面向殿。
2CHR|3|14|他又用蓝色、紫色、朱红色线和细麻织幔子，在其上绣基路伯。
2CHR|3|15|他在殿前造了两根柱子，高三十五肘；柱子上面的柱顶高五肘。
2CHR|3|16|他造链子在内殿里，安在柱顶上，又做一百个石榴，安在链子上。
2CHR|3|17|他把两根柱子立在殿前，一根在右边，一根在左边；右边的起名叫 雅斤 ，左边的起名叫 波阿斯 。
2CHR|4|1|他造一座铜坛，长二十肘，宽二十肘，高十肘。
2CHR|4|2|他又铸一个铜海，周围是圆的，直径十肘，高五肘，用绳子量周围是三十肘。
2CHR|4|3|铜海下面的周围有牛的样式，有十肘，绕着铜海；牛有两行，是造铜海的时候铸上去的。
2CHR|4|4|铜海安在十二头铜牛上：三头向北，三头向西，三头向南，三头向东。铜海安在牛上，牛尾都向内。
2CHR|4|5|铜海厚一掌，边如杯边，像百合花，容量是三千罢特。
2CHR|4|6|他又造十个盆：五个放在右边，五个放在左边，作洗涤之用。献燔祭所用之物都洗在盆内；但铜海是为祭司洗涤用的。
2CHR|4|7|他照所定的样式造十个金灯台，放在殿里：五个在右边，五个在左边。
2CHR|4|8|他造十张桌子，放在殿里：五张在右边，五张在左边。他又造一百个金碗。
2CHR|4|9|他建造祭司院和大院，以及院门，门扇包上铜。
2CHR|4|10|他把铜海安在殿的右边，就是东南边。
2CHR|4|11|户兰 又造了盆、铲子和盘子。这样， 户兰 为 所罗门 王做完了上帝殿的工：
2CHR|4|12|两根柱子和柱子顶上两个如碗的柱顶，以及盖着如碗柱顶的两个网子；
2CHR|4|13|四百个石榴，安在两个网子上，每网两行石榴，盖着柱子上面两个如碗的柱顶。
2CHR|4|14|他造盆座，又造其上的盆；
2CHR|4|15|铜海和其下的十二头牛；
2CHR|4|16|盆、铲子、肉叉。巧匠 户兰 给 所罗门 王为耶和华殿造的这一切器皿都是用磨亮的铜，
2CHR|4|17|是王在 约旦 平原、 疏割 和 撒利但 中间的泥巴地铸成的。
2CHR|4|18|所罗门 造这一切器皿，数量很多，铜的重量无法计算。
2CHR|4|19|所罗门 又为上帝的殿造了各样的器皿：金坛和献供饼的供桌；
2CHR|4|20|纯金的灯台和灯盏，可以照定例点在内殿前；
2CHR|4|21|灯台上的花和灯盏，以及灯剪，都是金的，而且是纯金的；
2CHR|4|22|纯金的钳子、盘子、勺子、火盆。至于殿门和至圣所的门扇，以及殿的门扇，都是金的。
2CHR|5|1|所罗门 王做完了耶和华殿一切的工，就把他父亲 大卫 分别为圣的金银和一切器皿都带来，放在上帝殿的库房里。
2CHR|5|2|于是， 所罗门 召集 以色列 的长老、各支派的领袖和 以色列 人的族长到 耶路撒冷 ，要把耶和华的约柜从 大卫城 ，就是 锡安 ，接上来。
2CHR|5|3|在七月节期的时候，所有的 以色列 人都聚集到王那里。
2CHR|5|4|以色列 众长老一来到， 利未 人就抬起约柜。
2CHR|5|5|祭司和 利未 人将约柜请上来，又把会幕和会幕一切的圣器皿都带上来。
2CHR|5|6|所罗门 王和聚集到他那里的 以色列 全会众都在约柜前献牛羊为祭，多得不可胜数，无法计算。
2CHR|5|7|祭司将耶和华的约柜请进内殿，就是至圣所，安置在两个基路伯的翅膀底下约柜自己的地方。
2CHR|5|8|基路伯张开翅膀在约柜上面的地方，从上面遮住约柜和抬柜的杠。
2CHR|5|9|这杠很长，从内殿前的约柜可以看见杠头，从外面却看不见。这杠直到今日还在那里。
2CHR|5|10|约柜里没有别的，只有两块石版，就是 以色列 人出 埃及 ，耶和华与他们立约的时候， 摩西 在 何烈山 所放的。
2CHR|5|11|当时，所有在那里的祭司，不论哪个班次供职的，都使自己分别为圣。祭司从圣所出来的时候，
2CHR|5|12|所有歌唱的 利未 人， 亚萨 、 希幔 、 耶杜顿 ，和他们的众儿子、众弟兄都穿细麻布衣服，站在祭坛的东边敲钹，鼓瑟，弹琴，和他们一起的还有一百二十个吹号的祭司。
2CHR|5|13|吹号的、歌唱的都合一齐声，赞美称谢耶和华。他们配合号筒、铙钹和其他乐器，扬声赞美耶和华： “耶和华本为善， 他的慈爱永远长存！” 那时，耶和华的殿充满了云彩。
2CHR|5|14|祭司因云彩的缘故不能站立供职，因为耶和华的荣光充满了上帝的殿。
2CHR|6|1|那时， 所罗门 说： “耶和华曾说要住在幽暗之处。
2CHR|6|2|我为你建了一座雄伟的殿宇， 作为你永远居住的地方。”
2CHR|6|3|王转过脸来为 以色列 全会众祝福， 以色列 全会众都站立。
2CHR|6|4|所罗门 说：“耶和华－ 以色列 的上帝是应当称颂的！因他亲口向我父 大卫 应许的，也亲手成就了；他曾说：
2CHR|6|5|‘自从那日我领我百姓出 埃及 地以来，我未曾在 以色列 各支派中选择一城，在那里为我的名建造殿宇，也未曾拣选一人作我百姓 以色列 的君王。
2CHR|6|6|但我选择 耶路撒冷 ，使我的名留在那里，又拣选 大卫 治理我的百姓 以色列 。’
2CHR|6|7|我父 大卫 的心意是要为耶和华－ 以色列 上帝的名建殿。
2CHR|6|8|耶和华却对我父 大卫 说：‘你有心为我的名建殿，这心意是好的；
2CHR|6|9|但你不可建殿，惟有你亲生的儿子才可为我的名建殿。’
2CHR|6|10|现在耶和华实现了他所应许的话，使我接续我父 大卫 坐 以色列 的王位，正如耶和华所说的，我也为耶和华－ 以色列 上帝的名建造了这殿。
2CHR|6|11|我将约柜安置在那里，柜内有耶和华的约，就是他与 以色列 人所立的约。”
2CHR|6|12|所罗门 当着 以色列 全会众，站在耶和华的坛前，举起手来。
2CHR|6|13|所罗门 曾造一个铜台，长五肘，宽五肘，高三肘，放在院中。他站在台上，当着 以色列 全会众双膝跪下，向天举手，
2CHR|6|14|说：“耶和华－ 以色列 的上帝啊，天上地下没有神明可与你相比！你向那些尽心行在你面前的仆人守约施慈爱，
2CHR|6|15|这约是你向你仆人 大卫 守的，是你应许他的。你亲口应许，亲手成就，正如今日一样。
2CHR|6|16|耶和华－ 以色列 的上帝啊，你向你仆人我父 大卫 应许说：‘你的子孙若谨慎自己的行为，遵行我的律法，像你在我面前所行的，就不断有人在我面前坐 以色列 的王位。’现在求你信守这话。
2CHR|6|17|耶和华－ 以色列 的上帝啊，现在求你成就向你仆人 大卫 所应许的话。
2CHR|6|18|“上帝果真与世人同住在地上吗？看哪，天和天上的天尚且不足容纳你，何况我所建的这殿呢？
2CHR|6|19|惟求耶和华－我的上帝垂顾仆人的祷告祈求，俯听仆人在你面前的祈祷呼求。
2CHR|6|20|愿你的眼目昼夜看顾这殿，就是你应许立为你名的居所；求你垂听祷告，你仆人向此处的祷告。
2CHR|6|21|你仆人和你百姓 以色列 向此处祈祷的时候，求你从天上你的居所垂听，垂听而赦免。
2CHR|6|22|“人若得罪邻舍，有人强迫他，要他起誓，他来到这殿，在你的坛前起誓，
2CHR|6|23|求你从天上垂听、处理，向你的仆人施行审判，定恶人有罪，照他所行的报应在他头上；定义人为义，照他的义赏赐他。
2CHR|6|24|“你的百姓 以色列 若得罪你，败在仇敌面前，却又归向你，宣认你的名，在这殿里向你祈求祷告，
2CHR|6|25|求你从天上垂听，赦免你百姓 以色列 的罪，使他们归回你赐给他们和他们列祖之地。
2CHR|6|26|“你的百姓若得罪了你，你使天闭塞不下雨；他们若向此处祷告，宣认你的名，因你的惩罚而离开他们的罪，
2CHR|6|27|求你在天上垂听，赦免你仆人你百姓 以色列 的罪，将当行的善道教导他们，并降雨在你的地，就是你赐给你百姓为业之地。
2CHR|6|28|“这地若有饥荒、瘟疫、焚风 、霉烂、蝗虫、蚂蚱，或有仇敌围困这地的城门，无论遭遇什么灾祸疾病，
2CHR|6|29|你的百姓 以色列 ，或众人或一人，自觉灾祸困苦，向这殿举手，无论祈求什么，祷告什么，
2CHR|6|30|求你从天上你的居所垂听赦免。因为你知道人心，惟有你知道世人的心，求你照各人所行的一切待他们，
2CHR|6|31|使他们在你赐给我们列祖的土地上一生一世敬畏你，遵行你的道。
2CHR|6|32|“论到不属你百姓 以色列 的外邦人，若为你的大名和大能的手，以及伸出来的膀臂，从远方而来，来向这殿祷告，
2CHR|6|33|求你从天上你的居所垂听，照着外邦人向你所求的一切而行，使地上万民都认识你的名，敬畏你，像你的百姓 以色列 一样，又使他们知道我所建造的是称为你名下的殿。
2CHR|6|34|“你的百姓若奉你的派遣出去，无论往何处与仇敌争战，他们若向你所选择的这城和我为你名所建造的殿祷告，
2CHR|6|35|求你从天上垂听他们的祷告祈求，为他们伸张正义。
2CHR|6|36|“你的百姓若得罪你，因为没有人不犯罪，你向他们发怒，把他们交在仇敌面前，掳他们的人把他们带到或远或近之地；
2CHR|6|37|他们若在被掳之地那里回心转意，在被掳之地悔改，向你恳求说：‘我们有罪了，我们悖逆了，我们作恶了’；
2CHR|6|38|他们若在被掳之地尽心尽性归向你，又向自己的地，就是你赐给他们列祖的地和你所选择的城，以及我为你名所建造的这殿祷告，
2CHR|6|39|求你从天上你的居所垂听他们的祷告祈求，为他们伸张正义，赦免你的百姓向你犯的罪。
2CHR|6|40|我的上帝啊，现在求你睁眼看，侧耳听在此处所献的祷告。
2CHR|6|41|“耶和华上帝啊，现在求你兴起， 与你有能力的约柜同入安歇之所。 耶和华上帝啊，愿你的祭司披上救恩， 愿你的圣民蒙福欢乐。
2CHR|6|42|耶和华上帝啊，求你不要厌弃你的受膏者， 要记得向你仆人 大卫 所施的慈爱。”
2CHR|7|1|所罗门 祈祷完毕，就有火从天降下来，烧尽燔祭和祭物。耶和华的荣光充满了殿；
2CHR|7|2|因耶和华的荣光充满了耶和华的殿，所以祭司不能进耶和华的殿。
2CHR|7|3|那火降下、耶和华的荣光在殿上的时候， 以色列 众人看见，就在石板地俯伏敬拜，称谢耶和华： “耶和华本为善， 他的慈爱永远长存！”
2CHR|7|4|王和众百姓在耶和华面前献祭。
2CHR|7|5|所罗门 王献二万二千头牛，十二万只羊为祭。这样，王和众百姓为上帝的殿行了奉献之礼。
2CHR|7|6|祭司各供其职侍立， 利未 人拿着耶和华的乐器，就是 大卫 王所造、为要颂赞耶和华的乐器，因他的慈爱永远长存；他们为 大卫 的赞美诗奏乐；祭司在众人面前吹号， 以色列 众人都站立。
2CHR|7|7|所罗门 因他所造的铜坛容不下燔祭、素祭和脂肪，就将耶和华殿前院子的中间分别为圣，在那里献燔祭和平安祭牲的脂肪。
2CHR|7|8|那时 所罗门 守节七日，从 哈马口 直到 埃及 溪谷的 以色列 众人都与他同在一起，成了一个极其盛大的会。
2CHR|7|9|第八日他们举行严肃会，行奉献坛的礼七日，守节七日。
2CHR|7|10|七月二十三日，王差遣百姓回自己的帐棚去；他们为耶和华向 大卫 和 所罗门 ，以及他百姓 以色列 所施的恩惠，心里都欢喜快乐。
2CHR|7|11|所罗门 建完了耶和华的殿和王宫；在耶和华的殿和王宫的工程上，凡他心中所要做的，都顺利做成了。
2CHR|7|12|夜间耶和华向 所罗门 显现，对他说：“我已听了你的祷告，也选择这地方归我作献祭的殿宇。
2CHR|7|13|我若使天闭塞不下雨，或使蝗虫吃这地的出产，或降瘟疫在我子民中，
2CHR|7|14|这称为我名下的子民，若是谦卑自己，祷告，寻求我的面，转离他们的恶行，我必从天上垂听，赦免他们的罪，医治他们的地。
2CHR|7|15|我必睁眼看，侧耳听在此处所献的祷告。
2CHR|7|16|现在我已选择这殿，分别为圣，使我的名永在其中；我的眼、我的心也必时常在那里。
2CHR|7|17|你若行在我面前，效法你父 大卫 所行的，遵行我一切所吩咐你的，谨守我的律例典章，
2CHR|7|18|我就必坚固你国度的王位，正如我与你父 大卫 所立的约，说：‘你的子孙必不断有人治理 以色列 。’
2CHR|7|19|“倘若你们转去，离弃我摆在你们面前的律例诫命，去事奉别神，敬拜它们，
2CHR|7|20|我就必把 以色列 人从我赐给他们的地上连根拔起，也必从我面前舍弃那为我名所分别为圣的殿，使它在万民中成为笑柄，被人讥诮。
2CHR|7|21|这殿虽然崇高，将来凡经过的人必惊讶说：‘耶和华为何向这地和这殿如此行呢？’
2CHR|7|22|人必说：‘因为此地的人离弃领他们祖先出 埃及 地的耶和华－他们的上帝，去亲近别神，敬拜事奉它们，所以耶和华使这一切灾祸临到他们。’”
2CHR|8|1|所罗门 建造耶和华的殿和王宫，用了二十年才完成。
2CHR|8|2|所罗门 修筑 希兰 送给他的城镇，使 以色列 人住在那里。
2CHR|8|3|所罗门 往 哈马．琐巴 去，攻取了那地方。
2CHR|8|4|所罗门 建造旷野的 达莫 ，建造 哈马 一切的储货城，
2CHR|8|5|又建造 上伯．和仑 、 下伯．和仑 ，成为有墙、门、闩的堡垒城。
2CHR|8|6|所罗门 建造 巴拉 和一切的储货城、战车城、战马城，以及他所想要建造的，在 耶路撒冷 、 黎巴嫩 ，和自己所治理全国中的一切建设。
2CHR|8|7|至于所有剩下的百姓，不属 以色列 的 赫 人、 亚摩利 人、 比利洗 人、 希未 人、 耶布斯 人，
2CHR|8|8|那些 以色列 人在当地不能灭尽的人， 所罗门 征召他们剩下的后代服劳役，直到今日。
2CHR|8|9|惟有 以色列 人， 所罗门 不使他们当奴仆做工，而是作他的战士、军官、战车长、骑兵长。
2CHR|8|10|这些是 所罗门 王的监工，共有二百五十名百姓的监工。
2CHR|8|11|所罗门 把法老的女儿迁出 大卫城 ，上到他为她建造的宫里，因 所罗门 说：“耶和华约柜所到之处都是圣地，所以我的妻子不可住在 以色列 王 大卫 的宫里。”
2CHR|8|12|那时， 所罗门 在走廊前他所筑的耶和华的坛上，向耶和华献燔祭，
2CHR|8|13|又遵照 摩西 的吩咐，在安息日、初一，以及每年在除酵节、七七节、住棚节三个节期，献每日所当献上的祭。
2CHR|8|14|所罗门 照着他父亲 大卫 所定的条例，分派祭司的班次，担任他们的职务，又分派 利未 人的任务，负责颂赞，并在祭司面前做每日当做的事，又派门口的守卫按着班次看守各门，因为神人 大卫 是这样吩咐的。
2CHR|8|15|王对众祭司和 利未 人的吩咐，无论是管理库房或任何事务，他们都不违背。
2CHR|8|16|所罗门 所有的工作都准备就绪，从立耶和华殿的根基直到完工的日子。耶和华的殿就完成了。
2CHR|8|17|那时， 所罗门 往 以东 地海岸的 以旬．迦别 和 以禄 去。
2CHR|8|18|希兰 派他的臣仆，把船只和熟悉航海的仆人送到 所罗门 那里。他们同 所罗门 的仆人到了 俄斐 ，从那里得了四百五十他连得金子，运到 所罗门 王那里。
2CHR|9|1|示巴 女王听见 所罗门 的名声，就来到 耶路撒冷 ，要用难题考问 所罗门 。她带着很多的随从，有骆驼驮着香料、许多金子和宝石。她来到 所罗门 那里，向他提出心中所有的问题。
2CHR|9|2|所罗门 回答了她所有的问题，没有一个问题太难，是 所罗门 不能向她解答的。
2CHR|9|3|示巴 女王看见 所罗门 的智慧和他所建造的宫殿，
2CHR|9|4|席上的食物，坐着的群臣，侍立的仆人和他们的服装，司酒长和他们的服装，以及他上耶和华殿的台阶 ，就诧异得神不守舍。
2CHR|9|5|她对王说：“我在本国所听到的话，论到你的事和你的智慧是真的！
2CHR|9|6|我本来不信那些话，及至我来亲眼看见了，看哪，人所告诉我的，还不及你丰富智慧的一半，超过我所听见的传闻。
2CHR|9|7|你的人是有福的！你这些常侍立在你面前、听你智慧话的仆人是有福的！
2CHR|9|8|耶和华－你的上帝是应当称颂的！他喜爱你，使你坐他的王位，为耶和华－你的上帝作王；因为你的上帝爱 以色列 ，要永远坚立它，所以立你作他们的王，使你秉公行义。”
2CHR|9|9|于是 示巴 女王把一百二十他连得金子、极多的香料和宝石送给 所罗门 王；从来没有像 示巴 女王送给 所罗门 王那么多的香料。
2CHR|9|10|希兰 的仆人和 所罗门 的仆人也从 俄斐 运了金子来，又运了檀香木和宝石来。
2CHR|9|11|王用檀香木为耶和华的殿和王宫做阶梯，又为歌唱的人做琴瑟； 犹大 地从来没有见过这样的。
2CHR|9|12|所罗门 王除了回赠 示巴 女王所带来的，凡她所提出的一切要求， 所罗门 王都送给她。于是女王和她臣仆转回，到本国去了。
2CHR|9|13|所罗门 每年所得的金子，重六百六十六他连得，
2CHR|9|14|另外还有从商人和贸易所收到的，以及 阿拉伯 诸王和各地的省长进贡给 所罗门 的金银。
2CHR|9|15|所罗门 王用锤出来的金子打成二百面盾牌，每面盾牌用六百舍客勒锤出来的金子；
2CHR|9|16|又用锤出来的金子打成三百面小盾牌，每面小盾牌用三百舍客勒金子。王把它们放在 黎巴嫩林宫 里。
2CHR|9|17|王又制造一个大的象牙宝座，包上纯金。
2CHR|9|18|宝座有六层台阶，又有金脚凳，与宝座相连。座位之处两旁有扶手，靠近扶手有两只狮子站立。
2CHR|9|19|六层台阶上有十二只狮子站立，分站左边和右边；任何国度都没有这样做的。
2CHR|9|20|所罗门 王一切的饮器都是金的， 黎巴嫩林宫 里所有的器皿都是纯金的。在 所罗门 的日子，银子算不了什么。
2CHR|9|21|因王的船只与 希兰 的仆人一同往 他施 去， 他施 船只每三年一次把金、银、象牙、猿猴、孔雀 运回来。
2CHR|9|22|所罗门 王的财宝与智慧胜过地上的众王。
2CHR|9|23|地上的众王都求见 所罗门 的面，要听上帝放在他心里的智慧。
2CHR|9|24|他们各带贡物，就是银器、金器、衣服、兵器、香料、马、骡子，每年都有一定的数量。
2CHR|9|25|所罗门 拥有给战车和马用的四千个棚子，还有一万二千名骑兵，安置在屯车城，在 耶路撒冷 的王那里。
2CHR|9|26|所罗门 统管诸王，从 大河 到 非利士 人的地，直到 埃及 的边界。
2CHR|9|27|王在 耶路撒冷 使银子多如石头，香柏木多如 谢非拉 的桑树。
2CHR|9|28|有人从 埃及 和各国为 所罗门 把马匹运来。
2CHR|9|29|所罗门 其余的事，自始至终，不都写在 拿单 先知的书上和 示罗 人 亚希雅 的《预言书》上，以及 易多 先见论 尼八 儿子 耶罗波安 的《默示书》上吗？
2CHR|9|30|所罗门 在 耶路撒冷 作全 以色列 的王四十年。
2CHR|9|31|所罗门 与他祖先同睡，葬在他父亲 大卫 的城里，他儿子 罗波安 接续他作王。
2CHR|10|1|罗波安 往 示剑 去，因 以色列 众人都到了 示剑 ，要立他作王。
2CHR|10|2|尼八 的儿子 耶罗波安 先前躲避 所罗门 王，逃往 埃及 ，住在那里；他听见这事，就从 埃及 回来。
2CHR|10|3|以色列 人派人去请他来。 耶罗波安 就和 以色列 众人来，与 罗波安 谈话，说：
2CHR|10|4|“你父亲使我们负重轭，现在求你减轻你父亲所加给我们的苦工和重轭，我们就服事你。”
2CHR|10|5|罗波安 对他们说：“过三天再来见我吧！”百姓就走了。
2CHR|10|6|罗波安 的父亲 所罗门 在世的时候，有侍立在他面前的长者， 罗波安 王和他们商议，说：“你们出个主意，好把话带回给这百姓。”
2CHR|10|7|他们对他说：“王若恩待这百姓，使他们喜悦，跟他们说好话，他们就永远作王的仆人了。”
2CHR|10|8|王不采纳长者给他出的主意，却和那些与他一同长大、在他面前侍立的年轻人商议。
2CHR|10|9|他对他们说：“这百姓对我说：‘你父亲使我们负重轭，求你减轻一些。’你们出个什么主意，我们好把话带回给他们。”
2CHR|10|10|那些与他一同长大的年轻人对他说：“这些百姓对王说：‘你父亲使我们负重轭，求你给我们减轻一些。’王要对他们如此说：‘我的小指头比我父亲的腰还粗呢！
2CHR|10|11|我父亲使你们负重轭，现在我必使你们负更重的轭！我父亲用鞭子惩罚你们，我却要用蝎子！’”
2CHR|10|12|耶罗波安 和众百姓遵照王所说“你们第三天再来见我”的话，第三天来到 罗波安 那里。
2CHR|10|13|王严厉地回答他们。 罗波安 王不采纳长者所出的主意，
2CHR|10|14|却照着年轻人所出的主意对他们说：“我 使你们负重轭，我必使你们负更重的轭！我父亲用鞭子惩罚你们，我却要用蝎子！”
2CHR|10|15|王不依从百姓，因这事件是出于上帝，为要应验耶和华藉 示罗 人 亚希雅 对 尼八 的儿子 耶罗波安 所说的话。
2CHR|10|16|以色列 众人见王不依从他们，百姓就回覆王说： “我们在 大卫 中有什么分呢？ 我们在 耶西 的儿子中没有产业！ 以色列 啊，各回自己的帐棚去吧！ 大卫 啊，现在你顾自己的家吧！” 于是， 以色列 众人都回自己的帐棚去了；
2CHR|10|17|至于住 犹大 城镇的 以色列 人， 罗波安 仍作他们的王。
2CHR|10|18|罗波安 王派监管劳役的 哈多兰 去， 以色列 人用石头打他，他就死了。 罗波安 王急忙上车，逃回 耶路撒冷 去了。
2CHR|10|19|这样， 以色列 背叛 大卫 家，直到今日。
2CHR|11|1|罗波安 来到 耶路撒冷 ，召集 犹大 家和 便雅悯 家，共十八万人，都是精选的战士，要与 以色列 争战，好将国夺回再归自己。
2CHR|11|2|但耶和华的话临到神人 示玛雅 ，说：
2CHR|11|3|“你去告诉 所罗门 的儿子 犹大 王 罗波安 和住 犹大 、 便雅悯 的 以色列 众人，说：
2CHR|11|4|‘耶和华如此说：你们不可上去与你们的弟兄争战。各自回家去吧！因为这事是出于我。’”众人就听从耶和华的话回去，不去与 耶罗波安 争战。
2CHR|11|5|罗波安 住在 耶路撒冷 ，在 犹大 为防御修筑城镇，
2CHR|11|6|他修筑 伯利恒 、 以坦 、 提哥亚 、
2CHR|11|7|伯．夙 、 梭哥 、 亚杜兰 、
2CHR|11|8|迦特 、 玛利沙 、 西弗 、
2CHR|11|9|亚多莱音 、 拉吉 、 亚西加 、
2CHR|11|10|琐拉 、 亚雅仑 、 希伯仑 。这都是 犹大 和 便雅悯 的坚固城。
2CHR|11|11|罗波安 又巩固这些堡垒，在其中安置军官，储备粮食、油和酒。
2CHR|11|12|他在各城里预备盾牌和枪，使城极其坚固。 犹大 和 便雅悯 都归了他。
2CHR|11|13|全 以色列 的祭司和 利未 人都从四方来归 罗波安 。
2CHR|11|14|利未 人放弃他们的郊野和产业，来到 犹大 与 耶路撒冷 ，因为 耶罗波安 和他的儿子拒绝他们，不许他们担任祭司事奉耶和华。
2CHR|11|15|耶罗波安 为丘坛，为山羊鬼魔，为自己所造的牛犊设立祭司。
2CHR|11|16|以色列 各支派中，凡立定心意寻求耶和华－ 以色列 上帝的，都随从 利未 人来到 耶路撒冷 献祭给耶和华－他们列祖的上帝。
2CHR|11|17|这就巩固了 犹大 王国，使 所罗门 的儿子 罗波安 强盛三年，因为这三年他们遵行 大卫 和 所罗门 的道。
2CHR|11|18|罗波安 娶 大卫 儿子 耶利末 的女儿 玛哈拉 为妻，又娶 耶西 儿子 以利押 的女儿 亚比孩 为妻，
2CHR|11|19|从她生了几个儿子，就是 耶乌施 、 示玛利雅 和 撒罕 。
2CHR|11|20|后来他又娶 押沙龙 的女儿 玛迦 ，从她生了 亚比雅 、 亚太 、 细撒 和 示罗密 。
2CHR|11|21|罗波安 有十八个妻和六十个妾，生了二十八个儿子，六十个女儿；他却爱 押沙龙 的女儿 玛迦 ，过于爱其他的妻妾。
2CHR|11|22|罗波安 立 玛迦 的儿子 亚比雅 作太子，在他兄弟中为首，因为要立他作王。
2CHR|11|23|罗波安 办事精明，把他众儿子分散在 犹大 和 便雅悯 全地各坚固城里，赐他们大量的粮食，又给他们娶许多妻子。
2CHR|12|1|罗波安 的王国稳固，他强盛的时候就离弃耶和华的律法，全 以色列 都跟从他。
2CHR|12|2|罗波安 王第五年， 埃及 王 示撒 上来攻打 耶路撒冷 ，因为他们背叛了耶和华。
2CHR|12|3|示撒 带着一千二百辆战车，六万名骑兵，以及跟随他从 埃及 出来的 路比 人、 苏基 人和 古实 人的军队，多得不可胜数。
2CHR|12|4|他攻取了 犹大 的坚固城，来到 耶路撒冷 。
2CHR|12|5|那时， 犹大 的领袖因为 示撒 的缘故聚集在 耶路撒冷 ，有先知 示玛雅 去见 罗波安 和众领袖，对他们说：“耶和华如此说：‘你们离弃了我，所以我也离弃你们，把你们交在 示撒 手里。’”
2CHR|12|6|于是 以色列 的领袖和王都谦卑说：“耶和华是公义的。”
2CHR|12|7|耶和华见他们谦卑，耶和华的话就临到 示玛雅 ，说：“他们既谦卑，我必不灭绝他们；我要使他们暂时得拯救，不藉着 示撒 的手将我的怒气倒在 耶路撒冷 。
2CHR|12|8|然而他们必作 示撒 的仆人，好叫他们知道，服事我与服事地上邦国有何分别。”
2CHR|12|9|于是， 埃及 王 示撒 上来攻取 耶路撒冷 ，夺了耶和华殿和王宫里的宝物，尽都带走，又夺走 所罗门 制造的金盾牌。
2CHR|12|10|罗波安 王制造铜盾牌代替那些金盾牌，交给看守王宫宫门的护卫长看管。
2CHR|12|11|每逢王进耶和华的殿，护卫兵就来，举起这些盾牌；随后仍将盾牌送回护卫室。
2CHR|12|12|王谦卑的时候，耶和华的怒气就转消了，不全然灭尽，并且在 犹大 中，情况也有好转。
2CHR|12|13|罗波安 王自强，在 耶路撒冷 作王。他登基的时候年四十一岁，在 耶路撒冷 ，就是耶和华从 以色列 众支派中所选择立他名的城，作王十七年。 罗波安 的母亲名叫 拿玛 ，是 亚扪 人。
2CHR|12|14|罗波安 行恶，因他没有立定心意寻求耶和华。
2CHR|12|15|罗波安 的事迹，自始至终不都写在 示玛雅 先知和 易多 先见的《史记》上吗？ 罗波安 与 耶罗波安 时常交战。
2CHR|12|16|罗波安 与他祖先同睡，葬在 大卫城 ，他的儿子 亚比雅 接续他作王。
2CHR|13|1|耶罗波安 王十八年， 亚比雅 登基作 犹大 王，
2CHR|13|2|在 耶路撒冷 作王三年。他母亲名叫 米该亚 ，是 基比亚 人 乌列 的女儿 。 亚比雅 常与 耶罗波安 交战。
2CHR|13|3|有一次 亚比雅 率领四十万精选的士兵出战，他们都是勇敢的战士； 耶罗波安 也率领八十万精选的大能勇士，迎着 亚比雅 摆阵。
2CHR|13|4|亚比雅 站在 以法莲 山区中的 洗玛脸山 上，说：“ 耶罗波安 和 以色列 众人哪，要听我说！
2CHR|13|5|耶和华－ 以色列 的上帝曾立盐约，将 以色列 国永远赐给 大卫 和他的子孙，你们不知道吗？
2CHR|13|6|但 大卫 儿子 所罗门 的臣仆、 尼八 的儿子 耶罗波安 起来背叛他的主人。
2CHR|13|7|有些无赖的歹徒聚集跟从他，逞强攻击 所罗门 的儿子 罗波安 ；那时 罗波安 还年轻，心志软弱，不能抵挡他们。
2CHR|13|8|“现在你们说要抗拒 大卫 子孙手下所治理的耶和华的国，你们的人数众多，你们那里又有 耶罗波安 为你们所造当作神明的金牛犊。
2CHR|13|9|你们不是驱逐耶和华的祭司 亚伦 的后裔和 利未 人吗？不是照着外邦人的恶俗为自己立祭司吗？无论何人牵一头公牛犊、七只公绵羊将自己分别出来，就可作虚无神明的祭司。
2CHR|13|10|至于我们，耶和华是我们的上帝，我们并没有离弃他。我们有事奉耶和华的祭司，都是 亚伦 的后裔，并有 利未 人各尽其职。
2CHR|13|11|他们每日早晚向耶和华献燔祭，烧芬芳的香，又在纯金的 供桌上摆供饼，每晚点燃金灯台上的灯盏，因为我们遵守耶和华－我们上帝的命令，但你们却离弃了他。
2CHR|13|12|看哪，率领我们的是上帝，又有他的祭司拿号向你们吹出响声。 以色列 人哪，不要与耶和华－你们列祖的上帝争战，因你们必不能得胜。”
2CHR|13|13|耶罗波安 却在 犹大 人的后头设伏兵。这样， 以色列 人在 犹大 人的前头，伏兵在 犹大 人的后头。
2CHR|13|14|犹大 人转过来，看哪，前后都有战事，就呼求耶和华，祭司也吹号。
2CHR|13|15|于是 犹大 人呐喊。 犹大 人呐喊的时候，上帝就击打 耶罗波安 和 以色列 众人，使他们败在 亚比雅 与 犹大 人面前。
2CHR|13|16|以色列 人在 犹大 人面前逃跑，上帝将他们交在 犹大 人手里。
2CHR|13|17|亚比雅 和他的军兵大大击杀 以色列 人， 以色列 人被杀仆倒的精兵有五十万。
2CHR|13|18|那时， 以色列 人被制伏了。 犹大 人得胜，因为他们倚靠耶和华－他们列祖的上帝。
2CHR|13|19|亚比雅 追赶 耶罗波安 ，攻取了他的几座城，就是 伯特利 和所属的乡镇 ， 耶沙拿 和所属的乡镇， 以法拉音 和所属的乡镇。
2CHR|13|20|亚比雅 在世的时候， 耶罗波安 不再强盛；耶和华击打他，他就死了。
2CHR|13|21|亚比雅 却渐渐强盛。他娶了十四个妻妾，生了二十二个儿子，十六个女儿。
2CHR|13|22|亚比雅 其余的事和他的言行都写在 易多 先知的评传上。
2CHR|14|1|亚比雅 与他祖先同睡，葬在 大卫城 ，他的儿子 亚撒 接续他作王。 亚撒 在位期间，国中太平十年。
2CHR|14|2|亚撒 行耶和华－他上帝眼中看为善为正的事，
2CHR|14|3|除掉外邦的祭坛和丘坛，打碎柱像，砍下 亚舍拉 ，
2CHR|14|4|吩咐 犹大 人寻求耶和华－他们列祖的上帝，遵行他的律法和诫命，
2CHR|14|5|又在 犹大 各城镇除掉丘坛和香坛。在他治理下，国中太平。
2CHR|14|6|他在 犹大 建造了几座坚固城。那些年间，国中太平，没有战争，因为耶和华赐他平安。
2CHR|14|7|他对 犹大 人说：“我们要建造这些城镇，四围筑墙，盖城楼，安门，做闩；地仍属于我们，因为我们寻求耶和华－我们的上帝；我们寻求他，他就赐我们四境平安。”于是他们建造城镇，诸事亨通。
2CHR|14|8|亚撒 的军兵，出自 犹大 拿盾牌拿枪的三十万人，出自 便雅悯 拿小盾牌拉弓的二十八万人；这些全都是大能的勇士。
2CHR|14|9|古实 人 谢拉 率领一百万军兵，三百辆战车，出来攻击 犹大 人，到了 玛利沙 。
2CHR|14|10|亚撒 出去迎战，在 玛利沙 的 洗法谷 彼此摆阵。
2CHR|14|11|亚撒 呼求耶和华－他的上帝说：“耶和华啊，在强弱之间，惟有你能帮助。耶和华－我们的上帝啊，求你帮助我们，因为我们仰赖你，奉你的名来抵挡这大军。耶和华啊，你是我们的上帝，不要让人胜过你。”
2CHR|14|12|于是耶和华击打 古实 人，使他们败在 亚撒 和 犹大 人面前， 古实 人就逃跑了。
2CHR|14|13|亚撒 和跟随他的军兵追赶他们，直到 基拉耳 。 古实 人被杀的很多，无法复原，因为他们在耶和华与他军兵面前被击溃。 犹大 人夺了许多财物，
2CHR|14|14|又攻打 基拉耳 四围一切的城镇；城中的人都惧怕耶和华。 犹大 人掳掠了一切的城镇，因其中的财物很多，
2CHR|14|15|又毁坏了群畜的圈，夺取许多的羊和骆驼，就回 耶路撒冷 去了。
2CHR|15|1|上帝的灵临到 俄德 的儿子 亚撒利雅 。
2CHR|15|2|他出来迎接 亚撒 ，对他说：“ 亚撒 ， 犹大 和 便雅悯 众人哪，要听我说：你们若顺从耶和华，耶和华必与你们同在；你们若寻求他，就必寻见；你们若离弃他，他必离弃你们。
2CHR|15|3|以色列 人不信真神，没有训诲的祭司，也没有律法，已经许多日子了。
2CHR|15|4|但他们在急难的时候归向耶和华－ 以色列 的上帝，寻求他，他就被他们寻见。
2CHR|15|5|那时，出入的人不得平安，各地的居民都遭大乱；
2CHR|15|6|他们被破坏殆尽，这国攻击那国，这城攻击那城，因为上帝用各样灾难扰乱他们。
2CHR|15|7|现在你们要刚强，不要手软，因你们所行的必得赏赐。”
2CHR|15|8|亚撒 听见这些话和 俄德 先知的预言，就壮起胆来，在 犹大 和 便雅悯 全地，以及 以法莲 山区所夺的各城，把其中的可憎之物尽都除掉，又在耶和华殿的走廊前重新修筑耶和华的坛。
2CHR|15|9|他又召集 犹大 和 便雅悯 众人，以及他们中间寄居的 以法莲 人、 玛拿西 人、 西缅 人。有许多 以色列 人归顺 亚撒 ，因为他们看见耶和华－他的上帝与他同在。
2CHR|15|10|亚撒 作王第十五年三月，他们都聚集在 耶路撒冷 。
2CHR|15|11|那日他们从所取的掳物中，将七百头牛和七千只羊献给耶和华。
2CHR|15|12|他们立约，要尽心尽性寻求耶和华－他们列祖的上帝。
2CHR|15|13|凡不寻求耶和华－ 以色列 上帝的，无论大小、男女，必被处死。
2CHR|15|14|他们就大声欢呼，吹号吹角，向耶和华起誓。
2CHR|15|15|犹大 众人为所起的誓欢喜，因他们尽心起誓，尽意寻求耶和华，耶和华就被他们寻见，且赐他们四境平安。
2CHR|15|16|亚撒 王甚至废了他祖母 玛迦 太后的位，因 玛迦 造了可憎的 亚舍拉 。 亚撒 砍下她的偶像，捣得粉碎，在 汲沦溪 边烧了，
2CHR|15|17|只是丘坛还没有从 以色列 中废去，然而 亚撒 一生有纯正的心。
2CHR|15|18|亚撒 将他父亲所分别为圣与自己所分别为圣的金银和器皿都奉到上帝的殿里。
2CHR|15|19|亚撒 作王直到第三十五年，都没有战事。
2CHR|16|1|亚撒 作王第三十六年， 以色列 王 巴沙 上来攻击 犹大 ，修筑 拉玛 ，不许人从 犹大 王 亚撒 那里出入。
2CHR|16|2|于是 亚撒 从耶和华殿和王宫的府库里拿出金银来，送给住在 大马士革 的 亚兰 王 便．哈达 ，说：
2CHR|16|3|“你父曾与我父立约，我与你也要这样立约。看哪，我把金银送给你，请你废掉你与 以色列 王 巴沙 所立的约，使他从我这里撤退。”
2CHR|16|4|便．哈达 听从了 亚撒 王，就派遣他的军官去攻打 以色列 的城镇。他们攻下了 以云 、 但 、 亚伯．玛音 和 拿弗他利 一切的储货城。
2CHR|16|5|巴沙 听见了，就停工不修筑 拉玛 ，任由他的工程停止。
2CHR|16|6|于是 亚撒 王率领 犹大 众人，运走 巴沙 修筑 拉玛 所用的石头和木料，用以修筑 迦巴 和 米斯巴 。
2CHR|16|7|那时， 哈拿尼 先见来见 犹大 王 亚撒 ，对他说：“因你仰赖 亚兰 王，没有仰赖耶和华－你的上帝，所以 亚兰 王的军兵逃脱了你的手。
2CHR|16|8|古实 人和 路比 人的军队不是非常强大吗？他们的战车骑兵不是极多吗？只因你仰赖耶和华，他就将他们交在你手里。
2CHR|16|9|因为耶和华的眼目遍察全地，要坚固向他存纯正之心的人。你在这事上行得愚昧；因此，以后你必有战争。”
2CHR|16|10|亚撒 恼恨先见，为了这事向他发怒，将他囚在监里。那时 亚撒 也虐待一些百姓。
2CHR|16|11|亚撒 自始至终的事迹，看哪，都写在《犹大和以色列诸王记》上。
2CHR|16|12|亚撒 作王三十九年的时候患了脚疾，非常严重。他生病的时候没有求耶和华，只求医生。
2CHR|16|13|他作王四十一年死了，与他祖先同睡，
2CHR|16|14|葬在 大卫城 自己所凿的坟墓里。人把他放在床上，床上堆满各样馨香的香料，就是按做香的作法调和的香料，又为他生一堆大火志哀。
2CHR|17|1|亚撒 的儿子 约沙法 接续他作王，奋勇自强，防备 以色列 。
2CHR|17|2|他安置军兵在 犹大 一切坚固城里，又安置驻军在 犹大 地和他父亲 亚撒 所得 以法莲 的城镇中。
2CHR|17|3|耶和华与 约沙法 同在，因为他行他祖先 大卫 从前所行的道，不去寻求诸 巴力 ，
2CHR|17|4|只寻求他父亲的上帝，遵行他的诫命，不效法 以色列 人的行为。
2CHR|17|5|所以耶和华坚定 约沙法 手中的国， 犹大 众人给他进贡； 约沙法 大有财富和尊荣。
2CHR|17|6|他乐意遵行耶和华的道，并且从 犹大 再次除掉一切丘坛和 亚舍拉 。
2CHR|17|7|他作王第三年，差遣官员 便．亥伊勒 、 俄巴底 、 撒迦利雅 、 拿坦业 、 米该亚 往 犹大 各城去教导百姓。
2CHR|17|8|跟他们一同去的有 利未 人 示玛雅 、 尼探雅 、 西巴第雅 、 亚撒黑 、 示米拉末 、 约拿单 、 亚多尼雅 、 多比雅 、 驼．巴多尼雅 ；跟他们一同的又有 以利沙玛 和 约兰 二位祭司。
2CHR|17|9|他们在 犹大 教导，带着耶和华的律法书，走遍 犹大 各城教导百姓。
2CHR|17|10|犹大 四围地上的邦国都惧怕耶和华，不敢与 约沙法 争战。
2CHR|17|11|有些 非利士 人送礼物，进贡银子给 约沙法 。 阿拉伯 人也送他七千七百只公绵羊，七千七百只公山羊。
2CHR|17|12|约沙法 日渐强大，他在 犹大 建造堡垒和储货城。
2CHR|17|13|他在 犹大 城镇中有许多工程，在 耶路撒冷 又有战士，就是大能的勇士。
2CHR|17|14|他们按着父家的数目如下： 犹大 族的千夫长以 押拿 为首，率领三十万大能的勇士；
2CHR|17|15|其次是 约哈难 千夫长，率领二十八万；
2CHR|17|16|其次是 细基利 的儿子 亚玛斯雅 ，他是一个自愿奉献给耶和华的人，率领二十万大能的勇士。
2CHR|17|17|便雅悯 族有大能的勇士 以利雅大 ，率领二十万拿弓箭和盾牌的人；
2CHR|17|18|其次是 约萨拔 ，率领十八万预备打仗的人。
2CHR|17|19|这些都是伺候王的，还有王在全 犹大 的坚固城所安置的不在其内。
2CHR|18|1|约沙法 大有财富和尊荣，他与 亚哈 结亲。
2CHR|18|2|过了几年，他下到 撒玛利亚 去见 亚哈 ； 亚哈 为他和跟从他的人宰了许多牛羊，劝他一同上去攻打 基列 的 拉末 。
2CHR|18|3|以色列 王 亚哈 问 犹大 王 约沙法 说：“你肯同我去攻打 基列 的 拉末 吗？”他回答说：“你我不分彼此，我的军队就是你的军队，我们必与你一同去争战。”
2CHR|18|4|约沙法 对 以色列 王说：“请你先求问耶和华的话。”
2CHR|18|5|于是 以色列 王召集先知四百人，问他们说：“我可以上去攻打 基列 的 拉末 吗？还是不要上去呢？”他们说：“可以上去，因为上帝必将那城交在王的手里。”
2CHR|18|6|约沙法 说：“这里还有没有耶和华的先知，我们好求问他呢？”
2CHR|18|7|以色列 王对 约沙法 说：“还有一个人，是 音拉 的儿子 米该雅 ，我们可以托他求问耶和华。只是我真的很恨他，因为他对我说预言，从不说吉言，总是说凶信。” 约沙法 说：“请王不要这么说。”
2CHR|18|8|以色列 王就召了一个官员来，说：“你快去，把 音拉 的儿子 米该雅 召来。”
2CHR|18|9|以色列 王和 犹大 王 约沙法 在 撒玛利亚 城门前的禾场，各穿朝服，坐在宝座上，所有的先知都在他们面前说预言。
2CHR|18|10|基拿拿 的儿子 西底家 为自己造了铁角，说：“耶和华如此说：‘你要用这些角抵触 亚兰 人，直到将他们灭尽。’”
2CHR|18|11|所有的先知也都这样预言说：“可以上 基列 的 拉末 去，必然得胜，因为耶和华必将那城交在王的手中。”
2CHR|18|12|那去召 米该雅 的使者对他说：“看哪，众先知都异口同声向王说吉言，你也跟他们说一样的话，说吉言吧！”
2CHR|18|13|米该雅 说：“我指着永生的耶和华起誓，我的上帝说什么，我就说什么。”
2CHR|18|14|米该雅 来到王那里，王问他：“ 米该雅 啊，我们可以上去攻打 基列 的 拉末 吗？还是不要上去呢？”他说：“可以上去，必然得胜，敌人必交在你们手里。”
2CHR|18|15|王对他说：“我要你发誓多少次，你才会奉耶和华的名向我说实话呢？”
2CHR|18|16|米该雅 说：“我看见 以色列 众人散布在山上，如同没有牧人的羊群一般。耶和华说：‘这些人没有主人，他们可以平安地各自回家去。’”
2CHR|18|17|以色列 王对 约沙法 说：“我岂没有告诉你，这人对我说预言，从不说吉言，只说凶信吗？”
2CHR|18|18|米该雅 说：“因此你们要听耶和华的话！我看见耶和华坐在宝座上，天上的万军侍立在他左右。
2CHR|18|19|耶和华 说：‘谁去引诱 以色列 王 亚哈 上 基列 的 拉末 去阵亡呢？’这个这样说，那个那样说。
2CHR|18|20|随后有一个灵出来，站在耶和华面前，说：‘我去引诱他。’耶和华问他：‘用什么方法呢？’
2CHR|18|21|他说：‘我要出去，在他众先知的口中成为谎言的灵。’耶和华说：‘这样，你去引诱他，必能成功。你出去，照样做吧！’
2CHR|18|22|现在，看哪，耶和华使谎言的灵入了你的这些先知的口，并且耶和华已经宣告要降祸于你。”
2CHR|18|23|基拿拿 的儿子 西底家 前来打 米该雅 一巴掌，说：“耶和华的灵从哪里离开我向你说话呢？”
2CHR|18|24|米该雅 说：“看哪，你进入严密的内室躲藏的那日，就必看见。”
2CHR|18|25|以色列 王说：“把 米该雅 带走，交回给 亚们 市长和 约阿施 王子。
2CHR|18|26|你们要说：‘王如此说：把这个人关在监狱里，使他受苦，吃不饱喝不足，直等到我平安回来。’”
2CHR|18|27|米该雅 说：“你若真的能平安回来，那就是耶和华没有藉我说话了。”他又说：“众百姓啊，你们都要听！”
2CHR|18|28|以色列 王和 犹大 王 约沙法 上 基列 的 拉末 去。
2CHR|18|29|以色列 王对 约沙法 说：“我要改装上阵，你可以仍穿王服。”于是 以色列 王改装，他们上阵去了。
2CHR|18|30|亚兰 王吩咐他的战车长说：“你们不要与他们的大将或小兵交战，只要单单攻击 以色列 王。”
2CHR|18|31|那些战车长看见 约沙法 就说：“这一定是 以色列 王！”他们转过去与他交战。 约沙法 一呼喊，耶和华就帮助他，上帝使他们转离他。
2CHR|18|32|战车长见他不是 以色列 王，就转身不追他了。
2CHR|18|33|有一人开弓，并不知情，箭恰巧射入 以色列 王铠甲的缝里。王对驾车的说：“我受重伤了，你掉过车来，载我离开战场！”
2CHR|18|34|那日，战况越来越猛， 以色列 王勉强站在战车上，面对 亚兰 人，直到傍晚。日落的时候，王就死了。
2CHR|19|1|犹大 王 约沙法 平安回 耶路撒冷 ，到自己的宫里。
2CHR|19|2|哈拿尼 的儿子 耶户 先见出来迎接 约沙法 王，对他说：“你怎么可以帮助恶人，爱那恨耶和华的人呢？因此耶和华的愤怒临到你了。
2CHR|19|3|然而你还有善行，因你从国中除掉 亚舍拉 ，立定心意寻求上帝。”
2CHR|19|4|约沙法 住在 耶路撒冷 ，以后又出巡民间，从 别是巴 直到 以法莲 山区，引导百姓归向耶和华－他们列祖的上帝。
2CHR|19|5|他在国中，在 犹大 一切坚固城设立审判官，各城都是如此。
2CHR|19|6|他对审判官说：“你们应当谨慎所做的事，因为你们审判不是为人，而是为耶和华。在审判的事上，他必与你们同在。
2CHR|19|7|现在，你们应当敬畏耶和华，谨慎办事，因为耶和华－我们的上帝没有不义，不看人的情面，也不受贿赂。”
2CHR|19|8|约沙法 从 利未 人和祭司，以及 以色列 族长中，也委派人在 耶路撒冷 为耶和华施行审判，为 耶路撒冷 的居民听讼断案 。
2CHR|19|9|约沙法 吩咐他们说：“你们当这样，以敬畏耶和华、诚实和纯正的心办事。
2CHR|19|10|你们住在各城的弟兄，若有争讼的案件呈到你们这里，或为流血，或犯律法、诫命、律例、典章，你们要警戒他们，免得他们得罪耶和华，以致愤怒临到你们和你们的弟兄；你们当这样行，就没有罪了。
2CHR|19|11|看哪，凡属耶和华的事，有 亚玛利雅 祭司长管理你们；凡属王的事，有 犹大 家的领袖 以实玛利 的儿子 西巴第雅 管理你们；在你们面前有 利未 人作官长。你们应当壮胆办事，愿耶和华与善人同在。”
2CHR|20|1|此后， 摩押 人和 亚扪 人，连同一些 米乌尼 人 来攻击 约沙法 。
2CHR|20|2|有人来报告 约沙法 说：“从海的那边， 以东 有大军来攻击你，看哪，他们在 哈洗逊．他玛 ，就是 隐．基底 。”
2CHR|20|3|约沙法 惧怕，就定意寻求耶和华，在全 犹大 宣告禁食。
2CHR|20|4|于是 犹大 人聚集，求耶和华帮助，甚至他们从 犹大 各城前来寻求耶和华。
2CHR|20|5|约沙法 站在 犹大 和 耶路撒冷 的会众中，在耶和华殿新的院子前，
2CHR|20|6|说：“耶和华－我们列祖的上帝啊，你不是天上的上帝吗？你不是万邦万国的主宰吗？在你手中有大能大力，无人能抵挡你。
2CHR|20|7|我们的上帝啊，你不是曾在你百姓 以色列 面前驱逐这地的居民，将这地赐给你朋友 亚伯拉罕 的后裔永远为业吗？
2CHR|20|8|他们住在这地，又为你的名建造圣所，说：
2CHR|20|9|‘若有祸患临到我们，或刀兵的惩罚，或瘟疫饥荒，我们在急难的时候，站在这殿前向你呼求，你必垂听并且拯救，因为你的名在这殿里。’
2CHR|20|10|现在，看哪， 以色列 人出 埃及 地的时候，你不容许 以色列 人侵犯 亚扪 人、 摩押 人和 西珥山 人， 以色列 人就离开他们，不灭绝他们。
2CHR|20|11|看哪，他们这样回报我们，要来驱逐我们离开你赐给我们为业之地。
2CHR|20|12|我们的上帝啊，你不惩罚他们吗？因为我们无力抵挡这来攻击我们的大军。我们不知道该怎么做，我们的眼目单仰望你。”
2CHR|20|13|犹大 众人和他们的孩童、妻子、儿女都站在耶和华面前。
2CHR|20|14|那时，耶和华的灵在会众中临到 利未 人 亚萨 的后裔 雅哈悉 ，他是 玛探雅 的玄孙， 耶利 的曾孙， 比拿雅 的孙子， 撒迦利雅 的儿子。
2CHR|20|15|他说：“ 犹大 众人、 耶路撒冷 的居民和 约沙法 王啊，你们要留心听，耶和华对你们如此说：‘不要因这大军恐惧惊惶，因为胜败不在乎你们，而是在乎上帝。
2CHR|20|16|明日你们要下去迎敌；看哪，他们从 洗斯坡 上来，你们必在 耶鲁伊勒 旷野前的谷口遇见他们。
2CHR|20|17|犹大 和 耶路撒冷 人哪，这次你们不要争战，要摆阵站着，看耶和华为你们施行拯救。不要恐惧，也不要惊惶。明日当出去迎敌，因为耶和华与你们同在。’”
2CHR|20|18|约沙法 屈身，脸伏于地， 犹大 众人和 耶路撒冷 的居民也俯伏在耶和华面前，敬拜耶和华。
2CHR|20|19|哥辖 子孙和 可拉 子孙的 利未 人都起来，用极大的声音赞美耶和华－ 以色列 的上帝。
2CHR|20|20|清晨，众人早起往 提哥亚 的旷野去。出去的时候， 约沙法 站着说：“ 犹大 人和 耶路撒冷 的居民哪，要听我说：信靠耶和华－你们的上帝就必站立得稳；信赖他的先知就必亨通。”
2CHR|20|21|约沙法 与百姓商议，就设立歌唱的人，颂赞耶和华，使他们穿上圣洁的礼服，走在军队前赞美耶和华： “当称谢耶和华， 因他的慈爱永远长存！”
2CHR|20|22|他们开始唱歌赞美的时候，耶和华派伏兵击杀那来攻击 犹大 的 亚扪 人、 摩押 人和 西珥山 人，他们就被打败了。
2CHR|20|23|亚扪 人和 摩押 人起来，击杀住 西珥山 的人，把他们灭尽；灭尽住 西珥山 的人之后，他们又彼此自相击杀。
2CHR|20|24|犹大 人来到旷野的了望楼，向那大军观看，看哪，遍地都是尸体，没有一个逃脱的。
2CHR|20|25|约沙法 和他的百姓就来收取掠物，找到许多牲畜 、财物、衣服 和珍宝。他们取掠物归为己有，直到无法携带；因为掠物太多，他们足足收取了三日。
2CHR|20|26|第四日，众人聚集在 比拉迦谷 ，在那里称颂耶和华；因此那地方名叫 比拉迦谷 ，直到今日。
2CHR|20|27|在 约沙法 率领下， 犹大 人和 耶路撒冷 人都欢欢喜喜地回 耶路撒冷 ，耶和华使他们因战胜仇敌而喜乐。
2CHR|20|28|他们弹琴、鼓瑟、吹号来到 耶路撒冷 ，进了耶和华的殿。
2CHR|20|29|地上所有的邦国听见耶和华打败 以色列 的仇敌，就都惧怕上帝。
2CHR|20|30|这样， 约沙法 的国得享太平，因为上帝赐他四境平安。
2CHR|20|31|约沙法 作 犹大 王，登基的时候年三十五岁，在 耶路撒冷 作王二十五年。他母亲名叫 阿苏巴 ，是 示利希 的女儿。
2CHR|20|32|约沙法 效法他父亲 亚撒 所行的道，不偏离左右，行耶和华眼中看为正的事。
2CHR|20|33|只是丘坛还没有废去，百姓也没有立定心意归向他们列祖的上帝。
2CHR|20|34|约沙法 其余的事，看哪，自始至终都写在 哈拿尼 的儿子 耶户 的书上，这些事也记载在《以色列诸王记》上。
2CHR|20|35|此后， 犹大 王 约沙法 与 以色列 王 亚哈谢 结盟； 亚哈谢 多行恶事。
2CHR|20|36|他们合伙造船要往 他施 去，就在 以旬．迦别 造船。
2CHR|20|37|玛利沙 人 多大瓦 的儿子 以利以谢 向 约沙法 预言说：“因你与 亚哈谢 结盟，耶和华必破坏你所造的。”后来那些船果然毁坏，不能往 他施 去了。
2CHR|21|1|约沙法 与他祖先同睡，与他祖先同葬在 大卫城 ，他的儿子 约兰 接续他作王。
2CHR|21|2|约兰 有几个兄弟，就是 约沙法 的儿子 亚撒利雅 、 耶歇 、 撒迦利雅 、 亚撒列夫 、 米迦勒 、 示法提雅 ；这些都是 以色列 王 约沙法 的儿子。
2CHR|21|3|他们的父亲把许多礼物，金银财宝和 犹大 的坚固城赐给他们，却把国赐给 约兰 ，因为他是长子。
2CHR|21|4|约兰 起来治理他父亲的国，奋勇自强，用刀杀了他所有的兄弟和 以色列 的几个领袖。
2CHR|21|5|约兰 登基的时候年三十二岁，在 耶路撒冷 作王八年。
2CHR|21|6|他行 以色列 诸王的道，正如 亚哈 家所行的，因他娶了 亚哈 的女儿为妻，行耶和华眼中看为恶的事。
2CHR|21|7|耶和华却因自己与 大卫 所立的约，不肯灭绝 大卫 的家，要照他所应许的，永远赐灯光给 大卫 和他的子孙。
2CHR|21|8|约兰 在位期间， 以东 背叛，自己立王治理他们，脱离 犹大 的权势。
2CHR|21|9|约兰 就率领他的军官和所有的战车过去。他夜间起来，攻打围困他的 以东 人和战车长。
2CHR|21|10|这样， 以东 背叛，脱离 犹大 的权势，直到今日。那时， 立拿 也背叛了，脱离它的权势，因为 约兰 离弃耶和华－他列祖的上帝。
2CHR|21|11|他又在 犹大 山岭 建造丘坛，使 耶路撒冷 的居民行淫，诱惑 犹大 。
2CHR|21|12|以利亚 先知写信给 约兰 说：“耶和华－你祖先 大卫 的上帝如此说：‘因为你不行你父 约沙法 和 犹大 王 亚撒 的道，
2CHR|21|13|反而行 以色列 诸王的道，使 犹大 和 耶路撒冷 居民行淫，像 亚哈 家行淫一样，又杀了你父家比你好的那些兄弟。
2CHR|21|14|看哪，耶和华必降大灾于你的百姓和你的妻妾、儿女，以及你一切所有的。
2CHR|21|15|至于你，你必患许多的病 ，你的肠子也必生许多的病，日渐沉重，直到肠子坠落下来。’”
2CHR|21|16|耶和华激发 非利士 人和靠近 古实 人的 阿拉伯 人的心来攻击 约兰 。
2CHR|21|17|他们上来攻击 犹大 ，侵入境内，掳掠了王宫里所有的财物和他的妻妾、儿女，除了他的小儿子 约哈斯 之外，没有留下一个儿子。
2CHR|21|18|这一切事以后，耶和华击打 约兰 ，使他的肠子患不能医治的病。
2CHR|21|19|这病缠绵日久，过了二年，肠子坠落下来，他就病重而死。他的百姓没有为他生火志哀，像从前为他祖先生火一样。
2CHR|21|20|约兰 登基的时候年三十二岁，在 耶路撒冷 作王八年。他逝世无人思慕，众人把他葬在 大卫城 ，只是不在列王的坟墓里。
2CHR|22|1|耶路撒冷 的居民立 约兰 的小儿子 亚哈谢 接续他作王，因为跟随 阿拉伯 人来攻营的军兵把 亚哈谢 所有的兄长都杀了； 犹大 王 约兰 的儿子 亚哈谢 就作了王。
2CHR|22|2|亚哈谢 登基的时候年四十二岁 ，在 耶路撒冷 作王一年。他母亲名叫 亚她利雅 ，是 暗利 的孙女。
2CHR|22|3|亚哈谢 也行 亚哈 家的道，因为他母亲给他主谋，使他行恶。
2CHR|22|4|他行耶和华眼中看为恶的事，像 亚哈 家一样；因他父亲死后，他们给他主谋，使他败坏。
2CHR|22|5|他也听从他们的计谋，与 以色列 王 亚哈 的儿子 约兰 同往 基列 的 拉末 去，与 亚兰 王 哈薛 交战。 亚兰 人打伤了 约兰 ，
2CHR|22|6|他回到 耶斯列 ，医治在 拉末 与 亚兰 王 哈薛 打仗时被击打所受的伤。 约兰 的儿子 犹大 王 亚哈谢 因为 亚哈 的儿子 约兰 病了，就下到 耶斯列 看望他。
2CHR|22|7|亚哈谢 去见 约兰 而遇害，这是出乎上帝；因为他一到就同 约兰 出去攻击 宁示 的孙子 耶户 ；这 耶户 是耶和华所膏，使他剪除 亚哈 家的。
2CHR|22|8|耶户 向 亚哈 家施行惩罚的时候，遇见 犹大 的众领袖和 亚哈谢 的侄子们正服事 亚哈谢 ，就把他们都杀了。
2CHR|22|9|亚哈谢 躲在 撒玛利亚 ， 耶户 寻找他，众人把他拿住，送到 耶户 那里，就杀了他。他们把他埋葬，因他们说，他是那尽心寻求耶和华之 约沙法 的儿子。这样， 亚哈谢 的家无力保住国权。
2CHR|22|10|亚哈谢 的母亲 亚她利雅 见她儿子死了，就起来剿灭 犹大 王室所有的后裔。
2CHR|22|11|但王的女儿 约示巴 将 亚哈谢 的儿子 约阿施 从那被杀的王子中偷出来，把他和他的奶妈藏在卧房里。 约示巴 是 约兰 王的女儿， 亚哈谢 的妹妹，祭司 耶何耶大 的妻子。她藏了 约阿施 ，躲避 亚她利雅 ，免受杀害。
2CHR|22|12|亚她利雅 治理这地的时候， 约阿施 和他们一同在上帝殿里藏了六年。
2CHR|23|1|第七年， 耶何耶大 奋勇自强，叫了 耶罗罕 的儿子 亚撒利雅 、 约哈难 的儿子 以实玛利 、 俄备得 的儿子 亚撒利雅 、 亚大雅 的儿子 玛西雅 ，和 细基利 的儿子 以利沙法 等众百夫长，与他们立约。
2CHR|23|2|他们走遍 犹大 ，从 犹大 各城召集 利未 人和 以色列 的众族长到 耶路撒冷 来。
2CHR|23|3|全会众在上帝殿里与王立约。 耶何耶大 对他们说：“看哪，王的儿子必作王，正如耶和华指着 大卫 子孙所应许的。
2CHR|23|4|你们要这样做：在安息日值班的祭司和 利未 人，三分之一要把守各门，
2CHR|23|5|三分之一要在王宫，三分之一要在 根基门 ；众百姓都要在耶和华殿的院内。
2CHR|23|6|除了祭司和供职的 利未 人之外，不准别人进耶和华的殿；只有他们可以进去，因为他们是神圣的。众百姓都要遵守耶和华所吩咐的。
2CHR|23|7|利未 人要手中各拿兵器，四围保护王；凡擅自进殿的，要被处死。王出入的时候，你们当跟随他。”
2CHR|23|8|利未 人和 犹大 众人都照着 耶何耶大 祭司一切所吩咐的去做，各带自己的人，无论安息日值班或不值班的都来，因为 耶何耶大 祭司不许他们下班。
2CHR|23|9|耶何耶大 祭司就把上帝殿里所藏 大卫 王的枪和大小盾牌交给百夫长，
2CHR|23|10|又分派众百姓手中各拿兵器，在祭坛和殿那里，从殿南到殿北，站在王的四围；
2CHR|23|11|他们领 约阿施 出来，给他戴上冠冕，把律法书交给他，立他作王。 耶何耶大 和他的儿子们膏他，他们说：“愿王万岁！”
2CHR|23|12|亚她利雅 听见百姓奔走赞美王的声音，就进耶和华的殿，到百姓那里。
2CHR|23|13|她观看，看哪，王站在殿门的柱旁，百夫长和号手在王旁边，国中的众百姓都欢乐吹号，又有歌唱的人用乐器领人歌唱赞美。 亚她利雅 就撕裂衣服，喊着说：“反了！反了！”
2CHR|23|14|耶何耶大 祭司带领管军兵的百夫长出来，对他们说：“把她从行列之间赶出去，凡跟随她的必用刀杀死！”因为祭司说：“不可在耶和华殿里杀她。”
2CHR|23|15|他们就下手拿住她；她进入通往王宫的 马门 ，他们就在那里把她杀了。
2CHR|23|16|耶何耶大 与众百姓，又与王立约，要作耶和华的子民。
2CHR|23|17|于是众百姓到 巴力 庙去，拆毁了庙，打碎祭坛和偶像，又在坛前把 巴力 的祭司 玛坦 杀了。
2CHR|23|18|耶何耶大 派官员在 利未 家的祭司手下看守耶和华的殿，他们是 大卫 所分派的，在耶和华殿中照 摩西 律法上所写，献燔祭给耶和华，又按 大卫 所定的，欢乐歌唱。
2CHR|23|19|耶何耶大 又设立守卫把守耶和华殿的各门，无论因何事而不洁净的人，都不准进去。
2CHR|23|20|他又率领百夫长和贵族，与民间的官长，以及国中的众百姓，请王从耶和华的殿下来，由 上门 正中进入王宫，使王坐在国度的王位上。
2CHR|23|21|国中的众百姓都欢乐，合城也都平静。他们已将 亚她利雅 用刀杀了。
2CHR|24|1|约阿施 登基的时候年方七岁，在 耶路撒冷 作王四十年。他母亲名叫 西比亚 ，是 别是巴 人。
2CHR|24|2|耶何耶大 祭司在世的日子， 约阿施 行耶和华眼中看为正的事。
2CHR|24|3|耶何耶大 为他娶了两个妻子，他生儿育女。
2CHR|24|4|此后， 约阿施 有心重修耶和华的殿，
2CHR|24|5|就召集祭司和 利未 人，吩咐他们说：“你们要往 犹大 各城去，向 以色列 众人征收银子，按每年的需要整修你们上帝的殿；你们要急速办理这事。”但 利未 人没有急速办理。
2CHR|24|6|王召了 耶何耶大 祭司长来，对他说：“从前耶和华的仆人 摩西 ，为法柜的帐幕与 以色列 会众所定的捐献，你为何不叫 利未 人照这例向 犹大 和 耶路撒冷 征收呢？”
2CHR|24|7|因为那恶妇 亚她利雅 的儿子们曾拆毁上帝的殿，又用耶和华殿中分别为圣的物供奉诸 巴力 。
2CHR|24|8|于是王下令造一个柜子，放在耶和华殿的门外，
2CHR|24|9|又通告 犹大 和 耶路撒冷 ，要将上帝仆人 摩西 在旷野所吩咐 以色列 的捐献送来给耶和华。
2CHR|24|10|众领袖和百姓都欢欢喜喜带捐献来，投入柜中，直到投满。
2CHR|24|11|利未 人见银子多了，把柜子抬到王所派的官长面前；这时王的书记和祭司长的助手就会来把柜子倒空，然后放回原处。日日都是这样做，积蓄的银子很多。
2CHR|24|12|王与 耶何耶大 把银子交给耶和华殿里办事的人，他们就雇了石匠、木匠重修耶和华的殿，又雇了铁匠、铜匠整修耶和华的殿。
2CHR|24|13|工人做工，修理工程在他们手中渐渐完成，他们将上帝的殿修理得如同从前一样，非常坚固。
2CHR|24|14|他们做完了，就把多余的银子拿到王与 耶何耶大 面前，用以制造耶和华殿供奉所用的器皿和调羹，以及金银的器皿。 耶何耶大 在世的日子，众人经常在耶和华殿里献燔祭。
2CHR|24|15|耶何耶大 年纪老迈，日子满足而死，死的时候年一百三十岁。
2CHR|24|16|众人把他与列王同葬在 大卫城 ，因为他在 以色列 中为上帝和他的殿做了美善的事。
2CHR|24|17|耶何耶大 死后， 犹大 的众领袖来叩拜王，那时王就听了他们。
2CHR|24|18|他们离弃耶和华－他们列祖上帝的殿，去事奉 亚舍拉 和偶像；因他们这罪，就有愤怒临到 犹大 和 耶路撒冷 。
2CHR|24|19|但上帝仍差遣先知到他们那里，引导他们归向耶和华。先知警戒他们，他们却不肯听。
2CHR|24|20|那时，上帝的灵感动 耶何耶大 的儿子 撒迦利亚 祭司，他就站在上面，对百姓说：“上帝如此说：‘你们为何干犯耶和华的诫命，以致不得亨通呢？因为你们离弃耶和华，所以他也离弃你们。’”
2CHR|24|21|众人谋害 撒迦利亚 ，照着王的吩咐，在耶和华殿的院内用石头打死他。
2CHR|24|22|这样， 约阿施 王不记念 撒迦利亚 的父亲 耶何耶大 向自己所施的恩，杀了他的儿子。 撒迦利亚 临死的时候说：“愿耶和华鉴察伸冤！”
2CHR|24|23|年底的时候， 亚兰 的军兵上来攻击 约阿施 ，来到 犹大 和 耶路撒冷 ，杀了百姓中的众领袖，把所掠取的财物全送到 大马士革 王那里。
2CHR|24|24|亚兰 的军兵虽只来了一小队人，耶和华却将极大的军队交在他们手里；因为 犹大 人离弃耶和华－他们列祖的上帝，所以 亚兰 人惩罚 约阿施 。
2CHR|24|25|亚兰 人离开 约阿施 的时候，他患重病 ；他的臣仆背叛他，要报 耶何耶大 祭司儿子 的流血之仇，在床上杀了他。他就死了，葬在 大卫城 ，只是不葬在列王的坟墓里。
2CHR|24|26|背叛他的是 亚扪 妇人 示米押 的儿子 撒拔 和 摩押 妇人 示米利 的儿子 约萨拔 。
2CHR|24|27|至于他的儿子们和他所受的众多警戒，以及他重修上帝殿的事，看哪，都写在《列王评传》上。他的儿子 亚玛谢 接续他作王。
2CHR|25|1|亚玛谢 登基的时候年二十五岁，在 耶路撒冷 作王二十九年。他母亲名叫 约耶但 ，是 耶路撒冷 人。
2CHR|25|2|亚玛谢 行耶和华眼中看为正的事，只是没有纯正的心。
2CHR|25|3|他的王国一巩固，就把杀他父王的臣仆杀了，
2CHR|25|4|却没有处死他们的儿子，这是照 摩西 律法书上耶和华所吩咐的说：“不可因子杀父，也不可因父杀子，各人要为自己的罪而死。”
2CHR|25|5|亚玛谢 召集 犹大 人，按着父家为全 犹大 和 便雅悯 设立千夫长、百夫长，又数点人数，从二十岁以上，能拿枪拿盾牌出去打仗的精兵共有三十万；
2CHR|25|6|又用一百他连得银子，从 以色列 招募了十万大能的勇士。
2CHR|25|7|有一个神人来见 亚玛谢 ，对他说：“王啊，不要带领 以色列 的军兵与你同去，因为耶和华不和 以色列 ，和任何 以法莲 的子孙同在。
2CHR|25|8|你若一定要去，就奋勇作战吧！但上帝必使你败在敌人面前，因为上帝能助人得胜，也能使人落败。”
2CHR|25|9|亚玛谢 问神人：“我给了 以色列 军队的那一百他连得银子怎么样呢？”神人回答：“耶和华会把比这些更多的赐给你。”
2CHR|25|10|于是 亚玛谢 把那从 以法莲 来的军兵分别出来，叫他们到自己的地方去。他们非常恼怒 犹大 ，气愤地回自己的地方去了。
2CHR|25|11|亚玛谢 壮起胆来，率领他的军队到 盐谷 ，杀了一万 西珥 人。
2CHR|25|12|犹大 人又生擒了一万人，把他们带到 西拉 山顶上，从 西拉 山顶扔下去，把他们全都摔碎了。
2CHR|25|13|但 亚玛谢 所打发回去、不许一同出征的那些军兵劫掠 犹大 各城，从 撒玛利亚 直到 伯．和仑 ，杀了三千人，抢了许多财物。
2CHR|25|14|亚玛谢 击杀 以东 人回来以后，他把 西珥 人的神像带回，立为自己的神明，在它们面前叩拜烧香。
2CHR|25|15|耶和华的怒气向 亚玛谢 发作，差派一个先知去见他，对他说：“这些神明不能救自己的百姓脱离你的手，你为何寻求它们呢？”
2CHR|25|16|先知与王说话的时候，王对他说：“难道我们立你作王的谋士吗？你住口吧！为何要挨打呢？”先知就止住了，却说：“我知道上帝已定意要消灭你，因为你行这事，不听从我的劝戒。”
2CHR|25|17|犹大 王 亚玛谢 经商议后，就派人去见 耶户 的孙子， 约哈斯 的儿子 以色列 王 约阿施 ，说：“来，让我们面对面较量吧！”
2CHR|25|18|以色列 王 约阿施 派人去见 犹大 王 亚玛谢 ，说：“ 黎巴嫩 的蒺藜派人去见 黎巴嫩 的香柏树，说：‘将你的女儿嫁给我的儿子。’但有一只野兽经过 黎巴嫩 ，把蒺藜践踏了。
2CHR|25|19|你说，看哪，你打败了 以东 ，就心高气傲，以此为荣。现在，你待在家里算了吧，为何要惹祸使自己和 犹大 一同败亡呢？”
2CHR|25|20|亚玛谢 却不肯听从。这是出乎上帝，好将他们交在敌人手里，因为他们寻求 以东 的神明。
2CHR|25|21|于是 以色列 王 约阿施 上来，在 犹大 的 伯．示麦 与 犹大 王 亚玛谢 面对面较量。
2CHR|25|22|犹大 败在 以色列 面前，他们逃跑，各人逃回自己的帐棚去了。
2CHR|25|23|以色列 王 约阿施 在 伯．示麦 擒住 约哈斯 的孙子， 约阿施 的儿子 犹大 王 亚玛谢 ，把他带到 耶路撒冷 ，又拆毁 耶路撒冷 的城墙，从 以法莲门 直到 角门 共四百肘。
2CHR|25|24|他带着 俄别．以东 所看守上帝殿里的一切金银和器皿，与王宫里的财宝，又带着人质，回 撒玛利亚 去了。
2CHR|25|25|约哈斯 的儿子 以色列 王 约阿施 死后， 犹大 王 约阿施 的儿子 亚玛谢 又活了十五年。
2CHR|25|26|亚玛谢 其余的事，自始至终，看哪，不都写在《犹大和以色列诸王记》上吗？
2CHR|25|27|自从 亚玛谢 离弃耶和华之后，在 耶路撒冷 有人背叛他，他就逃往 拉吉 ；他们却派人追到 拉吉 ，在那里杀了他。
2CHR|25|28|有人用马将他驮回，把他与祖先一同葬在 犹大 的城 。
2CHR|26|1|犹大 众百姓立 乌西雅 接续他父亲 亚玛谢 作王，那时他年十六岁。
2CHR|26|2|亚玛谢 王与他祖先同睡之后， 乌西雅 收复 以禄 回归 犹大 ，又重新修建。
2CHR|26|3|乌西雅 登基的时候年十六岁，在 耶路撒冷 作王五十二年。他母亲名叫 耶可利雅 ，是 耶路撒冷 人。
2CHR|26|4|乌西雅 行耶和华眼中看为正的事，效法他父亲 亚玛谢 一切所行的。
2CHR|26|5|撒迦利亚 是一个通晓上帝默示的人 ，他在世的日子， 乌西雅 定意寻求上帝； 乌西雅 寻求耶和华的日子，上帝使他亨通。
2CHR|26|6|他出去攻击 非利士 人，拆毁了 迦特 、 雅比尼 和 亚实突 的城墙，又在 非利士 人中，在 亚实突 境内建筑城镇。
2CHR|26|7|上帝帮助他攻击 非利士 人和住在 姑珥．巴力 的 阿拉伯 人，以及 米乌尼 人。
2CHR|26|8|米乌尼 人 向 乌西雅 进贡。他的名声传到 埃及 ，因他非常强盛。
2CHR|26|9|乌西雅 在 耶路撒冷 的 角门 和 谷门 ，以及城墙转角之处建筑城楼，非常坚固。
2CHR|26|10|他在旷野建筑了望楼，又挖了许多井，因为他在 谢非拉 和平原有很多牲畜。他在山区和肥沃的土地雇用耕种田地和修整葡萄园的人，因为他喜爱土地。
2CHR|26|11|乌西雅 又有军兵，照书记 耶利 和官长 玛西雅 所数点的，在王的一个将军 哈拿尼雅 手下，分队出战。
2CHR|26|12|族长和大能勇士的总数共二千六百人，
2CHR|26|13|他们手下的军兵共三十万七千五百人，都大有能力，善于作战，帮助王攻击仇敌。
2CHR|26|14|乌西雅 为全军预备盾牌、头盔、铠甲、枪、弓和甩石的机弦，
2CHR|26|15|又在 耶路撒冷 叫巧匠设计机器，安在城楼和角楼上，用以射箭，投掷大石。 乌西雅 的名声传到远方，因为他得了非凡的帮助，极其强盛。
2CHR|26|16|乌西雅 既强盛，就心高气傲，以致败坏。他干犯耶和华－他的上帝，进耶和华的殿，要在香坛上烧香。
2CHR|26|17|亚撒利雅 祭司率领八十名勇敢的耶和华的祭司，跟随他进去。
2CHR|26|18|他们阻止 乌西雅 王，对他说：“ 乌西雅 啊，给耶和华烧香不是你的事，而是 亚伦 子孙的事，他们是分别为圣来烧香的祭司。你出圣殿吧！因为你犯了罪，耶和华上帝必不使你得尊荣。”
2CHR|26|19|乌西雅 发怒，手拿香炉要烧香。他在耶和华殿中香坛旁向众祭司发怒的时候，他的额头在众祭司面前忽然长出痲疯 。
2CHR|26|20|亚撒利雅 祭司长和众祭司转向他，看哪，他的额头长出痲疯，就催他离开那里；他自己也急速出去，因为耶和华降灾于他。
2CHR|26|21|乌西雅 王患痲疯直到死的那日；他因为染上痲疯，就住在隔离的行宫里，与耶和华的殿隔绝。他儿子 约坦 管理王的家，治理这地的百姓。
2CHR|26|22|乌西雅 其余的事，自始至终， 亚摩斯 的儿子 以赛亚 先知都记录下来。
2CHR|26|23|乌西雅 与他祖先同睡，与他祖先同葬在田间的王陵；因为人说，他是长痲疯的。他的儿子 约坦 接续他作王。
2CHR|27|1|约坦 登基的时候年二十五岁，在 耶路撒冷 作王十六年。他母亲名叫 耶路沙 ，是 撒督 的女儿。
2CHR|27|2|约坦 行耶和华眼中看为正的事，效法他父亲 乌西雅 一切所行的，只是他不入耶和华的殿。百姓仍旧行败坏的事。
2CHR|27|3|约坦 建造耶和华殿的 上门 ，在 俄斐勒 城墙上有很多建设，
2CHR|27|4|又在 犹大 山区建造城镇，在树林中建筑营寨和了望楼。
2CHR|27|5|约坦 与 亚扪 人的王打仗，胜了他们。那年 亚扪 人向他进贡一百他连得银子，一万歌珥小麦，一万歌珥大麦；第二年、第三年 亚扪 人也这样做。
2CHR|27|6|约坦 日渐强盛，因为他在耶和华－他上帝面前行正道。
2CHR|27|7|约坦 其余的事和一切战役，以及他的行为，看哪，都写在《以色列和犹大列王记》上。
2CHR|27|8|他登基的时候年二十五岁，在 耶路撒冷 作王十六年。
2CHR|27|9|约坦 与他祖先同睡，葬在 大卫城 ，他儿子 亚哈斯 接续他作王。
2CHR|28|1|亚哈斯 登基的时候年二十岁，在 耶路撒冷 作王十六年。他不像他祖先 大卫 行耶和华眼中看为正的事，
2CHR|28|2|却行 以色列 诸王的道，又铸造诸 巴力 的像，
2CHR|28|3|照着耶和华从 以色列 人面前赶出的外邦人所行可憎的事，在 欣嫩子谷 烧香，用火焚烧他的儿女，
2CHR|28|4|又在丘坛上、山冈上、各青翠树下献祭烧香。
2CHR|28|5|耶和华－他的上帝将他交在 亚兰 王手里。 亚兰 王打败他，从他掳走了许多人，带到 大马士革 去。上帝又将他交在 以色列 王手里， 以色列 王向他大行杀戮。
2CHR|28|6|利玛利 的儿子 比加 一日之内在 犹大 杀了十二万人，都是勇士，因为他们离弃了耶和华－他们列祖的上帝。
2CHR|28|7|有一个叫 细基利 的 以法莲 勇士，杀了 玛西雅 王子、 押斯利甘 宫廷总管和 以利加拿 宰相。
2CHR|28|8|以色列 人掳了他们的弟兄，连妇人带儿女共二十万，又掠取了许多财物，把这些掠物带到 撒玛利亚 去。
2CHR|28|9|但那里有耶和华的一个先知，名叫 俄德 ，出来迎接往 撒玛利亚 去的军兵，对他们说：“看哪，耶和华－你们列祖的上帝恼怒 犹大 人，将他们交在你们手里，你们竟怒气冲天，向他们大行杀戮。
2CHR|28|10|如今你们又有意强逼 犹大 人和 耶路撒冷 人作你们的奴婢，你们岂不是也得罪了耶和华－你们的上帝吗？
2CHR|28|11|现在你们当听我说，要将从你们弟兄中掳来的释放回去，因耶和华的烈怒已临到你们了。”
2CHR|28|12|于是， 以法莲 人的几个领袖，就是 约哈难 的儿子 亚撒利雅 、 米实利末 的儿子 比利家 、 沙龙 的儿子 耶希西家 、 哈得莱 的儿子 亚玛撒 ，起来拦阻从战场上回来的人，
2CHR|28|13|对他们说：“你们不可把这些被掳的人带到这里，因我们已经得罪耶和华了。你们还想加增我们的罪恶过犯吗？因为我们的罪过深重，已经有烈怒临到 以色列 了。”
2CHR|28|14|于是带兵器的人将掳来的人口和掠取的财物都留在众领袖和全会众面前。
2CHR|28|15|以上提名的那些人就起来，照顾被掳的人；其中凡赤身的，就从所掠取的财物中拿出衣服和鞋来，给他们穿，又给他们吃喝，用膏抹他们；其中凡软弱的，就使他们骑驴，送到棕树城 耶利哥 他们弟兄那里。然后，他们就回 撒玛利亚 去了。
2CHR|28|16|那时， 亚哈斯 王派人去求 亚述 诸王 来帮助他，
2CHR|28|17|因为 以东 人又来攻击 犹大 ，掳掠俘虏。
2CHR|28|18|非利士 人也来侵占 谢非拉 和 犹大 的 尼革夫 的城镇，攻取了 伯．示麦 、 亚雅仑 、 基低罗 、 梭哥 和所属的乡镇、 亭拿 和所属的乡镇、 瑾锁 和所属的乡镇，就住在那里。
2CHR|28|19|因为 以色列 王 亚哈斯 在 犹大 放肆，大大干犯耶和华，所以耶和华使 犹大 卑微。
2CHR|28|20|亚述 王 提革拉．毗列色 来攻击他，不帮助他，反倒欺负他。
2CHR|28|21|亚哈斯 从耶和华殿里和王宫中，以及众领袖家中取财宝送给 亚述 王，也无济于事。
2CHR|28|22|这 亚哈斯 王在急难的时候，越发得罪耶和华。
2CHR|28|23|他向那攻击他的 大马士革 的神明献祭，说：“因为 亚兰 王的神明帮助他们，我也要向这些神明献祭，好让它们帮助我。”但那些神明却使他和全 以色列 败亡。
2CHR|28|24|亚哈斯 聚集上帝殿里的器皿，把上帝殿里的器皿都打碎了，并且封锁耶和华殿的门，又在 耶路撒冷 各处的转角为自己建筑祭坛。
2CHR|28|25|他在 犹大 各城建立丘坛，向别神烧香，惹耶和华－他列祖的上帝发怒。
2CHR|28|26|亚哈斯 其余的事和他一切的行为，自始至终，看哪，都写在《犹大和以色列诸王记》上。
2CHR|28|27|亚哈斯 与他祖先同睡，葬在 耶路撒冷 城里，却没有送入 以色列 诸王的坟墓。他的儿子 希西家 接续他作王。
2CHR|29|1|希西家 登基的时候年二十五岁，在 耶路撒冷 作王二十九年。他母亲名叫 亚比雅 ，是 撒迦利雅 的女儿。
2CHR|29|2|希西家 行耶和华眼中看为正的事，效法他祖先 大卫 一切所行的。
2CHR|29|3|元年正月，他开了耶和华殿的门，重新整修。
2CHR|29|4|他召祭司和 利未 人来，聚集在东边的广场，
2CHR|29|5|对他们说：“ 利未 人哪，当听我说：现在你们要将自己分别为圣，又将耶和华－你们列祖上帝的殿分别为圣，从圣所中除去污秽之物。
2CHR|29|6|因我们的祖先犯了罪，行耶和华－我们上帝眼中看为恶的事，离弃他，转脸背向耶和华的居所。
2CHR|29|7|他们又封锁走廊的门，吹灭灯火，不在圣所中向 以色列 的上帝烧香，或献燔祭。
2CHR|29|8|耶和华的愤怒临到 犹大 和 耶路撒冷 ，使他们恐惧，令人惊骇，使人嗤笑，正如你们亲眼所见的。
2CHR|29|9|看哪，我们的祖宗倒在刀下，我们的妻子儿女也为此被掳掠。
2CHR|29|10|现在我心中有意与耶和华－ 以色列 的上帝立约，好使他的烈怒转离我们。
2CHR|29|11|我的众子啊，现在不要懈怠；因为耶和华拣选你们站在他面前事奉他，作他的仆人，向他烧香。”
2CHR|29|12|于是， 利未 人起来，当中有 哥辖 的子孙， 亚玛赛 的儿子 玛哈 、 亚撒利雅 的儿子 约珥 ； 米拉利 的子孙， 亚伯底 的儿子 基士 、 耶哈利勒 的儿子 亚撒利雅 ； 革顺 人， 薪玛 的儿子 约亚 、 约亚 的儿子 伊甸 ；
2CHR|29|13|以利撒反 的子孙 申利 和 耶利 ； 亚萨 的子孙， 撒迦利雅 和 玛探雅 ；
2CHR|29|14|希幔 的子孙 耶歇 和 示每 ； 耶杜顿 的子孙 示玛雅 和 乌薛 。
2CHR|29|15|他们聚集他们的弟兄，将自己分别为圣，照着耶和华的话和王的吩咐，进去洁净耶和华的殿。
2CHR|29|16|祭司进入耶和华的内殿要洁净殿，把耶和华殿中所发现一切污秽之物都搬出去，搬到耶和华殿的院子，由 利未 人接走，搬出去到外头的 汲沦溪 。
2CHR|29|17|从正月初一开始分别为圣，初八就来到耶和华殿的走廊。他们又用了八日使耶和华的殿分别为圣，到正月十六日才完成。
2CHR|29|18|于是，他们到里面去见 希西家 王，说：“我们已将耶和华的全殿和燔祭坛，以及坛的一切器皿、供饼的供桌，与供桌的一切器皿都洁净了；
2CHR|29|19|并且连 亚哈斯 王在位犯罪的时候所废弃的器皿，我们也都预备齐全，分别为圣，看哪，它们都在耶和华的祭坛前。”
2CHR|29|20|希西家 王清早起来，召集城里的领袖都上耶和华的殿。
2CHR|29|21|他们牵了七头公牛，七只公羊，七只羔羊，七只公山羊，要为国、为殿、为 犹大 作赎罪祭。王吩咐 亚伦 的子孙众祭司在耶和华的坛上献祭。
2CHR|29|22|他们宰了公牛，祭司将血接来，洒在坛上；他们宰了公羊，把血洒在坛上，又宰了羔羊，也把血洒在坛上。
2CHR|29|23|他们把那些作赎罪祭的公山羊牵到王和会众面前，按手在公山羊上。
2CHR|29|24|祭司宰了羊，将血献在坛上作赎罪祭，为全 以色列 赎罪，因为王吩咐要为全 以色列 献上燔祭和赎罪祭。
2CHR|29|25|王又派 利未 人在耶和华殿中敲钹，鼓瑟，弹琴，正如 大卫 和王的先见 迦得 ，以及 拿单 先知所吩咐的，就是耶和华藉先知所吩咐的。
2CHR|29|26|利未 人拿 大卫 的乐器，祭司拿号，一同站立。
2CHR|29|27|希西家 吩咐在坛上献燔祭，开始献燔祭的时候，他们就唱赞美耶和华的歌，吹号，并用 以色列 王 大卫 的乐器伴奏。
2CHR|29|28|全会众都敬拜，歌唱的歌唱，吹号的吹号，如此直到燔祭献完了。
2CHR|29|29|献完了祭，王和所有在场跟随他的人都俯伏敬拜。
2CHR|29|30|希西家 王与众领袖吩咐 利未 人用 大卫 和 亚萨 先见的诗词颂赞耶和华，他们欢欢喜喜地颂赞，低头敬拜。
2CHR|29|31|希西家 回应说：“如今你们既承接圣职归耶和华，就要前来把祭物和感谢祭奉到耶和华的殿里。”会众就奉上祭物和感谢祭，凡甘心乐意的也奉上燔祭。
2CHR|29|32|会众所奉的燔祭数目如下：七十头公牛，一百只公羊，二百只羔羊，这些全都是要作燔祭献给耶和华的；
2CHR|29|33|又有分别为圣之物，就是六百头公牛，三千只绵羊。
2CHR|29|34|但祭司太少，不能剥尽所有燔祭牲的皮，所以他们的弟兄 利未 人帮助他们，直等献祭的事完毕，直到其他的祭司也分别为圣了；因 利未 人以正直的心分别为圣，胜过祭司。
2CHR|29|35|燔祭和平安祭牲的脂肪，以及与燔祭同献的浇酒祭很多。这样，耶和华殿中的事务俱都齐备了。
2CHR|29|36|希西家 和众百姓都因上帝为百姓所预备的而喜乐，因为这事办得很迅速。
2CHR|30|1|希西家 派人去见 以色列 和 犹大 众人，又写信给 以法莲 和 玛拿西 人，要他们到 耶路撒冷 耶和华的殿，向耶和华－ 以色列 的上帝守逾越节，
2CHR|30|2|因为王和众领袖，以及 耶路撒冷 全会众已经商议，要在二月份守逾越节。
2CHR|30|3|那时他们不能守，因为分别为圣的祭司不够，百姓也还没有聚集在 耶路撒冷 。
2CHR|30|4|这事在王与全会众眼中都看为合宜。
2CHR|30|5|于是他们下令，通告全 以色列 ，从 别是巴 直到 但 ，吩咐百姓都来，在 耶路撒冷 向耶和华－ 以色列 的上帝守逾越节，因为他们已经许久没有照所写的守这节了 。
2CHR|30|6|信差遵着王命，拿着王和众领袖所发的信，送达全 以色列 和 犹大 ，说：“ 以色列 人哪，当转向耶和华－ 亚伯拉罕 、 以撒 、 以色列 的上帝，好叫他转向你们这些脱离 亚述 诸王之手的余民。
2CHR|30|7|不要效法你们的祖先和你们的弟兄；他们干犯耶和华－他们列祖的上帝，以致耶和华使他们令人惊骇，正如你们所见的。
2CHR|30|8|现在，不要像你们祖先硬着颈项，只要归顺耶和华，进入他的圣所，就是永远成圣的居所，又要事奉耶和华－你们的上帝，好使他的烈怒转离你们。
2CHR|30|9|你们若转向耶和华，你们的弟兄和儿女必在掳掠他们的人面前蒙怜悯，得以归回这地，因为耶和华－你们的上帝有恩惠，有怜悯。你们若转向他，他必不会转脸不顾你们。”
2CHR|30|10|信差从这城跑到那城，传遍了 以法莲 和 玛拿西 之地，直到 西布伦 ；那里的人却戏笑他们，讥诮他们。
2CHR|30|11|然而 亚设 、 玛拿西 、 西布伦 中也有人谦卑自己，来到 耶路撒冷 。
2CHR|30|12|上帝也按手在 犹大 人身上，使他们一心遵行王与众领袖照着耶和华的话所发的命令。
2CHR|30|13|二月时，许多百姓聚集在 耶路撒冷 ，成为一个盛大的会，要守除酵节。
2CHR|30|14|他们起来，把 耶路撒冷 的祭坛和烧香的坛尽都除去，扔在 汲沦溪 中。
2CHR|30|15|二月十四日，他们宰了逾越节的羔羊。祭司与 利未 人觉得惭愧，就使自己分别为圣，把燔祭奉到耶和华的殿中。
2CHR|30|16|他们遵照神人 摩西 的律法，按定例站在自己的地方；祭司从 利未 人手里接过血来，洒出去。
2CHR|30|17|会众中有许多人尚未分别为圣，所以 利未 人为所有不洁的人宰逾越节的羔羊，使他们归耶和华为圣。
2CHR|30|18|从 以法莲 、 玛拿西 、 以萨迦 、 西布伦 来的许多百姓尚未自洁，他们却吃逾越节的羔羊，不合所写的条例。 希西家 为他们祷告说：“求至善的耶和华饶恕
2CHR|30|19|那凡专心寻求上帝耶和华－他列祖的上帝，却未照圣所洁净礼自洁的人。”
2CHR|30|20|耶和华应允 希西家 ，医治了百姓。
2CHR|30|21|在 耶路撒冷 的 以色列 人守除酵节七日，大大喜乐。 利未 人和祭司为耶和华演奏响亮的乐器，天天颂赞耶和华。
2CHR|30|22|希西家 慰劳所有精通礼仪，事奉耶和华的 利未 人。于是众人吃节期的筵席七日，又献平安祭，并且称谢耶和华－他们列祖的上帝。
2CHR|30|23|全会众商议，要再守节七日；于是他们欢欢喜喜地又守节七日。
2CHR|30|24|犹大 王 希西家 赐给会众一千头公牛，七千只羊；众领袖也赐给会众一千头公牛，一万只羊，并有许多祭司将自己分别为圣。
2CHR|30|25|犹大 全会众、祭司、 利未 人和从 以色列 来的全会众，以及那些从 以色列 地来的和住在 犹大 的寄居的人，尽都喜乐。
2CHR|30|26|这样，在 耶路撒冷 大有喜乐，因自从 以色列 王 大卫 的儿子 所罗门 以来，在 耶路撒冷 从未有过这样的喜乐。
2CHR|30|27|那时，祭司和 利未 人起来，为百姓祝福。他们的声音蒙上帝垂听，他们的祷告达到他天上的圣所。
2CHR|31|1|这一切事都完毕以后，在那里的 以色列 众人就到 犹大 的城镇，打碎柱像，砍断 亚舍拉 ，又在 犹大 、 便雅悯 、 以法莲 、 玛拿西 遍地把丘坛和祭坛完全拆毁。于是 以色列 众人各回各城，各归自己产业的地去了。
2CHR|31|2|希西家 分派祭司和 利未 人的班次，使祭司和 利未 人照各自的班次，按各自的职分献燔祭和平安祭，又在耶和华殿 的门内事奉，称谢颂赞耶和华。
2CHR|31|3|王又从自己的产业中分出一份来作燔祭，就是早晚的燔祭，和安息日、初一，以及节期的燔祭，都是按耶和华律法上所记载的。
2CHR|31|4|他又吩咐住 耶路撒冷 的百姓将祭司和 利未 人所应得的份给他们，使他们坚守耶和华的律法。
2CHR|31|5|命令一出， 以色列 人就把初熟的五谷、新酒、新油、蜜和田地的出产多多送来；他们把各样出产的十分之一大量送来。
2CHR|31|6|住 犹大 各城的 以色列 人和 犹大 人也将牛羊的十分之一，以及分别为圣归耶和华－他们上帝之物，就是十分取一之物，尽都送来，积成一堆一堆；
2CHR|31|7|他们从三月开始堆积，到七月才完成。
2CHR|31|8|希西家 和众领袖来，看见这些堆积物，就称颂耶和华，又为耶和华的百姓 以色列 祝福。
2CHR|31|9|希西家 向祭司和 利未 人查问这些堆积物。
2CHR|31|10|撒督 家的 亚撒利雅 祭司长告诉他说：“自从礼物开始送到耶和华的殿以来，我们不但吃饱，而且剩下的很多；因为耶和华赐福给他的百姓，所剩下的才这样丰盛。”
2CHR|31|11|希西家 吩咐要在耶和华殿里预备仓房，他们就预备了。
2CHR|31|12|他们诚心将礼物，十分取一之物，就是分别为圣之物，都搬入仓内。 利未 人 歌楠雅 主管这事，他的兄弟 示每 是副主管。
2CHR|31|13|耶歇 、 亚撒细雅 、 拿哈 、 亚撒黑 、 耶利摩 、 约撒拔 、 以列 、 伊斯玛基雅 、 玛哈 、 比拿雅 都是督办，在 歌楠雅 和他兄弟 示每 的手下，是 希西家 王和管理上帝殿的 亚撒利雅 所委派的。
2CHR|31|14|守东门的 利未 人 音拿 的儿子 可利 ，掌管献给上帝的甘心祭，发放献给耶和华的礼物和至圣的物。
2CHR|31|15|在祭司的各城里，在他手下忠心协助他的有 伊甸 、 (王民)雅(王民) 、 耶书亚 、 示玛雅 、 亚玛利雅 、 示迦尼雅 ，都按着班次分给他们的弟兄，无论大小，
2CHR|31|16|不论是否登录在家谱，凡三岁以上的男丁，每日进耶和华殿、按班次供职事奉的，都分给他，
2CHR|31|17|也发放给按父家登录在家谱的祭司；又按班次职任分给二十岁以上的 利未 人，
2CHR|31|18|又按家谱的登记，分给他们的小孩、妻子、儿女，给全体会众；因为他们忠诚，将自己分别为圣。
2CHR|31|19|住在各城郊野 亚伦 的子孙、按名受委任的人，要把应得的份给祭司中所有的男丁和载入家谱的 利未 人。
2CHR|31|20|希西家 在全 犹大 都这样办理，在耶和华－他上帝面前行良善、正直、忠诚的事。
2CHR|31|21|凡他所行的，无论是开始办上帝殿的事，是遵律法守诫命，是寻求他的上帝，他都尽心去做，无不亨通。
2CHR|32|1|在这些虔诚的事以后， 亚述 王 西拿基立 来侵犯 犹大 ，围困坚固城，想要攻破它们。
2CHR|32|2|希西家 见 西拿基立 来，定意要攻打 耶路撒冷 ，
2CHR|32|3|就与领袖和勇士商议，塞住城外的泉源；他们都帮助他。
2CHR|32|4|于是许多百姓聚集，塞住一切泉源，以及国中流通的小河，说：“ 亚述 诸王来，为何让他们得着许多水呢？”
2CHR|32|5|希西家 奋勇自强，修筑所有毁坏的城墙，升高城楼，又在城外筑另一片城墙，坚固 大卫城 的 米罗 ，制造许多兵器和盾牌。
2CHR|32|6|他设立军事将领管理百姓，召集他们在城门的广场，勉励他们，说：
2CHR|32|7|“你们当刚强壮胆，不要因 亚述 王和跟随他的大军恐惧惊慌，因为与我们同在的，比与他们同在的更大。
2CHR|32|8|与他们同在的是血肉之臂，但与我们同在的是耶和华－我们的上帝，他必帮助我们，为我们争战。”百姓因 犹大 王 希西家 的话就得到鼓励。
2CHR|32|9|此后， 亚述 王 西拿基立 和跟随他的全军攻打 拉吉 ，派臣仆到 耶路撒冷 见 犹大 王 希西家 和所有在 耶路撒冷 的 犹大 人，说：
2CHR|32|10|“ 亚述 王 西拿基立 如此说：‘你们倚靠什么，还留在 耶路撒冷 受困吗？
2CHR|32|11|希西家 说：耶和华－我们的上帝必救我们脱离 亚述 王的手，这不是诱惑你们，使你们受饥渴而死吗？
2CHR|32|12|希西家 岂不是将耶和华的丘坛和祭坛废去，并且吩咐 犹大 与 耶路撒冷 的人说：你们当在一个坛前敬拜，在其上烧香吗？
2CHR|32|13|我与我祖先向列邦民族所行的，你们岂不知道吗？列邦的神明何尝能救自己的国脱离我的手呢？
2CHR|32|14|我祖先所灭的那些国的神明，有谁能救自己的百姓脱离我的手呢？难道你们的上帝能救你们脱离我的手吗？
2CHR|32|15|现在，不要让 希西家 这样欺骗你们，诱惑你们，也不要相信他，因为没有一国一邦的神明能救自己的百姓脱离我的手和我祖先的手，你们的上帝也绝不能救你们脱离我的手。’”
2CHR|32|16|西拿基立 的臣仆还说了一些话来毁谤耶和华上帝和他的仆人 希西家 。
2CHR|32|17|西拿基立 也写信毁谤耶和华－ 以色列 的上帝，说：“列邦的神明既不能救自己的百姓脱离我的手， 希西家 的上帝也不能救他的百姓脱离我的手。”
2CHR|32|18|亚述 王的臣仆用 犹大 话向 耶路撒冷 城墙上的百姓大声呼喊，要恐吓他们，扰乱他们，以便取城。
2CHR|32|19|他们谈论 耶路撒冷 的上帝，如同谈论世上人手所造的神明一样。
2CHR|32|20|希西家 王和 亚摩斯 的儿子 以赛亚 先知为此祷告，向天呼求。
2CHR|32|21|耶和华就差遣一个使者进入 亚述 王的营中，把所有大能的勇士、官长和将领尽都灭了。 亚述 王满面羞愧地回到本国，进了他神明的庙中，他几个亲生的儿子在那里用刀杀了他。
2CHR|32|22|这样，耶和华救 希西家 和 耶路撒冷 的居民脱离 亚述 王 西拿基立 的手，也脱离一切仇敌的手，又赐他们四境平安 。
2CHR|32|23|有许多人到 耶路撒冷 将供物献与耶和华，又将宝物送给 犹大 王 希西家 。自此之后， 希西家 在列国人的眼中受人尊崇。
2CHR|32|24|那些日子， 希西家 病得要死，就向耶和华祷告，耶和华应允他，赐他一个预兆。
2CHR|32|25|希西家 却没有照他所蒙的恩回报，因他心里骄傲，所以愤怒要临到他，临到 犹大 和 耶路撒冷 。
2CHR|32|26|但 希西家 和 耶路撒冷 的居民为了心里骄傲，就一同谦卑，以致耶和华的愤怒在 希西家 的日子没有临到他们。
2CHR|32|27|希西家 大有财富和尊荣，他为自己建造府库，收藏金银、宝石、香料、盾牌和各样的宝器，
2CHR|32|28|又建造仓房，收藏五谷、新酒和新的油，又为各类牲畜盖棚立圈，
2CHR|32|29|并且为自己建立城镇，也拥有许多的羊群牛群，因为上帝赐他极多的财产。
2CHR|32|30|这 希西家 也塞住 基训 的上源，引水直下，流在 大卫城 的西边。 希西家 所行的事尽都亨通。
2CHR|32|31|但当 巴比伦 诸侯差遣使者来见 希西家 ，询问国中所发生的奇事时，上帝离开他，要考验他，好知道他心里的一切。
2CHR|32|32|希西家 其余的事和他的善行，看哪，都写在 亚摩斯 的儿子 以赛亚 先知的《默示书》上和《犹大和以色列诸王记》上。
2CHR|32|33|希西家 与他祖先同睡，葬在 大卫 子孙陵墓的斜坡上。他死的时候， 犹大 众人和 耶路撒冷 的居民都向他致敬。他的儿子 玛拿西 接续他作王。
2CHR|33|1|玛拿西 登基的时候年十二岁，在 耶路撒冷 作王五十五年。
2CHR|33|2|他行耶和华眼中看为恶的事，效法耶和华在 以色列 人面前赶出的列国那些可憎的事。
2CHR|33|3|他重新建筑他父亲 希西家 所拆毁的丘坛，为诸 巴力 筑坛，造 亚舍拉 ，又敬拜天上的万象，事奉它们。
2CHR|33|4|他在耶和华殿中筑坛，耶和华曾指着这殿说：“我的名必永远在 耶路撒冷 。”
2CHR|33|5|他在耶和华殿的两个院子为天上的万象筑坛，
2CHR|33|6|并在 欣嫩子谷 使他的儿子经火，又观星象，行法术，行邪术，求问招魂的和行巫术的，多行耶和华眼中看为恶的事，惹他发怒。
2CHR|33|7|他在上帝殿内立雕刻的偶像；上帝曾对 大卫 和他儿子 所罗门 说：“我在 以色列 众支派中所选择的 耶路撒冷 和这殿，必立我的名，直到永远。
2CHR|33|8|只要 以色列 人谨守遵行我藉 摩西 吩咐他们的一切律法、律例、典章，我就不再使他们的脚挪移，离开我所赐给他们列祖之土地。”
2CHR|33|9|玛拿西 引诱 犹大 和 耶路撒冷 的居民行恶，比耶和华在 以色列 人面前所灭的列国更严重。
2CHR|33|10|耶和华警戒 玛拿西 和他的百姓，他们却不听。
2CHR|33|11|所以耶和华使 亚述 王的将领来攻击他们，用手铐铐住 玛拿西 ，用铜链锁住他，把他带到 巴比伦 去。
2CHR|33|12|他在急难的时候恳求耶和华－他的上帝，并在他列祖的上帝面前极其谦卑。
2CHR|33|13|他祈祷耶和华，耶和华就应允他，垂听他的祷告，使他归回 耶路撒冷 ，仍坐王位。 玛拿西 这才知道惟独耶和华是上帝。
2CHR|33|14|此后， 玛拿西 在 大卫城 外，从谷内 基训 西边直到 鱼门 口，建筑城墙，环绕 俄斐勒 ；这墙建得很高。他又在 犹大 各坚固城内设立将领。
2CHR|33|15|他除掉外邦人的神像与耶和华殿中的偶像，又将他在耶和华殿的山上和 耶路撒冷 所筑的各坛都拆毁，抛在城外。
2CHR|33|16|他重修耶和华的祭坛，在坛上献平安祭和感谢祭，并吩咐 犹大 人事奉耶和华－ 以色列 的上帝。
2CHR|33|17|百姓却仍在丘坛上献祭，不过，他们只献给耶和华－他们的上帝。
2CHR|33|18|玛拿西 其余的事和他向上帝的祷告，以及先见奉耶和华－ 以色列 上帝的名警戒他的话，看哪，都在《以色列诸王记》上。
2CHR|33|19|他的祷告，上帝怎样应允他，他未谦卑以前的一切罪愆过犯，以及在何处建筑丘坛，设立 亚舍拉 和雕刻的偶像，看哪，都写在 何赛 的书上。
2CHR|33|20|玛拿西 与他祖先同睡，葬在自己的宫中，他儿子 亚们 接续他作王。
2CHR|33|21|亚们 登基的时候年二十二岁，在 耶路撒冷 作王二年。
2CHR|33|22|他行耶和华眼中看为恶的事，效法他父亲 玛拿西 所行的，祭祀他父亲 玛拿西 所雕刻的一切偶像，事奉它们，
2CHR|33|23|但他不像他父亲 玛拿西 在耶和华面前那样谦卑下来。这 亚们 的罪越犯越大。
2CHR|33|24|他的臣仆背叛他，在宫里杀了他。
2CHR|33|25|但这地的百姓杀了所有背叛 亚们 王的人；这地的百姓立他儿子 约西亚 接续他作王。
2CHR|34|1|约西亚 登基的时候年八岁，在 耶路撒冷 作王三十一年。
2CHR|34|2|他行耶和华眼中看为正的事，行他祖先 大卫 所行的道，不偏左右。
2CHR|34|3|他作王第八年，尚且年轻，就寻求他祖先 大卫 的上帝。到了十二年，他开始洁净 犹大 和 耶路撒冷 ，除掉丘坛、 亚舍拉 、雕刻的像和铸造的像。
2CHR|34|4|众人在他面前拆毁诸 巴力 的坛，砍断坛上高高的香坛，又把 亚舍拉 和雕刻的像，以及铸造的像打碎成灰，撒在向偶像献祭之人的坟上，
2CHR|34|5|把祭司的骸骨烧在他们的坛上，洁净了 犹大 和 耶路撒冷 。
2CHR|34|6|他又在 玛拿西 、 以法莲 、 西缅 、 拿弗他利 各城和四围的废墟 ，
2CHR|34|7|拆毁祭坛，把 亚舍拉 和雕刻的像打碎成灰，砍断 以色列 全地所有的香坛。于是他回 耶路撒冷 去了。
2CHR|34|8|约西亚 王十八年，这地和殿洁净了之后，他派 亚萨利雅 的儿子 沙番 、 玛西雅 市长、 约哈斯 的儿子 约亚 史官去整修耶和华－他上帝的殿。
2CHR|34|9|他们去见 希勒家 大祭司，把奉到上帝殿的银子交给他；这银子是看守殿门的 利未 人从 玛拿西 、 以法莲 ，和 以色列 所有幸存的人，以及 犹大 、 便雅悯 众人和 耶路撒冷 的居民收来的。
2CHR|34|10|他们把这银子交给耶和华殿里督工的，由他们转交整修耶和华殿的工匠，
2CHR|34|11|就是交给木匠和石匠，好为 犹大 王所毁坏的殿，买凿成的石头和作钩子与栋梁的木料。
2CHR|34|12|这些人办事诚实，管理他们的是 利未 人 米拉利 的子孙 雅哈 和 俄巴底 ，又有 哥辖 人 撒迦利亚 和 米书兰 ；还有所有善于奏乐的 利未 人。
2CHR|34|13|他们监督扛抬的人，督导一切做各样工的人。 利未 人中也有作书记、官员、守卫的。
2CHR|34|14|他们把奉到耶和华殿的银子运出来的时候， 希勒家 祭司发现了耶和华藉 摩西 所传的律法书。
2CHR|34|15|希勒家 对 沙番 书记说：“我在耶和华殿里发现了律法书。” 希勒家 把书递给 沙番 。
2CHR|34|16|沙番 把书拿到王那里，又把这事回覆王说：“凡交给仆人的手所办的事，他们都办好了。
2CHR|34|17|耶和华殿里所发现的银子已经倒出来，交在督工和工匠的手里了。”
2CHR|34|18|沙番 书记又向王报告说：“ 希勒家 祭司递给我一卷书。” 沙番 就在王面前朗读那书。
2CHR|34|19|王听见律法的话，就撕裂衣服。
2CHR|34|20|王吩咐 希勒家 与 沙番 的儿子 亚希甘 、 米迦 的儿子 亚比顿 、 沙番 书记和王的臣仆 亚撒雅 ，说：
2CHR|34|21|“你们去，以所发现这书上的话，为我、为 以色列 和 犹大 幸存的人求问耶和华；因为我们的祖先没有遵守耶和华的话，没有照这书上所记的一切去做，耶和华的烈怒就倒在我们身上。”
2CHR|34|22|于是， 希勒家 和王的人 都去见 户勒大 女先知，她是掌管礼服的 沙龙 的妻子， 沙龙 是 哈斯拉 的孙子， 特瓦 的儿子。 户勒大 住在 耶路撒冷 第二区。他们向她说明来意。
2CHR|34|23|她对他们说：“耶和华－ 以色列 的上帝如此说：‘你们可以回覆那派你们来见我的人说，
2CHR|34|24|耶和华如此说：看哪，我必照着在 犹大 王面前所读那书上记载的一切诅咒，降祸于这地方和其上的居民。
2CHR|34|25|因为他们离弃我，向别神烧香，用他们手所做的一切惹我发怒，所以我的愤怒必倒在这地方，总不止息。’
2CHR|34|26|然而，派你们来求问耶和华的 犹大 王，你们要这样回覆他：‘耶和华－ 以色列 的上帝如此说：至于你所听见的话，
2CHR|34|27|就是听见我指着这地方和其上居民所说的话，你的心就软化，在我面前谦卑下来，撕裂衣服，向我哭泣，因此我应允你。这是耶和华说的。
2CHR|34|28|看哪，我必使你归到你祖先那里，平安地进入坟墓，我要降于这地方和其上居民的一切灾祸，你不会亲眼看见。’”他们就去把这话回覆王。
2CHR|34|29|王派人召集 犹大 和 耶路撒冷 的众长老来。
2CHR|34|30|王和 犹大 众人、 耶路撒冷 的居民、祭司、 利未 人，以及所有的百姓，无论大小，都一同上到耶和华的殿去；王把殿里所发现的约书上面一切的话读给他们听。
2CHR|34|31|王站在自己的位上，在耶和华面前立约，要尽心尽性跟从耶和华，遵守他的诫命、法度、律例，实行这书上所记这约的话；
2CHR|34|32|又使所有住 耶路撒冷 和 便雅悯 的人都服从这约。于是 耶路撒冷 的居民都遵行上帝，就是他们列祖之上帝的约。
2CHR|34|33|约西亚 从 以色列 各处把一切可憎之物尽都除掉，使 以色列 境内的人都事奉耶和华－他们的上帝。 约西亚 在世的日子，众人都跟从耶和华－他们列祖的上帝，总不离开。
2CHR|35|1|约西亚 在 耶路撒冷 向耶和华守逾越节。正月十四日，他们宰了逾越节的羔羊。
2CHR|35|2|王分派祭司各尽其职，又勉励他们办耶和华殿中的事。
2CHR|35|3|他对那归耶和华为圣、教导 以色列 众人的 利未 人说：“你们将圣约柜安放在 以色列 王 大卫 儿子 所罗门 建造的殿里，不必再用肩扛抬。现在你们要服事耶和华－你们的上帝和他的百姓 以色列 。
2CHR|35|4|你们应当按着父家，照着班次，遵照 以色列 王 大卫 和他儿子 所罗门 所写的，预备自己。
2CHR|35|5|要按着你们百姓的弟兄、父家的班次，侍立在圣所；每父家的班次中要有几个 利未 人。
2CHR|35|6|要宰逾越节的羔羊，将自己分别为圣，为你们的弟兄预备，好遵守耶和华藉 摩西 所吩咐的话。”
2CHR|35|7|约西亚 从群畜中赐给所有在场的百姓，三万只小绵羊和小山羊，三千头牛，作逾越节的祭物；这些都是出自王的产业。
2CHR|35|8|约西亚 的众领袖也乐意把祭牲给百姓、祭司和 利未 人；管理上帝殿的 希勒家 、 撒迦利亚 、 耶歇 ，把二千六百只羔羊和三百头牛给祭司作逾越节的祭物。
2CHR|35|9|利未 人的族长 歌楠雅 和他两个兄弟 示玛雅 、 拿坦业 ，与 哈沙比雅 、 耶利 、 约撒拔 ，把五千只羔羊和五百头牛给 利未 人作逾越节的祭物。
2CHR|35|10|这样，事奉的工作都安排好了，照王所吩咐的，祭司站在自己的位上， 利未 人按着班次侍立。
2CHR|35|11|他们宰了逾越节的羔羊，祭司从他们手里接过血来 洒出去； 利未 人剥皮，
2CHR|35|12|把燔祭拿走，再按着父家的班次分给众百姓，照 摩西 书上所写的献给耶和华；献牛也是这样。
2CHR|35|13|他们按着常例，用火烤逾越节的羔羊。至于其他的圣物，他们用盆，用锅，用釜煮了，速速地送给众百姓。
2CHR|35|14|然后他们为自己和祭司预备祭物，因为作祭司的 亚伦 子孙献燔祭和脂肪，直到晚上。所以 利未 人为自己和作祭司的 亚伦 子孙预备。
2CHR|35|15|歌唱的 亚萨 子孙，照着 大卫 、 亚萨 、 希幔 和王的先见 耶杜顿 所吩咐的，站在自己的位上。守门的看守各门，不用离开他们的职守，因为他们的弟兄 利未 人给他们预备。
2CHR|35|16|当日，一切供奉耶和华、守逾越节，以及在耶和华坛上献燔祭的事，都照 约西亚 王的吩咐预备好了。
2CHR|35|17|那时，在场的 以色列 人都守逾越节，又守除酵节七日。
2CHR|35|18|自从 撒母耳 先知的日子以来，在 以色列 中没有守过这样的逾越节， 以色列 诸王也没有守过像 约西亚 、祭司、 利未 人、所有住 犹大 和 以色列 的人，以及 耶路撒冷 居民所守的逾越节。
2CHR|35|19|这逾越节是 约西亚 作王十八年时守的。
2CHR|35|20|约西亚 为殿做完这一切事以后， 埃及 王 尼哥 上来，要攻打靠近 幼发拉底河 的 迦基米施 ； 约西亚 出去迎击他。
2CHR|35|21|他派使者来见 约西亚 ，说：“ 犹大 王啊，我跟你有什么相干呢？我今日来不是要攻打你，而是要攻打与我争战之家，并且上帝吩咐我从速行事。你不要干预与我同在的上帝，免得他毁灭你。”
2CHR|35|22|约西亚 却不转脸离开他，反而改装要与他打仗。他不听从上帝藉 尼哥 的口所说的话，就来到 米吉多 平原争战。
2CHR|35|23|弓箭手射中 约西亚 王。王对他的臣仆说：“我受了重伤，你们载我离开战场吧！”
2CHR|35|24|他的臣仆扶他下了战车，上了他的副座车，送他到 耶路撒冷 。他就死了，葬在他祖先的坟墓里。全 犹大 和 耶路撒冷 都哀悼 约西亚 。
2CHR|35|25|耶利米 为 约西亚 作哀歌，所有歌唱的男女也唱哀歌，追悼 约西亚 ，直到今日。他们在 以色列 中以此为定例；看哪，这些哀歌写在《哀歌书》上。
2CHR|35|26|约西亚 其余的事和他遵照耶和华律法上所记而行的善事，
2CHR|35|27|以及他自始至终所行的，看哪，都写在《以色列和犹大列王记》上。
2CHR|36|1|这地的百姓立 约西亚 的儿子 约哈斯 在 耶路撒冷 接续他父亲作王。
2CHR|36|2|约哈斯 登基的时候年二十三岁，在 耶路撒冷 作王三个月。
2CHR|36|3|埃及 王在 耶路撒冷 废了他，又罚这地一百他连得银子，一他连得金子。
2CHR|36|4|埃及 王 尼哥 立 约哈斯 的哥哥 以利雅敬 作 犹大 和 耶路撒冷 的王，给他改名叫 约雅敬 。 尼哥 却将他的弟弟 约哈斯 带到 埃及 去。
2CHR|36|5|约雅敬 登基的时候年二十五岁，在 耶路撒冷 作王十一年。他行耶和华－他上帝眼中看为恶的事。
2CHR|36|6|巴比伦 王 尼布甲尼撒 上来攻击他，用铜链锁着他，要把他带到 巴比伦 去。
2CHR|36|7|尼布甲尼撒 又将耶和华殿里的一些器皿带到 巴比伦 ，放在 巴比伦 自己的宫里 。
2CHR|36|8|约雅敬 其余的事和他所行可憎的事，以及发生在他身上的事，看哪，都写在《以色列和犹大列王记》上，他儿子 约雅斤 接续他作王。
2CHR|36|9|约雅斤 登基的时候年八岁 ，在 耶路撒冷 作王三个月十天，他行耶和华眼中看为恶的事。
2CHR|36|10|过了一年， 尼布甲尼撒 王差遣人将 约雅斤 和耶和华殿里宝贵的器皿带到 巴比伦 ，然后立 约雅斤 的叔父 西底家 作 犹大 和 耶路撒冷 的王。
2CHR|36|11|西底家 登基的时候年二十一岁，在 耶路撒冷 作王十一年。
2CHR|36|12|他行耶和华－他上帝眼中看为恶的事，没有谦卑听从 耶利米 先知所传达耶和华的话。
2CHR|36|13|尼布甲尼撒 王曾叫他指着上帝起誓，他却背叛，硬着颈项，内心顽固，不归向耶和华－ 以色列 的上帝。
2CHR|36|14|众祭司长和百姓也多多犯罪，效法列国一切可憎的事，玷污耶和华在 耶路撒冷 分别为圣的殿。
2CHR|36|15|耶和华－他们列祖的上帝因为爱惜自己的百姓和居所，一再差遣使者去警戒他们。
2CHR|36|16|他们却嘲笑上帝的使者，藐视他的话，讥诮他的先知，以致耶和华向他的百姓大发烈怒，甚至无法可救。
2CHR|36|17|所以，耶和华使 迦勒底 人的王来攻击他们，在他们圣殿里用刀杀了他们的壮丁，不怜悯他们的少男少女、老人长者。耶和华把所有的人都交在他手里。
2CHR|36|18|他把上帝殿里一切的大小器皿与耶和华殿里的财宝，以及王和众领袖的财宝，全都带到 巴比伦 去。
2CHR|36|19|迦勒底 人焚烧了上帝的殿，拆毁 耶路撒冷 的城墙，用火烧了城里所有的宫殿，毁坏了城里一切宝贵的器皿。
2CHR|36|20|凡脱离刀剑的幸存者， 迦勒底 王都掳到 巴比伦 去，作他和他子孙的仆婢，直到 波斯 国兴起。
2CHR|36|21|这就应验耶和华藉 耶利米 的口所说的话：地得享安息；在荒凉的日子，地就守安息，直到满了七十年。
2CHR|36|22|波斯 王 居鲁士 元年，耶和华为要应验藉 耶利米 的口所说的话，就激发 波斯 王 居鲁士 的心，使他下诏书通告全国，说：
2CHR|36|23|“ 波斯 王 居鲁士 如此说：耶和华－天上的上帝已将地上万国赐给我，又委派我在 犹大 的 耶路撒冷 为他建造殿宇。你们中间凡作他子民的可以上去，愿耶和华－他的上帝与他同在。”
EZRA|1|1|波斯 王 居鲁士 元年，耶和华为要应验藉 耶利米 的口所说的话，就激发 波斯 王 居鲁士 的心，使他下诏书通告全国，说：
EZRA|1|2|“ 波斯 王 居鲁士 如此说：耶和华天上的上帝已将地上万国赐给我，又委派我在 犹大 的 耶路撒冷 为他建造殿宇。
EZRA|1|3|你们中间凡作他子民的，可以上 犹大 的 耶路撒冷 去，重建耶和华－ 以色列 上帝的殿，他是在 耶路撒冷 的上帝；愿上帝与这人同在。
EZRA|1|4|凡存留的人，无论寄居何处，那地的人要用金银、财物、牲畜帮助他，还要为 耶路撒冷 上帝的殿甘心献上礼物。”
EZRA|1|5|于是， 犹大 和 便雅悯 的族长、祭司、 利未 人，凡是心被上帝感动的人都起来，要上 耶路撒冷 去建造耶和华的殿。
EZRA|1|6|四围所有的人都拿银器 、金子、财物、牲畜、珍宝支持他们 ，此外还有甘心献的一切礼物 。
EZRA|1|7|居鲁士 王也把耶和华殿的器皿拿出来，这些器皿是 尼布甲尼撒 从 耶路撒冷 掠取，放在自己神明庙中的。
EZRA|1|8|波斯 王 居鲁士 派 米提利达 司库把这些器皿拿出来，点交给 犹大 的领袖 设巴萨 。
EZRA|1|9|它们的数目如下：金盘三十个，银盘一千个，刀二十九把，
EZRA|1|10|金碗三十个，备用银碗四百一十个，其他器皿一千件。
EZRA|1|11|金银器皿共有五千四百件。被掳的人从 巴比伦 上 耶路撒冷 的时候， 设巴萨 把这一切都带了上来。
EZRA|2|1|这些是从被掳之地上来的省民， 巴比伦 王 尼布甲尼撒 把他们掳到 巴比伦 ，他们重返 耶路撒冷 和 犹大 ，各归本城。
EZRA|2|2|他们是同 所罗巴伯 、 耶书亚 、 尼希米 、 西莱雅 、 利来雅 、 末底改 、 必珊 、 米斯拔 、 比革瓦伊 、 利宏 、 巴拿 一起回来的。 以色列 百姓的人数如下：
EZRA|2|3|巴录 的子孙二千一百七十二名；
EZRA|2|4|示法提雅 的子孙三百七十二名；
EZRA|2|5|亚拉 的子孙七百七十五名；
EZRA|2|6|巴哈．摩押 的后裔，就是 耶书亚 和 约押 的子孙二千八百一十二名；
EZRA|2|7|以拦 的子孙一千二百五十四名；
EZRA|2|8|萨土 的子孙九百四十五名；
EZRA|2|9|萨改 的子孙七百六十名；
EZRA|2|10|巴尼 的子孙六百四十二名；
EZRA|2|11|比拜 的子孙六百二十三名；
EZRA|2|12|押甲 的子孙一千二百二十二名；
EZRA|2|13|亚多尼干 的子孙六百六十六名；
EZRA|2|14|比革瓦伊 的子孙二千零五十六名；
EZRA|2|15|亚丁 的子孙四百五十四名；
EZRA|2|16|亚特 的后裔，就是 希西家 的子孙九十八名；
EZRA|2|17|比赛 的子孙三百二十三名；
EZRA|2|18|约拉 的子孙一百一十二名；
EZRA|2|19|哈顺 的子孙二百二十三名；
EZRA|2|20|吉罢珥 人九十五名；
EZRA|2|21|伯利恒 人一百二十三名；
EZRA|2|22|尼陀法 人五十六名；
EZRA|2|23|亚拿突 人一百二十八名；
EZRA|2|24|亚斯玛弗 人四十二名；
EZRA|2|25|基列．耶琳 人、 基非拉 人、 比录 人共七百四十三名；
EZRA|2|26|拉玛 人和 迦巴 人共六百二十一名；
EZRA|2|27|默玛 人一百二十二名；
EZRA|2|28|伯特利 人和 艾 人共二百二十三名；
EZRA|2|29|尼波 人五十二名；
EZRA|2|30|末必 人一百五十六名；
EZRA|2|31|另一个 以拦 的子孙一千二百五十四名；
EZRA|2|32|哈琳 的子孙三百二十名；
EZRA|2|33|罗德 人、 哈第 人、 阿挪 人共七百二十五名；
EZRA|2|34|耶利哥 人三百四十五名；
EZRA|2|35|西拿 人三千六百三十名。
EZRA|2|36|祭司： 耶书亚 家 耶大雅 的子孙九百七十三名；
EZRA|2|37|音麦 的子孙一千零五十二名；
EZRA|2|38|巴施户珥 的子孙一千二百四十七名；
EZRA|2|39|哈琳 的子孙一千零一十七名。
EZRA|2|40|利未 人： 何达威雅 的后裔，就是 耶书亚 和 甲篾 的子孙七十四名。
EZRA|2|41|歌唱的： 亚萨 的子孙一百二十八名。
EZRA|2|42|门口的守卫： 沙龙 的子孙、 亚特 的子孙、 达们 的子孙、 亚谷 的子孙、 哈底大 的子孙、 朔拜 的子孙，共一百三十九名。
EZRA|2|43|殿役： 西哈 的子孙、 哈苏巴 的子孙、 答巴俄 的子孙、
EZRA|2|44|基绿 的子孙、 西亚 的子孙、 巴顿 的子孙、
EZRA|2|45|利巴拿 的子孙、 哈迦巴 的子孙、 亚谷 的子孙、
EZRA|2|46|哈甲 的子孙、 萨买 的子孙、 哈难 的子孙、
EZRA|2|47|吉德 的子孙、 迦哈 的子孙、 利亚雅 的子孙、
EZRA|2|48|利汛 的子孙、 尼哥大 的子孙、 迦散 的子孙、
EZRA|2|49|乌撒 的子孙、 巴西亚 的子孙、 比赛 的子孙、
EZRA|2|50|押拿 的子孙、 米乌宁 的子孙、 尼普心 的子孙、
EZRA|2|51|巴卜 的子孙、 哈古巴 的子孙、 哈忽 的子孙、
EZRA|2|52|巴洗律 的子孙、 米希大 的子孙、 哈沙 的子孙、
EZRA|2|53|巴柯 的子孙、 西西拉 的子孙、 答玛 的子孙、
EZRA|2|54|尼细亚 的子孙、 哈提法 的子孙。
EZRA|2|55|所罗门 仆人的后裔： 琐太 的子孙、 琐斐列 的子孙、 比路大 的子孙、
EZRA|2|56|雅拉 的子孙、 达昆 的子孙、 吉德 的子孙、
EZRA|2|57|示法提雅 的子孙、 哈替 的子孙、 玻黑列．哈斯巴音 的子孙、 亚米 的子孙。
EZRA|2|58|殿役和 所罗门 仆人的后裔共三百九十二名。
EZRA|2|59|从 特．米拉 、 特．哈萨 、 基绿 、 亚顿 、 音麦 上来，不能证明他们的父系家族和后裔是否属 以色列 的如下：
EZRA|2|60|第莱雅 的子孙、 多比雅 的子孙、 尼哥大 的子孙，共六百五十二名。
EZRA|2|61|祭司中， 哈巴雅 的子孙、 哈哥斯 的子孙、 巴西莱 的子孙， 巴西莱 因为娶了 基列 人 巴西莱 的女儿为妻，所以就以此为名。
EZRA|2|62|这些人在族谱之中寻查自己的谱系，却寻不着，因此算为不洁，不得作祭司。
EZRA|2|63|省长对他们说，不可吃至圣的物，直到有会用乌陵和土明的祭司兴起来。
EZRA|2|64|全会众共有四万二千三百六十名。
EZRA|2|65|此外，还有他们的仆婢七千三百三十七名，又有歌唱的男女二百名。
EZRA|2|66|他们有七百三十六匹马，二百四十五匹骡子，
EZRA|2|67|四百三十五匹骆驼，六千七百二十匹驴。
EZRA|2|68|有些族长到了 耶路撒冷 耶和华的殿，为上帝的殿甘心献上礼物，要在原有的根基上重新建造。
EZRA|2|69|他们量力捐入工程的库房，有六万一千达利克 金子，五千弥那银子，以及一百件祭司的礼服。
EZRA|2|70|于是祭司、 利未 人、百姓中的一些人、歌唱的、门口的守卫、殿役，各住在自己的城里； 以色列 众人都住在自己的城里。
EZRA|3|1|到了七月， 以色列 人住在自己的城里；那时他们如同一人，聚集在 耶路撒冷 。
EZRA|3|2|约萨达 的儿子 耶书亚 和他的弟兄众祭司，以及 撒拉铁 的儿子 所罗巴伯 和他的弟兄，都起来建筑 以色列 上帝的坛，要照神人 摩西 律法书上所写的，在坛上献燔祭。
EZRA|3|3|他们在原有的根基上筑坛，因为他们惧怕邻邦民族，又在其上向耶和华早晚献燔祭，
EZRA|3|4|并照律法书上所写的守住棚节，按数照例每日献所当献的燔祭。
EZRA|3|5|此后，他们献常献的燔祭，并在初一和耶和华一切分别为圣的节期献祭，又向耶和华献各人的甘心祭。
EZRA|3|6|从七月初一起，虽然耶和华殿的根基尚未立定，他们开始向耶和华献燔祭。
EZRA|3|7|他们把银子给石匠、木匠，把粮食、酒、油给 西顿 人、 推罗 人，好将香柏树从 黎巴嫩 浮海运到 约帕 ，是照 波斯 王 居鲁士 所允准他们的。
EZRA|3|8|他们到了 耶路撒冷 上帝殿的第二年，二月的时候， 撒拉铁 的儿子 所罗巴伯 ， 约萨达 的儿子 耶书亚 和其余的弟兄，就是祭司和 利未 人，以及所有被掳归回 耶路撒冷 的人，就开工建造；他们派二十岁以上的 利未 人，监督建造耶和华殿的工作。
EZRA|3|9|于是 何达威雅 的后裔，就是 耶书亚 和他的子孙与弟兄、 甲篾 和他的子孙，他们和 利未 人 希拿达 的子孙与弟兄，都起来如同一人，监督那些在上帝殿里做工的人。
EZRA|3|10|工匠立耶和华殿根基的时候，祭司穿礼服吹号， 利未 人 亚萨 的子孙敲钹，都照 以色列 王 大卫 亲手所定的，站着赞美耶和华。
EZRA|3|11|他们彼此唱和，赞美称谢耶和华： “他本为善， 他向 以色列 永施慈爱。” 他们赞美耶和华的时候，众百姓大声呼喊，因为耶和华殿的根基已经立定。
EZRA|3|12|然而有许多祭司、 利未 人和族长，就是见过先前那殿的老年人，现在亲眼看见这殿立了根基，就大声哭号，也有许多人大声欢呼，
EZRA|3|13|百姓不能分辨欢呼的声音或哭号的声音，因为百姓大声呼喊，声音连远处都可听到。
EZRA|4|1|犹大 和 便雅悯 的敌人听说被掳归回的人为耶和华－ 以色列 的上帝建造殿宇，
EZRA|4|2|就去见 所罗巴伯 和族长，对他们说：“请让我们与你们一同建造，因为我们也与你们一样寻求你们的上帝。自从 亚述 王 以撒．哈顿 带我们上这地的日子以来，我们常向上帝献祭。”
EZRA|4|3|但 所罗巴伯 、 耶书亚 和其余 以色列 的族长对他们说：“我们建造上帝的殿与你们无关，因为我们要照 波斯 王 居鲁士 所吩咐的，自己为耶和华－ 以色列 的上帝协力建造。”
EZRA|4|4|那地的人就在 犹大 百姓建造的时候，使他们的手发软，扰乱他们。
EZRA|4|5|从 波斯 王 居鲁士 年间，直到 波斯 王 大流士 在位的时候，那些人贿赂谋士，要破坏他们的计划。
EZRA|4|6|亚哈随鲁 在位，他的国度刚开始的时候，他们上书控告 犹大 和 耶路撒冷 的居民。
EZRA|4|7|亚达薛西 年间， 比施兰 、 米特利达 、 他别 和他们 的同僚上书奏告 波斯 王 亚达薛西 。奏文是用 亚兰 文写的，以 亚兰 文呈上。
EZRA|4|8|利宏 省长、 伸帅 书记也上奏 亚达薛西 王，控告 耶路撒冷 如下
EZRA|4|9|（那时， 利宏 省长、 伸帅 书记和他们其余的同僚，法官、官员、军官、 波斯 官员 、 亚基卫 人、 巴比伦 人，和 书珊迦 人，就是 以拦 人 ，
EZRA|4|10|以及被 亚斯那巴 大人迁移、安置在 撒玛利亚城 和 大河 西边一带地方其余的人。现在 ，
EZRA|4|11|这是他们上奏 亚达薛西 王奏文的抄本）：“ 河西 的臣仆上奏 亚达薛西 王，现在
EZRA|4|12|请王知道，从王那里上到我们这里的 犹太 人，已经抵达 耶路撒冷 。他们正在重建这反叛恶劣的城，已经完成了城墙，正要修复根基。
EZRA|4|13|如今请王知道，这城若再建造，城墙完工，他们就不再进贡、纳粮、缴税，王的国库必受亏损。
EZRA|4|14|如今，我们吃的盐既然全是宫廷的盐，就不忍见王吃亏，因此奏告于王，
EZRA|4|15|请王考察先王史籍，必会在史籍上查知这城是反叛的城，对列王和各省有害；自古以来，城中常有悖逆的事，因此这城曾被拆毁。
EZRA|4|16|我们谨奏王知，这城若再建造，城墙完工， 河西 之地王就无份了。”
EZRA|4|17|那时王谕覆 利宏 省长、 伸帅 书记和他们其余的同僚，就是住 撒玛利亚 和 河西 一带地方的人，说：“愿你们平安。现在
EZRA|4|18|你们所呈给我们的奏本，已经清楚地在我面前读了。
EZRA|4|19|我已下令考查，得知这城自古以来果然背叛列王，其中常有反叛悖逆的事。
EZRA|4|20|也曾有强大的君王治理 耶路撒冷 ，统管 河西 全地，人就给他们进贡、纳粮、缴税。
EZRA|4|21|现在你们要下令叫这些人停工，使这城不得建造，等到我再降旨。
EZRA|4|22|你们当谨慎办这事，不可迟延，何必让损害加重，使王受亏损呢？”
EZRA|4|23|亚达薛西 王上谕的抄本在 利宏 和 伸帅 书记，以及他们的同僚面前宣读，他们就急忙往 耶路撒冷 去见 犹太 人，用势力和强权叫他们停工。
EZRA|4|24|于是，在 耶路撒冷 上帝殿的工程就停止了，直停到 波斯 王 大流士 第二年。
EZRA|5|1|那时， 哈该 先知和 易多 的孙子 撒迦利亚 ，两个先知奉 以色列 上帝的名向 犹大 和 耶路撒冷 的 犹太 人说预言。
EZRA|5|2|于是 撒拉铁 的儿子 所罗巴伯 和 约萨达 的儿子 耶书亚 起来，开始建造 耶路撒冷 上帝的殿，有上帝的先知在那里帮助他们。
EZRA|5|3|当时 河西 的 达乃 总督和 示他．波斯乃 ，以及他们的同僚来对 犹太 人这样说：“谁降旨让你们建造这殿，完成这建筑呢？”
EZRA|5|4|于是我们告诉他们建造这建筑物的人叫什么名字。
EZRA|5|5|但上帝的眼目看顾 犹太 人的长老，以致没有人叫他们停工，直到奏文上告 大流士 ，得着他对这事的回谕。
EZRA|5|6|这是 河西 的 达乃 总督和 示他．波斯乃 ，以及他们的同僚，就是住 河西 的官员 ，上书奏告 大流士 王的抄本，
EZRA|5|7|他们上书给王的奏文，其中写着：“愿 大流士 王诸事平安。
EZRA|5|8|请王知道，我们往 犹大 省去，到了至大上帝的殿。这殿是用凿成的石头建造的，梁木插入墙内。这项工程进行迅速，在他们手中顺利。
EZRA|5|9|于是我们问那些长老，对他们这样说：‘谁降旨让你们建造这殿，完成这建筑呢？’
EZRA|5|10|我们又问他们的名字，要记下他们领袖的名字，奏告于王。
EZRA|5|11|他们这样回答我们说：‘我们是天和地之上帝的仆人，重建多年前所建造的殿，就是 以色列 一位伟大的君王建造完成的。
EZRA|5|12|但因我们祖先惹天上的上帝发怒，上帝把他们交在 迦勒底 人 巴比伦 王 尼布甲尼撒 的手中，他就拆毁这殿，又把百姓掳到 巴比伦 。
EZRA|5|13|然而 巴比伦 王 居鲁士 元年，他降旨允准建造上帝的这殿。
EZRA|5|14|上帝殿中的金银器皿，就是 尼布甲尼撒 从 耶路撒冷 殿中掠取带到 巴比伦 庙里的， 居鲁士 王从 巴比伦 庙里取出来，交给派为省长，名叫 设巴萨 的，
EZRA|5|15|对他说：可以将这些器皿带去，放在 耶路撒冷 的殿中，在原处建造上帝的殿。
EZRA|5|16|于是那位 设巴萨 来建立 耶路撒冷 上帝殿的根基。但从那时直到如今，这殿尚未修建完毕。’
EZRA|5|17|现在，王若以为好，请查阅 巴比伦 王的档案库，看 居鲁士 王有没有降旨允准在 耶路撒冷 建造上帝的殿。请降旨指示我们王对这件事的心意。”
EZRA|6|1|于是 大流士 王降旨，要寻察典籍库，就是在 巴比伦 藏档案之处；
EZRA|6|2|在 玛代 省 亚马他城 的宫内寻得一卷，其中这样写着，“纪录如下：
EZRA|6|3|居鲁士 王元年，王降旨论到在 耶路撒冷 上帝的殿，要建造这殿作为献祭之处，坚固它的根基。殿高六十肘，宽六十肘，
EZRA|6|4|要用三层凿成的石头，一层木头 ，经费可出于王的库房。
EZRA|6|5|至于上帝殿的金银器皿，就是 尼布甲尼撒 从 耶路撒冷 的殿中掠取带到 巴比伦 的，必须归还，带回 耶路撒冷 的殿中，各按原处放在上帝的殿里。”
EZRA|6|6|“现在， 河西 的 达乃 总督和 示他．波斯乃 ，以及他们的同僚，就是住 河西 的官员，你们当远离那里。
EZRA|6|7|不要拦阻这上帝殿的工作，任由 犹太 人的省长和长老在原处建造上帝的这殿。
EZRA|6|8|我又降旨，吩咐你们为建造上帝的殿当向 犹太 人的长老这样行：从王的财产中，由 河西 所缴纳的贡银，迅速支付这些人，免得工程停顿。
EZRA|6|9|他们向天上的上帝献燔祭所需用的公牛犊、公绵羊、小绵羊，以及麦子、盐、酒、油，都要照 耶路撒冷 祭司的话，每日供给他们，不得有误；
EZRA|6|10|好叫他们献馨香的祭给天上的上帝，又为王和王众子的寿命祈祷。
EZRA|6|11|我再降旨，无论谁更改这命令，必从他房屋中拆出一根梁木，把他举起，悬在其上，又使他的房屋为此成为粪堆。
EZRA|6|12|任何王或百姓若伸手更改这命令，拆毁在 耶路撒冷 上帝的这殿，愿那立他名在那里的上帝将他们灭绝。我 大流士 降这谕旨，你们要速速遵行。”
EZRA|6|13|于是， 河西 的 达乃 总督和 示他．波斯乃 ，以及他们的同僚，急速遵行 大流士 王所颁的命令。
EZRA|6|14|犹太 人的长老因 哈该 先知和 易多 的孙子 撒迦利亚 的预言，就建造这殿，凡事顺利。他们遵照 以色列 上帝的命令和 波斯 王 居鲁士 、 大流士 、 亚达薛西 的谕旨，建造完毕。
EZRA|6|15|大流士 王第六年，亚达月初三，这殿完工了。
EZRA|6|16|以色列 人、祭司和 利未 人，以及其余被掳归回的人都欢欢喜喜地为上帝的这殿行奉献礼。
EZRA|6|17|他们为这上帝殿的奉献礼献了一百头公牛，二百只公绵羊，四百只小绵羊，又照 以色列 支派的数目献十二只公山羊，作 以色列 众人的赎罪祭。
EZRA|6|18|他们派祭司按着班次， 利未 人也按着班次在 耶路撒冷 事奉上帝，正如 摩西 律法书上所写的。
EZRA|6|19|正月十四日，被掳归回的人守逾越节。
EZRA|6|20|祭司和 利未 人一同自洁，他们全都洁净了。 利未 人为被掳归回的众人和他们的弟兄众祭司，并为自己宰逾越节的羔羊。
EZRA|6|21|从被掳之地归回的 以色列 人，并所有归附他们、除掉这地外邦人的污秽、寻求耶和华－ 以色列 上帝的人，都吃这羔羊。
EZRA|6|22|他们欢欢喜喜地守除酵节七日，因为耶和华使他们欢喜。耶和华又使 亚述 王的心转向他们，坚固他们的手，去做上帝－ 以色列 上帝殿的工。
EZRA|7|1|这些事以后， 波斯 王 亚达薛西 在位的时候，有个人叫 以斯拉 ，他是 西莱雅 的儿子， 西莱雅 是 亚撒利雅 的儿子， 亚撒利雅 是 希勒家 的儿子，
EZRA|7|2|希勒家 是 沙龙 的儿子， 沙龙 是 撒督 的儿子， 撒督 是 亚希突 的儿子，
EZRA|7|3|亚希突 是 亚玛利雅 的儿子， 亚玛利雅 是 亚撒利雅 的儿子， 亚撒利雅 是 米拉约 的儿子，
EZRA|7|4|米拉约 是 西拉希雅 的儿子， 西拉希雅 是 乌西 的儿子， 乌西 是 布基 的儿子，
EZRA|7|5|布基 是 亚比书 的儿子， 亚比书 是 非尼哈 的儿子， 非尼哈 是 以利亚撒 的儿子， 以利亚撒 是 亚伦 大祭司的儿子。
EZRA|7|6|这 以斯拉 从 巴比伦 上来，他是一个文士，精通耶和华－ 以色列 上帝所赐 摩西 的律法。王允准他一切所求的，因为耶和华－他上帝的手帮助他。
EZRA|7|7|亚达薛西 王第七年，有些 以色列 人、一些祭司、 利未 人、歌唱的、门口的守卫、殿役，上 耶路撒冷 去。
EZRA|7|8|王第七年五月， 以斯拉 到了 耶路撒冷 。
EZRA|7|9|正月初一，他从 巴比伦 起程，五月初一就到了 耶路撒冷 ，因为他上帝施恩的手帮助他。
EZRA|7|10|以斯拉 立志考究遵行耶和华的律法，又将律例典章教导 以色列 人。
EZRA|7|11|亚达薛西 王赐给精通耶和华诫命和 以色列 律例的文士 以斯拉 祭司的谕旨，抄本如下：
EZRA|7|12|“诸王之王 亚达薛西 ，达于精通天上之上帝律法的 以斯拉 祭司文士等等：现在
EZRA|7|13|住在我国中的 以色列 百姓、祭司、 利未 人，凡愿意上 耶路撒冷 去的，我降旨准他们与你同去。
EZRA|7|14|既然王与七个谋士派你去，照你手中上帝的律法视察 犹大 和 耶路撒冷 的景况；
EZRA|7|15|你又带着王和谋士乐意献给住 耶路撒冷 、 以色列 上帝的金银，
EZRA|7|16|和你在 巴比伦 全省所得的一切金银，以及百姓、祭司甘心献给 耶路撒冷 他们上帝殿的礼物，
EZRA|7|17|那么，你就当用这银子急速买公牛、公绵羊、小绵羊，和同献的素祭、浇酒祭，献在 耶路撒冷 你们上帝殿的坛上。
EZRA|7|18|剩下的金银，你和你的弟兄看怎样好，就怎样用，但总要遵照你们上帝的旨意。
EZRA|7|19|你要带着交托给你、在上帝殿中事奉用的器皿，到 耶路撒冷 上帝面前。
EZRA|7|20|你上帝殿里若再有需用的经费，是你负责供应的，可以从王的宝库里支取。
EZRA|7|21|“我 亚达薛西 王又降旨达于 河西 所有的司库：‘精通天上之上帝律法的 以斯拉 祭司文士无论向你们要什么，你们要速速办理，
EZRA|7|22|直至一百他连得银子，一百柯珥 麦子，一百罢特酒，一百罢特油，盐不限其数。
EZRA|7|23|凡天上之上帝所吩咐的，当为天上之上帝的殿切实办理。何必使愤怒临到王和王众子的国呢？
EZRA|7|24|我再吩咐你们：至于任何祭司、 利未 人、歌唱的、门口的守卫和殿役，以及在上帝的这殿事奉的人，不可要求他们进贡，纳粮，缴税。’
EZRA|7|25|“你， 以斯拉 啊，要照着你上帝赐你的智慧，指派所有明白你上帝律法的人作官长、审判官，治理 河西 所有的百姓，教导不明白上帝律法的人。
EZRA|7|26|凡不遵行你上帝律法和王命令的人，当速速定他的罪，或处死，或充军，或抄家，或囚禁。”
EZRA|7|27|以斯拉 说：“耶和华－我们列祖的上帝是应当称颂的！因他使王起这心愿，使 耶路撒冷 耶和华的殿得荣耀，
EZRA|7|28|他又在王和谋士，以及王所有大能的军官面前施恩于我。我因耶和华－我上帝的手的帮助，得以坚强，从 以色列 中召集领袖，与我一同上来。”
EZRA|8|1|这些是 亚达薛西 王在位的时候，同我从 巴比伦 上来的族长和他们的家谱：
EZRA|8|2|属 非尼哈 的子孙有 革顺 ；属 以他玛 的子孙有 但以理 ；属 大卫 的子孙有 哈突 ；
EZRA|8|3|属 示迦尼 的子孙；属 巴录 的子孙有 撒迦利亚 ，同着他按家谱计算，男丁一百五十人；
EZRA|8|4|属 巴哈．摩押 的子孙有 西拉希雅 的儿子 以利约乃 ，同着他有男丁二百人；
EZRA|8|5|属 萨土 的子孙有 雅哈悉 的儿子 示迦尼 ，同着他有男丁三百人；
EZRA|8|6|属 亚丁 的子孙有 约拿单 的儿子 以别 ，同着他有男丁五十人；
EZRA|8|7|属 以拦 的子孙有 亚他利雅 的儿子 耶筛亚 ，同着他有男丁七十人；
EZRA|8|8|属 示法提雅 的子孙有 米迦勒 的儿子 西巴第雅 ，同着他有男丁八十人；
EZRA|8|9|属 约押 的子孙有 耶歇 的儿子 俄巴底亚 ，同着他有男丁二百一十八人；
EZRA|8|10|属 巴尼 的子孙有 约细斐 的儿子 示罗密 ，同着他有男丁一百六十人；
EZRA|8|11|属 比拜 的子孙有 比拜 的儿子 撒迦利亚 ，同着他有男丁二十八人；
EZRA|8|12|属 押甲 的子孙有 哈加坦 的儿子 约哈难 ，同着他有男丁一百一十人；
EZRA|8|13|属 亚多尼干 的子孙，就是晚到的，他们的名字是 以利法列 、 耶利 、 示玛雅 ，同着他们有男丁六十人；
EZRA|8|14|属 比革瓦伊 的子孙有 乌太 和 撒刻 ，同着他们有男丁七十人。
EZRA|8|15|我召集这些人在流入 亚哈瓦 的河旁边，我们在那里扎营三日。我查看百姓和祭司，发现并没有 利未 人在那里，
EZRA|8|16|就派人到 以利以谢 、 亚列 、 示玛雅 、 以利拿单 、 雅立 、 以利拿单 、 拿单 、 撒迦利亚 、 米书兰 等领袖，以及 约雅立 和 以利拿单 教师那里。
EZRA|8|17|我吩咐他们往 迦西斐雅 地方去见那里的领袖 易多 ，又告诉他们当向 易多 和他的弟兄，就是 迦西斐雅 那地方的殿役说什么话，好为我们上帝的殿带事奉的人来。
EZRA|8|18|蒙我们上帝施恩的手帮助我们，他们在 以色列 的曾孙， 利未 的孙子， 抹利 的后裔中带了一个精明的人来，就是 示利比 ，还有他的众子与兄弟共十八人。
EZRA|8|19|另外，还有 哈沙比雅 ，同着他有 米拉利 的子孙 耶筛亚 ，以及他的众子和兄弟共二十人。
EZRA|8|20|从前 大卫 和众领袖派殿役服事 利未 人，现在从这殿役中也带了二百二十人来，全都是按名指定的。
EZRA|8|21|那时，我在 亚哈瓦河 边宣告禁食，为要在我们上帝面前刻苦己心，求他使我们和我们的孩子，以及一切所有的，都得平坦的道路。
EZRA|8|22|我以求王拨步兵骑兵帮助我们抵挡路上的仇敌为羞愧，因我们曾对王说：“我们上帝施恩的手必帮助凡寻求他的，但他的能力和愤怒必攻击凡离弃他的。”
EZRA|8|23|我们为此禁食祈求我们的上帝，他就应允我们。
EZRA|8|24|我分派十二位祭司长，就是 示利比 、 哈沙比雅 和与他们一起的兄弟十人，
EZRA|8|25|把王和谋士、军官，并在那里的 以色列 众人为我们上帝殿所献的金银和器皿，都秤了交给他们。
EZRA|8|26|我秤了交在他们手中的有六百五十他连得银子，一百他连得银器，一百他连得金子，
EZRA|8|27|二十个金碗，值一千达利克，上等光亮的铜器皿两个，珍贵如金。
EZRA|8|28|我对他们说：“你们归耶和华为圣，器皿也归为圣；金银是甘心献给耶和华－你们列祖之上帝的。
EZRA|8|29|你们要警醒看守，直到你们在祭司长和 利未 族长，以及 以色列 的各族长面前，在 耶路撒冷 耶和华殿的库房内，把这些过了秤。”
EZRA|8|30|于是，祭司和 利未 人把秤过的金银和器皿接过来，要带到 耶路撒冷 我们上帝的殿里。
EZRA|8|31|正月十二日，我们从 亚哈瓦河 边起行，要往 耶路撒冷 去。我们上帝的手保佑我们，救我们脱离仇敌和路上埋伏之人的手。
EZRA|8|32|我们到了 耶路撒冷 ，在那里住了三日。
EZRA|8|33|第四日，金银和器皿都在我们上帝的殿里过了秤，交在 乌利亚 的儿子 米利末 祭司的手中。同着他的有 非尼哈 的儿子 以利亚撒 ，还有 利未 人 耶书亚 的儿子 约撒拔 和 宾内 的儿子 挪亚底 。
EZRA|8|34|那时，这一切都点过秤过了，重量全写在册上。
EZRA|8|35|从被掳之地归回的人向 以色列 的上帝献燔祭，为 以色列 众人献十二头公牛，九十六只公绵羊，七十七只小绵羊，又献十二只公山羊作赎罪祭，这些全都是献给耶和华的燔祭。
EZRA|8|36|被掳归回的人把王的谕旨交给王的总督与 河西 的省长，他们就支助百姓和上帝的殿。
EZRA|9|1|这些事完成以后，众领袖来接近我，说：“ 以色列 百姓、祭司和 利未 人没有弃绝 迦南 人、 赫 人、 比利洗 人、 耶布斯 人、 亚扪 人、 摩押 人、 埃及 人和 亚摩利 人等列邦民族所行可憎的事。
EZRA|9|2|因他们为自己和儿子娶了这些外邦女子，以致圣洁的种籽和列邦民族混杂，而且领袖和官长在这事上是罪魁。”
EZRA|9|3|我一听见这事，就撕裂衣服和外袍，拔了头发和胡须，惊惶地坐着。
EZRA|9|4|凡为 以色列 上帝言语战兢的人，都因被掳归回之人所犯的罪，聚集到我这里来。我惊惶地坐着，直到献晚祭的时候。
EZRA|9|5|献晚祭的时候我从愁烦中起来，穿着撕裂的衣服和外袍，双膝跪下，向耶和华－我的上帝举手，
EZRA|9|6|说： “我的上帝啊，我抱愧蒙羞，不敢向你－我的上帝仰面，因为我们的罪孽多到灭顶，我们的罪恶滔天。
EZRA|9|7|从我们祖先的日子直到今日，我们的罪恶深重；因我们的罪孽，我们和君王、祭司都交在邻国诸王的手中，被杀害，掳掠，抢夺，脸上蒙羞，正如今日的景况。
EZRA|9|8|现在耶和华－我们的上帝暂且向我们施恩，为我们留下一些残存之民，使我们如钉子钉在他的圣所，好让我们的上帝光照我们的眼目，使我们在受辖制之中稍微复兴。
EZRA|9|9|我们是奴仆，然而在受辖制之中，我们的上帝没有丢弃我们，在 波斯 诸王面前向我们施恩，叫我们复兴，能重建我们上帝的殿，修补毁坏之处，使我们在 犹大 和 耶路撒冷 有城墙。
EZRA|9|10|“我们的上帝啊，既然如此，现在我们还有什么话可说呢？因为我们离弃了你的诫命，
EZRA|9|11|就是你藉你仆人众先知所吩咐的，说：‘你们要去得为业之地是污秽之地，因列邦民族的污秽和可憎的事，叫这地从这边到那边都充满了污秽。
EZRA|9|12|现在，不可把你们的女儿嫁给他们的儿子，也不可为你们的儿子娶他们的女儿，永不可求他们的平安和他们的利益，这样你们就可以强盛，吃这地的美物，并把这地留给你们的子孙永远为业。’
EZRA|9|13|我们因自己的恶行和大罪，遭遇这一切的事，但你－我们的上帝惩罚我们轻于我们罪所当得的，又为我们留下这些残存之民。
EZRA|9|14|我们岂可再违背你的诫命，与行这些可憎之事的民族结亲呢？若我们这样行，你岂不向我们发怒，将我们灭绝，以致没有一个余民或残存之民吗？
EZRA|9|15|耶和华－ 以色列 的上帝啊，你是公义的，我们才能剩下这些残存之民，正如今日的景况。看哪，我们在你面前有罪恶，因此无人能在你面前站立得住。”
EZRA|10|1|以斯拉 祷告，认罪，哭泣，俯伏在上帝殿前的时候，有 以色列 中的男女和孩童聚集到 以斯拉 那里，成了一个盛大的会，百姓无不痛哭。
EZRA|10|2|以拦 的子孙， 耶歇 的儿子 示迦尼 对 以斯拉 说：“我们娶了这地的外邦女子，干犯了我们的上帝，然而现在 以色列 人在这事上还有指望。
EZRA|10|3|现在，我们要与我们的上帝立约，送走所有的妻子和她们所生的，照着主和那些因我们上帝诫命战兢之人所议定的，按律法去行。
EZRA|10|4|起来，这是你当办的事，我们必支持你，你当奋勇而行。”
EZRA|10|5|以斯拉 就起来，叫祭司长和 利未 人，以及 以色列 众人起誓，要照这话去做；他们就起了誓。
EZRA|10|6|以斯拉 从上帝殿前起来，进入 以利亚实 的儿子 约哈难 的屋里，到了那里不吃饭，也不喝水，为被掳归回之人所犯的罪悲伤。
EZRA|10|7|他们通告 犹大 和 耶路撒冷 ，叫所有被掳归回的人聚集在 耶路撒冷 。
EZRA|10|8|凡不遵照领袖和长老所议定，三日之内不来的，就必毁坏他所有的财产，把他从被掳归回之人的会中开除。
EZRA|10|9|于是， 犹大 和 便雅悯 众人三日之内都聚集在 耶路撒冷 。那时是九月，那月的二十日，众百姓坐在上帝殿前的广场，因这事，又因下大雨，就都战抖。
EZRA|10|10|以斯拉 祭司站起来，对他们说：“你们有罪了，因为你们娶了外邦女子，增添 以色列 的罪恶。
EZRA|10|11|现在当向耶和华－你们列祖的上帝认罪，遵行他的旨意，离开这地的百姓和外邦女子。”
EZRA|10|12|全会众大声回答说：“好！我们必照着你的话去做。
EZRA|10|13|只是百姓众多，又逢大雨的季节，我们没有气力站在外面；这也不是一两天可以办完的事，因我们在这事上犯了大罪。
EZRA|10|14|让我们的领袖代表全会众留在那里。我们城镇中凡娶外邦女子的，当按所定的日期，会同本城的长老和审判官前来，直到办完这事，上帝的烈怒转离我们 。”
EZRA|10|15|惟有 亚撒黑 的儿子 约拿单 ， 特瓦 的儿子 雅哈谢 反对这事，并有 米书兰 和 利未 人 沙比太 支持他们。
EZRA|10|16|被掳归回的人就如此做了。 以斯拉 祭司按着父家指名选派一些族长 。十月初一，他们一同坐下来查办这事，
EZRA|10|17|到正月初一，才查清所有娶外邦女子的人数。
EZRA|10|18|在祭司中查出娶外邦女子的： 耶书亚 的子孙中，有 约萨达 的儿子，和他兄弟 玛西雅 、 以利以谢 、 雅立 、 基大利 ，
EZRA|10|19|他们承诺要送走他们的妻子。他们因有罪，就献羊群中的一只公绵羊赎罪；
EZRA|10|20|音麦 的子孙中，有 哈拿尼 、 西巴第雅 ；
EZRA|10|21|哈琳 的子孙中，有 玛西雅 、 以利雅 、 示玛雅 、 耶歇 、 乌西雅 ；
EZRA|10|22|巴施户珥 的子孙中，有 以利约乃 、 玛西雅 、 以实玛利 、 拿坦业 、 约撒拔 、 以利亚萨 。
EZRA|10|23|利未 人中，有 约撒拔 、 示每 、 基拉雅 ， 基拉雅 就是 基利他 ，还有 毗他希雅 、 犹大 、 以利以谢 。
EZRA|10|24|歌唱的人中有 以利亚实 。门口的守卫中，有 沙龙 、 提联 、 乌利 。
EZRA|10|25|以色列 人 巴录 的子孙中，有 拉米 、 耶西雅 、 玛基雅 、 米雅民 、 以利亚撒 、 玛基雅 、 比拿雅 。
EZRA|10|26|以拦 的子孙中，有 玛他尼 、 撒迦利亚 、 耶歇 、 押底 、 耶列末 、 以利雅 。
EZRA|10|27|萨土 的子孙中，有 以利约乃 、 以利亚实 、 玛他尼 、 耶列末 、 撒拔 、 亚西撒 。
EZRA|10|28|比拜 的子孙中，有 约哈难 、 哈拿尼雅 、 萨拜 、 亚勒 。
EZRA|10|29|巴尼 的子孙中，有 米书兰 、 玛鹿 、 亚大雅 、 雅述 、 示押 、 拉末 。
EZRA|10|30|巴哈．摩押 的子孙中，有 阿底拿 、 基拉 、 比拿雅 、 玛西雅 、 玛他尼 、 比撒列 、 宾内 、 玛拿西 。
EZRA|10|31|哈琳 的子孙中，有 以利以谢 、 伊示雅 、 玛基雅 、 示玛雅 、 西缅 、
EZRA|10|32|便雅悯 、 玛鹿 、 示玛利雅 。
EZRA|10|33|哈顺 的子孙中，有 玛特乃 、 玛达他 、 撒拔 、 以利法列 、 耶利买 、 玛拿西 、 示每 。
EZRA|10|34|巴尼 的子孙中，有 玛玳 、 暗兰 、 乌益 、
EZRA|10|35|比拿雅 、 比底雅 、 基禄 、
EZRA|10|36|瓦尼雅 、 米利末 、 以利亚实 、
EZRA|10|37|玛他尼 、 玛特乃 、 雅扫 、
EZRA|10|38|巴尼 、 宾内 、 示每 、
EZRA|10|39|示利米雅 、 拿单 、 亚大雅 、
EZRA|10|40|玛拿底拜 、 沙赛 、 沙赖 、
EZRA|10|41|亚萨利 、 示利米雅 、 示玛利雅 、
EZRA|10|42|沙龙 、 亚玛利雅 、 约瑟 。
EZRA|10|43|尼波 的子孙中，有 耶利 、 玛他提雅 、 撒拔 、 西比拿 、 雅玳 、 约珥 、 比拿雅 。
EZRA|10|44|这些人全都娶了外邦女子，其中也有生了儿女的 。
NEH|1|1|哈迦利亚 的儿子 尼希米 的言语如下： 亚达薛西 王二十年基斯流月，我在 书珊 城堡中。
NEH|1|2|那时，我有一个兄弟 哈拿尼 ，同几个人从 犹大 来。我问他们那些被掳归回、剩下残存的 犹太 人和 耶路撒冷 的情况。
NEH|1|3|他们对我说：“那些被掳归回剩下的余民在 犹大 省那里遭大难，受凌辱； 耶路撒冷 的城墙被拆毁，城门被火焚烧。”
NEH|1|4|我听见这话，就坐下哭泣，悲哀几日，在天上的上帝面前禁食祈祷，
NEH|1|5|说：“唉，耶和华－天上大而可畏的上帝，向爱你、守你诫命的人守约施慈爱的上帝啊，
NEH|1|6|愿你睁眼看，侧耳听你仆人今日昼夜在你面前，为你众仆人 以色列 人的祈祷，承认我们 以色列 人向你所犯的罪；我与我父家都犯了罪。
NEH|1|7|我们向你所行的非常败坏，没有遵守你吩咐你仆人 摩西 的诫命、律例、典章。
NEH|1|8|求你记念所吩咐你仆人 摩西 的话，说：‘你们若犯罪，我就把你们分散在万民中；
NEH|1|9|但你们若归向我，谨守遵行我的诫命，你们被赶散的人虽在天涯，我也必从那里将他们召集回来，带到我所选择立为我名居所的地方。’
NEH|1|10|他们是你的仆人和你的百姓，是你用大力和大能的手所救赎的。
NEH|1|11|唉，主啊，求你侧耳听你仆人的祈祷，听喜爱敬畏你名众仆人的祈祷，使你仆人今日亨通，在这人面前蒙恩。” 我是王的酒政。
NEH|2|1|亚达薛西 王二十年尼散月，酒摆在王面前 ，我拿起酒来奉给王。我在王面前从来没有愁容。
NEH|2|2|王对我说：“你既没有病，为什么面带愁容呢？这不是别的，必是你心中愁烦。”于是我非常惧怕。
NEH|2|3|我对王说：“愿王万岁！我祖先坟墓所在的那城荒凉，城门被火焚烧，我岂能面无愁容呢？”
NEH|2|4|王对我说：“你想求什么？”于是我向天上的上帝祈祷。
NEH|2|5|我对王说：“王若以为好，仆人若在王面前蒙宠爱，求王差遣我往 犹大 ，到我祖先坟墓所在的那城去，我好重新建造。”
NEH|2|6|那时王后坐在王的旁边，王对我说：“你要去多久？几时回来？”王看这事为好，就派我去。我给王定了日期。
NEH|2|7|我又对王说：“王若以为好，求王赐我诏书，通知 河西 的省长准我经过，直到 犹大 ；
NEH|2|8|又赐诏书，通知管理王园林的 亚萨 ，叫他给我木材，作为殿的营楼之门、城墙，和我自己要住的房屋的横梁。”王就允准我，因为我上帝施恩的手帮助我。
NEH|2|9|王派了军官和骑兵护送我。我到了 河西 的省长那里，将王的诏书交给他们。
NEH|2|10|和伦 人 参巴拉 和作臣仆的 亚扪 人 多比雅 ，听见有人来为 以色列 人争取利益，就很恼怒。
NEH|2|11|我到了 耶路撒冷 ，在那里停留了三天。
NEH|2|12|夜间我和跟随我的几个人起来；但上帝感动我心要为 耶路撒冷 做的事，我并没有告诉人。只有我自己骑的牲口，没有别的牲口在我那里。
NEH|2|13|当夜，我出了 谷门 ，往 野狗泉 去，到了 粪厂门 ，察看 耶路撒冷 的城墙，城墙被拆毁，城门被火焚烧。
NEH|2|14|我又往前，到了 泉门 ，又到 王池 ，但所骑的牲口没有地方可以过去。
NEH|2|15|于是我夜间沿溪而上，察看城墙，又转身进入 谷门 ，就回来了。
NEH|2|16|我往哪里去，我做什么事，官长都不知道。我也没有告诉 犹大 人、祭司、贵族、官长和其余做工的人。
NEH|2|17|以后，我对他们说：“我们所遭的难， 耶路撒冷 怎样荒凉，城门被火焚烧，你们都看见了。来吧，让我们重建 耶路撒冷 的城墙，免得再受凌辱！”
NEH|2|18|我告诉他们我上帝施恩的手怎样帮助我，以及王向我所说的话。他们就说：“我们起来建造吧！”于是他们使自己的手坚强，做这美好的工作。
NEH|2|19|但 和伦 人 参巴拉 、作臣仆的 亚扪 人 多比雅 和 阿拉伯 人 基善 听见就嗤笑我们，藐视我们，说：“你们所做的这事是什么呢？要背叛王吗？”
NEH|2|20|我回答他们的话，对他们说：“天上的上帝必使我们亨通。我们作他仆人的，要起来建造；你们却在 耶路撒冷 无份、无权、无名号 。”
NEH|3|1|那时， 以利亚实 大祭司和他的弟兄众祭司起来建立 羊门 ，将门分别为圣，安立门扇，直到 哈米亚楼 。他们又将它分别为圣，直到 哈楠业楼 。
NEH|3|2|在他旁边建造的是 耶利哥 人。在他旁边建造的是 音利 的儿子 撒刻 。
NEH|3|3|哈西拿 的子孙建立 鱼门 ，架横梁、安门扇，装闩和锁。
NEH|3|4|在他们旁边修造的是 哈哥斯 的孙子， 乌利亚 的儿子 米利末 。在他们旁边修造的是 米示萨别 的孙子， 比利迦 的儿子 米书兰 。在他们旁边修造的是 巴拿 的儿子 撒督 。
NEH|3|5|在他们旁边修造的是 提哥亚 人；但是他们的贵族不用肩 扛他们主人的工作。
NEH|3|6|巴西亚 的儿子 耶何耶大 与 比所玳 的儿子 米书兰 修造 古门 ，架横梁，安门扇，装闩和锁。
NEH|3|7|在他们旁边修造的是 基遍 人 米拉提 、 米伦 人 雅顿 、 基遍 人，和 河西 总督所管的 米斯巴 人。
NEH|3|8|在他旁边修造的是 哈海雅 的儿子 乌薛 银匠。在他旁边修造的是做香料的 哈拿尼雅 。他们修复 耶路撒冷 ，直到 宽墙 。
NEH|3|9|在他们旁边修造的是管理 耶路撒冷 城区的一半、 户珥 的儿子 利法雅 。
NEH|3|10|在他们旁边的是 哈路抹 的儿子 耶大雅 在自己房屋的对面修造。在他旁边修造的是 哈沙尼 的儿子 哈突 。
NEH|3|11|哈琳 的儿子 玛基雅 和 巴哈．摩押 的儿子 哈述 修造下一段和 炉楼 。
NEH|3|12|在他旁边修造的是管理 耶路撒冷 城区的另一半、 哈罗黑 的儿子 沙龙 和他的女儿们。
NEH|3|13|哈嫩 和 撒挪亚 的居民修造 谷门 ；他们立门，安门扇，装闩和锁，又修造城墙一千肘，直到 粪厂门 。
NEH|3|14|管理 伯．哈基琳 区、 利甲 的儿子 玛基雅 修造 粪厂门 ；他立门，安门扇，装闩和锁。
NEH|3|15|管理 米斯巴 区、 各．荷西 的儿子 沙仑 修造 泉门 ；他立门，盖门顶，安门扇，装闩和锁，又修造靠近王的花园 西罗亚池 的城墙，直到那从 大卫城 下来的台阶。
NEH|3|16|接续他修造的是管理 伯．夙 区的一半、 押卜 的儿子 尼希米 ，直到 大卫 坟地的对面，又到人造池，到达勇士的房屋。
NEH|3|17|接续他修造的是 利未 人 巴尼 的儿子 利宏 。在他旁边的是管理 基伊拉 区一半的 哈沙比雅 为本区修造。
NEH|3|18|接续他修造的是他们弟兄中管理 基伊拉 区的另一半、 希拿达 的儿子 宾内 。
NEH|3|19|在他旁边的是管理 米斯巴 、 耶书亚 的儿子 以谢珥 修造武库的上坡对面、城墙转弯处的那一段。
NEH|3|20|接续他的是 萨拜 的儿子 巴录 竭力修造下一段，从转弯处，直到 以利亚实 大祭司的府门。
NEH|3|21|接续他的是 哈哥斯 的孙子， 乌利亚 的儿子 米利末 修造下一段，从 以利亚实 的府门，直到 以利亚实 府的尽头。
NEH|3|22|接续他修造的是住平原的祭司。
NEH|3|23|接续他的是 便雅悯 与 哈述 在自己房屋的对面修造。接续他的是 亚难尼 的孙子， 玛西雅 的儿子 亚撒利雅 在自己房屋的旁边修造。
NEH|3|24|接续他的是 希拿达 的儿子 宾内 修造下一段，从 亚撒利雅 的房屋直到转弯处，又到城角。
NEH|3|25|乌赛 的儿子 巴拉 修造转弯处的对面和靠近护卫院、王宫上层凸出来的城楼。接续他的是 巴录 的儿子 毗大雅 ，
NEH|3|26|（殿役住在 俄斐勒 ，直到朝东 水门 的对面和凸出来的城楼。）
NEH|3|27|接续他的是 提哥亚 人又修造一段，对着那凸出来的大城楼，直到 俄斐勒 的城墙。
NEH|3|28|从 马门 往上，祭司各在自己房屋的对面修造。
NEH|3|29|接续他的是 音麦 的儿子 撒督 在自己房屋的对面修造。接续他修造的是 东门 的守卫、 示迦尼 的儿子 示玛雅 。
NEH|3|30|接续他的是 示利米雅 的儿子 哈拿尼雅 和 萨拉 的第六个儿子 哈嫩 修造下一段。接续他的是 比利迦 的儿子 米书兰 在自己房屋的对面修造。
NEH|3|31|接续他的是 玛基雅 银匠修造，直到殿役和商人的房屋，对着 集合门 ，直到角楼。
NEH|3|32|银匠与商人在角楼和 羊门 之间修造。
NEH|4|1|参巴拉 听见我们建造城墙就发怒，非常恼恨，并嗤笑 犹太 人。
NEH|4|2|他对他的弟兄和 撒玛利亚 的军兵说：“这些软弱的 犹太 人做什么呢？要为自己重建吗 ？要献祭吗？要一日完工吗？要使土堆里火烧过的石头再有用吗？”
NEH|4|3|亚扪 人 多比雅 在一旁说：“他们所修造的石墙，就是狐狸上去也必崩裂。”
NEH|4|4|我们的上帝啊，求你垂听，因为我们被藐视。求你使他们的毁谤归于他们自己头上，使他们在被掳之地成为掠物。
NEH|4|5|不要遮掩他们的罪孽，不要使他们的罪恶从你面前涂去，因为他们在修造的人前面惹你发怒。
NEH|4|6|这样，我们修造城墙，整个城墙就连接起来，到一半高，因为百姓一心做工。
NEH|4|7|参巴拉 、 多比雅 、 阿拉伯 人、 亚扪 人和 亚实突 人听见 耶路撒冷 城墙正在修造，破裂的地方开始进行修补，就非常愤怒。
NEH|4|8|大家同谋要来攻打 耶路撒冷 ，使城混乱。
NEH|4|9|然而，我们向我们的上帝祷告，又因他们的缘故，就派人站岗，昼夜防备他们。
NEH|4|10|但 犹大 有话说： “扛抬的人力气衰弱， 瓦砾太多， 我们自己不可能 建造城墙。”
NEH|4|11|我们的敌人说：“趁他们不知道，看不见的时候，我们进入他们中间，杀了他们，使工作停止。”
NEH|4|12|那靠近敌人居住的 犹太 人十次从各处来见我们，说：“你们必须回到我们那里。”
NEH|4|13|我叫百姓站在城墙后边低洼的空处，使百姓各按宗族站着，拿刀、拿枪、拿弓。
NEH|4|14|我察看了，就起来对贵族、官长和其余的百姓说：“不要怕他们！当记得主是大而可畏的。你们要为你们的弟兄、儿女、妻子、家园争战。”
NEH|4|15|仇敌听见我们知道了他们的计谋，上帝也破坏他们的计谋，我们就都回到城墙那里，各做各的工。
NEH|4|16|从那日起，我的仆人一半做工，一半拿枪、拿盾牌、拿弓、穿铠甲，官长都站在 犹大 全家的后边。
NEH|4|17|他们建造城墙；扛抬材料的人扛抬的时候，一手做工，一手拿兵器。
NEH|4|18|建造的人都腰间佩刀建造，吹角的人在我旁边。
NEH|4|19|我对贵族、官长和其余的百姓说：“这工程浩大，范围辽阔，我们在城墙上彼此相离很远。
NEH|4|20|你们一听见角声在哪里，就聚集到我们那里去。我们的上帝必为我们争战。”
NEH|4|21|于是，我们做这工程，一半的人拿枪，从天亮直到星宿出现的时候。
NEH|4|22|那时，我又对百姓说：“各人和他的仆人当在 耶路撒冷 过夜，好为我们夜间守卫，白昼做工。”
NEH|4|23|这样，我和弟兄仆人，以及跟从我的卫兵都不脱衣服，各人打水时 也拿着自己的兵器。
NEH|5|1|百姓和他们的妻子大大呼号，埋怨他们的弟兄 犹太 人。
NEH|5|2|有的说：“我们和儿女人口众多，必须得粮食吃，才能活下去。”
NEH|5|3|有的说：“我们典押了田地、葡萄园、房屋，才得粮食充饥。”
NEH|5|4|有的说：“我们借了钱付田地和葡萄园的税给王。
NEH|5|5|现在，我们的身体与我们弟兄的身体是一样的，我们的儿女与他们的儿女没有差别。看哪，我们却要迫使儿女作人的奴婢。我们有些女儿已被抢走了，我们却无能为力，因为我们的田地和葡萄园已经归了别人。”
NEH|5|6|我听见他们的呼号和这些话，就非常愤怒。
NEH|5|7|我心里作了决定，就斥责贵族和官长，对他们说：“你们各人借钱给弟兄，竟然索取利息！”于是我召开大会攻击他们。
NEH|5|8|我对他们说：“我们已尽力赎回我们的弟兄，就是卖到列国的 犹太 人；你们还要卖弟兄，让我们去买回来吗？”他们就静默不语，无话可答。
NEH|5|9|我又说：“你们做的这事不对！你们行事不是应该敬畏我们的上帝，免得列国我们的仇敌毁谤我们吗？
NEH|5|10|我和我的弟兄仆人也要把银钱粮食借给百姓，大家都当免除利息。
NEH|5|11|就在今日，你们要把他们的田地、葡萄园、橄榄园、房屋，以及向他们所取银钱的利息 、粮食、新酒和新油都归还他们。”
NEH|5|12|贵族和官长说：“我们必归还，不再向他们索取，必照你所说的去做。”我就召了祭司来，叫贵族和官长起誓，必照这话去做。
NEH|5|13|我也抖着胸前的衣袋，说：“凡不实行这话的，愿上帝照样抖他离开他的家和他劳碌得来的，直到抖空了。”全会众都说：“阿们！”又赞美耶和华。百姓就照着这话去做。
NEH|5|14|自从我奉派作 犹大 地省长的那日，就是从 亚达薛西 王二十年直到三十二年，共十二年之久，我与我弟兄都没有吃省长的俸禄。
NEH|5|15|在我以前的省长加重百姓的负担，向百姓索取粮食和酒，以及四十舍客勒银子 ，甚至他们的仆人也辖制百姓，但我因敬畏上帝不这样做。
NEH|5|16|我也努力修造城墙。我们并没有购置田地，我所有的仆人也都聚集在那里做工。
NEH|5|17|除了从四围列国来的人以外，有 犹太 人和官长一百五十人与我同席。
NEH|5|18|每日预备一头公牛，六只肥羊，又为我预备飞禽；每十日一次多多预备各样的酒。虽然如此，我并不索取省长的俸禄，因为这百姓负的劳役很重。
NEH|5|19|我的上帝啊，求你记念我为这百姓所做的一切，施恩于我。
NEH|6|1|参巴拉 、 多比雅 、 阿拉伯 人 基善 和我们其余的仇敌听见我已经建造了城墙，没有破裂之处在其中，那时我还没有在城门安门扇；
NEH|6|2|参巴拉 和 基善 就派人来见我，说：“请你来，我们在 阿挪 平原的村庄见面。”其实，他们想要害我。
NEH|6|3|于是我派使者到他们那里，说：“我正在进行大的工程，不能下去。我怎么能离开，下去见你们，而让工程停顿呢？”
NEH|6|4|他们这样派人来见我四次，我都用这话回答他们。
NEH|6|5|参巴拉 第五次同样派仆人来见我，手里拿着未封的信，
NEH|6|6|信上写着：“列国中有风声， 基善 也说，你和 犹太 人谋反，所以你建造城墙。据说，你要作他们的王，
NEH|6|7|并且你派先知在 耶路撒冷 指着你宣讲说，‘在 犹大 有王。’如今这些话必传给王知，现在请你来，我们一起商议。”
NEH|6|8|我就派人到他那里，说：“你所说的这些事，一概没有，是你心里捏造的。”
NEH|6|9|他们全都要使我们惧怕，说：“他们的手必软弱，不能工作，以致不能完工。”现在，求你坚固我的手。
NEH|6|10|我到了 米希大别 的孙子， 第来雅 的儿子 示玛雅 家里；那时，他闭门不出。他说：“我们可以在上帝的殿里，就在殿的中间会面，锁住殿门，因为他们要来杀你，要在夜里来杀你。”
NEH|6|11|我说：“像我这样的人岂会逃跑呢？像我这样的人岂能进入殿里保全生命呢？我不进去！”
NEH|6|12|我看清楚了，看哪，上帝并没有派他，是他自己说预言攻击我，是 多比雅 和 参巴拉 收买了他；
NEH|6|13|收买他的目的是要叫我惧怕，依从他犯罪，留下一个坏名声，好让他们毁谤我。
NEH|6|14|我的上帝啊，求你记得 多比雅 、 参巴拉 、 挪亚底 女先知和其余的先知，因他们行这些事，要叫我惧怕。
NEH|6|15|以禄月二十五日，城墙修完了，共修了五十二天。
NEH|6|16|我们所有的仇敌听见了，四围的列国就惧怕，愁眉不展，因为他们知道这工作得以完成，是出于我们的上帝。
NEH|6|17|而且，在那些日子， 犹大 的贵族屡次寄信给 多比雅 ， 多比雅 也回信给他们。
NEH|6|18|在 犹大 有许多人与 多比雅 结盟，因为他是 亚拉 的儿子 示迦尼 的女婿，并且他的儿子 约哈难 娶了 比利迦 的儿子 米书兰 的女儿。
NEH|6|19|他们也在我面前说 多比雅 的好话，又把我的话传给他。 多比雅 常寄信来，要叫我惧怕。
NEH|7|1|城墙修完，我安了门扇，门口的守卫、歌唱的和 利未 人都已派定。
NEH|7|2|我吩咐我的兄弟 哈拿尼 和城堡的官长 哈拿尼雅 管理 耶路撒冷 ，因为 哈拿尼雅 是一个忠信的人，敬畏上帝过于众人。
NEH|7|3|我对他们说：“等到太阳热的时候才可开 耶路撒冷 的城门；要派 耶路撒冷 的居民，各按班次在自己房屋的前面站岗。他们还在站岗的时候，就要关门上闩。”
NEH|7|4|城又宽又大，城中的百姓却稀少，房屋也还没有建造。
NEH|7|5|我的上帝感动我的心，我就召集贵族、官长和百姓，要登记家谱。我找到第一次上来之人的家谱，发现上面写着：
NEH|7|6|这些是从被掳之地上来的省民， 巴比伦 王 尼布甲尼撒 把他们掳去，他们重返 耶路撒冷 和 犹大 ，各归本城。
NEH|7|7|他们是同 所罗巴伯 、 耶书亚 、 尼希米 、 亚撒利雅 、 拉米 、 拿哈玛尼 、 末底改 、 必珊 、 米斯毗列 、 比革瓦伊 、 尼宏 、 巴拿 一起回来的。 以色列 百姓的人数如下：
NEH|7|8|巴录 的子孙二千一百七十二名；
NEH|7|9|示法提雅 的子孙三百七十二名；
NEH|7|10|亚拉 的子孙六百五十二名；
NEH|7|11|巴哈．摩押 的后裔，就是 耶书亚 和 约押 的子孙二千八百一十八名；
NEH|7|12|以拦 的子孙一千二百五十四名；
NEH|7|13|萨土 的子孙八百四十五名；
NEH|7|14|萨改 的子孙七百六十名；
NEH|7|15|宾内 的子孙六百四十八名；
NEH|7|16|比拜 的子孙六百二十八名；
NEH|7|17|押甲 的子孙二千三百二十二名；
NEH|7|18|亚多尼干 的子孙六百六十七名；
NEH|7|19|比革瓦伊 的子孙二千零六十七名；
NEH|7|20|亚丁 的子孙六百五十五名；
NEH|7|21|亚特 的后裔，就是 希西家 的子孙九十八名；
NEH|7|22|哈顺 的子孙三百二十八名；
NEH|7|23|比赛 的子孙三百二十四名；
NEH|7|24|哈拉 的子孙一百一十二名；
NEH|7|25|基遍 人九十五名；
NEH|7|26|伯利恒 人和 尼陀法 人共一百八十八名；
NEH|7|27|亚拿突 人一百二十八名；
NEH|7|28|伯．亚斯玛弗 人四十二名；
NEH|7|29|基列．耶琳 人、 基非拉 人、 比录 人共七百四十三名；
NEH|7|30|拉玛 人和 迦巴 人共六百二十一名；
NEH|7|31|默玛 人一百二十二名；
NEH|7|32|伯特利 人和 艾 人共一百二十三名；
NEH|7|33|别的 尼波 人五十二名；
NEH|7|34|另一个 以拦 子孙一千二百五十四名；
NEH|7|35|哈琳 的子孙三百二十名；
NEH|7|36|耶利哥 人三百四十五名；
NEH|7|37|罗德 人、 哈第 人、 阿挪 人共七百二十一名；
NEH|7|38|西拿 人三千九百三十名。
NEH|7|39|祭司： 耶书亚 家， 耶大雅 的子孙九百七十三名；
NEH|7|40|音麦 的子孙一千零五十二名；
NEH|7|41|巴施户珥 的子孙一千二百四十七名；
NEH|7|42|哈琳 的子孙一千零一十七名。
NEH|7|43|利未 人： 何达威 的后裔，就是 耶书亚 和 甲篾 的子孙七十四名。
NEH|7|44|歌唱的： 亚萨 的子孙一百四十八名。
NEH|7|45|门口的守卫： 沙龙 的子孙、 亚特 的子孙、 达们 的子孙、 亚谷 的子孙、 哈底大 的子孙、 朔拜 的子孙，共一百三十八名。
NEH|7|46|殿役： 西哈 的子孙、 哈苏巴 的子孙、 答巴俄 的子孙、
NEH|7|47|基绿 的子孙、 西亚 的子孙、 巴顿 的子孙、
NEH|7|48|利巴拿 的子孙、 哈迦巴 的子孙、 萨买 的子孙、
NEH|7|49|哈难 的子孙、 吉德 的子孙、 迦哈 的子孙、
NEH|7|50|利亚雅 的子孙、 利汛 的子孙、 尼哥大 的子孙、
NEH|7|51|迦散 的子孙、 乌撒 的子孙、 巴西亚 的子孙、
NEH|7|52|比赛 的子孙、 米乌宁 的子孙、 尼普心 的子孙、
NEH|7|53|巴卜 的子孙、 哈古巴 的子孙、 哈忽 的子孙、
NEH|7|54|巴洗律 的子孙、 米希大 的子孙、 哈沙 的子孙、
NEH|7|55|巴柯 的子孙、 西西拉 的子孙、 答玛 的子孙、
NEH|7|56|尼细亚 的子孙、 哈提法 的子孙。
NEH|7|57|所罗门 仆人的后裔： 琐太 的子孙、 琐斐列 的子孙、 比路大 的子孙、
NEH|7|58|雅拉 的子孙、 达昆 的子孙、 吉德 的子孙、
NEH|7|59|示法提雅 的子孙、 哈替 的子孙、 玻黑列．哈斯巴音 的子孙、 亚们 的子孙。
NEH|7|60|殿役和 所罗门 仆人的后裔共三百九十二名。
NEH|7|61|从 特．米拉 、 特．哈萨 、 基绿 、 亚顿 、 音麦 上来，不能证明他们的父系家族和后裔是否属 以色列 的如下：
NEH|7|62|第莱雅 的子孙、 多比雅 的子孙、 尼哥大 的子孙，共六百四十二名。
NEH|7|63|祭司中， 哈巴雅 的子孙、 哈哥斯 的子孙、 巴西莱 的子孙， 巴西莱 因为娶了 基列 人 巴西莱 的女儿为妻，所以就以此为名。
NEH|7|64|这些人在族谱之中寻查自己的谱系，却寻不着，因此算为不洁，不得作祭司。
NEH|7|65|省长对他们说，不可吃至圣的物，直到有会用乌陵和土明的祭司兴起来。
NEH|7|66|全会众共有四万二千三百六十名。
NEH|7|67|此外，还有他们的仆婢七千三百三十七名，又有歌唱的男女二百四十五名。
NEH|7|68|他们有七百三十六匹马，二百四十五匹骡子，
NEH|7|69|四百三十五匹骆驼，六千七百二十匹驴。
NEH|7|70|有些族长为工程捐助。省长捐入库房中的有一千达利克 金子，五十个碗，五百三十件祭司的礼服。
NEH|7|71|有些族长捐入工程的库房，有二万达利克金子，二千二百弥那银子。
NEH|7|72|其余百姓所捐的有二万达利克金子，二千弥那银子，六十七件祭司的礼服。
NEH|7|73|于是祭司、 利未 人、门口的守卫、歌唱的、百姓中的一些人、殿役，并 以色列 众人，都住在自己的城里。 到了七月， 以色列 人住在自己的城里。
NEH|8|1|那时，众百姓如同一人聚集在 水门 前的广场，请 以斯拉 文士将耶和华吩咐 以色列 的 摩西 的律法书带来。
NEH|8|2|七月初一， 以斯拉 祭司将律法书带到听了能明白的男女会众面前。
NEH|8|3|他在 水门 前的广场，从清早到中午，在男女和能明白的人面前读这律法书，众百姓都侧耳而听。
NEH|8|4|以斯拉 文士站在为这事特制的木台上。站在他旁边的有 玛他提雅 、 示玛 、 亚奈雅 、 乌利亚 和 希勒家 ；站在他右边的有 玛西雅 ；站在他左边的有 毗大雅 、 米沙利 、 玛基雅 、 哈顺 、 哈拔大拿 、 撒迦利亚 和 米书兰 。
NEH|8|5|以斯拉 站在上面，在众百姓眼前展开这书。他一展开，众百姓都站起来。
NEH|8|6|以斯拉 称颂耶和华至大的上帝，众百姓都举手应声说：“阿们！阿们！”他们低头，俯伏在地，敬拜耶和华。
NEH|8|7|耶书亚 、 巴尼 、 示利比 、 雅悯 、 亚谷 、 沙比太 、 荷第雅 、 玛西雅 、 基利他 、 亚撒利雅 、 约撒拔 、 哈难 、 毗莱雅 和 利未 人使百姓明白律法；百姓都站在自己的地方。
NEH|8|8|他们清清楚楚地念上帝的律法书，讲明意思，使百姓明白所念的。
NEH|8|9|尼希米 省长、 以斯拉 祭司文士，和教导百姓的 利未 人对众百姓说：“今日是耶和华－你们上帝的圣日，不要悲哀，也不要哭泣。”这是因为众百姓听见律法书上的话都哭了。
NEH|8|10|尼希米 对他们说：“你们去吃肥美的，喝甘甜的，有不能预备的就分给他，因为今日是我们主的圣日。你们不要忧愁，因靠耶和华而得的喜乐是你们的力量。”
NEH|8|11|于是 利未 人叫众百姓安静，说：“安静，因今日是圣日，不要忧愁。”
NEH|8|12|众百姓去吃喝，也分给别人，都大大喜乐，因为他们明白所教导他们的话。
NEH|8|13|次日，众百姓的族长、祭司和 利未 人都聚集到 以斯拉 文士那里，要明白律法书上的话。
NEH|8|14|他们发现律法书上写着，耶和华藉 摩西 吩咐 以色列 人要在七月的节期中住在棚里，
NEH|8|15|并要在各城和 耶路撒冷 传扬宣告说：“你们当出去，上山，把橄榄树、野橄榄树、番石榴树、棕树和各样茂密树的枝子取来，照着所写的搭棚。”
NEH|8|16|于是百姓出去，取了树枝来，各人在自己的房顶上，院子里，上帝殿的院内， 水门 的广场，和 以法莲门 的广场搭棚。
NEH|8|17|从被掳之地归回的全会众就搭棚，住在棚里。从 嫩 的儿子 约书亚 的时候直到这日， 以色列 人没有这样行。他们都大大喜乐。
NEH|8|18|从第一天直到末一天， 以斯拉 天天朗读上帝的律法书。他们守节七日，第八日照例有严肃会。
NEH|9|1|这月二十四日， 以色列 人聚集禁食，他们披麻蒙灰。
NEH|9|2|以色列 的后裔与所有的外邦人分别出来，站着承认自己的罪和祖先的罪孽。
NEH|9|3|那日的四分之一，他们站在自己的地方念耶和华－他们上帝的律法书，又在那日的四分之一认罪，敬拜耶和华－他们的上帝。
NEH|9|4|耶书亚 、 巴尼 、 甲篾 、 示巴尼 、 布尼 、 示利比 、 巴尼 、 基拿尼 站在 利未 人的台阶上，大声哀求耶和华－他们的上帝。
NEH|9|5|利未 人 耶书亚 、 甲篾 、 巴尼 、 哈沙尼 、 示利比 、 荷第雅 、 示巴尼 、 毗他希雅 说：“起来，称颂耶和华－你们的上帝，永世无尽：‘你荣耀之名是应当称颂的，超乎一切称颂和赞美。
NEH|9|6|“‘你，惟独你是耶和华！你造了天和天上的天，以及天上的万象，地和地上的万物，海和海中所有的；一切的生命全都是你赏赐的。天军都敬拜你。
NEH|9|7|你是耶和华上帝，曾拣选 亚伯兰 ，领他出 迦勒底 的 吾珥 ，给他改名叫 亚伯拉罕 。
NEH|9|8|你发现他在你面前心里忠诚，就与他立约，要把 迦南 人、 赫 人、 亚摩利 人、 比利洗 人、 耶布斯 人、 革迦撒 人之地赐给他的后裔，并且你也实现了你的话，因为你是公义的。
NEH|9|9|“‘你曾看见我们祖先在 埃及 所受的困苦，垂听他们在 红海 边的哀求，
NEH|9|10|施行神迹奇事在法老和他所有臣仆，以及他国中众百姓身上，因为你知道他们向我们祖先行事狂傲。你也得了名声，正如今日一样。
NEH|9|11|你在我们祖先面前把海分开，使他们走过海中干地，将追赶他们的人抛在深海，如石头抛在大水中。
NEH|9|12|白昼你用云柱引导他们，黑夜你用火柱照亮他们当行的路。
NEH|9|13|你降临在 西奈山 ，从天上与他们说话，赐给他们正直的典章、真实的律法、美好的律例与诫命，
NEH|9|14|又使他们知道你的圣安息日，并藉你仆人 摩西 传给他们诫命、律例、律法。
NEH|9|15|你从天上赐下粮食给他们充饥，使水从磐石流出给他们解渴。你吩咐他们进去，得你起誓应许要赐给他们的地。
NEH|9|16|“‘但我们的祖先行事狂傲，硬着颈项不听从你的诫命。
NEH|9|17|他们不肯顺从，也不记念你在他们中间所行的奇事，竟硬着颈项，居心悖逆，自立领袖，要回 埃及 他们为奴之地 。但你是乐意饶恕人，有恩惠，有怜悯，不轻易发怒，有丰盛慈爱的上帝，并没有丢弃他们。
NEH|9|18|他们虽然为自己铸了一头牛犊，说，这就是领你出 埃及 的神明，因而犯了亵渎的大罪，
NEH|9|19|你还是有丰富的怜悯，不把他们丢弃在旷野。白昼，云柱不离开他们，仍引导他们行路；黑夜，火柱仍照亮他们当行的路。
NEH|9|20|你赐下你良善的灵教导他们，没有收回吗哪不给他们吃，仍赐水给他们解渴。
NEH|9|21|在旷野四十年，你养育他们，他们一无所缺，衣服没有穿破，脚也没有肿。
NEH|9|22|你将列国和诸民族交给他们，把那些角落分给他们，他们就得了 西宏 之地，就是 希实本 王之地，和 巴珊 王 噩 之地。
NEH|9|23|你使他们的子孙多如天上的星，带他们到你对他们祖先说要进去得为业之地。
NEH|9|24|这样，这些子孙进去得了那地。你在他们面前制伏那地的居民 迦南 人，把 迦南 人和他们的君王，以及那地的民族，都交在他们手里，让他们任意处置。
NEH|9|25|他们得了坚固的城镇、肥沃的土地，取了装满各样美物的房屋、挖成的水井、葡萄园、橄榄园，以及许多果树。他们就吃了，而且饱足，身体肥胖，因你的大恩活得快乐。
NEH|9|26|“‘然而，他们不顺从，竟背叛你，将你的律法丢在背后，又杀害那些劝他们回转归向你的众先知，犯了亵渎的大罪。
NEH|9|27|所以你将他们交在敌人的手中，敌人就折磨他们。他们遭难的时候哀求你，你就从天上垂听，照你丰富的怜悯赐给他们拯救者，救他们脱离敌人的手。
NEH|9|28|但他们得享太平之后，又在你面前行恶，所以你丢弃他们，交在仇敌的手中，仇敌就辖制他们；然而他们转回哀求你，你就从天上垂听，屡次照你的怜悯拯救他们，
NEH|9|29|你警戒他们，要使他们归顺你的律法。他们却行事狂傲，不听从你的诫命，干犯你的典章，人若遵行就必因此存活。他们顽梗地扭转肩头，硬着颈项，不肯听从。
NEH|9|30|但你多年宽容他们，又以你的灵藉众先知劝戒他们，他们仍不侧耳而听，所以你将他们交在列邦民族的手中。
NEH|9|31|然而因你丰富的怜悯，你不全然灭绝他们，也不丢弃他们，因为你是有恩惠、有怜悯的上帝。
NEH|9|32|“‘现在，我们的上帝啊，你是至大、至能、至可畏、守约施慈爱的上帝；我们的君王、官长、祭司、先知、祖先和你的众百姓，从 亚述 诸王的时候直到今日所遭遇的一切苦难，求你不要看为小事。
NEH|9|33|在一切临到我们的事上，你是公义的，因为你所行的是信实，我们所做的是邪恶。
NEH|9|34|我们的君王、官长、祭司、祖先都不遵守你的律法，不听从你的诫命和你警戒他们的话。
NEH|9|35|他们在本国领受你大恩的时候，在你所赐给他们这广大肥沃之地不事奉你，也不转离他们的恶行。
NEH|9|36|看哪，我们今日成了奴仆！你赐给我们祖先享受土产和美物的地，看哪，我们在这地上竟作了奴仆！
NEH|9|37|这地许多的出产都归了诸王，就是你因我们的罪派来辖制我们的。他们任意辖制我们的身体和牲畜，我们遭了大难。’”
NEH|9|38|因这一切，我们立确实的约，写在册上。我们的领袖、 利未 人和祭司都用了印。
NEH|10|1|用印的是 哈迦利亚 的儿子 尼希米 省长、 西底家 ；
NEH|10|2|还有 西莱雅 、 亚撒利雅 、 耶利米 、
NEH|10|3|巴施户珥 、 亚玛利雅 、 玛基雅 、
NEH|10|4|哈突 、 示巴尼 、 玛鹿 、
NEH|10|5|哈琳 、 米利末 、 俄巴底亚 、
NEH|10|6|但以理 、 近顿 、 巴录 、
NEH|10|7|米书兰 、 亚比雅 、 米雅民 、
NEH|10|8|玛西亚 、 璧该 、 示玛雅 等祭司；
NEH|10|9|又有 利未 人 亚散尼 的儿子 耶书亚 、 希拿达 的子孙 宾内 、 甲篾 ，
NEH|10|10|他们的弟兄 示巴尼 、 荷第雅 、 基利他 、 毗莱雅 、 哈难 、
NEH|10|11|米迦 、 利合 、 哈沙比雅 、
NEH|10|12|撒刻 、 示利比 、 示巴尼 、
NEH|10|13|荷第雅 、 巴尼 、 比尼努 ；
NEH|10|14|还有百姓中的领袖 巴录 、 巴哈．摩押 、 以拦 、 萨土 、 巴尼 、
NEH|10|15|布尼 、 押甲 、 比拜 、
NEH|10|16|亚多尼雅 、 比革瓦伊 、 亚丁 、
NEH|10|17|亚特 、 希西家 、 押朔 、
NEH|10|18|荷第雅 、 哈顺 、 比赛 、
NEH|10|19|哈拉 、 亚拿突 、 尼拜 、
NEH|10|20|抹比押 、 米书兰 、 希悉 、
NEH|10|21|米示萨别 、 撒督 、 押杜亚 、
NEH|10|22|毗拉提 、 哈难 、 亚奈雅 、
NEH|10|23|何细亚 、 哈拿尼雅 、 哈述 、
NEH|10|24|哈罗黑 、 毗利哈 、 朔百 、
NEH|10|25|利宏 、 哈沙拿 、 玛西雅 、
NEH|10|26|亚希雅 、 哈难 、 亚难 、
NEH|10|27|玛鹿 、 哈琳 、 巴拿 。
NEH|10|28|其余的百姓、祭司、 利未 人、门口的守卫、歌唱的、殿役，所有与邻邦民族分别出来、归服上帝律法的，以及他们的妻子、儿女，凡有知识、能明白的，
NEH|10|29|都随从他们贵族的弟兄发咒起誓，要遵行上帝藉他仆人 摩西 所赐的律法，谨守遵行耶和华－我们主的一切诫命、典章、律例。
NEH|10|30|我们不把我们的女儿嫁给这地的居民，也不为我们的儿子娶他们的女儿。
NEH|10|31|这地的民族若在安息日，或什么圣日，带了货物或粮食来卖，我们必不买。每逢第七年必不耕种，凡欠我们债的必不追讨。
NEH|10|32|我们又为自己定例，每年各人捐献三分之一舍客勒，作为我们上帝殿之用：
NEH|10|33|为供饼、常献的素祭和燔祭，安息日、初一、节期所献的祭和圣物， 以色列 的赎罪祭，以及我们上帝殿里一切工作之用。
NEH|10|34|我们的祭司、 利未 人和百姓都抽签，每年按父家定期将奉献的木柴带到我们上帝的殿里，照着律法上所写的，烧在耶和华－我们上帝的坛上。
NEH|10|35|每年我们又将地上初熟的土产和各样树上初熟的果子，都奉到耶和华的殿里。
NEH|10|36|我们又照律法上所写的，将我们头胎的儿子和首生的牛羊都奉到我们上帝的殿，交给在上帝殿里供职的祭司；
NEH|10|37|并将初熟麦子所磨的面和举祭、各样树上的果子、新酒与新油奉给祭司，收在我们上帝殿的库房里，又把我们土地所产的十分之一奉给 利未 人，因 利未 人在我们一切城镇的土产中当取十分之一。
NEH|10|38|利未 人取十分之一的时候， 亚伦 的子孙中当有一个祭司与 利未 人同在。 利未 人也当从十分之一中取十分之一，奉到我们上帝的殿，收在库房的仓里。
NEH|10|39|因 以色列 人和 利未 人要把礼物，就是五谷、新酒和新油，带到收存圣所器皿的仓里，供职的祭司、门口的守卫、歌唱的都在那里。我们绝不会不顾我们上帝的殿。
NEH|11|1|百姓的领袖住在 耶路撒冷 。其余的百姓抽签，每十人中选一人来住在圣城 耶路撒冷 ，另外九人住在别的城镇。
NEH|11|2|凡甘心乐意住在 耶路撒冷 的，百姓都为他们祝福。
NEH|11|3|以色列 人、祭司、 利未 人、殿役和 所罗门 仆人的后裔都住在 犹大 的城镇，各在自己城内的地业中。本省的领袖住在 耶路撒冷 的如下：
NEH|11|4|住在 耶路撒冷 的有一些 犹大 人和 便雅悯 人。 犹大 人中有 法勒斯 的子孙 亚他雅 ； 亚他雅 是 乌西雅 的儿子， 乌西雅 是 撒迦利雅 的儿子， 撒迦利雅 是 亚玛利雅 的儿子， 亚玛利雅 是 示法提雅 的儿子， 示法提雅 是 玛勒列 的儿子；
NEH|11|5|又有 玛西雅 ； 玛西雅 是 巴录 的儿子， 巴录 是 谷．何西 的儿子， 谷．何西 是 哈赛雅 的儿子， 哈赛雅 是 亚大雅 的儿子， 亚大雅 是 约雅立 的儿子， 约雅立 是 撒迦利雅 的儿子， 撒迦利雅 是 示罗尼 的儿子；
NEH|11|6|住在 耶路撒冷 所有 法勒斯 的子孙共四百六十八名，都是勇士。
NEH|11|7|便雅悯 人中有 撒路 ； 撒路 是 米书兰 的儿子， 米书兰 是 约叶 的儿子， 约叶 是 毗大雅 的儿子， 毗大雅 是 哥赖雅 的儿子， 哥赖雅 是 玛西雅 的儿子， 玛西雅 是 以铁 的儿子， 以铁 是 耶筛亚 的儿子；
NEH|11|8|其次有 迦拜 、 撒来 ，共九百二十八名。
NEH|11|9|细基利 的儿子 约珥 是他们的长官； 哈西努亚 的儿子 犹大 是 耶路撒冷 的副长官。
NEH|11|10|祭司中有 约雅立 的儿子 耶大雅 ，又有 雅斤 ，
NEH|11|11|还有管理上帝殿的 西莱雅 ； 西莱雅 是 希勒家 的儿子， 希勒家 是 米书兰 的儿子， 米书兰 是 撒督 的儿子， 撒督 是 米拉约 的儿子， 米拉约 是 亚希突 的儿子；
NEH|11|12|还有他们的弟兄在殿里供职的，共八百二十二名；又有 亚大雅 ； 亚大雅 是 耶罗罕 的儿子， 耶罗罕 是 毗拉利 的儿子， 毗拉利 是 暗洗 的儿子， 暗洗 是 撒迦利亚 的儿子， 撒迦利亚 是 巴施户珥 的儿子， 巴施户珥 是 玛基雅 的儿子；
NEH|11|13|还有他的弟兄作族长的，共二百四十二名；又有 亚玛帅 ； 亚玛帅 是 亚萨列 的儿子， 亚萨列 是 亚哈赛 的儿子， 亚哈赛 是 米实利末 的儿子， 米实利末 是 音麦 的儿子；
NEH|11|14|还有他们的弟兄，大能的勇士共一百二十八名； 哈基多琳 的儿子 撒巴第业 是他们的长官。
NEH|11|15|利未 人中有 示玛雅 ； 示玛雅 是 哈述 的儿子， 哈述 是 押利甘 的儿子， 押利甘 是 哈沙比雅 的儿子， 哈沙比雅 是 布尼 的儿子；
NEH|11|16|又有 利未 人的族长 沙比太 和 约撒拔 管理上帝殿外面的事务；
NEH|11|17|祈祷的时候， 玛他尼 是主礼，开始称谢； 玛他尼 是 米迦 的儿子， 米迦 是 撒底 的儿子， 撒底 是 亚萨 的儿子；又有 玛他尼 弟兄中的 八布迦 为副；还有 押大 ； 押大 是 沙母亚 的儿子， 沙母亚 是 加拉 的儿子， 加拉 是 耶杜顿 的儿子；
NEH|11|18|在圣城所有的 利未 人共二百八十四名。
NEH|11|19|门口的守卫是 亚谷 和 达们 ，以及他们的弟兄，看守各门，共一百七十二名。
NEH|11|20|其余的 以色列 人、祭司、 利未 人都住在 犹大 一切的城镇，各在自己的地业中。
NEH|11|21|殿役却住在 俄斐勒 ； 西哈 和 基斯帕 管理他们。
NEH|11|22|在 耶路撒冷 ， 利未 人的长官，管理上帝殿事务的是歌唱者 亚萨 的子孙 乌西 ； 乌西 是 巴尼 的儿子， 巴尼 是 哈沙比雅 的儿子， 哈沙比雅 是 玛他尼 的儿子， 玛他尼 是 米迦 的儿子。
NEH|11|23|王为歌唱者下命令，确定他们每日当办的事 。
NEH|11|24|犹大 的儿子 谢拉 的子孙， 米示萨别 的儿子 毗他希雅 辅助王办理百姓一切的事。
NEH|11|25|至于村庄和所属的田地，有 犹大 人住在 基列．亚巴 和所属的乡镇 、 底本 和所属的乡镇、 叶甲薛 和所属的村庄、
NEH|11|26|耶书亚 、 摩拉大 、 伯．帕列 、
NEH|11|27|哈萨．书亚 、 别是巴 和所属的乡镇、
NEH|11|28|洗革拉 、 米哥拿 和所属的乡镇、
NEH|11|29|隐．临门 、 琐拉 、 耶末 、
NEH|11|30|撒挪亚 、 亚杜兰 和属它们的村庄、 拉吉 和所属的田地、 亚西加 和所属的乡镇；他们所住的地方是从 别是巴 直到 欣嫩谷 。
NEH|11|31|便雅悯 人从 迦巴 起，住在 密抹 、 亚雅 、 伯特利 和所属的乡镇、
NEH|11|32|亚拿突 、 挪伯 、 亚难雅 、
NEH|11|33|夏琐 、 拉玛 、 基他音 、
NEH|11|34|哈第 、 洗编 、 尼八拉 、
NEH|11|35|罗德 、 阿挪 、 革．夏纳欣 。
NEH|11|36|在 犹大 地区的 利未 人中，有些已归属 便雅悯 。
NEH|12|1|这些是同 撒拉铁 的儿子 所罗巴伯 以及 耶书亚 一起上来的祭司和 利未 人： 西莱雅 、 耶利米 、 以斯拉 、
NEH|12|2|亚玛利雅 、 玛鹿 、 哈突 、
NEH|12|3|示迦尼 、 利宏 、 米利末 、
NEH|12|4|易多 、 近顿 、 亚比雅 、
NEH|12|5|米雅民 、 玛底雅 、 璧迦 、
NEH|12|6|示玛雅 、 约雅立 、 耶大雅 、
NEH|12|7|撒路 、 亚木 、 希勒家 、 耶大雅 ；这些人在 耶书亚 的时代作祭司和他们弟兄的领袖。
NEH|12|8|利未 人有 耶书亚 、 宾内 、 甲篾 、 示利比 、 犹大 、 玛他尼 ； 玛他尼 和他的弟兄负责赞美诗歌。
NEH|12|9|他们的弟兄 八布迦 和 乌尼 按照班次站在他们的对面。
NEH|12|10|耶书亚 生 约雅金 ， 约雅金 生 以利亚实 ， 以利亚实 生 耶何耶大 ，
NEH|12|11|耶何耶大 生 约拿单 ， 约拿单 生 押杜亚 。
NEH|12|12|在 约雅金 的时代，祭司作族长的， 西莱雅 族有 米拉雅 ， 耶利米 族有 哈拿尼雅 ，
NEH|12|13|以斯拉 族有 米书兰 ， 亚玛利雅 族有 约哈难 ，
NEH|12|14|米利古 族有 约拿单 ， 示巴尼 族有 约瑟 ，
NEH|12|15|哈琳 族有 押拿 ， 米拉约 族有 希勒恺 ，
NEH|12|16|易多 族有 撒迦利亚 ， 近顿 族有 米书兰 ，
NEH|12|17|亚比雅 族有 细基利 ， 米拿民 族， 摩亚底 族有 毗勒太 ，
NEH|12|18|璧迦 族有 沙母亚 ， 示玛雅 族有 约拿单 ，
NEH|12|19|约雅立 族有 玛特乃 ， 耶大雅 族有 乌西 ，
NEH|12|20|撒来 族有 加莱 ， 亚木 族有 希伯 ，
NEH|12|21|希勒家 族有 哈沙比雅 ， 耶大雅 族有 拿坦业 。
NEH|12|22|在 以利亚实 、 耶何耶大 、 约哈难 、 押杜亚 的时代， 利未 人的族长都记在册上，祭司也一样，直到 波斯 王 大流士 在位的时候。
NEH|12|23|利未 人作族长的记在史籍上，一直记到 以利亚实 的儿子 约哈难 的时代。
NEH|12|24|利未 人的族长是 哈沙比雅 、 示利比 、 甲篾 的儿子 耶书亚 ，他们的弟兄站在他们的对面，照神人 大卫 的命令按着班次赞美称谢。
NEH|12|25|玛他尼 、 八布迦 、 俄巴底亚 、 米书兰 、 达们 、 亚谷 是门口的守卫，在库房的门口站岗。
NEH|12|26|这些人都在 约撒达 的孙子， 耶书亚 的儿子 约雅金 和 尼希米 省长，以及 以斯拉 祭司文士的时代供职。
NEH|12|27|为 耶路撒冷 城墙行奉献礼的时候，众人把各处的 利未 人召到 耶路撒冷 ，要以称谢、歌唱、敲钹、鼓瑟、弹琴，喜乐地行奉献礼。
NEH|12|28|歌唱的人从 耶路撒冷 的周围聚集，从 尼陀法 人的村庄、
NEH|12|29|伯．吉甲 ，以及 迦巴 和 亚斯玛弗 的田地而来；因为歌唱的人在 耶路撒冷 四围为自己建立了村庄。
NEH|12|30|祭司和 利未 人就洁净自己，也洁净百姓，以及城门和城墙。
NEH|12|31|我带 犹大 的领袖上城墙，把称谢的人分为两大队，在城墙上往右边的 粪厂门 行进，
NEH|12|32|在他们后面行进的有 何沙雅 与 犹大 一半的领袖，
NEH|12|33|又有 亚撒利雅 、 以斯拉 、 米书兰 、
NEH|12|34|犹大 、 便雅悯 、 示玛雅 、 耶利米 。
NEH|12|35|还有祭司的子孙，吹号的有 撒迦利亚 ； 撒迦利亚 是 约拿单 的儿子， 约拿单 是 示玛雅 的儿子， 示玛雅 是 玛他尼 的儿子， 玛他尼 是 米该亚 的儿子， 米该亚 是 撒刻 的儿子， 撒刻 是 亚萨 的儿子；
NEH|12|36|又有 撒迦利亚 的弟兄 示玛雅 、 亚撒利 、 米拉莱 、 基拉莱 、 玛艾 、 拿坦业 、 犹大 、 哈拿尼 ，各拿着神人 大卫 的乐器，由 以斯拉 文士在前面引领。
NEH|12|37|他们经过 泉门 往前，登 大卫城 的台阶，上城墙的斜坡，从 大卫 宫殿之上，直到朝东的 水门 。
NEH|12|38|第二队称谢的人要往反方向而行。我和一半的百姓在城墙上跟随他们，从 炉楼 之上，直到 宽墙 ；
NEH|12|39|又过了 以法莲门 、 古门 、 鱼门 、 哈楠业楼 、 哈米亚楼 ，直到 羊门 ，就在 护卫门 站住。
NEH|12|40|于是，这两队称谢的人连同我和一半跟随我的官长，站在上帝的殿里。
NEH|12|41|还有 以利亚金 、 玛西雅 、 米拿民 、 米该亚 、 以利约乃 、 撒迦利亚 、 哈楠尼亚 等吹号的祭司；
NEH|12|42|又有 玛西雅 、 示玛雅 、 以利亚撒 、 乌西 、 约哈难 、 玛基雅 、 以拦 和 以谢 。歌唱的大声唱歌，有 伊斯拉希雅 作指挥。
NEH|12|43|那日，众人献上丰盛的祭物，并且欢乐，因为上帝使他们大大欢乐，连妇女带孩童也都欢乐，甚至从远处都可听到 耶路撒冷 的欢声。
NEH|12|44|当日，有些人受派管理库房，把举祭、初熟之物，和所取的十一奉献，按各城的田地，照律法所定，归给祭司和 利未 人的份，都收在库房里。 犹大 人因祭司和 利未 人供职就欢乐。
NEH|12|45|祭司和 利未 人遵守上帝所吩咐的，守洁净礼。歌唱的和门口的守卫照着 大卫 和他儿子 所罗门 的命令也如此行。
NEH|12|46|古时，在 大卫 和 亚萨 的日子，有歌唱者的指挥，也有赞美称谢上帝的诗歌。
NEH|12|47|在 所罗巴伯 和 尼希米 的时代， 以色列 众人把歌唱者和门口的守卫每日当得的份供给他们，又把给 利未 人的分别出来； 利未 人又把给 亚伦 子孙的分别出来。
NEH|13|1|在那日，百姓听到人朗读 摩西 的律法书，发现书上写着， 亚扪 人和 摩押 人永不可入上帝的会；
NEH|13|2|因为他们没有拿食物和水来迎接 以色列 人，却雇了 巴兰 诅咒他们，但我们的上帝使那诅咒变为祝福。
NEH|13|3|以色列 人听见这律法，就与所有不同族群的人分别出来。
NEH|13|4|在这之前，与 多比雅 结亲的 以利亚实 祭司，受派管理我们上帝殿中的库房，
NEH|13|5|为 多比雅 预备了一间大屋子，就是从前收存素祭、乳香、器皿，和照例供给 利未 人、歌唱者、门口守卫的五谷、新酒和新油的十分之一，以及归祭司之举祭的屋子。
NEH|13|6|当这一切事发生的时候，我不在 耶路撒冷 ，因为 巴比伦 王 亚达薛西 三十二年，我回到王那里。过了多日，我又向王告假。
NEH|13|7|我来到 耶路撒冷 ，才知道 以利亚实 为 多比雅 所做、在上帝殿的院内为他预备屋子的那件恶事。
NEH|13|8|我非常愤怒，就把 多比雅 的一切家具都从屋子里抛出去。
NEH|13|9|我又吩咐人洁净这屋子，然后将上帝殿的器皿、素祭和乳香搬回那里。
NEH|13|10|我发现 利未 人当得的份无人供给他们，甚至供职的 利未 人与歌唱的都各奔回自己的田地去了。
NEH|13|11|我就斥责官长说：“你们为何不顾上帝的殿呢？”于是我召集 利未 人，使他们在自己的岗位上供职。
NEH|13|12|犹大 众人就把五谷、新酒和新油的十分之一送入库房。
NEH|13|13|我派 示利米雅 祭司、 撒督 文士和 利未 人 毗大雅 作司库管理库房，副手是 哈难 ； 哈难 是 撒刻 的儿子， 撒刻 是 玛他尼 的儿子；这些人都是忠实的，他们的职务是分派他们弟兄所当得的份。
NEH|13|14|我的上帝啊，求你因这事记念我，不要涂去我为上帝的殿与其中的礼仪所献的忠心。
NEH|13|15|那些日子，我在 犹大 见有人在安息日踹醡酒池，搬运禾捆驮在驴上，又把酒、葡萄、无花果和各样的担子在安息日扛入 耶路撒冷 ，我就在他们卖食物的那日警戒他们。
NEH|13|16|有一些住在城里的 推罗 人也把鱼和各样货物运进来，甚至在 耶路撒冷 ，在安息日卖给 犹大 人。
NEH|13|17|我就斥责 犹大 的贵族，对他们说：“你们怎么会做这恶事干犯安息日呢！
NEH|13|18|你们祖先岂不是这样做，以致我们的上帝使一切灾祸临到我们和这城吗？你们竟干犯安息日，使愤怒越发临到 以色列 ！”
NEH|13|19|安息日前一日黄昏的时候，我吩咐人把 耶路撒冷 城门锁上；我又吩咐，不过安息日不准开门。我也派几个仆人在城门口站岗，免得有人在安息日挑担子进城。
NEH|13|20|于是商人和贩卖各样货物的人，有一两次在 耶路撒冷 城外过夜。
NEH|13|21|我警告他们说：“你们为何在城墙前过夜呢？若再这样，我必下手办你们。”从此以后，他们在安息日就不再来了。
NEH|13|22|我吩咐 利未 人洁净自己来守城门，使安息日分别为圣。我的上帝啊，求你因这事记念我，照你丰盛的慈爱怜悯我。
NEH|13|23|那些日子，我又看见 犹太 人娶了 亚实突 、 亚扪 和 摩押 的女子为妻。
NEH|13|24|他们的儿女，一半说 亚实突 话，或其他种族的方言，不会说 犹大 话。
NEH|13|25|我就斥责他们，诅咒他们，打了他们几个人，拔下他们的胡须，叫他们指着上帝起誓：“你们不可把自己的女儿嫁给外邦人的儿子，也不可为自己和儿子娶他们的女儿。
NEH|13|26|以色列 王 所罗门 不也在这样的事上犯罪吗？在许多国家中并没有一位王像他，蒙他上帝喜爱，上帝立他作王治理全 以色列 。然而，连他也被外邦女子引诱犯罪。
NEH|13|27|我们岂能听凭你们行这一切大恶，娶外邦女子干犯我们的上帝呢？”
NEH|13|28|以利亚实 大祭司的孙子， 耶何耶大 的一个儿子是 和伦 人 参巴拉 的女婿，我就把他从我这里赶出去。
NEH|13|29|我的上帝啊，求你记得他们的罪，因为他们玷污了祭司的职分，违背祭司和 利未 人的约。
NEH|13|30|这样，我洁净他们，使他们脱离属外邦人的一切；我又分派祭司和 利未 人的班次，使他们各尽其职，
NEH|13|31|按定期奉献木柴和初熟的土产。我的上帝啊，求你记念我，施恩于我。
ESTH|1|1|这事发生在 亚哈随鲁 的时代， 亚哈随鲁 从 印度 直到 古实 统治一百二十七个省，
ESTH|1|2|就是 亚哈随鲁 王在 书珊 城堡中坐国度王位的那些日子。
ESTH|1|3|他在位第三年，为所有官员和臣仆摆设宴席，有 波斯 和 玛代 的权贵，各省的贵族与领袖在他面前。
ESTH|1|4|他把他荣耀国度的丰富和他伟大威严的尊贵给他们看了许多日子，共一百八十天。
ESTH|1|5|这些日子满了，王又为所有住 书珊 城堡的百姓，无论大小，在御花园的院子里摆设宴席七日。
ESTH|1|6|院子里有白色棉和蓝色线，用细麻绳、紫色绳系在白玉石柱的银环上，又有金银的床榻摆在红、白、黄、黑大理石镶嵌的地上。
ESTH|1|7|用金器皿盛酒，有很多不同的器皿，照王的厚意提供丰富的御酒。
ESTH|1|8|饮酒有规定，不准勉强人 ，因为王吩咐宫里所有的臣宰，让人各随己意。
ESTH|1|9|瓦实提 王后在 亚哈随鲁 王的宫内也为妇女摆设宴席。
ESTH|1|10|第七日， 亚哈随鲁 王饮酒，心中快乐，就吩咐在他面前侍立的七个太监 米户幔 、 比斯他 、 哈波拿 、 比革他 、 亚拔他 、 西达 、 甲迦 ，
ESTH|1|11|请 瓦实提 王后头戴王后的冠冕到王面前，让各民族和官员观看她的美貌，因为她容貌美丽。
ESTH|1|12|瓦实提 王后却不肯遵照太监所传的王命前来，所以王非常愤怒，怒火中烧。
ESTH|1|13|按王的常规，办事必先询问知例明法的人。那时，王询问通达时务的智慧人，
ESTH|1|14|就是在王左右常见王面、在国中坐高位的 波斯 和 玛代 的七个大臣， 甲示拿 、 示达 、 押玛他 、 他施斯 、 米力 、 玛西拿 、 米慕干 ：
ESTH|1|15|“ 瓦实提 王后不遵照太监所传的王命，照例应当怎样办理呢？”
ESTH|1|16|米慕干 在王和众官长面前回答说：“ 瓦实提 王后这事，不但得罪王，并且有害于 亚哈随鲁 王各省的臣民。
ESTH|1|17|因为王后这事必传到众妇人那里，她们就会藐视自己的丈夫，说：‘ 亚哈随鲁 王吩咐 瓦实提 王后到王面前，她却不来。’
ESTH|1|18|今日 波斯 和 玛代 的众夫人听见王后这事，必向王所有的官长照样说，如此必造成无数的藐视和愤怒。
ESTH|1|19|王若以为好，请降谕旨，写在 波斯 和 玛代 人的条例中，永不更改，不准 瓦实提 再到 亚哈随鲁 王面前，把她王后的位分赐给比她更好的妃子。
ESTH|1|20|王的谕旨一传遍全国，国土纵然辽阔，凡作妻子的，无论丈夫是尊贵或卑贱，都必尊敬他。”
ESTH|1|21|王和众官长都以这话为美，王就照 米慕干 的建议去做。
ESTH|1|22|王下诏书，用各省的文字、各族的语言通知各省，使凡作丈夫的在家中作主，各说本地的语言 。
ESTH|2|1|这些事以后， 亚哈随鲁 王的愤怒平息，就想起 瓦实提 和她所做的，以及自己怎样降旨办她。
ESTH|2|2|于是王的侍臣对王说：“请派人为王寻找美貌的少女；
ESTH|2|3|请王派官员在国中各省招聚所有美貌的少女到 书珊 城堡的女院，交给王所派掌管女子的太监 希该 ，给她们香膏涂抹。
ESTH|2|4|王眼中看为好的女子可以立为王后，代替 瓦实提 。”王以这话为美，就照样做。
ESTH|2|5|书珊 城堡中有一个 犹太 人名叫 末底改 ，是 便雅悯 人 基士 的曾孙， 示每 的孙子， 睚珥 的儿子。
ESTH|2|6|从前 巴比伦 王 尼布甲尼撒 把 犹大 王 耶哥尼雅 和百姓从 耶路撒冷 掳来， 末底改 也在被掳的人当中。
ESTH|2|7|末底改 抚养他叔叔的女儿 哈大沙 ，就是 以斯帖 ，因为她没有父母。这女子容貌美丽；她父母死了， 末底改 收她为自己的女儿。
ESTH|2|8|王的谕旨和敕令传出之后，许多女子被招聚到 书珊 城堡，交给掌管女子的 希该 ； 以斯帖 也被送入王宫，交给 希该 。
ESTH|2|9|希该 眼中宠爱 以斯帖 ，就恩待她，急忙给她涂抹的香膏和当得的份，又从王宫里挑选七个宫女来服事她，使她和她的宫女搬入女院上好的房屋。
ESTH|2|10|以斯帖 未曾将自己的籍贯宗族告诉人，因为 末底改 嘱咐她不可叫人知道。
ESTH|2|11|末底改 天天在女院前徘徊，要知道 以斯帖 是否平安，过得如何。
ESTH|2|12|众女子照例先涂抹身体十二个月：六个月用没药油，六个月用香料和涂抹的香膏。满了日期，每个女子挨次进去朝见 亚哈随鲁 王。
ESTH|2|13|女子进去朝见王是这样：从女院到王宫的时候，凡她所要的都必给她带进去。
ESTH|2|14|晚上她进去，次日回到另一个女院，交给掌管妃嫔的太监 沙甲 。除非王喜爱她，再提名召她，她就不再进去见王。
ESTH|2|15|末底改 的叔叔 亚比孩 的女儿，就是 末底改 收为自己女儿的 以斯帖 ，按次序要进去朝见王的时候，除了掌管女子的太监 希该 所分派给她的，她别无所求。凡看见 以斯帖 的都喜欢她。
ESTH|2|16|亚哈随鲁 王第七年十月，就是提别月， 以斯帖 被引入宫中朝见王。
ESTH|2|17|王爱 以斯帖 过于众女子，她在王面前蒙宠爱胜过众少女。王把王后的冠冕戴在她头上，立她为王后，代替 瓦实提 。
ESTH|2|18|王为所有的官长和臣仆摆设大宴席，称为 以斯帖 的宴席，又豁免各省的租税，并照王的厚意大颁赏赐。
ESTH|2|19|第二次招聚少女的时候， 末底改 坐在朝门。
ESTH|2|20|以斯帖 遵照 末底改 所嘱咐的，没有将籍贯宗族告诉人； 以斯帖 照 末底改 的吩咐去做，正如受他抚养的时候一样。
ESTH|2|21|那时候， 末底改 坐在朝门，王有两个守门的太监， 辟探 和 提列 ，恼恨 亚哈随鲁 王，想要下手害他。
ESTH|2|22|末底改 知道了这件事，就告诉 以斯帖 王后。 以斯帖 以 末底改 的名向王报告。
ESTH|2|23|这事经过查究后发现是真的，二人就被挂在木头上。这事在王面前记录在史籍上。
ESTH|3|1|这些事以后， 亚哈随鲁 王使 亚甲 人 哈米大他 的儿子 哈曼 尊大，提升了他，叫他的爵位超过所有与他同朝的官长。
ESTH|3|2|在朝门，王所有的臣仆都跪拜 哈曼 ，因为王如此吩咐，但 末底改 不跪不拜。
ESTH|3|3|在朝门，王的臣仆对 末底改 说：“你为何违背王的命令呢？”
ESTH|3|4|他们天天劝他，他还是不听，他们就告诉 哈曼 ，要看 末底改 的事是否站得住，因他已经告诉他们自己是 犹太 人。
ESTH|3|5|哈曼 见 末底改 不跪不拜，就非常愤怒。
ESTH|3|6|有人把 末底改 的宗族告诉 哈曼 。 哈曼 看下手只害 末底改 一人是小事，还图谋要灭绝 亚哈随鲁 王全国所有的 犹太 人，就是 末底改 的宗族。
ESTH|3|7|亚哈随鲁 王十二年正月，就是尼散月，人在 哈曼 面前抽普珥，普珥即签，要定何月何日；抽到了十二月，就是亚达月。
ESTH|3|8|哈曼 对 亚哈随鲁 王说：“有一民族散居在王国各省的民族中，与众不同；他们的律例与万民的律例不同，也不守王的律例，所以容留他们对王无益。
ESTH|3|9|王若以为好，请下谕旨灭绝他们，我就捐一万他连得银子交给管财政的人，纳入王的府库。”
ESTH|3|10|于是王从自己手上摘下戒指给 犹太 人的仇敌， 亚甲 人 哈米大他 的儿子 哈曼 。
ESTH|3|11|王对 哈曼 说：“这银子赐给你，这民族也交给你，可以照你眼中看为好的待他们。”
ESTH|3|12|正月十三日，王的一些书记受召而来，照着 哈曼 一切所吩咐的，用各省的文字、各族的语言，奉 亚哈随鲁 王的名写谕旨，又用王的戒指盖印，传给王的总督、各省的省长，以及各族的领袖。
ESTH|3|13|诏书由信差传到王的各省，限令一日之内，就是在十二月，亚达月十三日，把所有的 犹太 人，无论老少妇女孩子，全然剪除，杀戮灭绝，并抢夺他们的财产。
ESTH|3|14|这谕旨的抄本以敕令的方式在各省颁布，通知各族，预备等候那日。
ESTH|3|15|信差奉王的命令急忙起行，敕令传遍了 书珊 城堡。王同 哈曼 坐下饮酒， 书珊 城堡却陷入慌乱中。
ESTH|4|1|末底改 知道所发生的这一切事，就撕裂衣服，披麻蒙灰，在城中行走，痛哭哀号。
ESTH|4|2|他到了朝门前就停住脚步，因为穿麻衣的不可进朝门。
ESTH|4|3|王的谕旨和敕令所到的各省各处， 犹太 人都极其悲哀，禁食哭泣哀号，许多人躺在麻布和炉灰中。
ESTH|4|4|以斯帖 王后的宫女和太监来把这事告诉 以斯帖 ，她非常忧愁，就送衣服给 末底改 穿，要他脱下身上的麻衣，他却不肯接受。
ESTH|4|5|以斯帖 把王所派伺候她的一个太监 哈他革 召来，吩咐他去见 末底改 ，要知道到底发生了什么事，为何如此。
ESTH|4|6|于是 哈他革 出来，到朝门前的广场见 末底改 。
ESTH|4|7|末底改 把自己遭遇的一切，以及 哈曼 为灭绝 犹太 人答应捐入王库的银数都告诉了他；
ESTH|4|8|又把那传遍 书珊 、要灭绝 犹太 人的谕旨抄本交给 哈他革 ，要他给 以斯帖 看，并向她说明，嘱咐她去晋见王，向王恳求，为本族的人在王面前请命。
ESTH|4|9|哈他革 回来，把 末底改 的话告诉 以斯帖 。
ESTH|4|10|以斯帖 吩咐 哈他革 去见 末底改 ，说：
ESTH|4|11|“王所有的臣仆和各省的百姓都知道有一个定例，若未奉召见，擅入内院见王的，无论男女必被处死；除非王向他伸出金杖，不得存活。但我没有被召进去见王已经有三十天了。”
ESTH|4|12|他们把 以斯帖 的话告诉 末底改 。
ESTH|4|13|末底改 托人回覆 以斯帖 说：“你不要自己以为在王宫里强过任何 犹太 人，得以幸免。
ESTH|4|14|此时你若闭口不言， 犹太 人必从别处得解脱，蒙拯救；你和你父家必致灭亡。焉知你得了王后的位分不是为现今的机会吗？”
ESTH|4|15|以斯帖 吩咐人回覆 末底改 说：
ESTH|4|16|“你当去召集 书珊 所有的 犹太 人，为我禁食三昼三夜，不吃不喝；我和我的宫女也要这样禁食。然后我违例去晋见王，我若死就死吧！”
ESTH|4|17|于是 末底改 照 以斯帖 一切所吩咐的去做。
ESTH|5|1|第三日， 以斯帖 穿上朝服，站立在王宫的内院，对着王宫。王在殿里坐在宝座上，对着殿的门。
ESTH|5|2|王见 以斯帖 王后站在院内，她在王的眼中得恩宠，王向她伸出手中的金杖。 以斯帖 往前去摸杖头。
ESTH|5|3|王对她说：“ 以斯帖 王后啊，你要什么？无论你求什么，就是国的一半也必赐给你。”
ESTH|5|4|以斯帖 说：“王若以为好，请王带着 哈曼 今日赴我为王预备的宴席。”
ESTH|5|5|王说：“叫 哈曼 速速照 以斯帖 的话去做。”于是王带着 哈曼 赴 以斯帖 所预备的宴席。
ESTH|5|6|在宴席喝酒的时候，王又对 以斯帖 说：“你要什么，必赐给你；无论你求什么，就是国的一半也必给你。”
ESTH|5|7|以斯帖 回答说：“我所要的、我所求的，嗯......。
ESTH|5|8|我若在王眼前蒙恩，王若愿意赐我所要的，准我所求的，就请王和 哈曼 再赴我为你们预备的宴席。明日我必照王的话去做。”
ESTH|5|9|那日 哈曼 心中快乐，欢欢喜喜地出来。但是当他看见 末底改 在朝门不站起来，也不因他动一下，就满心恼怒 末底改 。
ESTH|5|10|哈曼 忍着气回家，叫人请他的一些朋友和他妻子 细利斯 来。
ESTH|5|11|哈曼 将他的荣华富贵、众多的儿女，和王使他尊大、提升他高过官长和臣仆的事，都述说给他们听。
ESTH|5|12|哈曼 又说：“ 以斯帖 王后预备宴席，除了我之外不许别人随王赴席。明日王后又请我随王赴席。
ESTH|5|13|只是每当我看见 犹太 人 末底改 坐在朝门，这一切对我就都毫无意义了。”
ESTH|5|14|他的妻子 细利斯 和他所有的朋友对他说：“叫人做一个五十肘高的木架，早晨求王把 末底改 挂在其上，然后你可以欢欢喜喜随王赴席。” 哈曼 认为这话很好，就叫人做了木架。
ESTH|6|1|那夜王睡不着觉，吩咐人取历史书，就是史籍，念给他听，
ESTH|6|2|发现书上写着：王有两个守门的太监 辟探 和 提列 ，想要下手害 亚哈随鲁 王， 末底改 告发了这件事。
ESTH|6|3|王说：“ 末底改 做了这事，有没有赐给他什么尊荣或高位呢？”伺候王的臣仆说：“没有赐给他什么。”
ESTH|6|4|王说：“谁在院子里？”那时 哈曼 正进入王宫的外院，要请王把 末底改 挂在他所预备的木架上。
ESTH|6|5|王的臣仆对他说：“看哪， 哈曼 站在院子里。”王说：“叫他进来。”
ESTH|6|6|哈曼 就进去。王对他说：“王所喜爱要赐尊荣的人，当如何待他呢？” 哈曼 心里说：“王所喜爱要赐尊荣的人，除了我，还有谁呢？”
ESTH|6|7|哈曼 就对王说：“王所喜爱要赐尊荣的人，
ESTH|6|8|当把王所穿的王袍拿来，牵了戴冠的御马，
ESTH|6|9|把王袍和御马都交给王一个极尊贵的大臣，吩咐人把王袍给王所喜爱要赐尊荣的人穿上，领他骑着御马走遍城里的广场，在他面前宣告：‘王所喜爱要赐尊荣的人，就是这样待他。’”
ESTH|6|10|王对 哈曼 说：“你速速把这王袍和御马，照你所说的，向坐在朝门的 犹太 人 末底改 去做。凡你所说的，一样都不可缺。”
ESTH|6|11|于是 哈曼 把王袍给 末底改 穿上，领他骑着御马走遍城里的广场，在他面前宣告：“王所喜爱要赐尊荣的人，就是这样待他。”
ESTH|6|12|末底改 仍回到朝门， 哈曼 却忧忧闷闷地蒙着头，急忙回家去了。
ESTH|6|13|哈曼 把所遭遇的一切都说给他妻子 细利斯 和他所有的朋友听。他的智囊团和他的妻子 细利斯 对他说：“你在 末底改 面前开始败落；他既是 犹太 人，你必不能胜过他，终必在他面前败落。”
ESTH|6|14|他们正跟 哈曼 说话的时候，王的几位太监来了，催 哈曼 快去赴 以斯帖 所预备的宴席。
ESTH|7|1|王带着 哈曼 来赴 以斯帖 王后的宴席。
ESTH|7|2|第二天在宴席喝酒的时候，王又对 以斯帖 说：“ 以斯帖 王后啊，你要什么，必赐给你；无论你求什么，就是国的一半也必给你。”
ESTH|7|3|以斯帖 王后回答说：“王啊，我若在你眼前蒙恩，王若以为好，我所要的，是王把我的性命赐给我；我所求的，是求我的本族。
ESTH|7|4|因为我和我的本族被出卖了，要被剪除，杀戮，灭绝。我们若被卖为奴为婢，我就闭口不言；但我们的痛苦比起王的损失，算不得什么 。”
ESTH|7|5|亚哈随鲁 王问 以斯帖 王后说：“擅敢起意如此行的是谁？这人在哪里呢？”
ESTH|7|6|以斯帖 说：“仇人敌人就是这恶人 哈曼 ！” 哈曼 在王和王后面前非常惊惶。
ESTH|7|7|王大怒，起来离开酒席往御花园去了。 哈曼 见王定意要加罪于他，就留下来求 以斯帖 王后救他的命。
ESTH|7|8|王从御花园回到酒席厅，见 哈曼 伏在 以斯帖 所靠的榻上；王说：“他竟敢在宫内、在我面前凌辱王后吗？”这话一出王口， 哈曼 的脸就被蒙住了。
ESTH|7|9|有一个伺候王名叫 哈波拿 的太监说：“看哪， 哈曼 还为那报告给王、救王有功的 末底改 做了一个五十肘高的木架，现今立在 哈曼 的家里。”王说：“把 哈曼 挂在木架上。”
ESTH|7|10|于是 哈曼 被挂在他为 末底改 所预备的木架上；王的愤怒才平息了。
ESTH|8|1|那日， 亚哈随鲁 王把 犹太 人的仇敌 哈曼 的家产赐给 以斯帖 王后。 末底改 也来到王面前，因为 以斯帖 已经告诉王， 末底改 跟她是什么关系。
ESTH|8|2|王摘下自己的戒指，就是从 哈曼 取回的，给了 末底改 。 以斯帖 派 末底改 管理 哈曼 的家产。
ESTH|8|3|以斯帖 又在王面前求情，俯伏在他脚前，流泪哀求他阻止 亚甲 人 哈曼 害 犹太 人的恶谋。
ESTH|8|4|王向 以斯帖 伸出金杖， 以斯帖 就起来，站在王面前，
ESTH|8|5|说：“王若以为好，我若在王面前蒙恩，王若认为合宜，我若在王眼前得喜悦，请王下谕旨，废除 亚甲 人 哈米大他 的儿子 哈曼 设谋，要杀灭王各省的 犹太 人所颁的诏书。
ESTH|8|6|我何忍见我本族的人受害？何忍见我同宗的人被灭呢？”
ESTH|8|7|亚哈随鲁 王对 以斯帖 王后和 犹太 人 末底改 说：“因为 哈曼 要下手害 犹太 人，看哪，我已把他的家产赐给 以斯帖 ，也把 哈曼 挂在木架上了。
ESTH|8|8|你们可以照你们看为好的，奉王的名写谕旨给 犹太 人，用王的戒指盖印；因为奉王的名所写、用王的戒指盖印的谕旨是不能废除的。”
ESTH|8|9|三月，就是西弯月二十三日，当时王的一些书记受召而来，按着 末底改 所吩咐的，用各省的文字、各族的语言，以及 犹太 人的文字语言写谕旨，传给那从 印度 直到 古实 一百二十七省的 犹太 人，以及总督、省长和领袖。
ESTH|8|10|末底改 奉 亚哈随鲁 王的名写谕旨，用王的戒指盖印，交给信差们骑上御用的王室快马去颁布。
ESTH|8|11|王准各城各镇的 犹太 人在一日之内，在十二月，就是亚达月的十三日聚集，在 亚哈随鲁 王的各省保护自己的性命，剪除，杀戮，灭绝那要攻击 犹太 人的各省各族所有的军队，以及他们的妻子儿女，夺取他们的财产为掠物。
ESTH|8|12|
ESTH|8|13|这谕旨的抄本以敕令的方式在各省颁布，通知各族，使 犹太 人预备等候那日，好在仇敌身上报仇。
ESTH|8|14|于是骑御用快马的信差奉王命催促，急忙起行；敕令传遍了 书珊 城堡。
ESTH|8|15|末底改 穿着蓝色白色的朝服，头戴大金冠冕，又穿紫色细麻布的外袍，从王面前出来； 书珊城 充满了欢乐的呼声。
ESTH|8|16|犹太 人有光荣，欢喜快乐，得享尊贵。
ESTH|8|17|王的谕旨和敕令所到的各省各城， 犹太 人都欢喜快乐，摆设宴席，以那日为吉日。国中许多民族的人因惧怕 犹太 人，就自称为 犹太 人。
ESTH|9|1|十二月，就是亚达月十三日，王的谕旨和敕令要执行的那一日， 犹太 人的仇敌盼望制伏他们，但 犹太 人反倒制伏了恨他们的人。
ESTH|9|2|犹太 人在 亚哈随鲁 王各省的城里聚集，下手击杀那些要害他们的人。没有人能在他们面前站立得住，因为各民族都惧怕他们。
ESTH|9|3|各省的领袖、总督、省长，和办理王事务的人，因惧怕 末底改 ，就都帮助 犹太 人。
ESTH|9|4|末底改 在朝中为大，名声传遍各省； 末底改 这人的权势日渐扩大。
ESTH|9|5|犹太 人用刀击杀所有的仇敌，杀灭他们，随意待那些恨他们的人。
ESTH|9|6|在 书珊 城堡中， 犹太 人杀灭了五百人。
ESTH|9|7|他们杀了 巴珊大他 、 达分 、 亚斯帕他 、
ESTH|9|8|破拉他 、 亚大利雅 、 亚利大他 、
ESTH|9|9|帕玛斯他 、 亚利赛 、 亚利代 、 瓦耶撒他 ；
ESTH|9|10|这十人都是 哈米大他 的孙子， 犹太 人的仇敌 哈曼 的儿子。 犹太 人却没有下手夺取财物。
ESTH|9|11|那日， 书珊 城堡中被杀的人数呈报到王面前。
ESTH|9|12|王对 以斯帖 王后说：“ 犹太 人在 书珊 城堡中杀灭了五百人，又杀了 哈曼 的十个儿子，在王其余的各省不知如何。你要什么，必赐给你；你还求什么，也必为你成就。”
ESTH|9|13|以斯帖 说：“王若以为好，求你允准 书珊 的 犹太 人，明日也照今日的谕旨去做，并把 哈曼 十个儿子的尸体挂在木架上。”
ESTH|9|14|王允准这么做。敕令传遍 书珊 ， 哈曼 十个儿子的尸体被挂了起来。
ESTH|9|15|亚达月十四日，在 书珊 的 犹太 人又聚集，在 书珊 杀了三百人，却没有下手夺取财物。
ESTH|9|16|亚达月十三日，在王各省其余的 犹太 人也都聚集，保护自己的性命，摆脱仇敌得享平安。他们杀了七万五千个恨他们的人，却没有下手夺取财物；十四日他们休息，以这日为设宴欢乐的日子。
ESTH|9|17|
ESTH|9|18|但 书珊 的 犹太 人却在十三日、十四日聚集；十五日休息，以这日为设宴欢乐的日子。
ESTH|9|19|所以住在无城墙的乡村的 犹太 人，都以亚达月十四日为设宴欢乐的吉日，彼此馈送礼物。
ESTH|9|20|末底改 记录这些事，写信给 亚哈随鲁 王各省远近所有的 犹太 人，
ESTH|9|21|吩咐他们每年守亚达月十四、十五两日，
ESTH|9|22|以这两日为 犹太 人摆脱仇敌得享平安、转忧为喜、转悲为乐的吉日，并在这两日设宴欢乐，彼此馈送礼物，赒济穷人。
ESTH|9|23|于是， 犹太 人照 末底改 所写给他们的，把开始所做的作为遵守的定例。
ESTH|9|24|因为 犹太 人的仇敌 亚甲 人 哈米大他 的儿子 哈曼 设谋要杀害 犹太 人，抽普珥，普珥即签，为要杀尽灭绝他们；
ESTH|9|25|但这阴谋 到了王面前，王却降旨使 哈曼 谋害 犹太 人的恶事归到他自己的头上，他和他的众子都被挂在木架上。
ESTH|9|26|所以 犹太 人照着普珥这名字称这两日为普珥日。他们因这信上一切的话，又因所看见所遇见的事，
ESTH|9|27|就规定自己与后裔，以及归化他们的人，每年按所写的、按时守这两日，永久不废。
ESTH|9|28|各省各城、世世代代、家家户户都记念并守这两日，使这普珥日在 犹太 人中不可废掉，在他们后裔中也永不遗忘。
ESTH|9|29|亚比孩 的女儿 以斯帖 王后和 犹太 人 末底改 以全权写第二封信，坚立这普珥日，
ESTH|9|30|送信给 亚哈随鲁 王国中一百二十七省所有的 犹太 人，祝他们平安和安稳，
ESTH|9|31|劝他们遵照 犹太 人 末底改 和 以斯帖 王后所规定的，按时守这普珥日，并照着 犹太 人为自己与后裔所规定的，禁食与哀求。
ESTH|9|32|以斯帖 规定了守普珥日的条例，这事也记录在书上。
ESTH|10|1|亚哈随鲁 王向国中和海岛的人征税。
ESTH|10|2|他以权柄能力所做的一切，以及他使 末底改 尊大、提升他的事，岂不都写在 玛代 和 波斯 王的史籍上吗？
ESTH|10|3|犹太 人 末底改 作 亚哈随鲁 王的宰相，在 犹太 人中为大，得许多弟兄的喜悦，为本族的人争取福利，为他所有的后代谋求幸福。
JOB|1|1|乌斯 地有一个人名叫 约伯 。这人完全、正直、敬畏上帝、远离恶事。
JOB|1|2|他生了七个儿子，三个女儿。
JOB|1|3|他的家产有七千只羊，三千匹骆驼，五百对牛，五百匹母驴，并有许多仆婢。这人在东方人中为至大。
JOB|1|4|他的儿子按着日子各在自己家里摆设宴席，派人去请他们的三个姊妹来，与他们一同吃喝。
JOB|1|5|宴席的日子过了， 约伯 派人去叫他们自洁。他清早起来，按着他们众人的数目献燔祭，因为他说：“恐怕我的儿子犯了罪，心中背弃 上帝。” 约伯 常常这样行。
JOB|1|6|有一天，上帝的众使者 来侍立在耶和华面前，撒但也来在其中。
JOB|1|7|耶和华对撒但说：“你从哪里来？”撒但回答耶和华说：“我从地上走来走去，在那里往返。”
JOB|1|8|耶和华对撒但说：“你曾用心察看我的仆人 约伯 没有？地上再没有人像他那样完全、正直、敬畏上帝、远离恶事。”
JOB|1|9|撒但回答耶和华说：“ 约伯 敬畏上帝，岂是无故呢？
JOB|1|10|你岂不是四面圈上篱笆围护他和他的家，以及他一切所有的吗？他手所做的都蒙你赐福，他的家产也在地上增多。
JOB|1|11|但你若伸手毁他一切所有的，他必当面背弃你。”
JOB|1|12|耶和华对撒但说：“看哪，凡他所有的都在你手中；只是不可伸手加害于他。”于是撒但从耶和华面前退出去。
JOB|1|13|有一天， 约伯 的儿女正在他们长兄的家里吃饭喝酒，
JOB|1|14|有报信的来见 约伯 ，说：“牛正耕地，母驴在旁边吃草，
JOB|1|15|示巴 人忽然闯来，把牲畜掳去，并用刀杀了仆人；惟有我一人逃脱，来报信给你。”
JOB|1|16|他还说话的时候，又有人来说：“上帝从天上降下火来，把羊群和仆人都吞灭了；惟有我一人逃脱，来报信给你。”
JOB|1|17|他还说话的时候，又有人来说：“ 迦勒底 人分成三队忽然闯来，把骆驼掳去，并用刀杀了仆人；惟有我一人逃脱，来报信给你。”
JOB|1|18|他还说话的时候，又有人来说：“你的儿女正在他们长兄的家里吃饭喝酒，
JOB|1|19|看哪，有狂风从旷野刮来，袭击房屋的四角，房屋倒塌在年轻人身上，他们就都死了；惟有我一人逃脱，来报信给你。”
JOB|1|20|约伯 就起来，撕裂外袍，剃了头，俯伏在地敬拜，
JOB|1|21|说：“我赤身出于母胎，也必赤身归回；赏赐的是耶和华，收取的也是耶和华。耶和华的名是应当称颂的。”
JOB|1|22|在这一切的事上， 约伯 并没有犯罪，也不以上帝为狂妄。
JOB|2|1|又有一天，上帝的众使者 来侍立在耶和华面前，撒但也来在其中。
JOB|2|2|耶和华问撒但说：“你从哪里来？”撒但回答说：“我从地上走来走去，在那里往返。”
JOB|2|3|耶和华对撒但说：“你曾用心察看我的仆人 约伯 没有？地上再没有人像他那样完全、正直、敬畏上帝、远离恶事。你虽激起我攻击他，无故吞灭他，他仍然持守他的纯正。”
JOB|2|4|撒但回答耶和华说：“人以皮代皮，情愿舍去一切所有的，来保全性命。
JOB|2|5|但你若伸手伤他的骨头和他的肉，他必当面背弃 你。”
JOB|2|6|耶和华对撒但说：“看哪，他在你手中，只要留下他的性命。”
JOB|2|7|于是撒但从耶和华面前退出去，击打 约伯 ，使他从脚掌到头顶长毒疮。
JOB|2|8|约伯 就坐在灰烬中，拿瓦片刮身体。
JOB|2|9|他的妻子对他说：“你仍然持守你的纯正吗？你背弃上帝，死了吧！”
JOB|2|10|约伯 却对她说：“你说话，正如愚顽的妇人。唉！难道我们从上帝手里得福，不也受祸吗？”在这一切的事上， 约伯 并没有以口犯罪。
JOB|2|11|约伯 的三个朋友， 提幔 人 以利法 、 书亚 人 比勒达 、 拿玛 人 琐法 ，听说这一切的灾祸临到他身上，各人就从自己的地方相约同来，为他悲伤，安慰他。
JOB|2|12|他们远远地举目观看，认不出他来，就放声大哭。各人撕裂外袍，向空中撒尘土，落在自己的头上。
JOB|2|13|他们同他七天七夜坐在地上，一句话也不对他说，因为他们见到了极大的痛苦。
JOB|3|1|此后， 约伯 开口诅咒自己的生日 。
JOB|3|2|约伯 说：
JOB|3|3|“愿我生的那日灭没， 说‘怀了男胎’的那夜也灭没。
JOB|3|4|愿那日变为黑暗， 愿上帝不从上面寻找它， 愿亮光不照于其上。
JOB|3|5|愿黑暗和死荫索取那日， 愿密云停在其上， 愿白天的昏暗 恐吓它。
JOB|3|6|愿那夜被幽暗夺取， 不在一年的日子中喜乐， 也不列入月中的数目。
JOB|3|7|看哪，愿那夜没有生育， 其间也没有欢乐的声音。
JOB|3|8|愿那些诅咒日子且能惹动 力威亚探 的， 诅咒那夜。
JOB|3|9|愿那夜黎明的星宿变为黑暗， 盼亮却不亮， 也不见晨曦破晓 ；
JOB|3|10|因它没有把怀我胎的门关闭， 也没有从我的眼中隐藏患难。
JOB|3|11|“我为何不出母胎而死？ 为何不出母腹就气绝呢？
JOB|3|12|为何有膝盖接收我？ 为何有奶哺养我呢？
JOB|3|13|不然，我现在已躺卧安睡， 而且，早已长眠安息；
JOB|3|14|与那些为自己重建荒凉之处， 地上的君王和谋士在一起；
JOB|3|15|或与把银子装满房屋， 拥有金子的王子在一起；
JOB|3|16|我为何不像流产的胎儿被埋藏， 如同未见光的婴孩？
JOB|3|17|在那里恶人止息搅扰， 在那里困乏人得享安息，
JOB|3|18|被囚的人同得安逸， 不再听见监工的声音。
JOB|3|19|大的小的都在那里， 奴仆脱离主人得自由。
JOB|3|20|“遭受患难的人为何有光赐给他呢？ 心中愁苦的人为何有生命赐给他呢？
JOB|3|21|他们等死，却不得死； 求死，胜于求隐藏的珍宝。
JOB|3|22|他们寻见坟墓， 就欢喜快乐，极其高兴。
JOB|3|23|这人的道路遮隐， 上帝又四面围困他。
JOB|3|24|我吃饭前就发出叹息， 我的唉哼涌出如水。
JOB|3|25|因我所恐惧的临到我， 我所惧怕的迎向我；
JOB|3|26|我不得安逸，不得平静， 也不得安息，却有患难来到。”
JOB|4|1|提幔 人 以利法 回答说：
JOB|4|2|“人想与你说话，你就厌烦吗？ 但谁能忍住不发言呢？
JOB|4|3|看哪，你素来教导许多人， 又坚固软弱的手。
JOB|4|4|你的言语曾扶助跌倒的人； 你使软弱的膝盖稳固。
JOB|4|5|但现在祸患临到 你，你就烦躁了； 它挨近你，你就惊惶。
JOB|4|6|你的倚靠不是在于你敬畏上帝吗？ 你的盼望不是在于你行事纯正吗？
JOB|4|7|“请你追想：无辜的人有谁灭亡？ 正直的人何处被剪除？
JOB|4|8|按我所见，耕罪孽的， 种毒害的，照样收割。
JOB|4|9|上帝一嘘气，他们就灭亡； 上帝一发怒，他们就消失。
JOB|4|10|狮子吼叫，猛狮咆哮， 少壮狮子的牙齿被敲断。
JOB|4|11|公狮因缺猎物而死， 母狮的幼狮都离散。
JOB|4|12|“有话暗中传递给我， 耳朵听其微小的声音。
JOB|4|13|世人沉睡的时候， 从夜间异象的杂念中，
JOB|4|14|恐惧战兢临到我身， 使我百骨战抖。
JOB|4|15|有灵从我面前经过， 我身上的毫毛竖立。
JOB|4|16|那灵停住， 我却不能辨其形状； 有形像在我眼前。 我在静默中听见有声音：
JOB|4|17|‘必死的人能比上帝公义吗？ 壮士能比造他的主纯洁吗？
JOB|4|18|看哪，主不信靠他的仆人， 尚且指他的使者为愚昧，
JOB|4|19|何况那些住在泥屋、 根基在尘土里、 被蛀虫所毁坏的人呢？
JOB|4|20|早晚之间，他们就被毁灭， 永归无有，无人理会。
JOB|4|21|他们帐棚的绳索岂不从中拔出来呢？ 他们死，且是无智慧而死。’”
JOB|5|1|“你呼求吧，有谁回答你呢？ 圣者之中，你转向哪一位呢？
JOB|5|2|愤怒害死愚妄人， 嫉妒杀死愚蠢的人。
JOB|5|3|我曾见愚妄人扎下根， 但我忽然诅咒他的住处。
JOB|5|4|他的儿女远离稳妥之地， 在城门口被欺压，无人搭救。
JOB|5|5|他的庄稼被饥饿的人吃尽了， 就是在荆棘里的也抢去了； 他的财宝被陷阱 张口吞没了。
JOB|5|6|因为祸患不是从尘土中出来， 患难也不是从土地里长出。
JOB|5|7|人生出来必遭遇患难， 如同火花 飞腾。
JOB|5|8|“至于我，我必寻求上帝， 把我的事情交托给他。
JOB|5|9|他行大事不可测度， 行奇事不可胜数。
JOB|5|10|他降雨在地面， 赐水于田野。
JOB|5|11|他将卑微的人安置在高处， 将哀痛的人举到稳妥之地。
JOB|5|12|他破坏通达人的计谋， 使他们手所做的不得成就。
JOB|5|13|他使有智慧的人中了自己的诡计， 叫狡诈人的计谋速速落空。
JOB|5|14|他们白昼遇见黑暗， 午间摸索如在夜间。
JOB|5|15|上帝拯救贫穷人脱离残暴人的手， 脱离他们口中的刀。
JOB|5|16|这样，贫寒人有指望， 不义的人闭口无言。
JOB|5|17|“看哪，上帝所惩治的人是有福的！ 所以你不可轻看全能者的管教。
JOB|5|18|因为他打伤，又包扎； 他击伤，又亲手医治。
JOB|5|19|你六次遭难，他必救你； 就是七次，灾祸也无法害你。
JOB|5|20|在饥荒中，他必救你脱离死亡； 在战争中，他必救你脱离刀剑的权势。
JOB|5|21|你必被隐藏，不受口舌之害； 灾害临到，你也不惧怕。
JOB|5|22|对于灾害饥馑，你必讥笑； 至于地上的野兽，你也不惧怕。
JOB|5|23|因为你必与田间的石头立约， 田里的野兽也必与你和好。
JOB|5|24|你必知道你的帐棚平安， 你查看你的羊圈，一无所失。
JOB|5|25|你也必知道你的后裔众多， 你的子孙像地上的青草。
JOB|5|26|你必寿高年迈才归坟墓， 好像禾捆按时收藏。
JOB|5|27|看哪，这道理我们已经考察，本是如此。 你须要听，要亲自明白。”
JOB|6|1|约伯 回答说：
JOB|6|2|“惟愿我的烦恼被秤一秤， 我一切的灾害放在天平里，
JOB|6|3|现今都比海沙更重， 所以我说话急躁。
JOB|6|4|因全能者的箭射中了我， 我的灵喝尽其毒； 上帝的惊吓摆阵攻击我。
JOB|6|5|野驴有草岂会叫唤？ 牛有饲料岂会吼叫？
JOB|6|6|食物淡而无盐岂可吃呢？ 蛋白有什么滋味呢？
JOB|6|7|那些可厌的食物， 我心不肯挨近。
JOB|6|8|“惟愿我得着所求的， 上帝赏赐我所切望的，
JOB|6|9|愿上帝把我压碎， 伸手将我剪除。
JOB|6|10|我因没有违弃那圣者的言语， 就仍以此为安慰， 在不止息的痛苦中还可欢跃。
JOB|6|11|我有什么气力使我等候？ 我有什么结局使我忍耐？
JOB|6|12|我的气力岂是石头的气力？ 我的肉身岂是铜呢？
JOB|6|13|在我里面岂不是无助吗？ 智慧岂不是从我心中被赶逐吗？
JOB|6|14|“灰心的人，他的朋友当以慈爱待他， 因为他将离弃敬畏全能者的心。
JOB|6|15|我的弟兄诡诈，好像河道， 像溪水流过的河床，
JOB|6|16|因结冰而混浊， 有雪藏在其中，
JOB|6|17|暖和的时候就溶化， 炎热时便从原处干涸。
JOB|6|18|商队偏离道路， 上到荒凉之地而死亡。
JOB|6|19|提玛 的商队瞻望， 示巴 的旅客等候。
JOB|6|20|他们因希望落空就抱愧， 来到那里便蒙羞。
JOB|6|21|现在你们正是这样 ， 看见惊吓的事就惧怕。
JOB|6|22|我岂说：‘请你们供给我， 从你们的财物中送礼给我’？
JOB|6|23|或说：‘请你们拯救我脱离敌人的手， 救赎我脱离残暴人的手’吗？
JOB|6|24|“请你们指教我，我就不作声； 我在何事上有错，请使我明白。
JOB|6|25|正直言语的力量何其大！ 但你们责备是责备什么呢？
JOB|6|26|绝望人的讲论既然如风， 你们还计划批驳言语吗？
JOB|6|27|你们甚至为孤儿抽签， 把朋友当货物。
JOB|6|28|“现在，请你们看着我， 我绝不当面说谎。
JOB|6|29|请你们转意，不要不公义； 请再转意，正义在我这里。
JOB|6|30|我的舌头岂有不公义吗？ 我的上膛岂不辨奸恶吗？”
JOB|7|1|“人在世上岂无劳役呢？ 他的日子不像雇工的日子吗？
JOB|7|2|像奴仆切慕阴凉， 像雇工等待工钱，
JOB|7|3|我也照样度过虚空的岁月， 愁烦的夜晚指定给我。
JOB|7|4|我躺卧的时候就说： ‘我何时可以起来呢？’漫漫长夜， 我总是翻来覆去，直到天亮。
JOB|7|5|我的肉体以虫子和尘土为衣， 我的皮肤才收了口又流脓。
JOB|7|6|我的日子比织布的梭更快， 都消耗在没有指望之中。
JOB|7|7|“你要记得，我的生命不过是一口气， 我的眼睛必不再看见福乐。
JOB|7|8|观看我的人，他的眼必不看见我； 你的眼目投向我，我却不在了。
JOB|7|9|云彩消散而去； 照样，人下阴间也不再上来。
JOB|7|10|他不再回自己的家， 他自己的地方也不再认得他。
JOB|7|11|“我甚至不封我的口； 我灵愁苦，要发出言语； 我心苦恼，要吐露哀情。
JOB|7|12|我岂是海洋，岂是大鱼， 你竟防守着我呢？
JOB|7|13|我若说：‘我的床必安慰我， 我的榻必分担我的苦情’，
JOB|7|14|你就用梦惊扰我， 用异象恐吓我。
JOB|7|15|甚至我宁可窒息死亡， 胜似留我这副骨头。
JOB|7|16|我厌弃生命，不愿永远活着。 你任凭我吧，因我的日子都是虚空。
JOB|7|17|人算什么，你竟看他为大， 将他放在心上，
JOB|7|18|每早晨鉴察他， 每时刻考验他？
JOB|7|19|你到何时才转眼不看我， 任凭我咽下唾沫呢？
JOB|7|20|鉴察人的主啊，我若有罪，于你何妨？ 为何以我当你的箭靶， 使我成为你的重担呢？
JOB|7|21|为何不赦免我的过犯， 除掉我的罪孽呢？ 我现今要躺卧在尘土中； 你要切切寻找我，我却不在了。”
JOB|8|1|书亚 人 比勒达 回答说：
JOB|8|2|“这些话你要说到几时？ 你口中的言语如狂风要到几时呢？
JOB|8|3|上帝岂能偏离公平？ 全能者岂能偏离公义？
JOB|8|4|或者你的儿女得罪了他， 他就把他们交在过犯的掌控中。
JOB|8|5|你若切切寻求上帝， 向全能者恳求；
JOB|8|6|你若纯洁正直， 他必定为你兴起， 使你公义的居所兴旺。
JOB|8|7|你起初虽然微小， 日后必非常强盛。
JOB|8|8|“请你询问上代， 思念他们祖先所查究的。
JOB|8|9|我们不过从昨日才有，一无所知， 因我们在世的日子好像影子。
JOB|8|10|他们岂不指教你，告诉你， 说出发自内心的言语呢？
JOB|8|11|“蒲草没有泥岂能生长？ 芦荻没有水岂能长大？
JOB|8|12|它还青翠，没有割下的时候， 比百样的草先枯槁。
JOB|8|13|凡忘记上帝的人，路途也是这样； 不虔敬人的指望要灭没。
JOB|8|14|他所仰赖的必折断， 他所倚靠的是蜘蛛网。
JOB|8|15|他要倚靠房屋，房屋却站立不住； 他要抓住房屋，房屋却不能存留。
JOB|8|16|他在日光之下茂盛， 嫩枝在园中蔓延；
JOB|8|17|他的根盘绕石堆， 钻入石缝 。
JOB|8|18|他若从本地被拔出， 那地就不认识他，说：‘我没有见过你。’
JOB|8|19|看哪，这就是他道路中的喜乐， 以后必另有人从尘土而生。
JOB|8|20|看哪，上帝必不丢弃完全人， 也不扶助邪恶人的手。
JOB|8|21|他还要以喜笑充满你的口， 以欢呼充满你的嘴唇。
JOB|8|22|恨恶你的要披戴羞愧， 恶人的帐棚必归于无有。”
JOB|9|1|约伯 回答说：
JOB|9|2|“我真的知道是这样， 但人在上帝前怎能成为义呢？
JOB|9|3|人若想要与他争辩， 千次中也不能回答一次。
JOB|9|4|他心里有智慧，且大有能力。 谁向上帝刚硬而得平安呢？
JOB|9|5|他把山挪移，山却不知， 他在怒气中，把山翻倒。
JOB|9|6|他使地震动，离其本位， 地的柱子就摇撼。
JOB|9|7|他吩咐太阳，太阳就不出来， 又封住众星。
JOB|9|8|他独自铺张诸天， 步行在海浪之上。
JOB|9|9|他造北斗、参星、昴星， 以及南方的星宿 ；
JOB|9|10|他行大事不可测度， 行奇事不可胜数。
JOB|9|11|看哪，他从我旁边经过，我看不见； 他走过，我没有察觉他。
JOB|9|12|看哪，他夺去，谁能阻挡他？ 谁敢对他说：‘你做什么呢？’
JOB|9|13|“上帝必不收回他的怒气， 扶助 拉哈伯 的，屈身在上帝以下。
JOB|9|14|既是这样，我怎敢回答他， 怎敢在他之前选择辩词呢？
JOB|9|15|我虽有义，也不能回答， 我要向那审判我的恳求。
JOB|9|16|我若呼求，纵然他应允我， 我仍不信他会侧耳听我的声音。
JOB|9|17|他用暴风 摧折我， 无故加增我的损伤。
JOB|9|18|他不容我喘一口气， 倒使我饱受苦恼。
JOB|9|19|若论力量，看哪，他真有能力！ 若论审判，‘谁能传我呢？’
JOB|9|20|我虽有义，我的口要定我有罪； 我虽完全，他必证明我为弯曲。
JOB|9|21|我虽完全，不顾自己； 我厌弃我的性命。
JOB|9|22|所以我说，都是一样； 完全人和恶人，他都灭绝。
JOB|9|23|若灾祸忽然带来死亡， 他必戏笑无辜人的苦难。
JOB|9|24|世界交在恶人手中； 他蒙蔽世界审判官的脸， 若不是他，那么是谁呢？
JOB|9|25|“我的日子比奔跑者更快， 急速过去，不见福乐。
JOB|9|26|我的日子如蒲草船掠过， 如鹰俯冲抓食。
JOB|9|27|我若说：‘我要忘记我的苦情， 强颜欢笑’，
JOB|9|28|我就因一切的愁苦而惧怕； 我知道你必不以我为无辜。
JOB|9|29|我必被定罪， 我何必徒然劳苦呢？
JOB|9|30|我若用雪水洗身， 用碱洁净我的手掌，
JOB|9|31|你还要把我扔在坑里， 我的衣服都憎恶我。
JOB|9|32|他不像我是个人，使我可以回答他， 使我们可以一同受审判。
JOB|9|33|我们中间没有仲裁者， 可以按手在我们两造之间。
JOB|9|34|愿他使他的杖离开我， 不使他的威严恐吓我，
JOB|9|35|我就说话，不惧怕他； 但对我来说，我却不是这样。”
JOB|10|1|“我厌恶自己的性命， 任由我述说自己的苦情； 因心里苦恼，我要说话。
JOB|10|2|我对上帝说，不要定我有罪， 要指示我，你为何与我争辩？
JOB|10|3|你手所造的，你又欺压，又藐视， 却光照恶人的计谋。 这事你以为美吗？
JOB|10|4|你的眼岂是肉眼？ 你察看岂像人察看吗？
JOB|10|5|你的日子岂像人的日子， 你的年岁岂像壮士的年岁，
JOB|10|6|你就追问我的罪孽， 寻察我的罪过吗？
JOB|10|7|其实，你知道我没有行恶， 也无人能施行拯救，脱离你的手。
JOB|10|8|你的手塑造我，造了我， 但我整个人却要一起被你吞灭。
JOB|10|9|求你记得，你制造我如泥土， 你还要使我归回尘土吗？
JOB|10|10|你不是倒出我来好像奶， 使我凝结如同奶酪吗？
JOB|10|11|你以皮和肉给我穿上， 用骨与筋把我联结起来。
JOB|10|12|你将生命和慈爱赐给我， 你也眷顾保全我的灵。
JOB|10|13|然而，你把这些事藏在你心里， 我知道这是你的旨意。
JOB|10|14|我若犯罪，你就察看我， 并不赦免我的罪。
JOB|10|15|我若行恶，我就有祸了； 我若行义，也不敢抬头， 而是饱受羞辱， 看见我的痛苦。
JOB|10|16|你如狮子昂首追捕我 ， 又在我身上显出奇事。
JOB|10|17|你更新你的见证对付我， 向我加增恼怒， 调遣军队攻击我。
JOB|10|18|“你为何使我出母胎呢？ 甚愿我当时气绝，没有眼睛看见我。
JOB|10|19|这样，就如从未有过我， 我一出母胎就被送入坟墓。
JOB|10|20|我的日子不是短少吗？求你停止， 求你放过我 ，使我可以稍得喜乐，
JOB|10|21|就是在我去而不返， 往黑暗和死荫之地以先。
JOB|10|22|那是乌黑之地， 犹如幽暗的死荫， 毫无秩序； 发出的光辉也像幽暗。”
JOB|11|1|拿玛 人 琐法 回答说：
JOB|11|2|“这许多的话岂不该回答吗？ 多嘴多舌的人岂可成为义呢？
JOB|11|3|你夸大的话岂能使人不作声吗？ 你戏笑的时候岂没有人使你受辱吗？
JOB|11|4|你说：‘我的教导纯全， 我在你眼前是清洁的。’
JOB|11|5|但是，惟愿上帝说话， 愿他张开嘴唇攻击你。
JOB|11|6|愿他将智慧的奥秘指示你， 因为健全的知识是两面的。 你当知道，上帝使你忘记你的一些罪孽。
JOB|11|7|你能寻见上帝的奥秘吗？ 你能寻见全能者的极限吗？
JOB|11|8|高如诸天，你能做什么？ 比阴间深，你能知道什么？
JOB|11|9|其量度比地长， 比海更宽。
JOB|11|10|他若经过，把人拘禁， 召集会众，谁能阻挡他呢？
JOB|11|11|因为他知道虚妄的人； 当他看见罪恶，岂不留意吗？
JOB|11|12|空虚的人若获得知识， 野驴生下的驹子也成了人。
JOB|11|13|“至于你，若坚固己心， 又向主举手；
JOB|11|14|你若远远脱离你手中的罪孽， 不容许不义住在你帐棚之中；
JOB|11|15|这样，你必仰起脸来，毫无瑕疵； 你也必安稳，无所惧怕。
JOB|11|16|你必忘记你的苦楚， 就是想起来，也如流过的水。
JOB|11|17|你在世要升高，比正午更明， 虽有黑暗，仍像早晨。
JOB|11|18|你因有指望就必稳固， 也必四围察看 ，安然躺下。
JOB|11|19|你躺卧，无人惊吓， 并有许多人向你求恩。
JOB|11|20|但恶人的眼睛要失明； 他们无路可逃， 他们的指望就是气绝身亡。”
JOB|12|1|约伯 回答说：
JOB|12|2|“你们果真是人物啊！ 智慧要与你们一同去死。
JOB|12|3|但我也有聪明，跟你们一样， 并非不及你们。 这些事，谁不知道呢？
JOB|12|4|我这求告上帝、蒙他应允的人 竟成了朋友所讥笑的； 又公义又完全的人竟遭受讥笑。
JOB|12|5|安逸的人心里藐视灾祸， 这灾祸在等待失足滑跌的人。
JOB|12|6|强盗的帐棚安宁， 惹上帝发怒的人稳固， 他们把上帝 握在自己手中 。
JOB|12|7|“你问走兽，走兽必指教你； 你问空中的飞鸟，飞鸟必告诉你；
JOB|12|8|或者你与地说话，地必指教你 ； 海中的鱼也必向你说明。
JOB|12|9|在这一切当中， 有谁不知道这是耶和华的手做成的呢？
JOB|12|10|凡动物的生命 和人类的气息都在他手中。
JOB|12|11|耳朵岂不辨别言语， 正如上膛品尝食物吗？
JOB|12|12|年老的有智慧， 寿高的有知识。
JOB|12|13|“在上帝有智慧和能力， 他有谋略和知识。
JOB|12|14|看哪，他拆毁，就不能重建； 他拘禁人，人就不得释放。
JOB|12|15|看哪，他使水止住，水就干了； 他把水放出，水就淹没大地。
JOB|12|16|在他有能力和智慧， 走迷的和使人迷路的都属他。
JOB|12|17|他把谋士剥衣掳去， 使审判官变为愚妄。
JOB|12|18|他解除君王的权势 ， 用带子捆住他们的腰。
JOB|12|19|他把祭司剥衣掳去， 使有权能的人倾覆。
JOB|12|20|他废去忠信者的言论， 夺去长者的见识。
JOB|12|21|他使贵族蒙羞受辱， 放松勇士的腰带。
JOB|12|22|他从黑暗中彰显深奥的事， 使死荫显出光明。
JOB|12|23|他使邦国兴旺而又毁灭， 使邦国扩展又被掠夺。
JOB|12|24|他将地上百姓中领袖的聪明夺去， 使他们迷失在荒凉无路之地。
JOB|12|25|他们在无光的黑暗中摸索； 他使他们摇晃像醉酒的人一样。”
JOB|13|1|“看哪，这一切，我眼都见过； 我耳都听过，而且明白。
JOB|13|2|你们所知道的，我也知道， 并非不及你们。
JOB|13|3|然而我要对全能者说话， 我愿与上帝理论。
JOB|13|4|但你们是编造谎言的， 全都是无用的医生。
JOB|13|5|惟愿你们全然不作声， 这就是你们的智慧！
JOB|13|6|请你们听我的答辩， 留心听我嘴唇的诉求。
JOB|13|7|你们要为上帝说不义的话吗？ 要为他说诡诈的言语吗？
JOB|13|8|你们要看上帝的情面吗？ 要为他争辩吗？
JOB|13|9|他查究你们，这岂是好事吗？ 人欺骗人，你们也要照样欺骗他吗？
JOB|13|10|你们若暗中看人的情面， 他必定要责备你们。
JOB|13|11|他的尊荣岂不叫你们惧怕吗？ 他岂不使惊吓临到你们吗？
JOB|13|12|你们可记念的谚语是灰烬的箴言； 你们的后盾是泥土的后盾。
JOB|13|13|“你们不要向我作声， 让我说话，无论如何我都承当。
JOB|13|14|我为何把我的肉挂在我的牙上， 将我的命放在我的手掌中呢？
JOB|13|15|看哪，他要杀我，我毫无指望 ， 然而我还要在他面前辩明我所行的。
JOB|13|16|这要成为我的拯救， 因为不虔诚的人不可到他面前。
JOB|13|17|你们要细听我的言语， 让我的申辩入你们耳中。
JOB|13|18|看哪，我已陈明我的案， 知道自己有义。
JOB|13|19|还有谁要和我争辩， 我现在就缄默不言，气绝而死。
JOB|13|20|惟有两件事不要向我施行， 我就不躲开你的面：
JOB|13|21|就是把你的手缩回，远离我身； 又不使你的威严恐吓我。
JOB|13|22|这样，你呼叫，我就回答； 或是让我说话，你回答我。
JOB|13|23|我的罪孽和我的罪有多少呢？ 求你叫我知道我的过犯与我的罪。
JOB|13|24|你为何转脸， 拿我当仇敌呢？
JOB|13|25|你要惊动被风吹的叶子吗？ 要追赶枯干的碎秸吗？
JOB|13|26|你写下苦楚对付我， 又使我担当幼年的罪孽。
JOB|13|27|你把我的脚锁上木枷， 察看我一切的道路， 为我的脚掌划定界限。
JOB|13|28|人像灭绝的烂物， 像虫蛀的衣裳。”
JOB|14|1|“人为妇人所生， 日子短少，多有患难。
JOB|14|2|他出来如花，凋谢而去； 他飞逝如影，不能存留。
JOB|14|3|这样的人你岂会睁眼看他， 又叫我 来，在你那里受审吗？
JOB|14|4|谁能使洁净出于污秽呢？ 谁也不能！
JOB|14|5|既然人的日子限定， 他的月数在于你， 你划定他的界限，他不能越过；
JOB|14|6|求你转眼不看他，使他得歇息， 直到他像雇工享受他的一天。
JOB|14|7|“因树有指望， 若被砍下，还可发芽， 嫩枝生长不息。
JOB|14|8|树根若衰老在地里， 树干也死在土中，
JOB|14|9|及至得了水气，还会发芽， 长出枝条，像新栽的树一样。
JOB|14|10|但壮士一死就消逝了； 人一气绝，他在何处呢？
JOB|14|11|海中的水枯竭， 江河消散干涸。
JOB|14|12|人一躺下就不再起来， 等到诸天没有了 ，仍不复醒， 也不能从睡中唤醒。
JOB|14|13|惟愿你把我藏在阴间， 把我隐藏，直到你的愤怒过去； 愿你为我定下期限，并记得我。
JOB|14|14|壮士若死了能再活吗？ 我在一切服役的日子中等待， 直到我退伍的时候来到。
JOB|14|15|你呼叫，我就回答你； 你手所做的，你必期待。
JOB|14|16|但如今你数点我的脚步， 不察看我的罪。
JOB|14|17|我的过犯被你密封在囊中， 你遮掩了我的罪孽。
JOB|14|18|“然而，山崩变为无有， 磐石从原处挪移。
JOB|14|19|流水冲蚀石头， 急流洗去地上的尘土； 你也照样灭绝人的指望。
JOB|14|20|你终必胜过人，使他消逝； 你改变他的容貌，把他送走。
JOB|14|21|他的儿子得尊荣，他不知道； 他们降为卑，他也不晓得。
JOB|14|22|他只觉得身上疼痛， 心中为自己悲哀。”
JOB|15|1|提幔 人 以利法 回答说：
JOB|15|2|“智慧人岂可用虚空的知识回答， 用东风充满自己的肚腹呢？
JOB|15|3|他岂可用无益的话， 用无济于事的言语理论呢？
JOB|15|4|你诚然废弃敬畏， 不在上帝面前默想。
JOB|15|5|你的罪孽指教你的口； 你选用诡诈人的舌头。
JOB|15|6|你自己的口定你有罪，并非是我； 你自己的嘴唇见证你的不是。
JOB|15|7|“你是头一个生下来的人吗？ 你受造在诸山之先吗？
JOB|15|8|你曾听见上帝的密旨吗？ 你要独自得尽智慧吗？
JOB|15|9|什么是你知道，我们不知道的呢？ 什么是你明白，我们不明白的呢？
JOB|15|10|我们这里有白发的和年老的， 比你父亲还年长。
JOB|15|11|上帝的安慰和对你温和的话， 你以为太小吗？
JOB|15|12|你的心为何失控， 你的眼为何冒火，
JOB|15|13|以致你的灵反对上帝， 你的口说出这样的言语呢？
JOB|15|14|人是什么，竟算为洁净呢？ 妇人所生的是什么，竟算为义呢？
JOB|15|15|看哪，上帝不信任他的众圣者； 在他眼前，天也不洁净，
JOB|15|16|何况那污秽可憎， 喝罪孽如水的世人呢！
JOB|15|17|“我指示你，你要听我； 我要陈述我所看见的，
JOB|15|18|就是智慧人从列祖所受， 传讲而不隐瞒的事。
JOB|15|19|这地惟独赐给他们， 并没有外人从他们中间经过。
JOB|15|20|恶人一生的日子绞痛难熬， 残暴人存留的年数也是如此。
JOB|15|21|惊吓的声音常在他耳中； 在平安时，毁灭者必临到他。
JOB|15|22|他不信自己能从黑暗中转回； 他被刀剑看守。
JOB|15|23|他飘流在外求食：‘哪里有食物呢？’ 他知道黑暗的日子在他手边预备好了。
JOB|15|24|急难困苦叫他害怕， 而且胜过他，好像君王预备上阵。
JOB|15|25|因他伸手攻击上帝， 逞强对抗全能者，
JOB|15|26|挺着颈项， 用盾牌坚厚的凸面向全能者直闯；
JOB|15|27|又因他的脸蒙上油脂， 腰上积满肥肉。
JOB|15|28|他住在荒凉的城镇， 房屋无人居住， 将成为废墟。
JOB|15|29|他不得富足， 财物不得常存， 产业在地上也不加增。
JOB|15|30|他不得脱离黑暗， 火焰要把他的嫩枝烧干； 因上帝口中的气，他要离去。
JOB|15|31|不要让他倚靠虚假，欺骗自己， 因虚假必成为他的报应。
JOB|15|32|他的日期未到之先，这事必实现； 他的枝子不得青绿。
JOB|15|33|他必像葡萄树，葡萄未熟就掉落； 又像橄榄树，一开花就凋谢。
JOB|15|34|因不敬虔之辈必不能生育， 受贿赂之人的帐棚必被火吞灭。
JOB|15|35|他们所怀的是毒害，所生的是罪孽， 肚腹里所预备的是诡诈。”
JOB|16|1|约伯 回答说：
JOB|16|2|“这样的话我听了许多； 你们全都是使人愁烦的安慰者。
JOB|16|3|如风的言语有穷尽吗？ 或者什么惹动你回答呢？
JOB|16|4|我也能说你们那样的话， 你们若处在我的景况， 我也可以堆砌言词攻击你们， 又可以向你们摇头。
JOB|16|5|但我必用口坚固你们， 颤动的嘴唇带来舒解。
JOB|16|6|“我若说话，痛苦仍不得缓解； 我若停止，痛苦就离开我吗？
JOB|16|7|但现在上帝使我困倦， 你使所有的亲友远离我，
JOB|16|8|你抓住我 ，成为见证起来攻击我； 我的枯瘦也当着我的面作证。
JOB|16|9|上帝发怒撕裂我，逼迫我， 向我咬牙切齿； 我的敌人怒目瞪我。
JOB|16|10|他们向我大大张口， 打我的耳光羞辱我， 聚在一起攻击我。
JOB|16|11|上帝把我交给不敬虔的人， 把我扔到恶人的手中。
JOB|16|12|我本是安逸，他折断我， 掐住我的颈项，把我摔碎， 又立我作他的箭靶。
JOB|16|13|他的弓箭手围绕我。 他刺破我的肾脏，并不留情， 把我的胆汁倾倒在地上。
JOB|16|14|他使我破裂，破裂又破裂， 如同勇士向我直闯。
JOB|16|15|“我把麻布缝在我的皮肤上， 把我的角放在尘土中。
JOB|16|16|我的脸因哭泣变红， 我的眼皮上有死荫。
JOB|16|17|我的手中却没有暴力， 我的祈祷也是纯洁的。
JOB|16|18|“地啊，不要遮盖我的血！ 不要让我的哀求有藏匿之处！
JOB|16|19|现今，看哪，在天有我的见证， 在上有我的保人。
JOB|16|20|我的朋友讥诮我， 我却向上帝眼泪汪汪。
JOB|16|21|愿人可与上帝理论， 如同人与朋友一样；
JOB|16|22|因为再过几年， 我必走那往而不返之路。”
JOB|17|1|“我的灵耗尽，我的日子消逝； 坟墓为我预备好了。
JOB|17|2|戏笑的人果真陪伴着我， 我的眼睛盯住他们的悖逆。
JOB|17|3|“愿你亲自为我付押担保。 谁还会与我击掌呢？
JOB|17|4|因你蒙蔽他们的心，使不明理， 所以你必不高举他们。
JOB|17|5|控告 朋友为了分享产业的， 他儿女的眼睛要失明。
JOB|17|6|“上帝使我成为人群中的笑谈， 他们吐唾沫在我脸上。
JOB|17|7|我的眼睛因忧愁昏花， 我的肢体全像影儿。
JOB|17|8|正直人因此必惊奇； 无辜的人要兴起攻击不敬虔之辈。
JOB|17|9|然而，义人要持守所行的道， 手洁的人要力上加力。
JOB|17|10|至于你们众人，再回来吧！ 你们中间，我找不到一个智慧人。
JOB|17|11|我的日子已经过去了， 我的谋算、我心的愿望已经断绝了。
JOB|17|12|他们以黑夜为白昼， 即使面临黑暗，以为亮光已近。
JOB|17|13|我若盼望阴间为我的家， 若下榻在黑暗中，
JOB|17|14|若对地府呼叫：‘你是我的父亲’， 若对虫呼叫：‘你是我的母亲、姊妹’，
JOB|17|15|这样，我的盼望在哪里呢？ 我所盼望的，谁能看见呢？
JOB|17|16|这盼望要下到阴间的门闩吗 ？ 要一起在尘土中安息吗 ？”
JOB|18|1|书亚 人 比勒达 回答说：
JOB|18|2|“你们寻索言语要到几时呢 ？ 你们要明白，然后我们才说话。
JOB|18|3|我们为何被视为畜生， 在你们眼中看为愚笨 呢？
JOB|18|4|在怒气中将自己撕裂的人哪， 难道大地要因你见弃、 磐石要挪开原处吗？
JOB|18|5|“恶人的亮光必要熄灭， 他的火焰必不照耀。
JOB|18|6|他帐棚中的亮光要变黑暗， 他上面的灯也必熄灭。
JOB|18|7|他强横的脚步必遭阻碍， 他的计谋必将自己绊倒。
JOB|18|8|他因自己的脚陷入网中， 走在缠人的网子上。
JOB|18|9|罗网必抓住他的脚跟， 陷阱必擒获他。
JOB|18|10|绳索为他藏在土里， 羁绊为他藏在路上。
JOB|18|11|四面的惊吓使他害怕， 在他脚跟后面追赶他。
JOB|18|12|他的力量必因饥饿衰败， 祸患要在他的旁边等候，
JOB|18|13|侵蚀他肢体的皮肤； 死亡的长子吞吃他的肢体。
JOB|18|14|他要从所倚靠的帐棚被拔出来， 带到使人惊恐的王那里。
JOB|18|15|不属他的必住在他的帐棚里， 硫磺必撒在他所住之处。
JOB|18|16|下边，他的根要枯干； 上边，他的枝子要剪除。
JOB|18|17|他的称号 从地上消失， 他的名字不在街上存留。
JOB|18|18|他必从光明中被驱逐到黑暗里， 他必被赶出世界。
JOB|18|19|他在自己百姓中必无子无孙， 在寄居之地也没有幸存者。
JOB|18|20|以后的人 要因他的日子惊讶， 以前的人 也被惊骇抓住。
JOB|18|21|不义之人的住处总是这样， 这就是不认识上帝之人的下场。”
JOB|19|1|约伯 回答说：
JOB|19|2|“你们搅扰我的心， 用言语压碎我要到几时呢？
JOB|19|3|你们这十次羞辱我， 苦待我也不以为耻。
JOB|19|4|果真我有错， 这错是在于我。
JOB|19|5|若你们真要向我夸大， 以我的羞辱来责备我，
JOB|19|6|就该知道是上帝倾覆我， 用罗网围绕我。
JOB|19|7|看哪，我喊冤叫屈，却不蒙应允； 我呼求，却没有公正。
JOB|19|8|上帝拦住我的道路，使我不得经过； 他使黑暗笼罩我的路径。
JOB|19|9|他剥去我的荣光， 摘去我头上的冠冕。
JOB|19|10|他在四围攻击我，我就走了； 他将我的指望如树拔出。
JOB|19|11|他向我发烈怒， 以我为他的敌人。
JOB|19|12|他的军队一齐上来， 修筑道路攻击我， 在我帐棚的四围安营。
JOB|19|13|“他把我的兄弟隔在远处， 使我认识的人全然与我生疏。
JOB|19|14|我的亲戚都离开了我； 我的密友都忘记了我。
JOB|19|15|在我家寄居的和我的使女， 都当我是陌生人； 我在他们眼中被视为外邦人。
JOB|19|16|我呼唤仆人，他却不回答； 我必须亲口求他。
JOB|19|17|我口的气味令我妻子厌恶， 我的同胞都憎恶我。
JOB|19|18|连小男孩也藐视我； 我起来，他们都嘲笑我。
JOB|19|19|我的知心朋友都憎恶我； 我平日所爱的人向我翻脸。
JOB|19|20|我的皮和肉紧贴骨头， 我得以逃脱，仅剩牙齿 。
JOB|19|21|我的朋友啊，可怜我！可怜我！ 因为上帝的手攻击我。
JOB|19|22|你们为什么仿佛上帝逼迫我， 吃我的肉还不满足呢？
JOB|19|23|“惟愿我的言语现在就写上， 都记录在书上；
JOB|19|24|用铁笔和铅， 刻在磐石上，存到永远。
JOB|19|25|我知道我的救赎主 活着， 末后他必站在尘土上。
JOB|19|26|我这皮肉灭绝之后 ， 我必在肉体之外 得见上帝。
JOB|19|27|我自己要见他， 亲眼要看他，并不像陌生人。 我的心肠在我里面耗尽了！
JOB|19|28|你们若说：‘我们怎么逼迫他呢？ 事情的根源是在于他 ’，
JOB|19|29|你们就当惧怕刀剑， 因为愤怒带来刀剑的刑罚。 这样，你们就知道有审判。”
JOB|20|1|拿玛 人 琐法 回答说：
JOB|20|2|“这样，我的思念叫我回答， 因为我心中急躁。
JOB|20|3|我听见那羞辱我的责备； 我悟性的灵回答我。
JOB|20|4|你岂不知道吗？亘古以来， 自从人被安置在地，
JOB|20|5|恶人欢乐的声音是暂时的， 不敬虔人的喜乐不过是转眼之间。
JOB|20|6|他的尊荣虽达到天上， 头虽顶到云中，
JOB|20|7|他必永远灭亡，像自己的粪一样。 看见他的人要说：‘他在哪里呢？’
JOB|20|8|他必如梦飞去，不再寻见； 他被赶走，如夜间的异象。
JOB|20|9|亲眼见过他的，必不再见他； 他自己的地方也不再见到他。
JOB|20|10|他的儿女要向穷人求恩； 他的手要赔还钱财。
JOB|20|11|他的骨头虽然满有年轻的活力， 却要和他一同躺卧在尘土之中。
JOB|20|12|“他口中以恶为甘甜， 把恶藏在舌头底下，
JOB|20|13|爱恋不舍， 含在口中。
JOB|20|14|他的食物在肚里却要翻转， 在他里面成为虺蛇的毒液。
JOB|20|15|他吞了财宝，还要吐出； 上帝要从他腹中掏出来。
JOB|20|16|他必吸饮虺蛇的毒汁， 毒蛇的舌头必杀他。
JOB|20|17|他不再看见溪流， 流奶与蜜之河。
JOB|20|18|他劳碌得来的要赔还，不得吞下； 赚取了财货，也不得欢乐。
JOB|20|19|他欺压穷人，弃之不顾， 强取非自己所盖的房屋 。
JOB|20|20|“他的肚腹不知安逸， 所贪恋的连一样也不放过，
JOB|20|21|剩余的没有一样他不吞吃， 所以他的福乐不能长久。
JOB|20|22|他在满足有余的时候，必有困苦临到； 凡受苦楚之人的手必加在他身上。
JOB|20|23|他的肚腹正要满足的时候， 上帝必将猛烈的愤怒降在他身上； 他正在吃饭的时候， 上帝要将这愤怒如雨降在他身上。
JOB|20|24|他要躲避铁的武器， 铜弓要将他射透。
JOB|20|25|箭一抽，就从他背上出来， 发亮的箭头从他胆中出来； 有惊惶临到他身上。
JOB|20|26|他的财宝隐藏在深沉的黑暗里； 有非人吹起的火要把他吞灭， 把他帐棚中所剩下的烧毁。
JOB|20|27|天要显明他的罪孽， 地要兴起去攻击他。
JOB|20|28|他家里出产的必消失， 在上帝愤怒的日子被冲走。
JOB|20|29|这是恶人从上帝所得的份， 是上帝为他所定的产业。”
JOB|21|1|约伯 回答说：
JOB|21|2|“你们要细心听我的言语， 这就算是你们的安慰。
JOB|21|3|请宽容我，我又要说话； 说了以后，任凭你嗤笑吧！
JOB|21|4|我岂是向人诉苦？ 我为何不是没有耐心呢？
JOB|21|5|你们要转向我而惊奇， 要用手捂口。
JOB|21|6|我每逢思想，心就惊惶， 战兢抓住我身。
JOB|21|7|恶人为何存活， 得享高寿，势力强盛呢？
JOB|21|8|他们的后裔与他们一起 ，坚立在他们面前， 他们得以眼见自己的子孙。
JOB|21|9|他们的家宅平安无惧， 上帝的杖不加在他们身上。
JOB|21|10|他们的公牛传种而不断绝， 母牛生牛犊而不掉胎。
JOB|21|11|他们打发小男孩出去，多如羊群， 他们的孩子踊跃跳舞。
JOB|21|12|他们随着琴鼓歌唱， 因箫声欢喜。
JOB|21|13|他们度日诸事亨通， 在平安中下到阴间。
JOB|21|14|他们对上帝说：‘离开我们吧！ 我们不想知道你的道路。
JOB|21|15|全能者是谁，我们何必事奉他呢？ 求告他有什么益处呢？’
JOB|21|16|看哪，他们亨通不是靠自己的手； 恶人的计谋离我好远。
JOB|21|17|“恶人的灯何尝熄灭？ 患难何尝临到他们呢？ 上帝何尝发怒，把灾祸分给他们呢？
JOB|21|18|他们何尝像风前的碎秸， 如暴风刮去的糠秕呢？
JOB|21|19|上帝为恶人的儿女积蓄罪孽， 不如本人遭报，好使他亲自知道。
JOB|21|20|愿他亲眼看见自己败亡， 亲自饮全能者的愤怒。
JOB|21|21|他的岁月既尽， 他身后还顾他的家吗？
JOB|21|22|谁能将知识教导上帝呢？ 是他审判那些居高位的。
JOB|21|23|有人至死身体强壮， 尽得平顺安逸；
JOB|21|24|他的肚腹充满奶汁 ， 他的骨髓滋润。
JOB|21|25|有人至死心中痛苦， 从未尝过福乐的滋味；
JOB|21|26|他们同样躺卧于尘土， 虫子覆盖他们。
JOB|21|27|“看哪，我知道你们的意念， 并残害我的计谋。
JOB|21|28|你们说：‘权贵的房屋在哪里？ 恶人住过的帐棚在哪里？’
JOB|21|29|你们没有询问那些过路的人吗？ 你们不承认他们的证据吗？
JOB|21|30|就是恶人在患难的日子得存留， 在愤怒的日子得逃脱。
JOB|21|31|他所行的，有谁当面给他说明？ 他所做的，有谁报应他呢？
JOB|21|32|然而他要被抬到坟地， 并有人看守墓穴。
JOB|21|33|他要以谷中的土块为甘甜； 人人要跟在他后面， 在他前面去的无数。
JOB|21|34|你们怎能以空话安慰我呢？ 你们的对答全都错谬！”
JOB|22|1|提幔 人 以利法 回答说：
JOB|22|2|“人能使上帝有益吗？ 智慧人能使他有益吗？
JOB|22|3|你为人公义，岂能叫全能者喜悦呢？ 你行为完全，岂能使他得利呢？
JOB|22|4|他岂是因你敬畏的心就责备你， 审判你吗？
JOB|22|5|你的罪恶岂不是大吗？ 你的罪孽不是没有穷尽吗？
JOB|22|6|因你无故强取弟兄的抵押， 剥去赤身者的衣服。
JOB|22|7|疲乏的人，你没有给他水喝； 饥饿的人，你没有给他食物。
JOB|22|8|有能力的人得土地； 尊贵的人住在其中。
JOB|22|9|你打发寡妇空手回去， 你折断孤儿的膀臂。
JOB|22|10|因此，有罗网环绕你， 有恐惧忽然使你惊惶；
JOB|22|11|或有黑暗使你看不见 ， 有洪水淹没你。
JOB|22|12|“上帝岂不是在高天吗？ 你看星宿的顶点何其高呢！
JOB|22|13|你说：‘上帝知道什么？ 他岂能透过幽暗施行审判呢？
JOB|22|14|密云将他遮盖，使他不能看见； 他周游穹苍。’
JOB|22|15|你要依从上古的道吗？ 这道是恶人行过的。
JOB|22|16|他们未到时候就被抓去 ； 他们的根基被江河冲去。
JOB|22|17|他们向上帝说：‘离开我们吧！’ 全能者能把他们怎么样呢？
JOB|22|18|然而，是上帝以美物充满他们的房屋； 恶人的计谋离我好远！
JOB|22|19|义人看见他们的结局 就欢喜； 无辜的人嗤笑他们：
JOB|22|20|‘攻击我们的果然被剪除， 剩余的都被火吞灭。’
JOB|22|21|“你要与上帝和好，要和平， 这样，福气必临到你。
JOB|22|22|你当领受他口中的教导， 将他的言语存在心里。
JOB|22|23|你若归向全能者，就必得建立。 你要从你帐棚中远离不义，
JOB|22|24|你要将黄金丢到尘土里， 将 俄斐 的金子丢在溪河石头之间；
JOB|22|25|全能者就必作你的黄金， 作你成堆的银子。
JOB|22|26|那时，你要以全能者为喜乐， 向上帝仰脸。
JOB|22|27|你要向他祷告，他就听你； 你也要还你的愿。
JOB|22|28|你定意要做何事，必然为你成就； 亮光也必照耀你的路。
JOB|22|29|当人降卑，你说：是因骄傲； 眼目谦卑的人，上帝必然拯救。
JOB|22|30|不是无辜的人，上帝尚且要搭救他 ； 他必因你手中的清洁得蒙拯救。”
JOB|23|1|约伯 回答说：
JOB|23|2|“如今我的哀告还算为悖逆； 我虽唉哼，他的手仍然重重责罚我 。
JOB|23|3|惟愿我知道哪里可以寻见上帝， 能到他的台前，
JOB|23|4|我就在他面前陈明我的案件， 满口辩诉。
JOB|23|5|我必知道他回答我的言语， 明白他向我所要说的。
JOB|23|6|他岂用大能与我争辩呢？ 不！他必理会我。
JOB|23|7|在那里正直人可以与他辩论， 我就必永远脱离那审判我的。
JOB|23|8|“看哪，我往前走，他不在那里； 往后退，也没有察觉他。
JOB|23|9|他在左边行事，我却看不见他； 他转向右边 ，我也见不到他。
JOB|23|10|然而他知道我所走的路； 他试炼我，我就如纯金。
JOB|23|11|我的脚紧跟他的步伐； 我谨守他的道，并不偏离。
JOB|23|12|他嘴唇的命令，我未曾背弃； 我看重他口中的言语，过于我需用的饮食 。
JOB|23|13|只是他心志已定，谁能使他转意呢？ 他心里所愿的，就行出来。
JOB|23|14|因此，为我所定的，他必做成， 这类的事他还有许多。
JOB|23|15|所以我在他面前惊惶； 我思想就惧怕他。
JOB|23|16|上帝使我丧胆， 全能者使我惊惶。
JOB|23|17|但我并非被黑暗剪除， 只是幽暗遮盖了我的脸。
JOB|24|1|“为何全能者不定下期限？ 为何认识他的人看不到那些日子呢？
JOB|24|2|有人挪移地界， 抢夺群畜去放牧。
JOB|24|3|他们拉走孤儿的驴， 强取寡妇的牛作抵押。
JOB|24|4|他们使贫穷人离开正道； 世上的困苦人尽都隐藏。
JOB|24|5|看哪，他们如同野驴出到旷野，殷勤寻找食物， 在野地给孩童糊口。
JOB|24|6|他们收割别人田间的庄稼， 摘取恶人剩余的葡萄。
JOB|24|7|他们终夜赤身无衣， 在寒冷中毫无遮盖。
JOB|24|8|他们在山上被大雨淋湿， 因没有避身之处就拥抱磐石。
JOB|24|9|又有人从母怀中抢走孤儿， 在困苦人身上强取抵押品 。
JOB|24|10|困苦人赤身无衣，到处流浪， 饿着肚子扛抬禾捆，
JOB|24|11|他们在围墙内榨油， 踹压酒池，自己却口渴。
JOB|24|12|在城内垂死的人呻吟， 受伤的人哀号； 上帝却不理会狂妄的事。
JOB|24|13|“又有人背弃光明， 不认识光明的道， 不留在光明的路上。
JOB|24|14|杀人者黎明起来， 杀害困苦人和贫穷人， 夜间又作盗贼。
JOB|24|15|奸夫的眼等候黄昏， 说：‘没有眼睛能见我’， 就把脸蒙住。
JOB|24|16|盗贼黑夜挖洞； 他们白日躲藏， 并不认识光明。
JOB|24|17|他们全都看早晨如死荫， 因为他们熟悉死荫的惊骇。
JOB|24|18|“恶人在水面上快速飘荡， 他们在地上所得的产业被诅咒； 无人再回到他们的葡萄园。
JOB|24|19|干旱炎热融化雪水； 阴间也如此吞没犯罪的人。
JOB|24|20|怀他的母胎忘记他； 虫子要吃他，觉得甘甜； 他不再被人记念； 不义的人必如树折断。
JOB|24|21|“他与不怀孕不生育的妇人交往 ， 却不善待寡妇。
JOB|24|22|然而上帝用能力保全有势力的人； 那性命难保的人仍然兴起。
JOB|24|23|上帝使他安稳，他就有所倚靠； 上帝的眼目看顾他们的道路。
JOB|24|24|他们高升，不过片刻就没有了； 他们降为卑，被除灭，与众人一样 ， 又如谷的穗子被割下。
JOB|24|25|若不是这样，谁能指证我是说谎的， 以我的言语为毫无根据呢？”
JOB|25|1|书亚 人 比勒达 回答说：
JOB|25|2|“上帝有统治之权，威严可畏； 他在高处施行和平。
JOB|25|3|他的军队岂能数算？ 他的光向谁不会升起呢 ？
JOB|25|4|这样，在上帝面前人怎能称义？ 妇人所生的怎能洁净？
JOB|25|5|看哪，在上帝眼前，月亮无光， 星宿也不皎洁，
JOB|25|6|更何况是如虫的人， 如蛆的世人呢！
JOB|26|1|约伯 回答说：
JOB|26|2|“无能的人蒙你何等的帮助！ 膀臂无力的人蒙你何等的拯救！
JOB|26|3|无智慧的人蒙你何等的指教！ 你向他显出丰富的知识。
JOB|26|4|你向谁发出言语？ 谁的灵从你而出？
JOB|26|5|在大水和水族以下， 阴魂战兢。
JOB|26|6|在上帝面前，阴间显露； 冥府 也不得遮掩。
JOB|26|7|上帝将北极铺在空中， 将大地悬在虚空。
JOB|26|8|他将水包在密云中， 盛水的云却不破裂。
JOB|26|9|他遮蔽宝座的正面， 把他的云彩铺在其上。
JOB|26|10|他在水面上划一圆圈， 直到光明与黑暗的交界。
JOB|26|11|天的柱子震动， 因他的斥责惊奇。
JOB|26|12|他以能力搅动 大海 ， 藉知识打伤 拉哈伯 。
JOB|26|13|他藉自己的灵使天空晴朗； 他的手刺杀爬得快的蛇。
JOB|26|14|看哪，这不过是上帝工作的些微； 我们听见他的话，是何等细微的声音！ 他大能的雷声谁能明白呢？”
JOB|27|1|约伯 继续发表他的言论说：
JOB|27|2|“我指着夺去我公道的永生上帝， 并使我心中愁苦的全能者起誓：
JOB|27|3|只要我的生命尚在我里面， 上帝所赐的气息仍在我鼻孔内，
JOB|27|4|我的唇绝不说不义， 我的舌也不说诡诈。
JOB|27|5|我断不以你们为义； 我至死不放弃自己的纯正！
JOB|27|6|我持定我的义，并不放松； 在世的日子，我的心不责备我。
JOB|27|7|“愿我的仇敌如恶人一样； 愿那起来攻击我的，如不义之人一般。
JOB|27|8|不敬虔的人有什么指望呢？ 上帝要剪除他，取他的性命。
JOB|27|9|患难临到他， 上帝岂听他的呼求？
JOB|27|10|他岂以全能者为乐， 随时求告上帝呢？
JOB|27|11|上帝手所做的，我要指教你们； 全能者所行的，我也不会隐瞒。
JOB|27|12|看哪，你们自己也都见过， 为何全变为这样虚妄呢？
JOB|27|13|“这是上帝为恶人所定的份， 残暴人从全能者所得的产业：
JOB|27|14|倘若他的儿女增多，仍被刀所杀； 他的子孙必不得饱食。
JOB|27|15|他遗留的人必死而埋葬， 他的寡妇也不哀哭。
JOB|27|16|他虽积蓄银子如尘沙， 堆积衣服如泥土，
JOB|27|17|他尽管堆积，义人却要穿上， 无辜的人却要分取银子。
JOB|27|18|他建造房屋如虫做窝， 又如守望者所搭的棚。
JOB|27|19|他虽富足躺卧，却不得收殓 ， 他张开眼睛，就不在了。
JOB|27|20|惊恐如洪水将他追上， 暴风在夜间将他刮去。
JOB|27|21|东风把他吹去，他就走了； 风将他刮离原地。
JOB|27|22|风 无情地击打他， 他试图逃脱风的手。
JOB|27|23|风要因他拍掌， 并要发叱声，使他离开原地。”
JOB|28|1|“银子有矿； 炼金有场。
JOB|28|2|铁从土里开采， 铜从矿石镕出。
JOB|28|3|人探索黑暗的尽头， 查究矿石直到极处， 那是幽暗和死荫；
JOB|28|4|他在无人居住之处开凿矿穴， 在无足迹之地被遗忘 ， 与人远离，悬空摇摆。
JOB|28|5|地出产粮食， 地底翻腾如火。
JOB|28|6|地的石头是蓝宝石之处， 那里还有金沙。
JOB|28|7|鸷鸟不知那条路， 鹰眼也未曾见过。
JOB|28|8|狂傲的野兽未曾踩踏， 猛烈的狮子也未曾经过。
JOB|28|9|“人动手凿开坚石， 翻倒山的根基，
JOB|28|10|在磐石中凿出水道， 亲眼看见各样宝物。
JOB|28|11|他封闭河川不得涓滴 ， 使隐藏之物显露出来。
JOB|28|12|“然而，智慧何处可寻？ 聪明之地在哪里？
JOB|28|13|智慧的价值 无人能知， 活人之地也无处可寻。
JOB|28|14|深渊说：‘不在我里面。’ 沧海说：‘不在我这里。’
JOB|28|15|智慧不可用黄金换取， 也不能用白银秤她的价值。
JOB|28|16|俄斐 的金子和贵重的红玛瑙， 以及蓝宝石，不足与她比拟；
JOB|28|17|黄金和玻璃不足与她比较； 纯金的器皿不足兑换她。
JOB|28|18|珊瑚、水晶都不值得提； 智慧的价值胜过宝石 。
JOB|28|19|古实 的红璧玺不足与她比较； 纯金也不足与她比拟。
JOB|28|20|“智慧从何处来呢？ 聪明之地在哪里？
JOB|28|21|她隐藏，远离众生的眼目， 她掩蔽，远离空中的飞鸟。
JOB|28|22|毁灭和死亡说： ‘我们风闻其名。’
JOB|28|23|“上帝明白智慧的道路， 知道智慧的所在。
JOB|28|24|因为他鉴察直到地极， 遍观普天之下，
JOB|28|25|要为风定轻重， 又度量诸水，
JOB|28|26|为雨定律例， 为雷电定道路。
JOB|28|27|那时他看见智慧，就谈论她， 坚定她，并且查究她。
JOB|28|28|他对人说：‘看哪，敬畏主就是智慧； 远离恶事就是聪明。’”
JOB|29|1|约伯 继续发表他的言论说：
JOB|29|2|“惟愿我如从前的岁月， 如上帝保护我的日子。
JOB|29|3|那时他的灯照在我头上， 我藉他的光行过黑暗。
JOB|29|4|在我壮年的时候， 上帝亲密的情谊临到我的帐棚中。
JOB|29|5|全能者仍与我同在， 我的儿女都环绕我。
JOB|29|6|我的脚洗在乳酪当中； 磐石为我流出油河。
JOB|29|7|我出到城门， 在广场安排座位，
JOB|29|8|年轻人见我而回避， 老年人起身站立。
JOB|29|9|王子都停止说话， 用手捂口；
JOB|29|10|领袖静默无声， 舌头贴住上膛。
JOB|29|11|耳朵听见了，称我有福； 眼睛看见了，就称赞我。
JOB|29|12|因我拯救了哀求的困苦人 和无人帮助的孤儿。
JOB|29|13|将要灭亡的为我祝福， 我使寡妇心中欢呼。
JOB|29|14|我穿上公义，它遮蔽我； 我的公平如外袍和冠冕。
JOB|29|15|我作瞎子的眼， 瘸子的脚。
JOB|29|16|我作贫穷人的父； 我不认识之人的案件，我也去查明。
JOB|29|17|我打破不义之人的大牙， 从他牙齿中夺走他所抢的。
JOB|29|18|我说：‘我要增添我的日子如尘沙， 我必死在自己家中 。
JOB|29|19|我的根伸展到水边， 露水夜宿我的枝上。
JOB|29|20|我的荣耀在我身上更新， 我的弓在我手中日新。’
JOB|29|21|“人听我说话而等候， 为我的教导而静默。
JOB|29|22|我说话之后，他们就不再说； 我的言语滴在他们身上。
JOB|29|23|他们等候我如等雨水， 又张口如切慕春雨。
JOB|29|24|我向他们微笑，他们不敢相信； 他们不使我脸上的光失色。
JOB|29|25|我为他们选择道路，又坐首位； 我如君王在军队中居住， 又如人安慰哀伤的人。”
JOB|30|1|“但如今，比我年轻的人讥笑我； 我曾藐视他们的父亲， 不放在我的牧羊犬中。
JOB|30|2|他们的精力既已衰败， 手中的气力于我何益？
JOB|30|3|他们因穷乏饥饿，没有生气， 在荒废凄凉的幽暗中啃干燥之地。
JOB|30|4|他们在草丛之中采咸草， 罗腾 树的根成为他们的食物。
JOB|30|5|他们从人群中被赶出， 人追喊他们如贼一般，
JOB|30|6|以致他们住在荒谷， 住在地洞和岩穴中。
JOB|30|7|他们在草丛中叫唤， 在荆棘下挤成一团。
JOB|30|8|这都是愚顽卑微人的儿女； 他们被鞭打，赶出境外。
JOB|30|9|“现在这些人以我为歌曲， 以我为笑谈。
JOB|30|10|他们厌恶我，躲避我， 不住地吐唾沫在我脸上。
JOB|30|11|上帝松开我的弓弦 使我受苦， 他们就在我面前脱去辔头。
JOB|30|12|这伙人在我右边起来， 他们推开我的脚， 筑灾难之路攻击我。
JOB|30|13|他们毁坏我的道， 加增我的灾害； 他们毋须人帮助。
JOB|30|14|他们来，如同闯进大缺口， 在暴风间滚动。
JOB|30|15|惊恐倾倒在我身上， 我的尊荣被逐如风； 我的福禄如云飘去。
JOB|30|16|“现在我的心极其悲伤， 困苦的日子将我抓住。
JOB|30|17|夜间，我里面的骨头刺痛， 啃着我的没有止息。
JOB|30|18|我的外衣因大力扭皱 ， 内衣的领子把我勒住。
JOB|30|19|上帝把我扔在淤泥之中， 我就像尘土和灰烬一样。
JOB|30|20|我呼求你，你不应允我； 我站起来，你只是望着我。
JOB|30|21|你对我变得残忍， 大能的手追逼我。
JOB|30|22|你把我提到风中，使我乘风而去， 使我消失在烈风之中。
JOB|30|23|我知道你要使我归于死亡， 到那为众生所定的阴宅。
JOB|30|24|“然而，人在废墟岂不伸手？ 遇灾难时一定呼救。
JOB|30|25|人遭难的日子，我岂不为他哭泣呢？ 人贫穷的时候，我岂不为他忧愁呢？
JOB|30|26|我仰望福气，灾祸就来到； 我等待光明，黑暗便来临。
JOB|30|27|我内心烦扰不安， 困苦的日子临到我身。
JOB|30|28|我在阴暗中行走，没有日光 ， 我在会众中站立求救。
JOB|30|29|我与野狗为弟兄， 我跟鸵鸟为同伴。
JOB|30|30|我的皮肤变黑脱落， 我的骨头因热烧焦。
JOB|30|31|我的琴音变为哀泣； 我的箫声变为哭声。”
JOB|31|1|“我与眼睛立约， 怎能凝望少女呢？
JOB|31|2|从至上的上帝所得之分， 从至高全能者所得之业是什么呢？
JOB|31|3|岂不是祸患临到不义的， 灾害临到作恶的吗？
JOB|31|4|上帝岂不察看我的道路， 数点我所有的脚步吗？
JOB|31|5|“我若与虚谎同行， 我脚若紧跟诡诈，
JOB|31|6|愿上帝用公道的天平秤我， 愿他知道我的纯正。
JOB|31|7|我的脚步若偏离正路， 我的心若随从我眼目， 我的手掌若粘有污秽；
JOB|31|8|愿我栽种，别人来吃， 我的农作物连根拔出。
JOB|31|9|“我心若因妇人受迷惑， 在邻舍的门外等候，
JOB|31|10|就愿我妻子给别人推磨， 别人与她同寝。
JOB|31|11|因为这是邪恶的事， 审判官裁定的罪孽。
JOB|31|12|这是一场火，直烧到毁灭 ， 必拔除我一切的家产。
JOB|31|13|“我的仆婢与我争辩， 我若藐视不听他们的冤情，
JOB|31|14|上帝兴起的时候，我怎样行呢？ 他察问的时候，我怎样回答他呢？
JOB|31|15|造我在母腹中的，不也是造了他吗？ 在母胎中使我们成形的，岂不是同一位吗？
JOB|31|16|“我若不让贫寒人遂其所愿， 或是叫寡妇眼中失望，
JOB|31|17|或独自吃自己的食物， 孤儿没有吃其中些许；
JOB|31|18|从我年轻时，孤儿就与我一同长大，我好像他的父亲， 我从出母腹就扶助寡妇 ；
JOB|31|19|我若见人因无衣死亡， 或见贫穷人毫无遮盖；
JOB|31|20|我若不使他真心为我祝福， 不使他因我羊的毛得暖；
JOB|31|21|我若举手攻击孤儿， 因为在城门口见有帮助我的；
JOB|31|22|情愿我的肩膀从肩胛骨脱落， 我的膀臂从肱骨折断。
JOB|31|23|因上帝降的灾祸使我恐惧 ， 因他的威严，我什么都不能。
JOB|31|24|“我若以黄金为我的指望， 对纯金说：你是我的倚靠；
JOB|31|25|我若因财物丰裕， 因手多得资财而欢喜；
JOB|31|26|我若见太阳发光， 明月运行，
JOB|31|27|心就暗暗被引诱， 口亲吻自己的手；
JOB|31|28|这也是审判官裁定的罪孽， 因为我背弃了至上的上帝。
JOB|31|29|“我若见恨我的遇难就欢喜， 见他遭灾就高兴；
JOB|31|30|其实我没有容许口犯罪， 以诅咒要他的性命；
JOB|31|31|若我帐棚中的人未曾说： ‘谁不以他的肉食吃饱呢？’
JOB|31|32|我未曾让旅客在街上过夜， 却开门迎接行路的人；
JOB|31|33|我若像 亚当 遮掩自己的过犯， 将罪孽藏在怀中；
JOB|31|34|我若因大大惧怕众人， 又因宗族的藐视而恐惧， 以致我缄默不言，闭门不出；
JOB|31|35|惟愿有一位肯听我！ 看哪，我的记号，愿全能者回答我！ 愿那与我争讼的写下状词！
JOB|31|36|我必把它带在肩上， 绑在头上为冠冕。
JOB|31|37|我必向上帝述说我脚步的数目， 如同王子进到他面前。
JOB|31|38|“若我的田地喊冤告我， 犁沟也一同哭泣；
JOB|31|39|我若吃地的出产不给银钱， 或叫地的原主丧命；
JOB|31|40|愿蒺藜生长代替麦子， 恶臭的草代替大麦。” 约伯 的话说完了。
JOB|32|1|于是这三个人因 约伯 看自己为义就停止，不再回答他。
JOB|32|2|那时 布西 人， 兰 族 巴拉迦 的儿子 以利户 发怒了。他向 约伯 发怒，因 约伯 自以为义，不以上帝为义。
JOB|32|3|他又向 约伯 的三个朋友发怒，因为他们想不出回答的话来，仍以 约伯 为有罪。
JOB|32|4|以利户 因为他们比自己年老，就等候要与 约伯 说话。
JOB|32|5|以利户 见这三个人口中无话回答，就发怒。
JOB|32|6|布西 人 巴拉迦 的儿子 以利户 回答说： “我年轻，你们年长， 因此我退让，不敢向你们陈述我的意见。
JOB|32|7|我说：‘年长的当先说话； 寿高的当以智慧教导人。’
JOB|32|8|其实，是人里面的灵， 全能者的气使人有聪明。
JOB|32|9|寿高的不都有智慧， 年老的不都明白公平。
JOB|32|10|因此我说：‘你们要听我， 我也要陈述我的意见。’
JOB|32|11|“看哪，我等候你们的话， 侧耳听你们的高见； 直到你们找到要说的言语。
JOB|32|12|我留心听你们， 看哪，你们中间无一人能折服 约伯 ， 回答他的话。
JOB|32|13|你们切不可说：‘我们寻得智慧； 上帝能胜他 ，人却不能。’
JOB|32|14|约伯 没有用言语与我争辩； 我也不用你们的话回答他。
JOB|32|15|“他们惊惶不再回答， 一言不发。
JOB|32|16|我岂因他们不说话， 因他们站住不再回答，仍旧等候呢？
JOB|32|17|我也要以我的一番话回答， 我也要陈述我的意见。
JOB|32|18|因为我满怀言语， 我里面的灵激动我。
JOB|32|19|看哪，我的肚腹如酒囊没有气孔， 又如新皮袋 快要破裂。
JOB|32|20|我要说话，使我舒畅； 我要张开嘴唇回答。
JOB|32|21|我必不看人的情面， 也不奉承人。
JOB|32|22|我不懂得奉承； 不然，造我的主必快快除灭我。”
JOB|33|1|“但是， 约伯 啊，请听我的言语， 侧耳听我一切的话。
JOB|33|2|看哪，我开口， 我的舌在上膛发言。
JOB|33|3|我的言语要表明心中的正直， 我嘴唇所知道的就诚实地说。
JOB|33|4|上帝的灵造了我， 全能者的气使我得生。
JOB|33|5|你若能够，就请回答我； 请你站起来，在我面前陈明。
JOB|33|6|看哪，我在上帝面前与你一样， 也是用泥土造成的。
JOB|33|7|看哪，我不用威严恐吓你， 也不用势力重压你。
JOB|33|8|“其实，你向我耳朵说话， 我听见你言语的声音：
JOB|33|9|‘我是纯洁无过的， 我是无辜的，在我里面没有罪孽。
JOB|33|10|看哪，上帝找机会攻击我， 以我为他的仇敌，
JOB|33|11|把我的脚锁上木枷， 察看我一切的道路。’
JOB|33|12|“看哪，你这话无理，我要回答你， 因上帝比世人更大。
JOB|33|13|你为何与他争论： ‘他任何事都不向人解答’？
JOB|33|14|上帝说一次、两次， 人却不理会。
JOB|33|15|世人在床上沉睡安眠时， 在梦中和夜间的异象里，
JOB|33|16|上帝就开通世人的耳朵， 把警告印在他们心上 ，
JOB|33|17|好叫人转离自己的行为， 叫壮士远离骄傲，
JOB|33|18|拦阻人不陷入地府， 不让他命丧刀下 。
JOB|33|19|“人在床上被疼痛惩治， 骨头不住地挣扎，
JOB|33|20|以致生命厌弃食物， 心中厌恶美味。
JOB|33|21|他的肉消瘦，难以看见； 先前看不见的骨头都凸出来。
JOB|33|22|他的性命临近地府， 他的生命挨近灭命者。
JOB|33|23|一千天使中， 若有一个作传话的临到他， 指示人所当行的事，
JOB|33|24|上帝就施恩给他，说： ‘要救赎他 免得下入地府， 我已经得了赎价。
JOB|33|25|他的肉要比孩童的肉更嫩； 他就返老还童。’
JOB|33|26|他向上帝祷告，上帝就悦纳他； 他必欢呼朝见上帝的面， 因上帝恢复他的义。
JOB|33|27|他在人前歌唱说： ‘我犯了罪，颠倒是非， 却没有受该得的报应。
JOB|33|28|上帝救赎我的性命免入地府， 我的生命也必见光。’
JOB|33|29|“看哪，上帝两次、三次 向人行这一切的事，
JOB|33|30|为要从地府救回人的性命， 使他被生命之光照耀。
JOB|33|31|约伯 啊，你当留心听我； 不要作声，我要说话。
JOB|33|32|你若有话说，可以回答我； 你只管说，因我愿以你为义。
JOB|33|33|若不然，你当听我； 不要作声，我要把智慧教导你。”
JOB|34|1|以利户 继续说：
JOB|34|2|“你们智慧人要听我的言语， 有知识的人要侧耳听我。
JOB|34|3|因为耳朵辨别言语， 好像上膛品尝食物。
JOB|34|4|我们当选择公理， 彼此知道何为善。
JOB|34|5|约伯 曾说：‘我是公义的， 上帝夺去我的公理。
JOB|34|6|我有理，岂能说谎呢？ 我无过，受的箭伤却不能医治。’
JOB|34|7|哪一个人像 约伯 ， 喝讥诮如同喝水呢？
JOB|34|8|他与作恶的结伴， 和恶人同行。
JOB|34|9|他说：‘人以上帝为乐， 总是无益。’
JOB|34|10|“所以，你们明理的人要听我， 上帝断不致行恶， 全能者断不致不义。
JOB|34|11|他必按人所做的报应人， 使各人照所行的得报。
JOB|34|12|确实地，上帝必不作恶， 全能者必不偏离公平。
JOB|34|13|谁派他治理大地？ 谁安定全世界呢？
JOB|34|14|他若专心为己， 将灵和气收归自己，
JOB|34|15|凡血肉之躯必一同死亡； 世人必归于尘土。
JOB|34|16|“你若明理，当听这话， 侧耳听我言语的声音。
JOB|34|17|难道恨恶公平的可以掌权吗？ 那有公义、有大能的，你岂可定他有罪呢？
JOB|34|18|你会对君王说：‘你是卑鄙的’； 对贵族说：‘你们是邪恶的’吗？
JOB|34|19|他待王子不徇情面， 也不看重富足的过于贫寒的， 因为他们都是他手所造的。
JOB|34|20|一瞬间他们就死亡。 百姓在半夜中被震动而去世； 有权力的被夺去，非藉人手。
JOB|34|21|“上帝的眼目观看人的道路， 察看他每一脚步。
JOB|34|22|没有黑暗，没有死荫， 能给作恶者在那里藏身。
JOB|34|23|上帝不必再三传人 到他面前受审判。
JOB|34|24|他毋须调查就粉碎有大能的人， 指定别人代替他们。
JOB|34|25|所以他知道他们的行为， 使他们在夜间倾倒压碎。
JOB|34|26|他在众目睽睽下击打他们， 如同击打恶人。
JOB|34|27|因为他们转离不跟从他， 不留心他一切的道，
JOB|34|28|甚至使贫寒人的哀声达到他那里； 他也听了困苦人的哀声。
JOB|34|29|他安静，谁能定罪呢？ 他转脸，谁能见他呢？ 无论一国或一人都是如此。
JOB|34|30|不虔敬的人不得作王， 免得百姓陷入圈套。
JOB|34|31|“有谁对上帝说： ‘我受了责罚，必不再犯罪；
JOB|34|32|我所看不明的，求你指教我； 我若行了不义，必不再行’？
JOB|34|33|他因你拒绝不接受， 就随你的心愿施行报应吗？ 选择的是你，不是我。 你所知道的，只管说吧！
JOB|34|34|明理的人必对我说， 听我的智慧人也说：
JOB|34|35|‘ 约伯 说话没有知识， 他的言语毫无智慧。’
JOB|34|36|愿 约伯 被考验到底， 因他回答像恶人一样。
JOB|34|37|他在罪上又加悖逆； 在我们中间引起疑惑 ， 用许多言语轻慢上帝。”
JOB|35|1|以利户 继续说：
JOB|35|2|“你以为这话有理， 说：‘我在上帝面前是公义的。’
JOB|35|3|你说：‘这对你有什么益处？ 我不犯罪有什么好处呢？’
JOB|35|4|至于我，我要用言语回答你 和跟你一起的朋友。
JOB|35|5|你要向天观看， 瞻望那高于你的穹苍。
JOB|35|6|你若犯罪，能使上帝受何害呢？ 你的过犯加增，能使上帝受何损呢？
JOB|35|7|你若是公义，能加增他什么呢？ 他从你手里还接受什么呢？
JOB|35|8|你的罪恶只影响像你这类的人； 你的公义也只影响世人。
JOB|35|9|“人因多受欺压就哀求， 因强权者的膀臂而求救。
JOB|35|10|但无人说：‘造我的上帝在哪里？ 他使人夜间歌唱，
JOB|35|11|教导我们多过地上的走兽， 使我们比空中的飞鸟更聪明。’
JOB|35|12|因为恶人骄傲， 他们在那里呼求，他却不回答。
JOB|35|13|虚妄的呼求，上帝必不垂听； 全能者必不留意。
JOB|35|14|何况你说，你不得见他。 案件就在他面前，你等候他吧。
JOB|35|15|但如今因他未曾发怒降罚， 也一点都不理会狂傲，
JOB|35|16|所以 约伯 开口说虚妄的话， 多多发表无知识的言语。”
JOB|36|1|以利户 继续说：
JOB|36|2|“你再给我片时，我就指示你， 因我还有话要为上帝说。
JOB|36|3|我要把我的知识从远处引来， 我要将公义归给造我的主。
JOB|36|4|我的言语绝不虚假， 有全备知识的与你同在。
JOB|36|5|“看哪，上帝有大能，并不藐视人； 他的心智能力广大。
JOB|36|6|他不让恶人活着， 却为困苦人伸冤。
JOB|36|7|他的眼目不远离义人， 却使他们和君王同坐宝座， 永远被高举 。
JOB|36|8|他们若被锁链捆住， 被苦难的绳索缠住，
JOB|36|9|他就向他们指示他们的作为和过犯， 以及他们的狂妄自大。
JOB|36|10|他也开通他们的耳朵来领受教导， 吩咐他们回转离开罪孽。
JOB|36|11|他们若听从事奉他， 就必度日亨通， 历年享福。
JOB|36|12|他们若不听从，就要被刀杀灭， 无知无识而死。
JOB|36|13|“那心中不敬虔的人积蓄怒气； 上帝捆绑他们，他们竟不求救。
JOB|36|14|他们必在青年时死亡， 与神庙娼妓一样丧命。
JOB|36|15|上帝藉着困苦救拔困苦人， 藉所受的欺压开通他们的耳朵。
JOB|36|16|上帝也必引你脱离患难， 进入宽阔不狭窄之地； 摆在你席上的必满有肥甘。
JOB|36|17|“但你充满着恶人的辩辞， 辩辞和审判抓住你。
JOB|36|18|不可让愤怒触动你，使你破口谩骂 ； 也不可因赎价大而偏行。
JOB|36|19|你的呼求 和一切的势力， 果真有用，使你不遭患难吗？
JOB|36|20|不要切慕黑夜， 就是众民在本处被除灭的时候。
JOB|36|21|你要谨慎，不可偏向罪孽， 因你选择罪孽过于苦难。
JOB|36|22|看哪，上帝因他的能力而崇高； 有谁像他那样作教师呢？
JOB|36|23|谁派定他的道路呢？ 谁能说：‘你行了不义’？
JOB|36|24|“你要记得颂赞他的作为， 就是人所歌颂的。
JOB|36|25|他的作为，万人都看见； 世人也从远处观看。
JOB|36|26|看哪，上帝崇高，我们不能知道； 他的年数，不能测度。
JOB|36|27|因他吸取水点， 水点就从云雾中变成雨；
JOB|36|28|云彩将雨落下， 沛然降于世人。
JOB|36|29|又有谁能明白密云如何铺张， 和上帝行宫的雷声呢？
JOB|36|30|看哪，他的亮光普照自己的四围； 他覆盖海的深处。
JOB|36|31|因他用这些审判 众民， 又赐丰富的粮食。
JOB|36|32|他以闪电遮手掌， 命令它击中靶子。
JOB|36|33|所发的雷声将他显明， 牲畜也指明要起暴风 。”
JOB|37|1|“因此我心战兢， 从原处移动。
JOB|37|2|听啊，听他轰轰的声音， 是上帝口中所发的响声。
JOB|37|3|他发响声震遍天下， 他的闪电直到地极。
JOB|37|4|随后，人听见他的声音， 是那轰轰的声音； 他发出威严的雷声， 而不加以遏止。
JOB|37|5|上帝发出奇妙的雷声； 他行大事，我们不能测透。
JOB|37|6|他对雪说：‘要降在地上’； 对大雨和暴雨也是这样说。
JOB|37|7|他封住各人的手， 叫所造的万人都知道他的作为。
JOB|37|8|野兽进入穴中， 卧在自己洞内。
JOB|37|9|暴风来自内宫， 寒冷出于狂风。
JOB|37|10|上帝嘘气成冰， 凝结宽阔之水，
JOB|37|11|使密云盛满水气， 乌云散布闪电。
JOB|37|12|云藉着他的指引游行旋转， 在世界的地面上行他一切所吩咐的，
JOB|37|13|或为责罚，或为他的地， 或为慈爱，都是他所行的。
JOB|37|14|“ 约伯 啊，侧耳听这话， 要站立，思想上帝奇妙的作为。
JOB|37|15|你知道上帝如何安排这些， 如何使云中的闪电照耀吗？
JOB|37|16|你知道云彩如何浮于空中， 知识全备者奇妙的作为吗？
JOB|37|17|你知道南风使地寂静， 你的衣服就变为热吗？
JOB|37|18|你岂能与上帝同铺穹苍， 坚固如同铸成的镜子吗？
JOB|37|19|我们因在黑暗中，不会陈说， 请你指教我们该对他说什么。
JOB|37|20|有人告诉他我要说话吗？ 岂有人说他愿被吞灭吗？
JOB|37|21|“现在，人不得见穹苍的亮光； 风一吹过，天色晴朗。
JOB|37|22|金色的光辉来自北方， 在上帝那里有可畏的威严。
JOB|37|23|全能者，我们不能测度； 他大有能力，又有公平， 满有公义，必不苦待人。
JOB|37|24|所以，世人敬畏他； 凡自以为 有智慧的，他都不看顾。”
JOB|38|1|那时，耶和华从旋风中回答 约伯 说：
JOB|38|2|“谁用无知的言语使我的旨意暗昧不明？
JOB|38|3|你要如勇士束腰； 我问你，你可以让我知道。
JOB|38|4|“我立大地根基的时候，你在哪里？ 你若明白事理，只管说吧！
JOB|38|5|你知道是谁定地的尺度， 是谁把准绳拉在其上吗？
JOB|38|6|地的根基安置在何处？ 地的角石是谁安放的？
JOB|38|7|那时，晨星一同歌唱； 上帝的众使者也都欢呼。
JOB|38|8|“当海水冲出，如出母胎， 谁用门将它关闭呢？
JOB|38|9|是我用云彩当海的衣服， 用幽暗当包裹它的布，
JOB|38|10|为它定界限， 又安门和闩，
JOB|38|11|说：‘你只可到这里，不可越过； 你狂傲的浪要到此止住。’
JOB|38|12|“你有生以来，曾命定晨光， 曾使黎明知道自己的地位，
JOB|38|13|抓住地的四极， 把恶人从其中驱逐出来吗？
JOB|38|14|地改变如泥上盖印， 万物出现如衣服一样。
JOB|38|15|亮光不照恶人， 高举的膀臂也必折断。
JOB|38|16|“你曾进到海之源， 或在深渊的隐密处行走吗？
JOB|38|17|死亡的门曾向你显露吗？ 死荫的门你曾见过吗？
JOB|38|18|地的广大，你能测透吗？ 你若全知道，只管说吧！
JOB|38|19|“往光明居所的路在哪里？ 黑暗的地方在何处？
JOB|38|20|你能将它带到其领域， 能辨明其居所之路吗？
JOB|38|21|你知道的，因为那时你已出生， 你活的日子数目也多。
JOB|38|22|“你曾进入雪之库， 或见过雹的仓吗？
JOB|38|23|雪雹是我为灾难的时候， 为打仗和战争的日子所预备。
JOB|38|24|光亮从何路分开？ 东风从何路分散遍地？
JOB|38|25|“谁为大雨分道， 谁为雷电开路，
JOB|38|26|使雨降在无人之地， 在无人居住的旷野，
JOB|38|27|使荒废凄凉之地得以丰足， 青草得以生长？
JOB|38|28|“雨有父亲吗？ 露珠是谁生的呢？
JOB|38|29|冰出于谁的胎？ 天上的霜是谁生的呢？
JOB|38|30|诸水坚硬如石头， 深渊之面凝结成冰。
JOB|38|31|“你能为昴星系结吗？ 你能为参星解带吗？
JOB|38|32|你能按时领出星宿吗？ 能引导北斗与其众星吗？
JOB|38|33|你知道天的定律吗？ 你能使地归其权下吗？
JOB|38|34|“你能向密云扬起声来， 使倾盆的雨遮盖你吗？
JOB|38|35|你能发出闪电，使它们 行走， 并对你说：‘我们在这里’吗？
JOB|38|36|谁将智慧放在朱鹭 中？ 谁将聪明赐给雄鸡 ？
JOB|38|37|谁能用智慧数算云彩？ 谁能倾倒天上的瓶呢？
JOB|38|38|那时，尘土聚集成团， 土块紧紧结连。
JOB|38|39|“你能为母狮抓取猎物， 使少壮的狮子饱足吗？
JOB|38|40|那时，它们在洞中蹲伏， 在隐密处埋伏。
JOB|38|41|谁能为乌鸦预备食物呢？ 那时，乌鸦之雏哀求上帝， 因无食物飞来飞去。”
JOB|39|1|“你知道岩石间的野山羊几时生产吗？ 你能观察母鹿下小鹿吗？
JOB|39|2|你能数算它们怀胎的月数吗？ 你知道它们几时生产吗？
JOB|39|3|它们屈身，生下幼儿， 就解除了阵痛。
JOB|39|4|其子渐渐肥壮，在荒野长大； 它们出去，不再归回。
JOB|39|5|“谁放野驴自由？ 谁解开快驴的绳索？
JOB|39|6|我使旷野作它的住处， 使盐地当它的居所。
JOB|39|7|它嘲笑城内的喧嚷， 不听赶牲口的喝声。
JOB|39|8|诸山是它漫游的草场， 它寻找各样青绿之物。
JOB|39|9|“野牛岂肯服事你？ 岂肯在你的槽旁过夜？
JOB|39|10|你岂能用套绳将野牛系于犁沟？ 它岂肯随你耙松山谷之地？
JOB|39|11|你岂可因它力大就倚靠它？ 岂可把你的工交给它做呢？
JOB|39|12|你岂能靠它把你的谷物运回， 又收聚在你的禾场上吗？
JOB|39|13|“鸵鸟的翅膀欢然拍动， 但岂是鹳的翎毛和羽毛吗 ？
JOB|39|14|因它把蛋留在地上， 使蛋在尘土中得温暖，
JOB|39|15|却忘记脚会把蛋踹碎， 野兽会践踏它。
JOB|39|16|它粗暴待雏，似乎不是自己生的； 虽徒然劳苦 ，也不惧怕。
JOB|39|17|因为上帝使它忘记智慧， 也未将悟性分给它。
JOB|39|18|它几时挺身展开翅膀， 就嘲笑马和骑马的人。
JOB|39|19|“马的力量是你所赐的吗？ 它颈项上的鬃是你披上的吗？
JOB|39|20|是你叫它跳跃像蝗虫吗？ 它喷气之威严使人惊惶。
JOB|39|21|它用蹄在谷中挖地 ，以能力欢跃； 它出去迎击仇敌 。
JOB|39|22|它嘲笑惧怕，并不惊惶， 也不因刀剑退却。
JOB|39|23|箭袋在它身上铮铮有声， 枪和短枪闪闪发亮。
JOB|39|24|它震颤激动，将地吞下 ； 一听角声就站不住。
JOB|39|25|每逢角声一响，它说：‘啊哈！’ 它从远处闻到战争的气息， 听见军官如雷的吼声和呐喊。
JOB|39|26|“鹰展开翅膀向南飞翔， 岂是藉着你的智慧吗？
JOB|39|27|大鹰上腾在高处搭窝， 岂是听你的指示吗？
JOB|39|28|它住在山岩， 以山峰和坚固之所为家，
JOB|39|29|从那里窥察食物， 眼睛自远方了望。
JOB|39|30|它的雏吸血； 被杀的人在哪里，它也在哪里。”
JOB|40|1|耶和华继续对 约伯 说：
JOB|40|2|“强辩的岂可与全能者争论？ 与上帝辩驳的可以回答吧！”
JOB|40|3|于是， 约伯 回答耶和华说：
JOB|40|4|“看哪，我是卑贱的！我用什么回答你呢？ 我只好用手捂住我的口。
JOB|40|5|我说了一次，就不回答； 说了两次，不再说了。”
JOB|40|6|于是，耶和华从旋风中回答 约伯 说：
JOB|40|7|“你要如勇士束腰； 我问你，你可以让我知道。
JOB|40|8|你岂可废弃我的判断？ 岂可定我有罪，好显自己为义吗？
JOB|40|9|你有上帝那样的膀臂吗？ 你能像他那样发雷声吗？
JOB|40|10|“你要以荣耀庄严为妆饰， 以尊荣威严为衣服。
JOB|40|11|你要发出你满溢的怒气， 见一切骄傲的人，使他降卑；
JOB|40|12|你见一切骄傲的人，将他制伏， 把恶人践踏在原来地方。
JOB|40|13|你将他们一同埋藏在尘土中， 把他们的脸遮蔽在隐密处 。
JOB|40|14|这样，我也向你承认， 你的右手能救你自己。
JOB|40|15|“看哪，我造河马， 也造了你； 它吃草像牛一样。
JOB|40|16|看哪，它的力气在腰间， 能力在肚腹的肌肉上。
JOB|40|17|它挺直 尾巴如香柏树， 它大腿的筋紧密结合。
JOB|40|18|它的骨头好像铜管； 它的肢体仿佛铁棍。
JOB|40|19|“它在上帝所造之物中为首， 只有创造它的能携刀临近它。
JOB|40|20|诸山为它产出食物， 百兽也在那里游玩。
JOB|40|21|它伏在莲叶之下， 在芦苇和沼泽的隐密处。
JOB|40|22|莲叶的阴影遮蔽它， 溪旁的柳树环绕它。
JOB|40|23|看哪，河水泛滥，它不慌张； 连 约旦河 涨到它口边，它也安然自若。
JOB|40|24|谁能在它眼前捉拿它呢？ 谁能以圈套穿它鼻子呢？”
JOB|41|1|“你能用鱼钩钓上 力威亚探 吗？ 能用绳子压下它的舌头吗？
JOB|41|2|你能用绳索穿它的鼻子吗？ 能用钩子穿它的腮骨吗？
JOB|41|3|它岂向你连连恳求， 向你说温柔的话吗？
JOB|41|4|它岂肯与你立约， 让你拿它永远作奴仆吗？
JOB|41|5|你岂可拿它当雀鸟玩耍？ 岂可将它系来给你幼女？
JOB|41|6|合伙的鱼贩岂可拿它当货物？ 他们岂可把它分给商人呢？
JOB|41|7|你能用倒钩扎满它的皮， 能用鱼叉叉满它的头吗？
JOB|41|8|把你的手掌按在它身上吧！ 想一想与它搏斗，你就不再这样做了！
JOB|41|9|看哪，对它有指望是徒然的； 一见它，岂不也丧胆吗？
JOB|41|10|没有那么凶猛的人敢惹它。 这样，谁能在我面前站立得住呢？
JOB|41|11|谁能与我对质，使我偿还呢？ 天下万物都是我的。
JOB|41|12|“我不能缄默不提 它的肢体和力量，以及健美的骨骼。
JOB|41|13|谁能剥它的外皮？ 谁能进它的铠甲之间 呢？
JOB|41|14|谁能开它的腮颊？ 它牙齿的四围是可畏的。
JOB|41|15|它的背上有一排排的鳞甲 ， 紧紧闭合，封得严密。
JOB|41|16|这鳞甲一一相连， 气不得透入其间，
JOB|41|17|互相连接， 胶结一起，不能分开。
JOB|41|18|它打喷嚏就发出光来， 它的眼睛好像晨曦 。
JOB|41|19|从它口中发出烧着的火把， 有火星飞迸出来；
JOB|41|20|从它鼻孔冒出烟来， 如烧开的锅在沸腾 。
JOB|41|21|它的气点着煤炭， 有火焰从它口中发出。
JOB|41|22|它颈项中存着劲力， 恐惧在它面前蹦跳。
JOB|41|23|它的肉块紧紧结连， 紧贴其身，不能摇动。
JOB|41|24|它的心结实如石头， 如下面的磨石那样结实。
JOB|41|25|它一起来，神明都恐惧， 因崩溃而惊慌失措。
JOB|41|26|人用刀剑扎它，是无用的， 枪、标枪、尖枪也一样。
JOB|41|27|它以铁为干草， 以铜为烂木。
JOB|41|28|箭不能使它逃走， 它看弹石如碎秸。
JOB|41|29|它当棍棒作碎秸， 它嘲笑短枪的飕飕声。
JOB|41|30|它肚腹下面是尖瓦片； 它如钉耙刮过淤泥。
JOB|41|31|它使深渊滚沸如锅， 使海洋如锅中膏油。
JOB|41|32|它使走过以后的路发光， 令人觉得深渊如同白发。
JOB|41|33|尘世上没有像它那样的受造物， 一无所惧。
JOB|41|34|凡高大的，它盯着看； 它在一切狂傲的野兽中作王。”
JOB|42|1|约伯 回答耶和华说：
JOB|42|2|“我知道，你万事都能做； 你的计划不能拦阻。
JOB|42|3|谁无知使你的旨意隐藏呢？ 因此我说的，我不明白； 这些事太奇妙，是我不知道的。
JOB|42|4|求你听我，我要说话； 我问你，求你让我知道。
JOB|42|5|我从前风闻有你， 现在亲眼看见你。
JOB|42|6|因此我撤回 ， 在尘土和炉灰中懊悔。”
JOB|42|7|耶和华对 约伯 说话以后，耶和华就对 提幔 人 以利法 说：“我的怒气向你和你两个朋友发作，因为你们议论我，不如我的仆人 约伯 说的正确。
JOB|42|8|现在你们要为自己取七头公牛，七只公羊，到我的仆人 约伯 那里去，为自己献上燔祭，我的仆人 约伯 就为你们祈祷。我必悦纳他，不按你们的愚妄处置你们。你们议论我，不如我的仆人 约伯 说的正确。”
JOB|42|9|于是 提幔 人 以利法 、 书亚 人 比勒达 、 拿玛 人 琐法 遵照耶和华所吩咐的去做，耶和华就悦纳 约伯 。
JOB|42|10|约伯 为他的朋友祈祷。耶和华就使 约伯 从苦境 中转回，并且耶和华赐给他的比他从前所有的加倍。
JOB|42|11|约伯 的兄弟、姊妹，和以前所认识的人都来到他那里，在他家里跟他一同吃饭。他们因耶和华所降于他的一切灾祸，都为他悲伤，安慰他。每人送他一块可锡塔 和一个金环。
JOB|42|12|这样，耶和华后来赐福给 约伯 比先前更多。他有一万四千只羊，六千匹骆驼，一千对牛，一千匹母驴。
JOB|42|13|他也有七个儿子，三个女儿。
JOB|42|14|他给长女起名叫 耶米玛 ，次女叫 基洗亚 ，三女叫 基连哈朴 。
JOB|42|15|在全地的妇女中找不着像 约伯 的女儿那样美貌的。她们的父亲使她们在兄弟中得产业。
JOB|42|16|此后， 约伯 又活了一百四十年，得见他的四代儿孙。
JOB|42|17|这样， 约伯 年纪老迈，日子满足而死。
PS|1|1|不从恶人的计谋， 不站罪人的道路， 不坐傲慢人的座位， 惟喜爱耶和华的律法， 昼夜思想 他的律法； 这人便为有福！
PS|1|2|
PS|1|3|他要像一棵树栽在溪水旁， 按时候结果子， 叶子也不枯干。 凡他所做的尽都顺利。
PS|1|4|恶人并不是这样， 却像糠秕被风吹散。
PS|1|5|因此，当审判的时候恶人必站立不住， 罪人在义人的会众中也是如此。
PS|1|6|因为耶和华知道义人的道路， 恶人的道路却必灭亡。
PS|2|1|列国为什么争闹？ 万民为什么图谋虚妄？
PS|2|2|世上的君王都站稳， 臣宰一同算计， 要对抗耶和华， 对抗他的受膏者：
PS|2|3|“我们要挣脱他们的捆绑， 脱去他们的绳索。”
PS|2|4|那坐在天上的必讥笑， 主必嗤笑他们。
PS|2|5|那时，他要在怒中责备他们， 在烈怒中惊吓他们：
PS|2|6|“我已经在 锡安 －我的圣山 膏立了我的君王。”
PS|2|7|我要传耶和华的圣旨， 他对我说：“你是我的儿子， 我今日生了你。
PS|2|8|你求我，我就将列国赐你为基业， 将地极赐你为田产。
PS|2|9|你必用铁杖打破他们， 把他们如同陶匠的瓦器摔碎。”
PS|2|10|现在，君王啊，应当谨慎！ 世上的审判官哪，要听劝戒！
PS|2|11|当存敬畏的心事奉耶和华， 又当战兢而快乐。
PS|2|12|当亲吻儿子，免得他发怒， 你们就在半途中灭亡， 因为他的怒气快要发作。 凡投靠他的，都是有福的。
PS|3|1|耶和华啊，我的敌人何其增多！ 许多人起来攻击我。
PS|3|2|许多人议论我： “他得不到上帝的帮助。”（细拉）
PS|3|3|但你－耶和华是我四围的盾牌， 是我的荣耀，又是令我抬起头来的。
PS|3|4|我用我的声音求告耶和华， 他就从他的圣山上应允我。（细拉）
PS|3|5|我躺下，我睡觉，我醒来， 耶和华都保佑我。
PS|3|6|虽有成万的百姓周围攻击我， 我也不惧怕。
PS|3|7|耶和华啊，求你兴起！ 我的上帝啊，求你救我！ 因为你打断我所有仇敌的腮骨， 敲碎了恶人的牙齿。
PS|3|8|救恩属于耶和华； 愿你赐福给你的百姓。（细拉）
PS|4|1|显我为义的上帝啊， 我呼求的时候，求你应允我！ 我在困境中，你曾使我宽畅； 求你怜悯我，听我的祷告！
PS|4|2|你们这些人哪，你们把我的尊荣变为羞辱，要到几时呢？ 你们喜爱虚妄，寻找虚假，要到几时呢？ （细拉）
PS|4|3|你们要知道，耶和华已将虔诚人分别出来归他自己； 我求告耶和华，他必垂听。
PS|4|4|应当畏惧，不可犯罪； 在床上的时候，要心里思想，并要安静。（细拉）
PS|4|5|当献上公义的祭， 又当倚靠耶和华。
PS|4|6|有许多人说：“谁能指示我们什么好处？ 耶和华啊，求你用你脸上的光照耀我们。”
PS|4|7|你使我心里喜乐， 胜过那丰收五谷新酒的人。
PS|4|8|我必平安地躺下睡觉， 因为独有你－耶和华使我安然居住。
PS|5|1|耶和华啊，求你侧耳听我的言语， 顾念我的心思！
PS|5|2|我的王，我的上帝啊，求你留心听我呼求的声音！ 因为我向你祈祷。
PS|5|3|耶和华啊，早晨你必听我的声音； 早晨我要向你陈明我的心思，并要警醒。
PS|5|4|因为你不是喜爱邪恶的上帝， 恶人不能与你同住。
PS|5|5|狂傲的人不能站在你眼前； 凡作恶的，都是你所恨恶的。
PS|5|6|说谎言的，你必灭绝； 好流人血、玩弄诡诈的，都为耶和华所憎恶。
PS|5|7|至于我，我必凭你丰盛的慈爱进入你的居所， 我要存敬畏你的心向你的圣殿下拜。
PS|5|8|耶和华啊，求你因我仇敌的缘故，凭你的公义引领我， 使你的道路在我面前正直。
PS|5|9|因为他们口中没有诚实， 心里充满邪恶， 他们的喉咙是敞开的坟墓； 他们用舌头谄媚人。
PS|5|10|上帝啊，求你定他们的罪！ 愿他们因自己的计谋跌倒； 求你因他们过犯众多赶逐他们， 因为他们背叛了你。
PS|5|11|凡投靠你的，愿他们喜乐，时常欢呼， 因为你庇护他们； 又愿那爱你名的人都靠你欢欣。
PS|5|12|耶和华啊，因为你必赐福给义人， 你必用恩惠如同盾牌四面护卫他。
PS|6|1|耶和华啊，求你不要在怒中责备我， 不要在烈怒中惩罚我！
PS|6|2|耶和华啊，求你怜悯我，因为我软弱。 耶和华啊，求你医治我，因为我的骨头战抖。
PS|6|3|我的心也大大惊惶。 耶和华啊，你要等到几时呢？
PS|6|4|耶和华啊，求你转回搭救我， 因你的慈爱拯救我。
PS|6|5|因为死了的人不会记念你， 在阴间有谁称谢你？
PS|6|6|我因呻吟而困乏； 我每夜流泪，使床铺漂起， 把褥子湿透。
PS|6|7|我的眼睛因忧愁而昏花， 因敌人的缘故，我的眼目模糊不清。
PS|6|8|你们所有作恶的人，离开我吧！ 因为耶和华听了我哀哭的声音。
PS|6|9|耶和华听了我的恳求， 耶和华必接纳我的祷告。
PS|6|10|我所有的仇敌都必羞愧，大大惊惶； 转眼之间，他们要羞愧撤退。
PS|7|1|耶和华－我的上帝啊，我投靠你！ 求你救我脱离所有追赶我的人，搭救我出来！
PS|7|2|免得他们像狮子撕裂我， 甚至撕碎，无人搭救。
PS|7|3|耶和华－我的上帝啊，我若行了这事， 若有罪孽在我手里，
PS|7|4|我若以恶回报我的朋友， 连那无故与我为敌的，我也救了他 ，
PS|7|5|就任凭仇敌追赶我，直到追上， 把我的性命踏在地上， 使我的荣耀归于灰尘。（细拉）
PS|7|6|耶和华啊，求你在怒中起来， 挺身而立，抵挡我敌人的烈怒！ 求你为我兴起！你已经发令施行审判。
PS|7|7|愿万民聚集环绕你！ 愿你居高位统治他们！
PS|7|8|耶和华向万民施行审判； 耶和华啊，求你按我的公义 和我心中的纯正判断我。
PS|7|9|愿恶人的恶断绝！ 愿你坚立义人！ 因为公义的上帝察验人的心肠肺腑。
PS|7|10|上帝是我的盾牌， 他拯救心里正直的人。
PS|7|11|上帝是公义的审判者， 又是天天向恶人发怒的上帝。
PS|7|12|若有人不回头，他的刀必磨快， 弓必上弦，预备妥当。
PS|7|13|他也预备了致死的兵器， 他所射的是火箭。
PS|7|14|看哪，恶人怀邪恶， 养毒害，生虚假。
PS|7|15|他掘了坑，挖得太深， 竟掉在自己所挖的陷阱里。
PS|7|16|他的毒害必回到自己头上， 他的残暴必落到自己的脑袋上。
PS|7|17|我要照着耶和华的公义称谢他， 要歌颂耶和华至高者的名。
PS|8|1|耶和华－我们的主啊， 你的名在全地何其美！ 你将你的荣耀彰显于天 。
PS|8|2|你因敌人的缘故， 从孩童和吃奶的口中建立了能力， 使仇敌和报仇的闭口无言。
PS|8|3|我观看你手指所造的天， 并你所陈设的月亮星宿。
PS|8|4|人算什么，你竟顾念他！ 世人算什么，你竟眷顾他！
PS|8|5|你使他比上帝 微小一点， 赐他荣耀尊贵为冠冕。
PS|8|6|你派他管理你手所造的， 使万物，就是一切的牛羊、 田野的牲畜、空中的鸟、海里的鱼， 凡游在水里的，都服在他的脚下。
PS|8|7|
PS|8|8|
PS|8|9|耶和华－我们的主啊， 你的名在全地何其美！
PS|9|1|我要一心称谢耶和华， 传扬你一切奇妙的作为。
PS|9|2|我要因你欢喜快乐； 至高者啊，我要歌颂你的名！
PS|9|3|我的仇敌回转撤退的时候， 他们在你面前跌倒灭亡。
PS|9|4|因你已经为我伸冤，为我辩护； 你坐在宝座上，按公义审判。
PS|9|5|你曾斥责列国，灭绝恶人； 你曾涂去他们的名，直到永永远远。
PS|9|6|仇敌到了尽头； 他们遭毁坏，直到永远。 你拆毁他们的城镇， 连他们的名字 也都消灭！
PS|9|7|惟耶和华坐在王位上，直到永远； 他已经为审判摆设宝座。
PS|9|8|他要按公义审判世界， 按正直判断万民。
PS|9|9|耶和华要作受欺压者的庇护所， 在患难时的庇护所。
PS|9|10|耶和华啊，认识你名的人要倚靠你， 因你没有离弃寻求你的人。
PS|9|11|应当歌颂居于 锡安 的耶和华， 将他所做的传扬在万民中。
PS|9|12|那位追讨流人血的， 他记念受屈的人， 不忘记困苦人的哀求。
PS|9|13|耶和华啊，求你怜悯我！ 你是从死门把我提升起来的， 求你看那恨我的人所加给我的苦难，
PS|9|14|好让我述说你一切的美德。 我要在 锡安 的城门因你的救恩欢乐。
PS|9|15|外邦人陷在自己所掘的坑中， 他们的脚被自己暗设的网罗缠住了。
PS|9|16|耶和华已将自己显明，他已施行审判； 恶人被自己手所做的缠住了 。（细拉）
PS|9|17|恶人，就是忘记上帝的外邦人， 都必归到阴间。
PS|9|18|贫穷人必不永久被忘， 困苦人的指望必不永远落空。
PS|9|19|耶和华啊，求你兴起，不容世人得胜！ 愿外邦人在你面前受审判！
PS|9|20|耶和华啊，求你使他们恐惧， 愿外邦人知道自己不过是人。（细拉）
PS|10|1|耶和华啊，你为什么站在远处？ 在患难的时候为什么隐藏？
PS|10|2|恶人骄横地追逼困苦人； 愿他们陷在自己所设的计谋里。
PS|10|3|因为恶人以自己的心愿自夸， 贪财的背弃耶和华，并且轻慢他 。
PS|10|4|恶人面带骄傲，不寻找耶和华； 他的思想中全无上帝。
PS|10|5|他的路时常亨通， 你的审判不在他眼里。 至于他所有的敌人，他都向他们发怒气。
PS|10|6|他心里说：“我必不动摇， 世世代代不遭灾难。”
PS|10|7|他满口咒骂、诡诈、欺压， 舌底尽是毒害、奸恶。
PS|10|8|他在村庄埋伏等候， 在隐密处杀害无辜的人， 他的眼睛窥探无倚无靠的人。
PS|10|9|他埋伏在暗地，如狮子蹲在洞中。 他埋伏，要俘掳困苦人； 他拉网，就把困苦人掳去。
PS|10|10|他屈身蹲伏， 无倚无靠的人就倒在他的暴力之下。
PS|10|11|他心里说：“上帝竟忘记了， 上帝转脸永不观看。”
PS|10|12|耶和华啊，求你兴起！ 上帝啊，求你举手！ 不要忘记困苦人！
PS|10|13|恶人为何轻慢上帝， 心里说“你必不追究”？
PS|10|14|你已经察看， 顾念人的忧患和愁苦， 放在你的手中。 无倚无靠的人把自己交托给你， 你向来是帮助孤儿的。
PS|10|15|求你打断恶人的膀臂， 至于坏人，求你追究他的恶，直到净尽。
PS|10|16|耶和华永永远远为王， 外邦人从他的地已经灭绝了。
PS|10|17|耶和华啊，困苦人的心愿你早已听见； 你必坚固他们的心，也必侧耳听他们的祈求，
PS|10|18|为要给孤儿和受欺压的人伸冤， 使世上的人不再威吓他们。
PS|11|1|我投靠耶和华； 你们怎么对我说：“你当像鸟逃到你们的山去；
PS|11|2|看哪，恶人弯弓，把箭搭在弦上， 要在暗中射那心里正直的人。
PS|11|3|根基若毁坏， 义人还能做什么呢？”
PS|11|4|耶和华在他的圣殿里， 耶和华在天上的宝座上； 他的眼睛察看， 他的眼目 察验世人。
PS|11|5|耶和华考验义人； 惟有恶人和喜爱暴力的人，他心里恨恶。
PS|11|6|他要向恶人密布罗网， 烈火、硫磺、热风作他们杯中的份。
PS|11|7|因为耶和华是公义的，他喜爱义行， 正直人必得见他的面。
PS|12|1|耶和华啊，求你帮助，因虔诚人断绝了， 世人中间忠信的人消失了。
PS|12|2|人人向邻舍说谎； 他们说话嘴唇油滑，心口不一。
PS|12|3|愿耶和华剪除一切油滑的嘴唇， 夸大的舌头。
PS|12|4|他们说：“我们必能以舌头取胜， 我们的嘴唇是自己的， 谁能作我们的主呢？”
PS|12|5|耶和华说：“因为困苦人的冤屈 和贫穷人的叹息， 我现在要起来， 把他安置在他所切慕的稳妥之地。”
PS|12|6|耶和华的言语是纯净的言语， 如同银子在泥做的炉中炼过七次。
PS|12|7|耶和华啊，你必保护他们， 你必保佑他们永远脱离这世代的人。
PS|12|8|卑鄙的人在世人中高升时， 就有恶人四处横行。
PS|13|1|耶和华啊，你忘记我要到几时呢？要到永远吗？ 你转脸不顾我要到几时呢？
PS|13|2|我心里筹算，终日愁苦，要到几时呢？ 我的仇敌升高压制我，要到几时呢？
PS|13|3|耶和华－我的上帝啊，求你看顾我，应允我！ 求你使我眼目明亮，免得我沉睡至死；
PS|13|4|免得我的仇敌说“我胜了他”； 免得我的敌人在我动摇的时候喜乐。
PS|13|5|但我倚靠你的慈爱， 我的心因你的救恩快乐。
PS|13|6|我要向耶和华歌唱， 因他厚厚地恩待我。
PS|14|1|愚顽人心里说：“没有上帝。” 他们都败坏，行了可憎恶的事， 没有一个人行善。
PS|14|2|耶和华从天上垂看世人， 要看有明白的没有， 有寻求上帝的没有。
PS|14|3|他们都偏离正路，一同变为污秽， 没有行善的， 连一个也没有。
PS|14|4|作恶的都没有知识吗？ 他们吞吃我的百姓如同吃饭一样， 并不求告耶和华。
PS|14|5|他们在那里大大害怕， 因为上帝在义人的族类中。
PS|14|6|你们叫困苦人的筹算变为羞辱， 然而耶和华是他的避难所。
PS|14|7|但愿 以色列 的救恩出自 锡安 。 当耶和华救回他被掳子民的时候， 雅各 要快乐， 以色列 要欢喜。
PS|15|1|耶和华啊，谁能寄居你的帐幕？ 谁能居住你的圣山？
PS|15|2|就是行为正直、做事公义、 心里说实话的人。
PS|15|3|他不以舌头谗害人， 不恶待朋友， 也不随伙毁谤邻舍。
PS|15|4|他眼中藐视匪类， 却尊重那敬畏耶和华的人。 他发了誓，虽然自己吃亏也不更改。
PS|15|5|他不放债取利， 不受贿赂以害无辜。 做这些事的人必永不动摇。
PS|16|1|上帝啊，求你保佑我， 因为我投靠你。
PS|16|2|我 曾对耶和华说：“你是我的主， 我的福气惟独从你而来。”
PS|16|3|论到世上的圣民，他们是尊贵的人， 是我最喜悦的。
PS|16|4|追逐 别神的， 他们的愁苦必增加； 他们所浇奠的血我不献上， 我嘴唇也不提别神的名号。
PS|16|5|耶和华是我的产业，是我杯中的福分； 我所得的，你为我持守。
PS|16|6|用绳量给我的地界，坐落在佳美之处； 我的产业实在美好。
PS|16|7|我要称颂那指引我的耶和华， 在夜间我的心肠也指教我。
PS|16|8|我让耶和华常在我面前， 因他在我右边，我就不致动摇。
PS|16|9|因此，我的心欢喜，我的灵 快乐； 我的肉身也要安然居住。
PS|16|10|因为你必不将我的灵魂 撇在阴间， 也不让你的圣者见地府 。
PS|16|11|你必将生命的道路指示我。 在你面前有满足的喜乐， 在你右手中有永远的福乐。
PS|17|1|耶和华啊，求你垂听公义的呼声， 留心听我的呼求！ 求你侧耳听我这没有诡诈的嘴唇的祈祷！
PS|17|2|愿判我公正的话从你面前发出， 愿你的眼睛察看正直。
PS|17|3|你已经考验我的心， 你在夜间鉴察我。 你熬炼我，却找不到错失， 我立志叫我口中没有过失。
PS|17|4|论到人的行为，我谨守你嘴唇的言语， 不走残暴人的道路。
PS|17|5|我的脚紧紧跟随你的脚踪， 我的两脚未曾滑跌。
PS|17|6|上帝啊，我求告你，因为你必应允我； 求你向我侧耳，听我的言语。
PS|17|7|求你显出你奇妙的慈爱， 你用右手拯救投靠你的人，脱离那起来攻击他们的人。
PS|17|8|求你保护我，如同保护眼中的瞳人， 把我隐藏在你翅膀的荫下，
PS|17|9|使我脱离欺压我的恶人， 脱离那围困我要害我命的仇敌。
PS|17|10|他们的心被油脂包裹， 用口说骄傲的话。
PS|17|11|他们追逼我 ，现在他们围困了我们， 瞪着眼，要把我们推倒在地。
PS|17|12|他像狮子要贪吃猎物， 又像少壮狮子蹲伏在暗处。
PS|17|13|耶和华啊，求你兴起，前去迎敌，把他打倒！ 求你用你的刀救我的命脱离恶人。
PS|17|14|耶和华啊，求你用手救我脱离世人， 脱离那只在今生有福分的世人！ 你以财宝充满他们的肚腹， 他们因有儿女就满足， 将其余的财物留给他们的孩子。
PS|17|15|至于我，我必因公正得见你的面； 我醒了的时候，你的形像使我满足。
PS|18|1|耶和华我的力量啊，我爱你！
PS|18|2|耶和华是我的岩石、我的山寨、我的救主、 我的上帝、我的磐石、我所投靠的。 他是我的盾牌， 是拯救我的角，是我的碉堡。
PS|18|3|我要求告当赞美的耶和华， 我必从仇敌手中被救出来。
PS|18|4|死亡的绳索勒住我， 毁灭的急流惊吓我，
PS|18|5|阴间的绳索缠绕我， 死亡的圈套临到我。
PS|18|6|我在急难中求告耶和华， 向我的上帝呼求。 他从殿中听了我的声音， 我在他面前的呼求必进入他耳中。
PS|18|7|那时，因他发怒地就震动战抖， 山的根基也震动挪移。
PS|18|8|他的鼻孔冒烟上腾， 他的口发火焚烧，连煤炭也烧着了。
PS|18|9|他使天垂下，亲自降临， 黑云在他脚下。
PS|18|10|他乘坐基路伯飞行， 藉着风的翅膀快飞，
PS|18|11|以黑暗为藏身之处， 以水的黑暗、天空的密云作四围的行宫。
PS|18|12|因他发出光辉， 冰雹和火炭穿透密云。
PS|18|13|耶和华在天上打雷， 至高者发出声音，就有冰雹和火炭 。
PS|18|14|他射出箭来，使仇敌四散； 发出连串的闪电，击溃他们。
PS|18|15|耶和华啊，你的斥责一发， 你鼻孔的气一出， 海底就显现， 大地的根基也暴露。
PS|18|16|他从高天伸手抓住我， 把我从大水中拉上来。
PS|18|17|他救我脱离强敌和那些恨我的人， 因为他们比我强盛。
PS|18|18|我遭遇灾难的日子，他们来攻击我； 但耶和华是我的倚靠。
PS|18|19|他领我到宽阔之处， 他救拔我，因他喜爱我。
PS|18|20|耶和华必按我的公义报答我， 按我手中的清洁赏赐我。
PS|18|21|因为我遵守耶和华的道， 未曾作恶离开我的上帝。
PS|18|22|他的一切典章常在我面前， 他的律例我也未曾丢弃。
PS|18|23|我在他面前作了完全人， 我也保护自己远离罪孽。
PS|18|24|所以耶和华按我的公义， 在他眼前按我手中的清洁赏赐我。
PS|18|25|慈爱的人，你以慈爱待他； 完全的人，你以完善待他。
PS|18|26|清洁的人，你以清洁待他； 歪曲的人，你以弯曲待他。
PS|18|27|困苦的百姓，你必拯救； 高傲的眼目，你使他降卑。
PS|18|28|你必点亮我的灯； 耶和华－我的上帝必照明我的黑暗。
PS|18|29|我藉着你冲入敌军， 藉着我的上帝跳过城墙。
PS|18|30|至于上帝，他的道是完全的； 耶和华的话是纯净的。 凡投靠他的，他就作他们的盾牌。
PS|18|31|除了耶和华，谁是上帝呢？ 除了我们的上帝，谁是磐石呢？
PS|18|32|惟有那以力量束我的腰、 使我行为完全的，他是上帝。
PS|18|33|他使我的脚快如母鹿， 使我站稳在高处。
PS|18|34|他教导我的手能争战， 我的膀臂能开铜造的弓。
PS|18|35|你赐救恩给我作盾牌， 你的右手扶持我， 你的庇护 使我为大。
PS|18|36|你使我脚步宽阔， 我的脚踝未曾滑跌。
PS|18|37|我要追赶我的仇敌，且要追上他们； 若不将他们灭绝，我总不归回。
PS|18|38|我要打伤他们，使他们站不起来； 他们必倒在我的脚下。
PS|18|39|你曾以力量束我的腰，使我能争战； 也曾使那起来攻击我的，都服在我以下。
PS|18|40|你又使我的仇敌在我面前转身逃跑， 使我剪除那恨我的人。
PS|18|41|他们呼求，却无人拯救； 就是呼求耶和华，他也不应允。
PS|18|42|我捣碎他们，如同风前的灰尘； 倾倒 他们，如同街上的泥土。
PS|18|43|你救我脱离百姓的纷争， 立我作列国的元首； 我素不认识的百姓必事奉我。
PS|18|44|他们一听见我的名声就必顺从我， 外邦人要投降我。
PS|18|45|外邦人要丧胆， 战战兢兢地出营寨。
PS|18|46|耶和华永远活着。 愿我的磐石被称颂， 愿救我的上帝受尊崇。
PS|18|47|这位上帝为我伸冤， 使万民服在我以下。
PS|18|48|他拯救我脱离仇敌， 又把我举起，高过那些起来攻击我的人， 救我脱离残暴的人。
PS|18|49|耶和华啊，因此我要在外邦中称谢你， 歌颂你的名。
PS|18|50|耶和华赐极大的救恩给他所立的王， 施慈爱给他的受膏者， 就是给 大卫 和他的后裔，直到永远。
PS|19|1|诸天述说上帝的荣耀， 穹苍传扬他手的作为。
PS|19|2|这日到那日发出言语， 这夜到那夜传出知识。
PS|19|3|无言无语， 也无声音可听。
PS|19|4|它们的声浪 传遍天下， 它们的言语传到地极。 上帝在其中为太阳安设帐幕，
PS|19|5|太阳如同新郎步出洞房， 又如勇士欢然奔路。
PS|19|6|它从天这边出来，绕到天那边， 没有一物可隐藏得不到它的热气。
PS|19|7|耶和华的律法全备，使人苏醒； 耶和华的法度确定，使愚蒙人有智慧。
PS|19|8|耶和华的训词正直，使人心快活； 耶和华的命令清洁，使人眼目明亮。
PS|19|9|耶和华的典章真实，全然公义， 敬畏耶和华是纯洁的，存到永远，
PS|19|10|比金子可羡慕，比极多的纯金可羡慕； 比蜜甘甜，比蜂房下滴的蜜甘甜。
PS|19|11|因此你的仆人受警戒， 遵守这些有极大的赏赐。
PS|19|12|谁能察觉自己的错失呢？ 求你赦免我隐藏的过犯。
PS|19|13|求你拦阻仆人不犯任意妄为的罪， 不容这罪辖制我， 我就完全，免犯大罪。
PS|19|14|耶和华－我的磐石，我的救赎主啊， 愿我口中的言语，心里的意念在你面前蒙悦纳。
PS|20|1|愿耶和华在你患难的日子应允你， 愿 雅各 的上帝的名保护你。
PS|20|2|愿他从圣所救助你， 从 锡安 坚固你，
PS|20|3|记念你的一切祭物， 悦纳你的燔祭，（细拉）
PS|20|4|将你心所愿的赐给你， 成就你的一切筹算。
PS|20|5|我们要因你的救恩夸胜， 要奉我们上帝的名竖立旌旗。 愿耶和华成就你一切所求的！
PS|20|6|现在我知道耶和华必救护他的受膏者， 从他神圣的天上应允他， 用右手的能力救护他。
PS|20|7|有人靠车，有人靠马， 但我们要提耶和华－我们上帝的名。
PS|20|8|他们都屈身仆倒， 我们却起来，坚立不移。
PS|20|9|耶和华啊，求你拯救； 我们呼求的时候，愿王应允我们！
PS|21|1|耶和华啊，王必因你的能力欢喜； 因你的救恩，他的快乐何其大！
PS|21|2|他心里所愿的，你已经赐给他； 他嘴唇所求的，你未尝不应允。（细拉）
PS|21|3|你以美善的福气迎接他， 把纯金的冠冕戴在他头上。
PS|21|4|他向你祈求长寿，你就赐给他， 就是日子长久，直到永远。
PS|21|5|他因你的救恩大有荣耀， 你将尊荣威严加在他身上。
PS|21|6|你使他有洪福，直到永远， 又使他在你面前欢喜快乐。
PS|21|7|王倚靠耶和华， 因至高者的慈爱，王必不动摇。
PS|21|8|你的手要搜出所有的仇敌， 你的右手要搜出那些恨你的人。
PS|21|9|你的脸出现的时候，要使他们如在炎热的火炉中。 耶和华要在他的震怒中吞灭他们， 那火要把他们烧尽。
PS|21|10|你必从世上灭绝他们的幼苗， 从人间灭绝他们的后裔。
PS|21|11|因为他们有意加害于你； 他们想出计谋，却不能做成。
PS|21|12|你必使他们转身逃跑， 向着他们的脸搭箭在弦。
PS|21|13|耶和华啊，愿你因自己的能力显为至高！ 这样，我们就唱诗，歌颂你的大能。
PS|22|1|我的上帝，我的上帝，为什么离弃我？ 为什么远离不救我，不听我的呻吟？
PS|22|2|我的上帝啊，我白日呼求，你不应允； 夜间呼求，也不得安宁。
PS|22|3|但你是神圣的， 用 以色列 的赞美为宝座。
PS|22|4|我们的祖宗倚靠你； 他们倚靠你，你解救他们。
PS|22|5|他们哀求你，就蒙解救； 他们倚靠你，就不羞愧。
PS|22|6|但我是虫，不是人， 被众人羞辱，被百姓藐视。
PS|22|7|凡看见我的都嗤笑我； 他们撇嘴摇头：
PS|22|8|“他把自己交托给耶和华，让耶和华救他吧！ 耶和华既喜爱他，可以搭救他吧！”
PS|22|9|但你是叫我出母腹的， 我在母怀里，你就使我有倚靠的心。
PS|22|10|我自出母胎就交在你手里， 自我出母腹，你就是我的上帝。
PS|22|11|求你不要远离我！ 因为灾难临头，无人帮助。
PS|22|12|许多公牛环绕我， 巴珊 大力的公牛四面围困我。
PS|22|13|它们向我张口， 好像猎食吼叫的狮子。
PS|22|14|我如水被倒出， 我的骨头都脱了节， 我的心如蜡，在我里面熔化。
PS|22|15|我的精力枯干，如同瓦片， 我的舌头紧贴上颚。 你将我安置在死灰中。
PS|22|16|犬类围着我，恶党环绕我； 他们扎了我的手、我的脚。
PS|22|17|我数遍我的骨头； 他们瞪着眼看我。
PS|22|18|他们分我的外衣， 为我的内衣抽签。
PS|22|19|耶和华啊，求你不要远离我！ 我的救主啊，求你快来帮助我！
PS|22|20|求你救我的性命脱离刀剑， 使我仅有的 脱离犬类，
PS|22|21|求你救我脱离狮子的口； 你已经应允我，使我脱离野牛的角。
PS|22|22|我要将你的名传给我的弟兄， 在会众中我要赞美你。
PS|22|23|敬畏耶和华的人哪，要赞美他！ 雅各 的后裔啊，要荣耀他！ 以色列 的后裔啊，要惧怕他！
PS|22|24|因为他没有藐视、憎恶受苦的人， 也没有转脸不顾他们； 那受苦之人呼求的时候，他就垂听。
PS|22|25|我在大会中赞美你的话是从你而来， 我要在敬畏耶和华的人面前还我的愿。
PS|22|26|愿困苦的人吃得饱足， 愿寻求耶和华的人赞美他。 愿你们的心永远活着！
PS|22|27|地的四极都要想念耶和华，并且归顺他， 列国的万族都要在你面前敬拜。
PS|22|28|因为国度属于耶和华， 他是管理列国的。
PS|22|29|地上富足的人都必吃喝而敬拜， 凡下到尘土中不能存活自己性命的人， 都要在他面前下拜 ；
PS|22|30|必有后裔事奉他， 主所做的事必传给后代。
PS|22|31|他们必来传他的公义给尚未出生的子民， 这是他的作为。
PS|23|1|耶和华是我的牧者， 我必不致缺乏。
PS|23|2|他使我躺卧在青草地上， 领我在可安歇的水边。
PS|23|3|他使我的灵魂苏醒 ， 为自己的名引导我走义路。
PS|23|4|我虽然行过死荫的幽谷， 也不怕遭害， 因为你与我同在； 你的杖、你的竿，都安慰我。
PS|23|5|在我敌人面前，你为我摆设筵席； 你用油膏了我的头，使我的福杯满溢。
PS|23|6|我一生一世必有恩惠慈爱随着我； 我且要住在 耶和华的殿中，直到永远。
PS|24|1|地和其中所充满的， 世界和住在其中的，都属耶和华。
PS|24|2|他把地建立在海上， 安定在江河之上。
PS|24|3|谁能登耶和华的山？ 谁能站在他的圣所？
PS|24|4|就是手洁心清，意念不向虚妄， 起誓不怀诡诈的人。
PS|24|5|他必蒙耶和华赐福， 又蒙救他的上帝使他成义。
PS|24|6|这是寻求耶和华的族类， 是寻求你面的 雅各 。（细拉）
PS|24|7|众城门哪，要抬起头来！ 永久的门户啊，你们要被举起！ 荣耀的王将要进来！
PS|24|8|这荣耀的王是谁呢？ 就是有力有能的耶和华， 在战场上大有能力的耶和华！
PS|24|9|众城门哪，要抬起头来！ 永久的门户啊，你们要高举！ 荣耀的王将要进来！
PS|24|10|这荣耀的王是谁呢？ 万军之耶和华是荣耀的王！（细拉）
PS|25|1|耶和华啊，我的心仰望你。
PS|25|2|我的上帝啊，我素来倚靠你； 求你不要叫我羞愧， 不要叫我的仇敌向我夸胜。
PS|25|3|凡等候你的必不羞愧， 惟有那无故行奸诈的必要羞愧。
PS|25|4|耶和华啊，求你将你的道指示我， 将你的路指教我！
PS|25|5|求你指教我，引导我进入你的真理， 因为你是救我的上帝。 我整日等候你。
PS|25|6|耶和华啊，求你记念你的怜悯和慈爱， 因为这是亘古以来所常有的。
PS|25|7|求你不要记得我幼年的罪愆和我的过犯； 耶和华啊，求你因你的良善，按你的慈爱记念我。
PS|25|8|耶和华是良善正直的， 因此，他必教导罪人走正路。
PS|25|9|他要按公平引领谦卑人， 将他的道指教他们。
PS|25|10|凡遵守他的约和他法度的人， 耶和华都以慈爱信实待他。
PS|25|11|耶和华啊，求你因你名的缘故赦免我的罪， 因我的罪重大。
PS|25|12|谁敬畏耶和华， 耶和华必教导他当选择的道路。
PS|25|13|他要安然居住， 他的后裔必承受土地。
PS|25|14|耶和华与敬畏他的人亲密， 他要将自己的约指示他们。
PS|25|15|我的眼目时常仰望耶和华， 因他必将我的脚从网里拉出来。
PS|25|16|求你转向我，怜悯我， 因我孤独困苦。
PS|25|17|我心里愁苦甚多， 求你救我脱离我的祸患。
PS|25|18|求你看顾我的困苦、我的艰难， 赦免我一切的罪。
PS|25|19|求你察看我的仇敌， 因为他们人数众多，并且痛恨我。
PS|25|20|求你保护我的性命，搭救我， 使我不致羞愧，因为我投靠你。
PS|25|21|愿纯全、正直保护我， 因为我等候你。
PS|25|22|上帝啊，求你救赎 以色列 脱离他一切的愁苦。
PS|26|1|耶和华啊，求你为我伸冤， 因我向来行事纯正； 我倚靠耶和华，必不动摇。
PS|26|2|耶和华啊，求你察看我，考验我， 熬炼我的肺腑心肠。
PS|26|3|因为你的慈爱常在我眼前， 我也按你的真理而行。
PS|26|4|我未曾与虚妄的人同坐， 也不与伪善的人来往。
PS|26|5|我痛恨恶人的集会， 必不与恶人同坐。
PS|26|6|耶和华啊，我要洗手表明无辜， 才环绕你的祭坛；
PS|26|7|我好发出称谢的声音， 述说你一切奇妙的作为。
PS|26|8|耶和华啊，我喜爱你所住的殿 和你显荣耀的居所。
PS|26|9|不要把我的性命和罪人一同除掉， 不要把我的生命和好流人血的一同除掉。
PS|26|10|他们的手中有奸恶， 他们的右手满有贿赂。
PS|26|11|至于我，却要行事纯正； 求你救赎我，怜悯我！
PS|26|12|我的脚站在平坦的地方， 在聚会中我要称颂耶和华！
PS|27|1|耶和华是我的亮光，是我的拯救， 我还怕谁呢？ 耶和华是我生命的保障， 我还惧谁呢？
PS|27|2|那作恶的就是我的仇敌， 前来吃我肉的时候就绊跌仆倒。
PS|27|3|虽有军队安营攻击我，我的心也不害怕； 虽然兴起战争攻击我，我仍旧安稳。
PS|27|4|有一件事，我曾求耶和华，我仍要寻求， 就是一生一世住在耶和华的殿中， 瞻仰他的荣美，在他的殿宇里求问。
PS|27|5|因为我遭遇患难，他必将我隐藏在他的帐棚里， 把我藏在他帐幕的隐密处， 将我高举在磐石上。
PS|27|6|现在我得以昂首，高过四面的仇敌。 我要在他的帐幕里欢然献祭， 我要唱诗歌颂耶和华。
PS|27|7|耶和华啊，我呼求的时候，求你垂听我的声音； 求你怜悯我，应允我。
PS|27|8|你说：“你们当寻求我的面。” 那时我的心向你说： “耶和华啊，你的面我正要寻求。”
PS|27|9|求你不要转脸不顾我， 不要发怒赶逐你的仆人， 你向来是帮助我的。 救我的上帝啊，不要离开我， 也不要撇弃我。
PS|27|10|即使我的父母撇弃我， 耶和华终必收留我。
PS|27|11|耶和华啊，求你将你的道指教我， 因我仇敌的缘故引导我走平坦的路。
PS|27|12|求你不要把我交给敌人，遂其所愿； 因为妄作见证的和口吐凶言的都起来攻击我。
PS|27|13|我深信在活人之地 必得见耶和华的恩惠。
PS|27|14|要等候耶和华， 当壮胆，坚固你的心， 要等候耶和华！
PS|28|1|耶和华啊，我要求告你！ 我的磐石啊，求你不要向我缄默！ 倘若你向我闭口， 我就如下入地府的人一样。
PS|28|2|我呼求你，向你至圣所举手的时候， 求你垂听我恳求的声音！
PS|28|3|不要把我和坏人并作恶的一同除掉； 他们跟邻舍说平安，心里却是奸恶。
PS|28|4|求你按着他们所做的， 按他们的恶行对待他们； 求你照着他们手所做的对待他们， 将他们应得的报应加给他们。
PS|28|5|他们既然不尊重耶和华的作为， 也不尊重他手所做的， 耶和华就必毁坏他们，不建立他们。
PS|28|6|耶和华是应当称颂的， 因为他听了我恳求的声音。
PS|28|7|耶和华是我的力量，是我的盾牌， 我心里倚靠他就得帮助。 我心中欢乐， 我要用诗歌称谢他。
PS|28|8|耶和华是他百姓的力量， 又是他受膏者得救的保障。
PS|28|9|求你拯救你的百姓，赐福给你的产业； 求你牧养他们，扶持他们，直到永远。
PS|29|1|上帝的子民 哪，你们要将荣耀、能力归给耶和华， 都归给耶和华！
PS|29|2|要将耶和华的名的荣耀归给他， 要敬拜神圣荣耀的耶和华 。
PS|29|3|耶和华的声音在众水上， 荣耀的上帝打雷； 耶和华打雷在大水之上。
PS|29|4|耶和华的声音大有能力， 耶和华的声音满有威严。
PS|29|5|耶和华的声音震碎香柏树， 耶和华震碎 黎巴嫩 的香柏树。
PS|29|6|他使 黎巴嫩 跳跃如牛犊， 使 西连 跳跃如野牛犊。
PS|29|7|耶和华的声音使火焰分岔。
PS|29|8|耶和华的声音震动旷野， 耶和华震动 加低斯 的旷野。
PS|29|9|耶和华的声音惊动母鹿落胎， 树林也脱落净光。 凡在他殿中的，都述说他的荣耀。
PS|29|10|耶和华坐在洪水之上为王； 耶和华坐着为王，直到永远。
PS|29|11|耶和华必赐力量给他的百姓， 耶和华必赐平安的福给他的百姓。
PS|30|1|耶和华啊，我要尊崇你， 因为你救了我，不让仇敌向我夸耀。
PS|30|2|耶和华－我的上帝啊， 我呼求你，你医治了我。
PS|30|3|耶和华啊，你救我的性命脱离阴间， 使我存活，不至于下入地府。
PS|30|4|耶和华的圣民哪，你们要歌颂他， 要颂扬他神圣的名字 。
PS|30|5|因为，他的怒气不过是转眼之间； 他的恩典乃是一生之久。 一宿虽然有哭泣， 早晨便必欢呼。
PS|30|6|至于我，我凡事顺利，就说： “我永不动摇。”
PS|30|7|耶和华啊，你曾施恩，使我稳固如山； 你转脸不顾，我就惊惶。
PS|30|8|耶和华啊，我曾求告你； 我向耶和华恳求：
PS|30|9|“我被害流血，下到地府，有何益处呢？ 尘土岂能称谢你、传扬你的信实吗？
PS|30|10|耶和华啊，求你应允我，怜悯我！ 耶和华啊，求你帮助我！”
PS|30|11|你将我的哀哭变为跳舞， 脱去我的麻衣，为我披上喜乐，
PS|30|12|使我的灵 歌颂你，不致缄默。 耶和华－我的上帝啊，我要称谢你，直到永远！
PS|31|1|耶和华啊，我投靠你， 求你使我永不羞愧， 凭你的公义搭救我！
PS|31|2|求你侧耳听我， 快快救我！ 求你作我坚固的磐石， 拯救我的保障！
PS|31|3|你真是我的岩石、我的山寨， 求你为你名的缘故引导我，指教我。
PS|31|4|求你救我脱离人为我暗设的网罗， 因为你是我的保障。
PS|31|5|我将我的灵交在你手里； 耶和华─信实的上帝啊，你救赎了我。
PS|31|6|我 恨恶那信奉虚无神明 的人； 我却倚靠耶和华。
PS|31|7|我要因你的慈爱欢喜快乐， 因为你见过我的困苦， 知道我心中的艰难。
PS|31|8|你未曾把我交在仇敌手里， 你使我的脚站在宽阔的地方。
PS|31|9|耶和华啊，求你怜悯我， 因为我在急难之中； 我的眼睛因忧愁而昏花， 我的身心也已耗尽。
PS|31|10|我的生命为愁苦所消耗， 我的年岁为叹息所荒废； 我的力量因我的罪孽 衰败， 我的骨头也枯干。
PS|31|11|我因所有的敌人成了羞辱， 在我邻舍跟前更加羞辱； 那认识我的都惧怕我， 在街上看见我的都躲避我。
PS|31|12|我被遗忘，如同死人，无人记念； 我好像破碎的器皿。
PS|31|13|我听见许多人的毁谤， 四围尽是惊吓； 他们一同商议攻击我， 图谋害我的性命。
PS|31|14|耶和华啊，我仍要倚靠你； 我说：“你是我的上帝。”
PS|31|15|我终生的事在你手中， 求你救我脱离仇敌的手和那些迫害我的人。
PS|31|16|求你使你的脸向仆人发光， 凭你的慈爱拯救我。
PS|31|17|耶和华啊，求你叫我不致羞愧， 因为我曾呼求你； 求你使恶人羞愧， 使他们在阴间缄默无声。
PS|31|18|那撒谎的人逞骄傲轻慢， 出狂妄的话攻击义人， 愿他的嘴哑而无言。
PS|31|19|在世人眼前， 你为敬畏你的人所积存的， 为投靠你的人所施行的， 是何等大的恩惠啊！
PS|31|20|你必将他们藏在你面前的隐密处， 免得遭人暗算； 你要隐藏他们在棚子里， 免受口舌的争闹。
PS|31|21|耶和华是应当称颂的， 因为我在围城里，他向我施展奇妙的慈爱。
PS|31|22|至于我，我曾惊惶地说： “我从你眼前被隔绝。” 然而，我呼求你的时候， 你仍听我恳求的声音。
PS|31|23|耶和华的圣民哪，你们都要爱他！ 耶和华保护诚实可靠的人， 却加倍报应行事骄傲的人。
PS|31|24|凡仰望耶和华的人， 你们都要壮胆，坚固你们的心！
PS|32|1|过犯得赦免， 罪恶蒙遮盖的人有福了！
PS|32|2|耶和华不算为有罪， 内心没有诡诈的人有福了！
PS|32|3|我闭口不认罪的时候， 因终日呻吟而骨头枯干。
PS|32|4|黑夜白日，你的手压在我身上沉重； 我的精力耗尽 ，如同夏天的干旱。（细拉）
PS|32|5|我向你陈明我的罪， 不隐瞒我的恶。 我说：“我要向耶和华承认我的过犯”； 你就赦免我的罪恶。（细拉）
PS|32|6|为此，凡虔诚人都当趁你可寻找 的时候向你祷告； 大水泛滥的时候，必不临到他。
PS|32|7|你是我藏身之处， 你必保佑我脱离苦难， 以得救的欢呼 四面环绕我。（细拉）
PS|32|8|我要教导你，指示你当行的路， 我要定睛在你身上劝戒你。
PS|32|9|你不可像那无知的骡马， 须用嚼环缰绳勒住， 不然，它就不会靠近你。
PS|32|10|恶人必多受苦楚； 惟独倚靠耶和华的，必有慈爱四面环绕他。
PS|32|11|义人哪，你们应当靠耶和华欢喜快乐， 心里正直的人哪，你们都当欢呼。
PS|33|1|义人哪，你们当因耶和华欢呼， 正直人理当赞美耶和华。
PS|33|2|你们要弹琴称谢耶和华， 用十弦瑟歌颂他。
PS|33|3|应当向他唱新歌， 弹得巧妙，声音洪亮。
PS|33|4|因为耶和华的言语正直， 他的作为尽都信实。
PS|33|5|他喜爱公义和公平， 遍地满了耶和华的慈爱。
PS|33|6|诸天藉耶和华的话而造， 万象藉他口中的气而成。
PS|33|7|他聚集海水如垒， 收藏深洋在仓库。
PS|33|8|愿全地都敬畏耶和华！ 愿世上的居民都惧怕他！
PS|33|9|因为他说有，就有， 命立，就立。
PS|33|10|耶和华使列国的筹算归于无有， 使万民的计谋全无功效。
PS|33|11|耶和华的筹算永远立定， 他心中的计划万代长存。
PS|33|12|以耶和华为上帝的，那国有福了！ 耶和华拣选为自己产业的，那民有福了！
PS|33|13|耶和华从天上观看， 看见所有的人，
PS|33|14|从他的居所察看地上每一个居民，
PS|33|15|他塑造他们的心， 洞察他们一切的作为。
PS|33|16|君王不能因兵多得胜， 勇士不能因力大得救。
PS|33|17|靠马得救是枉然的， 马也不能因力大救人。
PS|33|18|看哪，耶和华的眼目看顾敬畏他的人 和仰望他慈爱的人，
PS|33|19|要救他们的性命脱离死亡， 使他们在饥荒中存活。
PS|33|20|我们的心向来等候耶和华； 他是我们的帮助，是我们的盾牌。
PS|33|21|我们的心必靠他欢喜， 因为我们向来倚靠他的圣名。
PS|33|22|耶和华啊，求你照着我们所仰望你的， 向我们施行慈爱！
PS|34|1|我要时时称颂耶和华， 赞美他的话常在我口中。
PS|34|2|我的心必因耶和华夸耀， 谦卑的人听见就喜乐。
PS|34|3|你们要和我一同尊耶和华为大， 让我们一同高举他的名。
PS|34|4|我曾寻求耶和华，他就应允我， 救我脱离一切的恐惧。
PS|34|5|仰望他的人，就有光荣； 他们 的脸必不蒙羞。
PS|34|6|这困苦人呼求，耶和华就垂听， 救他脱离一切的患难。
PS|34|7|耶和华的使者在敬畏他的人四围安营， 要搭救他们。
PS|34|8|你们要尝尝主恩的滋味，便知道他是美善； 投靠他的人有福了！
PS|34|9|耶和华的圣民哪，你们当敬畏他， 因敬畏他的一无所缺。
PS|34|10|少壮狮子尚且缺食忍饿， 但寻求耶和华的什么好处都不缺。
PS|34|11|孩子们哪，来听我！ 我要将敬畏耶和华的道教导你们。
PS|34|12|有谁喜爱生命， 爱慕长寿，得享美福？
PS|34|13|你要禁止舌头不出恶言， 嘴唇不说诡诈的话。
PS|34|14|要弃恶行善， 寻求和睦，一心追求。
PS|34|15|耶和华的眼目看顾义人， 他的耳朵听他们的呼求。
PS|34|16|耶和华向行恶的人变脸， 要从地上除灭他们的名字 。
PS|34|17|义人呼求，耶和华听见了， 就拯救他们脱离一切患难。
PS|34|18|耶和华靠近伤心的人， 拯救心灵痛悔的人。
PS|34|19|义人多有苦难， 但耶和华救他脱离这一切，
PS|34|20|又保护他全身的骨头， 连一根也不折断。
PS|34|21|恶必害死恶人， 恨恶义人的，必被定罪。
PS|34|22|耶和华救赎他仆人的性命， 凡投靠他的，必不致定罪。
PS|35|1|耶和华啊，与我相争的，求你与他们相争！ 与我争战的，求你与他们争战！
PS|35|2|求你拿着大小盾牌， 起来帮助我；
PS|35|3|举起枪来，抵挡那追赶我的。 求你对我说：“我是拯救你的。”
PS|35|4|愿那寻索我命的，蒙羞受辱！ 愿那谋害我的，退后羞愧！
PS|35|5|愿他们像风前的糠秕， 有耶和华的使者赶逐他们。
PS|35|6|愿他们的道路又暗又滑， 有耶和华的使者追赶他们。
PS|35|7|因他们无故为我暗设网罗， 无故挖坑，要害我的命。
PS|35|8|愿灾祸忽然临到他身上！ 愿他暗设的网罗缠住自己！ 愿他落在其中遭灾祸！
PS|35|9|我的心必靠耶和华快乐， 靠他的救恩欢喜。
PS|35|10|我全身的骨头要说： “耶和华啊，谁能像你 救护困苦人脱离那比他强壮的， 救护困苦贫穷人脱离那抢夺他的？”
PS|35|11|凶恶的见证人起来， 盘问我所不知道的事。
PS|35|12|他们向我以恶报善， 使我丧失儿子。
PS|35|13|至于我，他们有病的时候， 我穿麻衣，禁食，刻苦己心； 我所求的都归到自己身上。
PS|35|14|我如此行，好像他是我的朋友，我的兄弟； 我屈身悲哀，如同哀悼自己的母亲。
PS|35|15|我在患难中，他们却欢喜，大家聚集， 我所不认识的卑贱人 聚集攻击我， 他们不住地撕裂我。
PS|35|16|他们试探我，不断嘲笑我 ， 向我咬牙切齿。
PS|35|17|主啊，你看着不理要到几时呢？ 求你救我的性命脱离他们的残害， 救我仅有的 脱离少壮狮子！
PS|35|18|我在大会中要称谢你， 在许多百姓中要赞美你。
PS|35|19|求你不容那无理与我为仇的向我夸耀！ 不容那无故恨我的向我瞪眼！
PS|35|20|因为他们不说平安， 倒想出诡诈的言语扰害地上安静的人。
PS|35|21|他们大大张口攻击我，说： “啊哈，啊哈，我们已经亲眼看见了！”
PS|35|22|耶和华啊，你已经看见了，求你不要沉默！ 主啊，求你不要远离我！
PS|35|23|我的上帝─我的主啊，求你醒来，求你奋起， 还我公正，伸明我冤！
PS|35|24|耶和华－我的上帝啊，求你按你的公义判断我， 不容他们向我夸耀！
PS|35|25|不容他们心里说：“啊哈，遂我们的心愿了！” 不容他们说：“我们已经把他吞了！”
PS|35|26|愿那喜欢我遭难的一同抱愧蒙羞！ 愿那向我妄自尊大的披戴惭愧，蒙受羞辱！
PS|35|27|愿那喜悦我被判为义 的欢呼快乐； 愿他们常说：“当尊耶和华为大！ 耶和华喜悦他的仆人平安。”
PS|35|28|我的舌头要论说你的公义， 要常常赞美你。
PS|36|1|过犯在恶人的心底向他说话 ， 他的眼中不怕上帝。
PS|36|2|他自夸自媚， 以致罪孽无法察觉，不被恨恶。
PS|36|3|他口中的言语尽是罪孽诡诈， 他不再有智慧，也不再行善。
PS|36|4|他在床上图谋罪孽， 定意行不善的道，不憎恶恶事。
PS|36|5|耶和华啊，你的慈爱上及诸天， 你的信实达到穹苍，
PS|36|6|你的公义好像高山， 你的判断如同深渊； 耶和华啊，人民、牲畜，你都救护。
PS|36|7|上帝啊，你的慈爱何其宝贵！ 世人投靠在你翅膀的荫下。
PS|36|8|他们必因你殿里的丰盛得以饱足， 你也必叫他们喝你那喜乐的泉水。
PS|36|9|因为在你那里有生命的泉源， 在你的光中，我们必得见光。
PS|36|10|愿你常施慈爱给认识你的人， 常以公义待心里正直的人。
PS|36|11|不容骄傲人的脚践踏我， 不容凶恶人的手赶逐我。
PS|36|12|在那里，作恶的人已经仆倒； 他们被推倒，不能再起来。
PS|37|1|不要为作恶的心怀不平， 也不要嫉妒那行不义的人。
PS|37|2|因为他们如草快被割下， 又如绿色的嫩草快要枯干。
PS|37|3|你当倚靠耶和华而行善， 安居地上，以他的信实为粮；
PS|37|4|又当以耶和华为乐， 他就将你心里所求的赐给你。
PS|37|5|当将你的道路交托耶和华， 并倚靠他，他就必成全。
PS|37|6|他要使你的公义如光发出， 使你的公平明如正午。
PS|37|7|你当安心倚靠耶和华，耐性等候他， 不要因那道路通达的和那恶谋成就的心怀不平。
PS|37|8|当止住怒气，离弃愤怒； 不要心怀不平，以致作恶。
PS|37|9|因为作恶的必被剪除； 惟有等候耶和华的必承受土地。
PS|37|10|还有片时，恶人要归于无有； 你就是细察他的住处，也不存在。
PS|37|11|但谦卑的人必承受土地， 以丰盛的平安为乐。
PS|37|12|恶人设谋要害义人， 向他咬牙。
PS|37|13|但主必笑他， 因见他受罚的日子将要来到。
PS|37|14|恶人刀已出鞘，弓已上弦， 要砍倒困苦贫穷的人， 要杀害行为正直的人。
PS|37|15|他们的刀必刺入自己的心， 他们的弓必折断。
PS|37|16|一个义人所有的虽少， 强过许多恶人的富余。
PS|37|17|因为恶人的膀臂必折断； 但耶和华扶持义人。
PS|37|18|耶和华知道完全人的日子， 他们的产业要存到永远。
PS|37|19|他们在患难的时候必不致羞愧， 在饥荒的日子必得饱足。
PS|37|20|恶人却要灭亡。 耶和华的仇敌要像草地的华美 ； 他们要毁灭，在烟中消失 。
PS|37|21|恶人借贷却不偿还； 义人恩待人，并且施舍。
PS|37|22|蒙耶和华赐福的必承受土地； 他所诅咒的必被剪除。
PS|37|23|义人的脚步为耶和华所稳定； 他的道路，耶和华也喜爱。
PS|37|24|他虽失脚也不致全身仆倒， 因为耶和华搀扶他的手。
PS|37|25|我从前年幼，现在年老， 却未见过义人被弃， 也未见过他的后裔求乞。
PS|37|26|他常常恩待人，借贷给人， 他的后裔也必蒙福。
PS|37|27|你当离恶行善， 就可永远安居。
PS|37|28|因为耶和华喜爱公平， 不撇弃他的圣民， 他们永蒙保佑； 但恶人的后裔必被剪除。
PS|37|29|义人必承受土地， 永居其上。
PS|37|30|义人的口发出智慧， 他的舌头讲说公平。
PS|37|31|上帝的律法在他心里， 他的步伐总不摇动。
PS|37|32|恶人窥探义人， 想要杀他。
PS|37|33|耶和华必不把他交在恶人手中， 当审判的时候，也不定他的罪。
PS|37|34|你当等候耶和华，遵守他的道， 他就抬举你，使你承受土地； 你必看到恶人被剪除。
PS|37|35|我见过恶人大有势力， 高耸如本地青翠的树木。
PS|37|36|有人 从那里经过，看哪，他已不存在， 我寻找他，却寻不着了。
PS|37|37|你要细察那完全人，观看那正直人， 因为和平的人有好结局。
PS|37|38|至于罪人，必一同灭绝， 恶人的结局必被剪除。
PS|37|39|义人得救是出于耶和华， 在患难时耶和华作他们的避难所。
PS|37|40|耶和华帮助他们，解救他们； 他解救他们脱离恶人，把他们救出来， 因为他们投靠他。
PS|38|1|耶和华啊，求你不要在怒中责备我， 不要在烈怒中惩罚我！
PS|38|2|因为你的箭射入我身， 你的手压住我。
PS|38|3|因你的恼怒，我的肉无一完全； 因我的罪过，我的骨头也不安宁。
PS|38|4|我的罪孽高过我的头， 如同重担叫我担当不起。
PS|38|5|因我的愚昧， 我的伤发臭流脓。
PS|38|6|我疼痛，大大蜷曲， 整日哀痛。
PS|38|7|我满腰灼热， 我的肉无一完全。
PS|38|8|我被压碎，身心虚弱； 因心里痛苦，我就呻吟。
PS|38|9|主啊，我的心愿都在你面前， 我的叹息不向你隐瞒。
PS|38|10|我心颤栗，体力衰微， 眼中无光。
PS|38|11|我遭遇灾病，良朋密友都袖手旁观， 我的亲戚本家也远远站立。
PS|38|12|那寻索我命的设下罗网， 那想要害我的口出恶言， 整日思想诡计。
PS|38|13|但我如聋子听不见， 像哑巴不能开口。
PS|38|14|我如听不见的人， 无法用口答辩。
PS|38|15|耶和华啊，我仰望你！ 主－我的上帝啊，你必应允我！
PS|38|16|我曾说：“恐怕他们向我夸耀， 我失脚的时候，他们向我夸口。”
PS|38|17|我就要跌倒， 我的痛苦常在我面前。
PS|38|18|我要承认我的罪孽， 要因我的罪忧愁。
PS|38|19|但我的仇敌又活泼又强壮， 无理恨我的增多了。
PS|38|20|以恶报善的与我作对， 但我追求良善。
PS|38|21|耶和华啊，求你不要撇弃我！ 我的上帝啊，求你不要远离我！
PS|38|22|拯救我的主啊， 求你快快帮助我！
PS|39|1|我曾说：“我要谨慎我的言行， 免得我的舌头犯罪； 恶人在我面前的时候， 我要用嚼环勒住我的口。”
PS|39|2|我默然无声，连好话也不出口， 我的愁苦就更加深。
PS|39|3|我的心在我里面发热； 我默想的时候，火就烧起， 我用舌头说话：
PS|39|4|“耶和华啊，求你让我晓得我的结局， 我的寿数几何， 使我知道我的生命何等短暂！
PS|39|5|看哪，你使我的年日窄如手掌， 我一生的年数，在你面前如同无有； 各人最稳妥的时候，真是全然虚幻。（细拉）
PS|39|6|世人行动实系幻影， 他们忙乱，真是枉然， 积蓄财宝，不知将来有谁收取。
PS|39|7|“主啊，如今我等什么呢？ 我的指望在乎你！
PS|39|8|求你救我脱离一切的过犯， 不要使我受愚顽人的羞辱。
PS|39|9|我保持沉默，闭口不言， 因为这一切都是你所做的。
PS|39|10|求你从我身上免去你的责罚； 因你手的责打，我就消灭。
PS|39|11|因人的罪恶你惩罚管教他的时候， 如蛀虫一般，吃掉他所喜爱的。 世人真是虚幻！（细拉）
PS|39|12|“耶和华啊，求你听我的祷告， 侧耳听我的呼求！ 我流泪，求你不要静默无声！ 因为在你面前我是客旅， 是寄居的，像我列祖一般。
PS|39|13|求你宽容我， 使我在去而不返之先可以喜乐。”
PS|40|1|我曾耐性等候耶和华， 他垂听我的呼求。
PS|40|2|他从泥坑里， 从淤泥中，把我拉上来， 使我的脚立在磐石上， 使我脚步稳健。
PS|40|3|他使我口唱新歌， 就是赞美我们上帝的话。 许多人必看见而惧怕， 并要倚靠耶和华。
PS|40|4|那倚靠耶和华、 不理会狂傲和偏向虚假的， 这人有福了！
PS|40|5|耶和华－我的上帝啊，你所行的奇事 和你为我们设想的计划，多到无法尽述； 若要述说陈明，不可胜数。
PS|40|6|祭物和礼物，你不喜爱， 你已经开通我的耳朵； 燔祭和赎罪祭非你所要。
PS|40|7|那时我说：“看哪，我来了！ 我的事在经卷上已经记载了。
PS|40|8|我的上帝啊，我乐意照你的旨意行， 你的律法在我心里。”
PS|40|9|我在大会中传讲公义的佳音， 看哪，必不制止我的嘴唇； 耶和华啊，这一切你都知道。
PS|40|10|我未曾把你的公义藏在心里， 我已陈明你的信实和你的救恩； 在大会中我未曾隐瞒你的慈爱和信实。
PS|40|11|耶和华啊，求你不要向我止住你的怜悯！ 愿你的慈爱和信实常常保佑我！
PS|40|12|因有无数的祸患围困我， 我的罪孽追上了我，使我不能看见， 这罪孽比我的头发还多， 我的胆量丧失了。
PS|40|13|耶和华啊，求你开恩搭救我！ 耶和华啊，求你速速帮助我！
PS|40|14|愿那些寻找我、要灭我命的，一同抱愧蒙羞！ 愿那些喜悦我遭害的，退后受辱！
PS|40|15|愿那些对我说“啊哈、啊哈”的， 因羞愧而败亡！
PS|40|16|愿一切寻求你的，因你欢喜快乐！ 愿那些喜爱你救恩的，常说：“当尊耶和华为大！”
PS|40|17|我本是困苦贫穷的，主却顾念我。 你是帮助我的，搭救我的； 我的上帝啊，求你不要耽延！
PS|41|1|眷顾贫寒人的有福了 ！ 在患难的日子，耶和华必搭救他。
PS|41|2|耶和华必保全他，使他存活， 他要在地上享福。 求你不要把他交给仇敌，遂其所愿。
PS|41|3|他病重在榻，耶和华必扶持他； 他在病中，你必使他离开病床。
PS|41|4|我曾说：“耶和华啊，求你怜悯我， 医治我，因为我得罪了你。”
PS|41|5|我的仇敌用恶言议论我： “他几时才会死，他的名几时才会消灭呢？”
PS|41|6|当他来看我的时候，说的是假话； 他心存奸恶，走到外边才说出来。
PS|41|7|所有恨我的，都一同交头接耳议论我， 他们设计要害我。
PS|41|8|他们说：“他有怪病缠身， 他已躺下，必不能再起来。”
PS|41|9|连我知己的朋友， 我所信赖、吃我饭的人也用脚踢我。
PS|41|10|耶和华啊，求你怜悯我， 使我起来，好报复他们！
PS|41|11|我因此就知道你喜爱我， 我的仇敌不得向我夸胜。
PS|41|12|你因我纯正就扶持我， 使我永远站立在你面前。
PS|41|13|耶和华－ 以色列 的上帝是应当称颂的， 从亘古直到永远。阿们！阿们！ 可拉后裔的诗。交给圣咏团长。
PS|42|1|上帝啊，我的心切慕你， 如鹿切慕溪水。
PS|42|2|我的心渴想上帝，就是永生上帝， 我几时得朝见上帝呢？
PS|42|3|我昼夜以眼泪当食物， 人不住地对我说：“你的上帝在哪里呢？”
PS|42|4|我从前与众人同往， 领他们到上帝的殿里， 大家用欢呼称颂的声音守节； 我追想这些事， 我的心极其悲伤。
PS|42|5|我的心哪，你为何忧闷？ 为何在我里面烦躁？ 应当仰望上帝， 因我还要称谢他，我当面的拯救，
PS|42|6|我的上帝。我的心在我里面忧闷， 所以我从 约旦 地， 从 黑门岭 ，从 米萨山 记念你。
PS|42|7|你的瀑布发声，深渊就与深渊响应， 你的波浪洪涛漫过我身。
PS|42|8|白昼，耶和华必施慈爱； 黑夜，我要歌颂祈祷赐我生命的上帝。
PS|42|9|我要对上帝－我的磐石说： “你为何忘记我呢？ 我为何因仇敌的欺压时常哀痛呢？”
PS|42|10|我的敌人辱骂我， 好像敲碎我的骨头， 他们不住地对我说： “你的上帝在哪里呢？”
PS|42|11|我的心哪，你为何忧闷？ 为何在我里面烦躁？ 应当仰望上帝， 因我还要称谢他，我当面的拯救，我的上帝。
PS|43|1|上帝啊，求你为我伸冤， 向不虔诚的国为我辩护； 求你救我脱离诡诈不义的人。
PS|43|2|你是作我保障 的上帝，为何丢弃我呢？ 我为何因仇敌的欺压时常哀痛呢？
PS|43|3|求你发出你的亮光和信实，好引导我， 带我到你的圣山，到你的居所！
PS|43|4|我就走到上帝的祭坛， 到赐我喜乐的上帝那里。 上帝，我的上帝啊， 我要弹琴称谢你！
PS|43|5|我的心哪，你为何忧闷？ 为何在我里面烦躁？ 应当仰望上帝， 我还要称谢他，我当面的拯救，我的上帝。
PS|44|1|上帝啊，你在古时， 我们列祖的日子所做的事， 我们亲耳听见了， 我们的列祖曾为我们述说。
PS|44|2|你曾用手赶出外邦人， 却栽培了我们的列祖； 你苦待万民， 却叫我们的列祖发达。
PS|44|3|因为他们不是靠自己的刀剑承受土地， 也不是靠自己的膀臂得胜， 而是靠你的右手、你的膀臂， 和你脸上的亮光， 因为你喜爱他们。
PS|44|4|上帝啊，你是我的君王， 求你发命令使 雅各 得胜。
PS|44|5|靠你，我们要推倒我们的敌人； 靠你的名，我们要践踏那兴起攻击我们的人。
PS|44|6|因为我必不倚靠我的弓， 我的刀也不能使我得胜。
PS|44|7|惟有你拯救我们脱离敌人， 使恨我们的人羞愧。
PS|44|8|我们要常常因上帝夸耀， 要永远颂扬你的名。（细拉）
PS|44|9|但如今你丢弃了我们，使我们受辱， 不和我们的军队同去。
PS|44|10|你使我们在敌人前转身撤退， 使那恨我们的人任意抢夺。
PS|44|11|你使我们如羊当作食物， 把我们分散在列国中。
PS|44|12|你卖了你的子民也不获利， 所得的并未加添你的资财。
PS|44|13|你使我们受邻国的羞辱， 被四围的人嗤笑讥讽。
PS|44|14|你使我们在列国中成了笑柄， 在万民中使人摇头。
PS|44|15|因辱骂者和毁谤者的声音， 因仇敌和报仇者的缘故， 我的凌辱常常在我面前， 我脸上的羞愧将我遮蔽，
PS|44|16|
PS|44|17|这些事都临到我们身上， 我们却没有忘记你， 也没有违背你的约；
PS|44|18|我们的心并未退缩， 我们的脚也没有偏离你的路。
PS|44|19|你在野狗出没之处压伤我们， 以死荫笼罩我们。
PS|44|20|倘若我们忘记上帝的名， 或向外邦神明举手，
PS|44|21|上帝岂不鉴察这事吗？ 因为他晓得人心里的隐秘。
PS|44|22|我们为你的缘故终日被杀， 人看我们如将宰的羊。
PS|44|23|主啊，求你睡醒，为何尽睡呢？ 求你醒来，不要永远丢弃我们！
PS|44|24|你为何转脸， 不顾我们所遭的苦难和所受的欺压呢？
PS|44|25|我们俯伏在尘土上， 我们的肚腹紧贴地面。
PS|44|26|求你兴起帮助我们！ 因你的慈爱救赎我们！
PS|45|1|我心里涌出美辞， 我为王朗诵我的诗章， 我的舌头是敏捷文士的手笔。
PS|45|2|你比世人更美， 你嘴里满有恩惠； 所以上帝赐福给你，直到永远。
PS|45|3|勇士啊，愿你腰间佩刀， 大展荣耀和威严，
PS|45|4|为真理、谦卑、公义威严地驾车前进，无不得胜； 愿你的右手显明可畏的事。
PS|45|5|你的箭锋快，射中王的仇敌的心， 万民仆倒在你之下。
PS|45|6|上帝啊，你的宝座是永永远远的， 你国度的权杖是正直的权杖。
PS|45|7|你喜爱公义，恨恶罪恶， 所以上帝，就是你的上帝，用喜乐油膏你， 胜过膏你的同伴。
PS|45|8|你的衣服散发没药、沉香、肉桂的香气， 象牙宫中丝弦乐器的声音使你欢喜。
PS|45|9|你的妃嫔之中有列王的女儿， 王后佩戴 俄斐 金饰站立在你右边。
PS|45|10|女子啊，要倾听，要思想，要侧耳而听！ 不要记念你本族和你父家，
PS|45|11|王就羡慕你的美貌； 因为他是你的主，你当向他下拜。
PS|45|12|推罗 必来送礼， 百姓中富足的人也必向你求恩。
PS|45|13|君王的女儿在宫里极其荣华， 她的衣服是金线绣的；
PS|45|14|她穿锦绣的衣服，引到王面前， 陪伴她的童女随从她，也被带到你面前。
PS|45|15|她们要欢喜快乐， 被引导进入王宫。
PS|45|16|你的子孙要接续你列祖， 你要立他们在各地作王。
PS|45|17|我必使万代记念你的名， 万民要永永远远称谢你。
PS|46|1|上帝是我们的避难所，是我们的力量， 是我们在患难中随时的帮助。
PS|46|2|所以，地虽改变， 山虽摇动到海心，
PS|46|3|其中的水虽澎湃翻腾， 山虽因海涨而战抖， 我们也不害怕。（细拉）
PS|46|4|有一道河，这河的分汊使上帝的城欢喜， 这城就是至高者居住的圣所。
PS|46|5|上帝在其中，城必不动摇； 到天一亮，上帝必帮助这城。
PS|46|6|万邦喧嚷，国度动摇； 上帝出声，地就熔化。
PS|46|7|万军之耶和华与我们同在， 雅各 的上帝是我们的避难所！（细拉）
PS|46|8|你们来看耶和华的作为， 看他使地怎样荒凉。
PS|46|9|他止息战争，直到地极； 他折弓、断枪，把战车焚烧在火中。
PS|46|10|你们要休息，要知道我是上帝！ 我必在列国中受尊崇，在全地也受尊崇。
PS|46|11|万军之耶和华与我们同在， 雅各 的上帝是我们的避难所！
PS|47|1|万民哪，你们都要鼓掌！ 用欢呼的声音向上帝呼喊！
PS|47|2|因为耶和华至高者是可畏的， 他是治理全地的大君王。
PS|47|3|他使万民服在我们以下， 又使万族服在我们脚下。
PS|47|4|他为我们选择产业， 就是他所爱之 雅各 的荣耀。（细拉）
PS|47|5|上帝上升，有喊声相送； 耶和华上升，有角声相送。
PS|47|6|你们要向上帝歌颂，歌颂！ 向我们的王歌颂，歌颂！
PS|47|7|因为上帝是全地的王， 你们要用圣诗歌颂！
PS|47|8|上帝作王治理列国， 上帝坐在他的圣宝座上。
PS|47|9|万民的君王聚集， 要作 亚伯拉罕 的上帝的子民， 因为地上的盾牌是属上帝的， 他为至高！
PS|48|1|耶和华本为大！ 在我们上帝的城中， 在他的圣山上， 当受大赞美。
PS|48|2|锡安山 －大君王的城， 在北面居高华美， 为全地所喜悦。
PS|48|3|上帝在城的宫殿中， 自显为避难所。
PS|48|4|看哪，诸王会合， 一同经过。
PS|48|5|他们见了这城就惊奇丧胆， 急忙逃跑。
PS|48|6|战兢在那里抓住他们， 他们好像临产的妇人一样阵痛。
PS|48|7|上帝啊，你用东风击破 他施 的船只。
PS|48|8|我们在万军之耶和华的城里， 就是我们上帝的城里， 所看见的正如我们所听见的。 上帝必坚立这城，直到永远。（细拉）
PS|48|9|上帝啊，我们在你的殿中 想念你的慈爱。
PS|48|10|上帝啊，你受的赞美正与你的名相称，直到地极！ 你的右手满了公义。
PS|48|11|因你的判断， 锡安山 应当欢喜， 犹大 的城镇 应当快乐。
PS|48|12|你们当周游 锡安 ， 四围环绕，数点城楼，
PS|48|13|细看它的城郭， 察看它的宫殿， 为要传扬给后代。
PS|48|14|因为这上帝永永远远为我们的上帝， 他必作我们引路的，直到死时 。
PS|49|1|万民哪，你们都当听这话！ 世上所有的居民， 无论贵贱贫富， 都当侧耳而听！
PS|49|2|
PS|49|3|我口要说智慧的言语， 我心思想通达的道理。
PS|49|4|我要侧耳听比喻， 用琴解谜语。
PS|49|5|在患难的日子，追逼我的人的奸恶 环绕我， 我何必惧怕？
PS|49|6|他们那些倚靠财货， 自夸钱财多的人，
PS|49|7|没有一个能赎自己的弟兄 ， 能将赎价给上帝，
PS|49|8|让他长远活着，不见地府 ； 因为赎生命的价值极贵， 只可永远罢休。
PS|49|9|
PS|49|10|他要见智慧人死， 愚昧人和畜牲一般的人一同灭亡， 把他们的财货留给别人。
PS|49|11|他们虽以自己的名叫自己的地， 坟墓却作他们永远的家， 作他们世世代代的居所。
PS|49|12|人居尊贵中不能长久， 如同死亡的畜类一样。
PS|49|13|他们所行之道本为自己的愚昧， 后来的人却还佩服他们的话语。（细拉）
PS|49|14|他们如同羊群注定要下阴间， 死亡必作他们的牧者； 到了早晨，正直人必管辖他们。 他们的形像必被阴间所灭，无处可容身。
PS|49|15|然而上帝必救赎我的命脱离阴间的掌控， 因他必收纳我。（细拉）
PS|49|16|见人发财、家室日益显赫的时候， 你不要惧怕；
PS|49|17|因为他死的时候什么也不能带去， 他的荣耀不能随他下去。
PS|49|18|他活着的时候，虽然自夸为有福 ─你若自己行得好，人必夸奖你─
PS|49|19|他仍必与历代的祖宗一样同归死亡， 永不见光。
PS|49|20|人在尊贵中而不醒悟， 就如死亡的畜类一样。
PS|50|1|大能者上帝－耶和华已经发言呼召天下， 从日出之地到日落之处。
PS|50|2|从全然美丽的 锡安 中， 上帝已经发光了。
PS|50|3|我们的上帝要来，绝不闭口； 有烈火在他面前吞灭， 有暴风在他四围刮起。
PS|50|4|他呼召上天下地， 为要审判他的子民：
PS|50|5|“召集我的圣民， 就是那些用祭物与我立约的人，到我这里来。”
PS|50|6|诸天必表明他的公义， 因为上帝是施行审判的。（细拉）
PS|50|7|“听啊，我的子民，我要说话！ 以色列 啊，我要审问你； 我是上帝，是你的上帝！
PS|50|8|我并不因你的祭物责备你； 你的燔祭常在我面前。
PS|50|9|我不从你家中取公牛， 也不从你圈内取公山羊；
PS|50|10|因为，林中的百兽是我的， 千山的牲畜也是我的。
PS|50|11|山中 的飞鸟，我都知道， 田野的走兽也都属我。
PS|50|12|“我若是饥饿，不用告诉你， 因为世界和其中所充满的都是我的。
PS|50|13|我岂吃公牛的肉呢？ 我岂喝公山羊的血呢？
PS|50|14|你们要以感谢为祭献给上帝， 又要向至高者还你的愿，
PS|50|15|并要在患难之日求告我， 我必搭救你，你也要荣耀我。”
PS|50|16|但上帝对恶人说：“你怎敢传讲我的律例， 口中提到我的约呢？
PS|50|17|其实你恨恶管教， 将我的言语抛在脑后。
PS|50|18|你见了盗贼就乐意与他同伙， 又和行奸淫的人同流合污。
PS|50|19|“你的口出恶言， 你的舌编造诡诈。
PS|50|20|你坐着，毁谤你的兄弟， 谗害你亲母的儿子。
PS|50|21|你做了这些事，我闭口不言， 你想我正如你一样； 其实我要责备你，将这些事摆在你眼前。
PS|50|22|“你们忘记上帝的，要思想这事， 免得我把你们撕碎，无人搭救。
PS|50|23|凡以感谢献祭的就是荣耀我； 那按正路而行的，我必使他得着上帝的救恩。”
PS|51|1|上帝啊，求你按你的慈爱恩待我！ 按你丰盛的怜悯涂去我的过犯！
PS|51|2|求你将我的罪孽洗涤净尽， 洁除我的罪！
PS|51|3|因为我知道我的过犯； 我的罪常在我面前。
PS|51|4|我向你犯罪，惟独得罪了你， 在你眼前行了这恶， 以致你责备的时候显为公义， 判断的时候显为清白。
PS|51|5|看哪，我是在罪孽里生的， 在我母亲怀胎的时候就有了罪。
PS|51|6|你所喜爱的是内心的诚实； 求你在我隐密处使我得智慧。
PS|51|7|求你用牛膝草洁净我，我就干净； 求你洗涤我，我就比雪更白。
PS|51|8|求你使我得听欢喜快乐的声音， 使你所压伤的骨头可以踊跃。
PS|51|9|求你转脸不看我的罪， 涂去我一切的罪孽。
PS|51|10|上帝啊，求你为我造清洁的心， 使我里面重新有正直 的灵。
PS|51|11|不要丢弃我，使我离开你的面； 不要从我收回你的圣灵。
PS|51|12|求你使我重得救恩之乐， 以乐意的灵来扶持我，
PS|51|13|我就把你的道指教有过犯的人， 罪人必归顺你。
PS|51|14|上帝啊，你是拯救我的上帝； 求你救我脱离流人血的罪！ 我的舌头就高唱你的公义。
PS|51|15|主啊，求你使我嘴唇张开， 我的口就传扬赞美你的话！
PS|51|16|你本不喜爱祭物，若喜爱，我就献上； 燔祭你也不喜悦。
PS|51|17|上帝所要的祭就是忧伤的灵； 上帝啊，忧伤痛悔的心，你必不轻看。
PS|51|18|求你随你的美意善待 锡安 ， 建造 耶路撒冷 的城墙。
PS|51|19|那时，你必喜爱公义的祭 和燔祭，全牲的燔祭； 那时，人必将公牛献在你坛上。
PS|52|1|勇士啊，你为何作恶自夸？ 上帝的慈爱是常存的。
PS|52|2|你这行诡诈的人哪， 你的舌头像快利的剃刀，图谋毁灭。
PS|52|3|你爱恶胜似爱善， 又爱说谎，胜于爱说公义。（细拉）
PS|52|4|诡诈的舌头啊， 你爱说一切毁灭的话！
PS|52|5|上帝也要毁灭你，直到永远。 他要抓住你，从帐棚中拉你出来， 从活人之地将你拔除。（细拉）
PS|52|6|义人要看见而惧怕， 并要笑他。
PS|52|7|看哪，这就是那不以上帝为保障的人， 他只倚靠丰富的财物，在邪恶上坚立自己。
PS|52|8|至于我，就像上帝殿中的青橄榄树， 我永永远远倚靠上帝的慈爱。
PS|52|9|我要称谢你，直到永远， 因为你做了这事。 我也要在你圣民面前仰望你的名， 这名本为美好。
PS|53|1|愚顽人心里说：“没有上帝。” 他们都败坏，行了可憎恶的罪孽， 没有一个人行善。
PS|53|2|上帝从天上垂看世人， 要看有明白的没有， 有寻求上帝的没有。
PS|53|3|他们全都退后，一同变为污秽， 没有行善的， 连一个也没有。
PS|53|4|作恶的都没有知识吗？ 他们吞吃我的百姓如同吃饭一样， 并不求告上帝。
PS|53|5|他们在无可惧怕之处就大大害怕， 因为上帝使那安营攻击你之人的骨头散开了。 你使他们蒙羞，因为上帝弃绝了他们。
PS|53|6|但愿 以色列 的救恩出自 锡安 。 当上帝救回他被掳子民的时候， 雅各 要快乐， 以色列 要欢喜。
PS|54|1|上帝啊，求你因你的名拯救我， 凭你的大能为我伸冤。
PS|54|2|上帝啊，求你听我的祷告， 侧耳听我口中的言语。
PS|54|3|因为陌生人兴起攻击我， 强横的人寻索我的性命； 他们眼中没有上帝。（细拉）
PS|54|4|看哪，上帝是帮助我的， 主是扶持我性命的，
PS|54|5|他要报应我仇敌所作的恶； 求你凭你的信实灭绝他们。
PS|54|6|我要把甘心祭献给你； 耶和华啊，我要颂扬你的名，这名本为美好。
PS|54|7|他从一切的急难中把我救出来， 我的眼睛也看见了我的仇敌遭报。
PS|55|1|上帝啊，求你侧耳听我的祷告， 不要隐藏不听我的恳求！
PS|55|2|求你留心听我，应允我。 我哀叹不安，发出呻吟，
PS|55|3|都因仇敌的声音，恶人的欺压； 他们将罪孽加在我身上，发怒气加害我。
PS|55|4|我的心在我里面阵痛， 死亡的恐怖落在我身。
PS|55|5|恐惧战兢临到了我， 惊恐笼罩我。
PS|55|6|我说：“但愿我有翅膀像鸽子， 我就飞去，得享安息。
PS|55|7|看哪，我要远走高飞， 宿在旷野。（细拉）
PS|55|8|我要速速逃到避难之所， 脱离狂风暴雨。”
PS|55|9|主啊，求你吞灭他们，变乱他们的言语！ 因为我在城中见了凶暴争吵的事。
PS|55|10|他们昼夜在城墙上绕行， 城内也有罪孽和奸恶。
PS|55|11|邪恶在其中， 欺压和诡诈不离街市。
PS|55|12|原来，不是仇敌辱骂我， 若是仇敌，还可忍受； 也不是恨我的人向我狂妄自大， 若是恨我的人，我必躲避他。
PS|55|13|不料是你；你原与我同等， 是我的朋友，是我的知己！
PS|55|14|我们素常彼此交谈，以为甘甜； 我们结伴在上帝的殿中同行。
PS|55|15|愿死亡忽然临到他们！ 愿他们活生生地下入阴间！ 因为他们的住处都是邪恶， 他们的内心充满奸恶。
PS|55|16|至于我，我要求告上帝， 耶和华必拯救我。
PS|55|17|晚上、早晨、中午我要哀声悲叹， 他就垂听我的声音。
PS|55|18|他救赎我的命脱离攻击我的人， 使我得享平安， 因为与我相争的人很多。
PS|55|19|那不愿改变、不敬畏上帝的人， 从太古常存的上帝必听见而使他受苦。（细拉）
PS|55|20|他背了约， 伸手攻击与他和好的人。
PS|55|21|他的口如奶油光滑， 他的心却怀着敌意； 他的话比油柔和， 其实是拔出的刀。
PS|55|22|你要把你的重担卸给耶和华， 他必扶持你， 他永不叫义人动摇。
PS|55|23|上帝啊，你必使恶人坠入灭亡的坑； 那好流人血、行诡诈的人必活不过半生， 但我要倚靠你。
PS|56|1|上帝啊，求你怜悯我，因为有人践踏我， 终日攻击欺压我。
PS|56|2|我的仇敌终日践踏我， 逞骄傲攻击我的人很多。
PS|56|3|我惧怕的时候要倚靠你。
PS|56|4|我倚靠上帝，我要赞美他的话语； 我倚靠上帝，必不惧怕。 血肉之躯能把我怎么样呢？
PS|56|5|他们终日扭曲我的话， 千方百计加害于我。
PS|56|6|他们聚集，埋伏，窥探我的脚踪， 等候要害我的命。
PS|56|7|他们岂能脱罪呢 ？ 上帝啊，求你在怒中使万民败落！
PS|56|8|我几次流离，你都数算； 求你把我的眼泪装在你的皮袋里。 这一切不都记在你的册子上吗？
PS|56|9|我呼求的日子，仇敌都要转身撤退。 上帝帮助我，这是我所知道的。
PS|56|10|我倚靠上帝，我要赞美他的话语； 我倚靠耶和华，我要赞美他的话语。
PS|56|11|我倚靠上帝，必不惧怕。 人能把我怎么样呢？
PS|56|12|上帝啊，我要向你还所许的愿， 我要以感谢祭回报你；
PS|56|13|因为你救我的命脱离死亡。 你保护我的脚不跌倒， 使我在生命的光中行在上帝面前。
PS|57|1|上帝啊，求你怜悯我，怜悯我， 因为我的心投靠你。 我要投靠在你翅膀荫下， 直等到灾害过去。
PS|57|2|我要求告至高的上帝， 就是为我成全万事的上帝。
PS|57|3|那践踏我的人辱骂我的时候， 上帝必从天上施恩救我，(细拉) 他必向我施行慈爱和信实。
PS|57|4|至于我的性命， 我好像躺卧在吞噬人的狮子当中； 他们的牙齿是枪、箭， 他们的舌头是快刀。
PS|57|5|上帝啊，愿你崇高过于诸天！ 愿你的荣耀高过全地！
PS|57|6|他们为我的脚设下网罗，压迫我； 他们在我面前掘了坑，自己反掉在其中。（细拉）
PS|57|7|上帝啊，我心坚定，我心坚定； 我要唱诗，我要歌颂！
PS|57|8|我的灵 啊，你当醒起！ 琴瑟啊，当醒起！ 我自己要极早醒起！
PS|57|9|主啊，我要在万民中称谢你， 在万族中歌颂你！
PS|57|10|因为你的慈爱高及诸天， 你的信实达到穹苍。
PS|57|11|上帝啊，愿你崇高过于诸天！ 愿你的荣耀高过全地！
PS|58|1|你们缄默不语，真合公义吗？ 你们审判世人，岂按正直吗？
PS|58|2|不然！你们心中作恶， 量出你们在地上手中的残暴。
PS|58|3|恶人一出母胎就与上帝疏远， 一离母腹就走错路，说谎话。
PS|58|4|他们的毒气好像蛇的毒气， 他们好像聋的毒蛇塞住耳朵，
PS|58|5|听不见弄蛇者的声音， 也听不见魔术师的咒语。
PS|58|6|上帝啊，求你敲碎他们口中的牙！ 耶和华啊，求你敲掉少壮狮子的大牙！
PS|58|7|愿他们消灭，如急流的水一般； 他们瞄准射箭的时候，箭头仿佛折断。
PS|58|8|愿他们像蜗牛腐烂消失， 又像妇人流掉的胎儿，未见天日。
PS|58|9|你们用荆棘烧火，锅还未热， 上帝就用旋风把未烧着的和已烧着的一齐刮去。
PS|58|10|义人见仇敌遭报就欢喜， 他要在恶人的血中洗脚。
PS|58|11|因此，人必说：“义人诚然有善报， 在地上果然有施行审判的上帝！”
PS|59|1|我的上帝啊，求你救我脱离仇敌， 把我安置在高处，脱离那些起来攻击我的人。
PS|59|2|求你救我脱离作恶的人， 救我脱离好流人血的人！
PS|59|3|因为他们埋伏要害我命， 强悍的人聚集攻击我， 耶和华啊，不是为我的过犯， 也不是为我的罪愆。
PS|59|4|我虽然无过，他们急忙摆阵攻击我。 求你兴起，来帮助我，来鉴察！
PS|59|5|万军之耶和华上帝－ 以色列 的上帝啊， 求你醒起，惩治万国！ 不要怜悯行诡诈的恶人！（细拉）
PS|59|6|他们晚上转回， 叫号如狗，围城绕行。
PS|59|7|看哪，他们口中喷吐恶言， 嘴里有刀： “有谁听见呢？”
PS|59|8|但你－耶和华必讥笑他们， 你要嗤笑万国。
PS|59|9|我 的力量啊，我要等候你， 因为上帝是我的庇护所。
PS|59|10|我的上帝要以慈爱 迎接我， 上帝要叫我看见我的仇敌遭报。
PS|59|11|主，我们的盾牌啊， 不要杀他们，免得我的子民遗忘； 求你用你的能力使他们四散， 使他们降为卑。
PS|59|12|愿他们因口中的罪和嘴唇的言语， 被自己的骄傲抓住， 他们所说的尽是咒骂和谎话。
PS|59|13|求你发怒，使他们消灭， 求你使他们消灭，归于无有， 使他们知道上帝在 雅各 中间掌权， 直到地极。（细拉）
PS|59|14|他们晚上转回， 叫号如狗，围城绕行。
PS|59|15|他们到处走动觅食， 若不饱足就咆哮不已。
PS|59|16|但我要歌颂你的能力， 早晨要高唱你的慈爱； 因为你是我的庇护所， 在急难的日子作过我的避难所。
PS|59|17|我的力量啊，我要歌颂你； 因为上帝是我的庇护所， 是赐恩给我的上帝。
PS|60|1|上帝啊，你丢弃了我们，破坏了我们； 你曾发怒，求你使我们复兴！
PS|60|2|你使地震动，崩裂； 求你将裂口补好，因为地在摇动。
PS|60|3|你让你的子民遇见艰难， 使我们喝那令人东倒西歪的酒。
PS|60|4|你把旌旗赐给敬畏你的人， 可以躲避弓箭 。（细拉）
PS|60|5|求你应允我们 ，用右手施行拯救， 好让你所亲爱的人得救。
PS|60|6|上帝在他的圣所 说： “我要欢乐； 要划分 示剑 ， 丈量 疏割谷 。
PS|60|7|基列 是我的， 玛拿西 是我的。 以法莲 是护卫我头的， 犹大 是我的权杖。
PS|60|8|摩押 是我的沐浴盆， 我要向 以东 扔鞋。 非利士 啊，你还能因我欢呼吗？”
PS|60|9|谁能领我进坚固城？ 谁能引我到 以东 地？
PS|60|10|上帝啊，你真的丢弃了我们吗？ 上帝啊，你不和我们的军队同去吗？
PS|60|11|求你帮助我们攻击敌人， 因为人的帮助是枉然的。
PS|60|12|我们倚靠上帝才得施展大能， 因为践踏我们敌人的就是他。
PS|61|1|上帝啊，求你听我的呼求， 留心听我的祷告！
PS|61|2|我心里发昏的时候， 要从地极求告你。 求你领我到那比我更高的磐石，
PS|61|3|因为你是我的避难所， 是我的坚固台，使我脱离仇敌。
PS|61|4|我要永远住在你的帐幕里！ 我要投靠在你翅膀下的隐密处！（细拉）
PS|61|5|上帝啊，你听了我所许的愿； 你将产业赐给敬畏你名的人。
PS|61|6|求你加添王的寿数， 使他的年岁存到世世代代。
PS|61|7|愿他在上帝面前永远坐在王位上， 求你预备慈爱和信实保佑他！
PS|61|8|这样，我要歌颂你的名，直到永远， 天天还我所许的愿。
PS|62|1|我的心默默无声，专等候上帝， 我的救恩从他而来。
PS|62|2|惟独他是我的磐石，我的拯救； 他是我的庇护所，我必不大大动摇。
PS|62|3|你们大家攻击一人，使他被杀， 如歪斜的墙、将倒的壁，要到几时呢？
PS|62|4|他们彼此商议，要把他从高位上拉下来； 他们喜爱谎话，口虽祝福，心却诅咒。（细拉）
PS|62|5|我的心哪，你当默默无声，专等候上帝， 因为我的盼望是从他而来。
PS|62|6|惟独他是我的磐石，我的拯救； 他是我的庇护所，我必不动摇。
PS|62|7|我的拯救、我的荣耀都在于上帝； 我力量的磐石、我的避难所都在于上帝。
PS|62|8|百姓啊，要时时倚靠他， 在他面前倾心吐意； 上帝是我们的避难所。（细拉）
PS|62|9|人真是虚空， 人真是虚假； 放在天平里就必浮起， 他们一共比空气还轻。
PS|62|10|不要仗势欺人， 也不要因抢夺而骄傲； 若财宝加增，不要放在心上。
PS|62|11|上帝说了一次、两次，我都听见了， 就是能力属乎上帝。
PS|62|12|主啊，慈爱也是属乎你， 因为你照着各人所做的报应他。
PS|63|1|上帝啊，你是我的上帝， 我要切切寻求你； 在干旱疲乏无水之地， 我的心灵渴想你，我的肉身切慕你。
PS|63|2|我在圣所中曾如此瞻仰你， 为要见你的能力和你的荣耀。
PS|63|3|因你的慈爱比生命更好， 我的嘴唇要颂赞你。
PS|63|4|我还活着的时候要这样称颂你， 我要奉你的名举手。
PS|63|5|我在床上记念你， 在夜更的时候思念你； 我的心像吃饱了骨髓肥油， 我也要以欢乐的嘴唇赞美你。
PS|63|6|
PS|63|7|因为你曾帮助了我， 我要在你翅膀的荫下欢呼。
PS|63|8|我的心紧紧跟随你； 你的右手扶持了我。
PS|63|9|但那些寻索要灭我命的人 必往地底下去；
PS|63|10|他们必被刀剑所杀， 成为野狗的食物。
PS|63|11|但是王必因上帝欢喜， 凡指着他发誓的都要夸耀， 因为说谎之人的口必被塞住。
PS|64|1|上帝啊，我哀叹的时候，求你听我的声音！ 求你保护我的性命，不受仇敌的惊吓！
PS|64|2|求你把我隐藏， 使我脱离作恶之人的暗谋， 脱离作孽之人的扰乱。
PS|64|3|他们磨舌如刀， 发出苦毒的言语，好像瞄准了的箭，
PS|64|4|要在暗地里射完全人； 他们忽然射他，并不惧怕。
PS|64|5|他们彼此勉励，设下恶计； 他们商量，暗设圈套， 说：“谁能看见呢？”
PS|64|6|他们图谋奸恶： “我们完成了精密的策划。” 各人的意念心思是深沉的。
PS|64|7|但上帝要用箭射他们， 他们忽然受了伤。
PS|64|8|他们必然绊跌，被自己的舌头所害； 凡看见他们的都必摇头。
PS|64|9|众人都要害怕， 要传扬上帝的工作， 并且明白他的作为。
PS|64|10|义人必因耶和华欢喜，并要投靠他； 凡心里正直的人都必夸耀。
PS|65|1|上帝啊，在 锡安 ，人都等候赞美你， 也要向你还所许的愿。
PS|65|2|听祷告的主啊， 凡有血肉之躯的都要来就你。
PS|65|3|罪孽胜了我； 至于我们的过犯，你都要赦免。
PS|65|4|你所拣选、使他亲近你、住在你院中的， 这人有福了！ 我们要因你居所、你圣殿的美福知足。
PS|65|5|拯救我们的上帝啊，你必以威严秉公义应允我们； 地极和海角远方的人都倚靠你。
PS|65|6|你既以大能束腰， 就用力量安定诸山，
PS|65|7|使诸海的响声和其中波浪的响声， 并万民的喧哗，都平静了。
PS|65|8|住在地极的人因你的神迹惧怕， 你使日出日落之地都欢呼。
PS|65|9|你眷顾地， 降雨使地大大肥沃。 上帝的河满了水； 你这样浇灌了地， 好为人预备五谷。
PS|65|10|你浇透地的犁沟，润泽犁脊， 降甘霖，使地松软； 其中生长的，蒙你赐福。
PS|65|11|你以恩惠为年岁的冠冕， 你的路径都滴下油脂，
PS|65|12|滴在旷野的草场上。 小山以欢乐束腰，
PS|65|13|草场以羊群为衣， 谷中也长满了五谷； 这一切都欢呼歌唱。
PS|66|1|全地都当向上帝欢呼！
PS|66|2|当歌颂他名的荣耀， 使赞美他的话大有荣耀！
PS|66|3|当对上帝说：“你的作为何等可畏！ 因你的大能，仇敌要向你投降。
PS|66|4|全地要敬拜你，歌颂你， 要歌颂你的名。”（细拉）
PS|66|5|你们来看上帝所做的， 他向世人所做之事是可畏的。
PS|66|6|他将海变成干地，使百姓步行过河； 我们在那里要因他欢喜。
PS|66|7|他用权能治理，直到永远。 他的眼睛鉴察万民； 悖逆的人不可自高。（细拉）
PS|66|8|万民哪，你们当称颂我们的上帝， 使人得听赞美他的声音。
PS|66|9|他使我们的性命存活， 不叫我们的脚摇动。
PS|66|10|上帝啊，你曾考验我们， 你熬炼我们，如炼银子一样。
PS|66|11|你使我们进入罗网， 把重担放在我们身上。
PS|66|12|你使人坐车轧我们的头； 我们经过水火， 你却使我们到丰富之地。
PS|66|13|我要带着燔祭进你的殿， 向你还我的愿，
PS|66|14|就是在急难时我嘴唇所发的、 口中所许的。
PS|66|15|我要将肥牛的燔祭 和公羊的香祭献给你， 又要把公牛和公山羊献上。（细拉）
PS|66|16|敬畏上帝的人哪，你们都来听！ 我要述说他为我所做的事。
PS|66|17|我曾用口求告他， 我的舌头也称他为高。
PS|66|18|我若心里注重罪孽， 主必不听。
PS|66|19|但上帝实在听见了， 他留心听了我祷告的声音。
PS|66|20|上帝是应当称颂的！ 他没有推却我的祷告， 也没有使他的慈爱离开我。
PS|67|1|愿上帝怜悯我们，赐福给我们， 使他的脸向我们发光，（细拉）
PS|67|2|好让全地得知你的道路， 万国得知你的救恩。
PS|67|3|上帝啊，愿万民称谢你！ 愿万民都称谢你！
PS|67|4|愿万族都快乐欢呼； 因为你必按公正审判万民， 引导地上的万族。（细拉）
PS|67|5|上帝啊，愿万民称谢你！ 愿万民都称谢你！
PS|67|6|地已经出了土产， 上帝，我们的上帝，要赐福给我们。
PS|67|7|上帝要赐福给我们， 地的四极都要敬畏他！
PS|68|1|愿上帝兴起，使他的仇敌四散， 使那恨他的人从他面前逃跑。
PS|68|2|你驱逐他们 ，如烟被吹散； 恶人见上帝的面就消灭，如蜡被火熔化。
PS|68|3|惟有义人必然欢喜， 在上帝面前快乐， 他们要在喜乐中欢欣。
PS|68|4|你们当向上帝唱诗，歌颂他的名； 为那驾车经过旷野的修平道路 。 他的名是耶和华， 你们要在他面前欢乐！
PS|68|5|上帝在他的圣所作孤儿的父， 作寡妇的伸冤者。
PS|68|6|上帝使孤独的有家， 使被囚的出来享福； 惟有悖逆的要住在干旱之地。
PS|68|7|上帝啊，当你走在百姓前头， 在旷野行进，（细拉）
PS|68|8|地见上帝的面就震动，天也降雨； 西奈山 见 以色列 上帝的面也震动。
PS|68|9|上帝啊，你降下大雨； 你的产业 以色列 疲乏的时候，你使他坚固。
PS|68|10|你的会众住在境内； 上帝啊，你在恩惠中为困苦人预备所需的。
PS|68|11|主发命令， 传好信息的妇女成了大群：
PS|68|12|“统领大军的君王逃跑了，逃跑了！” 在家等候的妇女也分得了掠物。
PS|68|13|你们躺卧在羊圈， 好像鸽子的翅膀镀银，翎毛镀金一般。
PS|68|14|全能者在境内赶散列王的时候， 势如飘雪在 撒们 。
PS|68|15|巴珊山 是极其宏伟 的山， 巴珊山 是多峰多岭的山。
PS|68|16|你们多峰多岭的山哪， 为何以妒忌的眼光看上帝所愿居住的山？ 耶和华必住这山，直到永远！
PS|68|17|上帝的车辇累万盈千； 主在其中，好像在 西奈 圣山一样。
PS|68|18|你已经升上高天，掳掠了俘虏； 你在人间，就是在悖逆的人中，受了供献， 使耶和华上帝可以与他们同住。
PS|68|19|天天背负我们重担的主， 就是拯救我们的上帝， 是应当称颂的！（细拉）
PS|68|20|上帝是为我们施行拯救的上帝； 人能脱离死亡是在乎主─耶和华。
PS|68|21|但上帝要打破他仇敌的头， 就是那常犯罪之人的头颅。
PS|68|22|主说：“我要使百姓从 巴珊 归来， 使他们从深海转回，
PS|68|23|好叫你打碎仇敌，使你的脚踹在血中， 使你狗的舌头也有份。”
PS|68|24|上帝啊，你是我的上帝，我的王； 人已经看见你行走，进入圣所。
PS|68|25|歌唱的行在前，作乐的随在后， 都在击鼓的童女中间：
PS|68|26|“从 以色列 源头而来的啊， 你们当在各会中称颂上帝─耶和华！”
PS|68|27|在那里，有统管他们的小 便雅悯 ， 有 犹大 的领袖和他们的一群人， 有 西布伦 的领袖， 有 拿弗他利 的领袖。
PS|68|28|你的上帝已赐给你力量 ； 上帝啊，求你坚固你为我们所成全的事！
PS|68|29|因你 耶路撒冷 的殿， 列王必带贡物献给你。
PS|68|30|求你斥责芦苇中的野兽和公牛群， 并万民中的牛犊。 直到他们带着银块来朝贡 ； 上帝已经赶散好战的万民 。
PS|68|31|埃及 的使臣要出来， 古实 人要急忙向上帝伸出手来。
PS|68|32|地上的国度啊， 你们要向上帝歌唱， 要歌颂主，（细拉）
PS|68|33|就是那驾行在亘古的诸天之上的主！ 听啊，他发出声音，是极大的声音。
PS|68|34|你们要将能力归给上帝； 他的威荣在 以色列 之上， 他的能力显在天上。
PS|68|35|上帝啊，你从圣所显为可畏， 以色列 的上帝是那将力量权能赐给他百姓的。 上帝是应当称颂的！
PS|69|1|上帝啊，求你救我！ 因为众水就要淹没我。
PS|69|2|我深陷在淤泥中，没有立脚之地； 我到了深水之中，波涛漫过我身。
PS|69|3|我因呼求困乏，喉咙发干； 我因等候上帝，眼睛失明。
PS|69|4|无故恨我的，比我的头发还多； 无理与我为仇、要把我剪除的，甚为强盛。 我没有抢夺，他们竟然要我偿还！
PS|69|5|上帝啊，我的愚昧，你原知道， 我的罪愆不能向你隐瞒。
PS|69|6|万军之主耶和华啊， 求你不要让那等候你的因我蒙羞！ 以色列 的上帝啊， 求你不要让那寻求你的因我受辱！
PS|69|7|因我为你的缘故受了辱骂， 满面羞愧。
PS|69|8|我的兄弟把我当陌生人， 我母亲的儿子把我当外邦人。
PS|69|9|因我为你的殿心里焦急，如同火烧， 并且辱骂你的人的辱骂都落在我身上。
PS|69|10|我哭泣，以禁食刻苦我心； 这倒成了我的羞辱。
PS|69|11|我拿麻布当衣裳， 却成了他们的笑柄。
PS|69|12|坐在城门口的谈论我， 酒徒也以我为歌曲。
PS|69|13|至于我，耶和华啊，在悦纳的时候我向你祈祷。 上帝啊，求你按你丰盛的慈爱， 凭你拯救的信实应允我！
PS|69|14|求你搭救我脱离淤泥， 不叫我陷在其中； 求你使我脱离那些恨我的人， 使我脱离深水。
PS|69|15|求你不容波涛漫过我， 不容深渊吞灭我， 不容深坑在我以上合口。
PS|69|16|耶和华啊，求你应允我！ 因为你的慈爱本为美好； 求你按你丰盛的怜悯转回眷顾我！
PS|69|17|不要转脸不顾你的仆人； 我在急难之中，求你速速应允我！
PS|69|18|求你亲近我，救赎我！ 求你因我仇敌的缘故将我赎回！
PS|69|19|你知道我所受的辱骂、欺凌、羞辱； 我的敌人都在你面前。
PS|69|20|辱骂刺伤我的心， 使我忧愁。 我指望有人体恤，却没有一个； 指望有人安慰，却找不着一个。
PS|69|21|他们拿苦胆给我当食物； 我渴了，他们拿醋给我喝。
PS|69|22|愿他们的筵席在他们面前变为罗网， 在他们平安的时候 变为圈套。
PS|69|23|愿他们的眼睛昏花，看不见； 求你使他们的腰常常战抖。
PS|69|24|求你将你的恼恨倒在他们身上， 使你的烈怒追上他们。
PS|69|25|愿他们的住处变为废墟， 他们的帐棚无人居住。
PS|69|26|因为你所击打的，他们就迫害； 你所击伤的，他们述说 他的愁苦。
PS|69|27|求你使他们罪上加罪， 不容他们在你面前称义。
PS|69|28|愿他们从生命册上被涂去， 不得名列在义人之中。
PS|69|29|但我困苦忧伤； 上帝啊，愿你的救恩将我安置在高处。
PS|69|30|我要以诗歌赞美上帝的名， 以感谢尊他为大！
PS|69|31|这就让耶和华喜悦，胜似献牛， 献有角有蹄的公牛。
PS|69|32|谦卑的人看见了就喜乐； 寻求上帝的人，愿你们的心苏醒。
PS|69|33|因为耶和华听了穷乏的人， 不藐视被囚的人。
PS|69|34|愿天和地、 海洋和其中一切的动物都赞美他！
PS|69|35|因为上帝要拯救 锡安 ，建造 犹大 的城镇； 他的子民要在那里居住，得地为业。
PS|69|36|他仆人的后裔要承受这地， 爱他名的人要住在其中。
PS|70|1|上帝啊，求你快快搭救我！ 耶和华啊，求你速速帮助我！
PS|70|2|愿那些寻索我命的，抱愧蒙羞； 愿那些喜悦我遭害的，退后受辱。
PS|70|3|愿那些对我说“啊哈、啊哈”的， 因羞愧退后。
PS|70|4|愿所有寻求你的，因你欢喜快乐； 愿那些喜爱你救恩的，常说：“当尊上帝为大！”
PS|70|5|但我是困苦贫穷的； 上帝啊，求你速速到我这里来！ 你是帮助我的，搭救我的； 耶和华啊，求你不要耽延！
PS|71|1|耶和华啊，我投靠你， 求你叫我永不羞愧！
PS|71|2|求你凭你的公义搭救我，救拔我； 侧耳听我，拯救我！
PS|71|3|求你作我常来栖身 的磐石， 你已经吩咐要救我， 因为你是我的岩石、我的山寨。
PS|71|4|我的上帝啊，求你救我脱离恶人的手， 脱离不义和残暴之人的手。
PS|71|5|主耶和华啊，你是我所盼望的； 自我年幼，你是我所倚靠的。
PS|71|6|我自出母胎被你扶持， 使我出母腹的是你。 我要常常赞美你！
PS|71|7|许多人看我为异类， 但你是我坚固的避难所。
PS|71|8|我要满口述说赞美你的话 终日荣耀你。
PS|71|9|我年老的时候，求你不要丢弃我！ 我体力衰弱时，求你不要离弃我！
PS|71|10|我的仇敌议论我， 那些窥探要害我命的一同商议，
PS|71|11|说：“上帝已经离弃他； 你们去追赶他，捉拿他吧！ 因为没有人搭救。”
PS|71|12|上帝啊，求你不要远离我！ 我的上帝啊，求你速速帮助我！
PS|71|13|愿那与我为敌的，羞愧灭亡； 愿那谋害我的，受辱蒙羞。
PS|71|14|我却要常常仰望， 并要越发赞美你。
PS|71|15|我的口要终日述说你的公义和你的救恩， 因我无从计算其数。
PS|71|16|我要述说主耶和华的大能， 我单要提说你的公义。
PS|71|17|上帝啊，自我年幼，你就教导我； 直到如今，我传扬你奇妙的作为。
PS|71|18|上帝啊，我年老发白的时候， 求你不要离弃我！ 等我宣扬你的能力给下一代， 宣扬你的大能给后世的人。
PS|71|19|上帝啊，你的公义极高； 行过大事的上帝啊，谁能像你？
PS|71|20|你是叫我多经历重大急难的， 必使我再活过来， 从地的深处救我上来。
PS|71|21|你必使我越发昌大， 又转来安慰我。
PS|71|22|我的上帝啊，我要鼓瑟称谢你， 称谢你的信实！ 以色列 的圣者啊，我要弹琴歌颂你！
PS|71|23|我歌颂你的时候，我的嘴唇要欢呼； 我的性命，就是你所救赎的，也要欢呼。
PS|71|24|我的舌头也必终日讲论你的公义， 因为那些谋害我的人已经蒙羞受辱了。
PS|72|1|上帝啊，求你将你的公平赐给王， 将你的公义赐给王的儿子。
PS|72|2|使他按公义审判你的子民， 按公平审判你的困苦人。
PS|72|3|大山小山都要因公义 使百姓得享平安。
PS|72|4|他必为百姓中困苦的人伸冤， 拯救贫穷之辈， 压碎那欺压人的人。
PS|72|5|太阳还存，月亮犹在， 人要敬畏你 ，直到万代！
PS|72|6|他必降临，像雨降在已割的草地上， 如甘霖滋润田地。
PS|72|7|在他的日子，公义 要兴旺， 大有平安，除非月亮不在。
PS|72|8|他要执掌权柄，从这海直到那海， 从 大河 直到地极。
PS|72|9|住在旷野的必在他面前下拜， 他的仇敌必要舔土。
PS|72|10|他施 和海岛的王要进贡， 示巴 和 西巴 的王要献礼物。
PS|72|11|众王都要叩拜他， 万国都要事奉他。
PS|72|12|贫穷人呼求，他要搭救， 无人帮助的困苦人，他也搭救。
PS|72|13|他要怜悯贫寒和贫穷的人， 拯救贫穷人的性命。
PS|72|14|他要救赎他们脱离欺压和残暴， 他们的血在他眼中看为宝贵。
PS|72|15|愿他永远活着， 示巴 的金子要献给他； 愿人常常为他祷告，终日祝福他。
PS|72|16|在地的山顶上，愿五谷茂盛， 所结的谷实响动，如 黎巴嫩 的树林； 愿城里的人兴旺，如地上的草。
PS|72|17|愿他的名存到永远， 他的名如太阳之长久 ； 愿人因他蒙福， 万国称他为有福。
PS|72|18|惟独耶和华－ 以色列 的上帝能行奇事， 他是应当称颂的！
PS|72|19|他荣耀的名也当称颂，直到永远。 愿他的荣耀充满全地！ 阿们！阿们！
PS|72|20|耶西 的儿子－ 大卫 的祈祷完毕。 亚萨的诗。
PS|73|1|上帝实在恩待 以色列 那些清心的人！
PS|73|2|至于我，我的脚几乎失闪， 我的步伐险些走偏；
PS|73|3|因为我嫉妒狂傲的人， 我看见恶人享平安。
PS|73|4|他们的力气强壮， 他们死的时候也没有疼痛。
PS|73|5|他们不像别人受苦， 也不像别人遭灾。
PS|73|6|所以，骄傲如链子戴在他们项上， 残暴像衣裳覆盖在他们身上。
PS|73|7|他们的眼睛 因体胖而凸出， 他们的内心放任不羁 。
PS|73|8|他们讥笑人，凭恶意说欺压人的话。 他们说话自高；
PS|73|9|他们的口亵渎上天， 他们的舌毁谤全地。
PS|73|10|所以他的百姓归到这里， 享受满杯的水 。
PS|73|11|他们说：“上帝怎能晓得？ 至高者哪会知道呢？”
PS|73|12|看哪，这就是恶人， 他们常享安逸，财宝增多。
PS|73|13|我实在徒然洁净了我的心， 徒然洗手表明我的无辜，
PS|73|14|因为我终日遭灾难， 每日早晨受惩治。
PS|73|15|我若说“我要这样讲”， 就是愧对这世代的众儿女了。
PS|73|16|我思索要明白这事， 眼看实系为难，
PS|73|17|直到我进了上帝的圣所， 思想他们的结局。
PS|73|18|你实在把他们安放在滑地， 使他们跌倒灭亡；
PS|73|19|他们转眼之间成了何等荒凉！ 他们被惊恐灭尽了。
PS|73|20|人睡醒了，怎样看梦， 主啊，你醒了也必照样轻看他们的影像。
PS|73|21|因此，我心里苦恼， 肺腑被刺。
PS|73|22|我这样愚昧无知， 在你面前如同畜牲。
PS|73|23|然而，我常与你同在； 你搀扶我的右手。
PS|73|24|你要以你的训言引导我， 以后你必接我到荣耀里。
PS|73|25|除你以外，在天上我有谁呢？ 除你以外，在地上我也没有所爱慕的。
PS|73|26|我的肉体和我的心肠衰残； 但上帝是我心里的力量， 又是我的福分，直到永远。
PS|73|27|看哪，远离你的，必要死亡； 凡离弃你行淫的，你都灭绝了。
PS|73|28|但我亲近上帝是于我有益； 我以主耶和华为我的避难所， 好叫我述说你一切的作为。
PS|74|1|上帝啊，你为何永远丢弃我们呢？ 为何向你草场的羊发怒，如烟冒出呢？
PS|74|2|求你记念你古时得来的会众， 就是你所赎、作你产业支派的， 并记念你向来居住的 锡安山 。
PS|74|3|求你举步去看那日久荒凉之地， 看仇敌在圣所中所做的一切恶事。
PS|74|4|你的敌人在你会中吼叫， 他们竖起自己的标帜为记号，
PS|74|5|好像人扬起斧子 对着林中的树，
PS|74|6|现在将圣所中的雕刻 ， 全都用斧子锤子打坏。
PS|74|7|他们用火焚烧你的圣所， 亵渎你名的居所于地。
PS|74|8|他们心里说“我们要尽行毁灭”； 就在遍地烧毁敬拜上帝聚会的所在。
PS|74|9|我们看不见自己的标帜，不再有先知， 我们当中也无人知道这灾祸要到几时。
PS|74|10|上帝啊，敌人辱骂要到几时呢？ 仇敌藐视你的名要到永远吗？
PS|74|11|你为什么缩回你的右手？ 求你从怀中伸出手来，毁灭他们。
PS|74|12|上帝自古以来是我的王， 在这地上施行拯救。
PS|74|13|你曾用能力将海分开， 你打破水里大鱼的头。
PS|74|14|你曾压碎 力威亚探 的头， 把它给旷野的禽兽作食物。
PS|74|15|你曾分裂泉源和溪流； 使长流的江河枯干。
PS|74|16|白昼属你，黑夜也属你； 亮光和太阳是你预备的。
PS|74|17|地的一切疆界是你立的， 夏天和冬天是你定的。
PS|74|18|耶和华啊，仇敌辱骂，愚顽之辈藐视你的名； 求你记念这事。
PS|74|19|不要将属你的斑鸠 交给野兽， 不要永远忘记你困苦人的性命。
PS|74|20|求你顾念所立的约， 因为地上黑暗之处遍满了凶暴。
PS|74|21|不要让受欺压的人蒙羞回去； 要使困苦贫穷的人赞美你的名。
PS|74|22|上帝啊，求你起来为自己辩护！ 求你记念愚顽人怎样终日辱骂你。
PS|74|23|不要忘记你敌人的喧闹， 就是那时常上升、起来对抗你之人的喧哗。
PS|75|1|上帝啊，我们称谢你，我们称谢你！ 你的名临近，人 都述说你奇妙的作为。
PS|75|2|我选定了日期， 必按正直施行审判。
PS|75|3|地和其上的居民都熔化了； 我亲自坚立地的柱子。（细拉）
PS|75|4|我对狂傲的人说：“不要狂傲！” 对凶恶的人说：“不要举角！”
PS|75|5|不要把你们的角高举， 不要挺着颈项 说话。
PS|75|6|因为高举非从东，非从西， 也非从南而来。
PS|75|7|惟有上帝断定， 他使这人降卑，使那人升高。
PS|75|8|耶和华的手里有杯， 杯内满了调和起沫的酒； 他倒出来， 地上的恶人都必喝，直到喝尽它的渣滓。
PS|75|9|但我要宣扬，直到永远！ 我要歌颂 雅各 的上帝！
PS|75|10|恶人一切的角，我要砍断； 惟有义人的角必被高举。
PS|76|1|在 犹大 ，上帝为人所认识； 在 以色列 ，他的名为大。
PS|76|2|在 撒冷 有他的住处， 在 锡安 有他的居所。
PS|76|3|他在那里折断弓上的火箭、 盾牌、刀剑和战争的兵器。（细拉）
PS|76|4|你是光荣的， 比猎物 之山更威严。
PS|76|5|心中勇敢的人都被掠夺； 他们睡了长觉，没有一个英雄能措手。
PS|76|6|雅各 的上帝啊，你的斥责一发， 战车和战马都沉睡了。
PS|76|7|你，惟独你是可畏的！ 你的怒气一发，谁能在你面前站得住呢？
PS|76|8|你从天上使人听判断。 上帝起来施行审判， 要救地上所有困苦的人； 那时地就惧怕而静默。（细拉）
PS|76|9|
PS|76|10|人的愤怒终必称谢你， 你要以人的余怒束腰。
PS|76|11|你们当向耶和华－你们的上帝许愿，还愿； 在他四围的人都当拿贡物献给那可畏的主。
PS|76|12|他要挫折王子的骄气， 向地上的君王显为可畏。
PS|77|1|我要向上帝发声呼求； 我向上帝发声，他必侧耳听我。
PS|77|2|我在患难之日寻求主， 在夜间不住地举手祷告 ， 我的心不肯受安慰。
PS|77|3|我想念上帝，就烦躁不安； 我沉思默想，心灵发昏。（细拉）
PS|77|4|你使我不能闭眼； 我心烦乱，甚至不能说话。
PS|77|5|我追想古时之日， 上古之年。
PS|77|6|夜间我想起我的歌曲 ， 我的心默想，我的灵仔细省察：
PS|77|7|“难道主要永远丢弃我， 不再施恩吗？
PS|77|8|难道他的慈爱永远穷尽， 他的应许世世废弃吗？
PS|77|9|难道上帝忘记施恩， 因发怒就止住他的怜悯吗？”（细拉）
PS|77|10|我说，至高者右手的能力已改变， 这是我的悲哀。
PS|77|11|我要记念耶和华所做的， 要记念你古时的奇事；
PS|77|12|我要思想你所做的， 默念你的作为。
PS|77|13|上帝啊，你的道是神圣的； 有何神明大如上帝呢？
PS|77|14|你是行奇事的上帝， 你曾在万民中彰显能力。
PS|77|15|你曾用膀臂赎了你的子民， 就是 雅各 和 约瑟 的子孙。（细拉）
PS|77|16|上帝啊，众水见你， 众水一见你就都惊惶， 深渊也都战抖。
PS|77|17|密云倒出水来， 天空发出响声， 你的箭也飞行四方。
PS|77|18|你的雷声在旋风之中， 闪电照亮世界， 大地战抖震动。
PS|77|19|你的道在海中， 你的路在大水之中， 你的脚踪无人知道。
PS|77|20|你曾藉 摩西 和 亚伦 的手引导你的百姓， 好像领羊群一般。
PS|78|1|我的子民哪，要侧耳听我的训诲， 竖起耳朵听我口中的言语。
PS|78|2|我要开口说比喻， 我要解开古时的谜语，
PS|78|3|是我们所听见、所知道， 我们的祖宗告诉我们的。
PS|78|4|我们不要向子孙隐瞒这些事， 而要将耶和华的美德和他的能力， 并他所行的奇事，述说给后代听。
PS|78|5|他在 雅各 中立法度， 在 以色列 中设律法； 他吩咐我们的祖宗要传给子孙，
PS|78|6|使将要生的后代子孙可以晓得。 他们也要起来告诉他们的子孙，
PS|78|7|好让他们仰望上帝， 不忘记上帝的作为， 惟遵守他的命令；
PS|78|8|不要像他们的祖宗， 是顽梗悖逆、心不坚定， 向上帝心不忠实之辈。
PS|78|9|以法莲 人带着兵器，拿着弓， 临阵之日转身退后。
PS|78|10|他们不遵守上帝的约， 不肯照他的律法行；
PS|78|11|又忘记他的作为 和他所彰显的奇事。
PS|78|12|他在 埃及 地，在 琐安 田， 在他们祖宗眼前施行奇事。
PS|78|13|他把海分开，使他们过去， 又叫水立起如垒。
PS|78|14|他白日用云彩， 终夜用火光引导他们。
PS|78|15|他在旷野使磐石裂开， 多多地给他们水喝，如从深渊而出。
PS|78|16|他使水从磐石涌出， 叫水如江河下流。
PS|78|17|他们却仍旧得罪他， 在干旱之地悖逆至高者。
PS|78|18|他们心中试探上帝， 随自己所欲的求食物，
PS|78|19|并且妄论上帝说： “上帝岂能在旷野摆设筵席吗？
PS|78|20|他虽曾击打磐石，使水涌出，如江河泛滥； 他还能赐粮食吗？ 还能为他的百姓预备吃的肉吗？”
PS|78|21|所以，耶和华听见就发怒， 有烈火向 雅各 点燃， 有怒气向 以色列 上腾；
PS|78|22|因为他们不信服上帝， 不倚赖他的拯救。
PS|78|23|然而他却吩咐天空， 又敞开天上的门，
PS|78|24|降吗哪像雨，给他们吃， 将天上的粮食赐给他们。
PS|78|25|各人就吃大能者的食物； 他赐下粮食，使他们饱足。
PS|78|26|他令东风吹在天空， 用能力引来南风。
PS|78|27|他降肉像雨，多如尘土， 降飞鸟，多如海沙，
PS|78|28|落在他自己的营中， 在他帐幕的四周围。
PS|78|29|他们吃了，而且饱足； 这样就随了他们所欲的。
PS|78|30|但在他们满足食欲以前， 食物还在他们口中的时候，
PS|78|31|上帝的怒气就向他们上腾， 杀了他们当中肥壮的人， 打倒 以色列 的青年。
PS|78|32|虽是这样，他们仍旧犯罪， 不信他奇妙的作为。
PS|78|33|因此，他使他们的日子全归虚空， 叫他们的年岁尽属惊恐。
PS|78|34|他杀他们的时候，他们才求问他， 回心转意，切切寻求上帝。
PS|78|35|他们追念上帝是他们的磐石， 至高的上帝是他们的救赎主。
PS|78|36|他们却用口谄媚他， 用舌向他说谎。
PS|78|37|他们的心向他不坚定， 不忠于他的约。
PS|78|38|但他有怜悯， 赦免他们的罪孽， 没有灭绝他们， 而且屡次撤销他的怒气， 不发尽他的愤怒。
PS|78|39|他想念他们不过是血肉之躯， 是一阵去而不返的风。
PS|78|40|他们在旷野悖逆他， 在荒地令他担忧，何其多呢！
PS|78|41|他们再三试探上帝， 惹动 以色列 的圣者。
PS|78|42|他们不追念他手的能力， 和他救赎他们脱离敌人的日子；
PS|78|43|他怎样在 埃及 显神迹， 在 琐安 田显奇事，
PS|78|44|把江河并河汊的水都变为血， 使他们不能喝。
PS|78|45|他使苍蝇成群落在他们当中，吃尽他们， 又叫青蛙灭了他们，
PS|78|46|将他们的果实交给蚂蚱， 把他们劳碌得来的交给蝗虫。
PS|78|47|他降冰雹打坏他们的葡萄树， 下寒霜打坏他们的桑树，
PS|78|48|将他们的牲畜交给冰雹， 把他们的群畜交给闪电。
PS|78|49|他使猛烈的怒气和愤怒、恼恨、苦难， 成了一群降灾的使者，临到他们。
PS|78|50|他为自己的怒气修平了路， 将他们的性命交给瘟疫， 使他们死亡，
PS|78|51|在 埃及 击杀所有的长子， 在 含 的帐棚中击杀他们壮年时头生的。
PS|78|52|他却领出自己的子民如羊， 在旷野引导他们如羊群。
PS|78|53|他领他们稳稳妥妥地，使他们不致害怕； 海却淹没他们的仇敌。
PS|78|54|他带他们到自己圣地的边界， 到他右手所得的这山地。
PS|78|55|他在他们面前赶出外邦人， 用绳子抽签量地给他们为业， 让 以色列 支派的人住在自己的帐棚里。
PS|78|56|他们仍旧试探，悖逆至高的上帝， 不遵守他的法度，
PS|78|57|反倒退后，行诡诈，像他们的祖宗一样， 他们翻转，如同松弛的弓，
PS|78|58|以丘坛惹他发怒， 以雕刻的偶像使他忌恨。
PS|78|59|上帝听见就发怒， 全然弃绝了 以色列 ，
PS|78|60|甚至离弃 示罗 的帐幕， 就是他在人间所搭的帐棚；
PS|78|61|又将他有能力的约柜 交给人掳去， 将他的荣耀交在敌人手中；
PS|78|62|并将他的百姓交给刀剑， 向他的产业发怒。
PS|78|63|壮丁被火烧灭， 童女也无婚礼颂歌。
PS|78|64|祭司倒在刀下， 寡妇却不哀哭。
PS|78|65|那时，主像睡觉的人醒来， 如勇士饮酒呼喊。
PS|78|66|他击退敌人， 叫他们永蒙羞辱。
PS|78|67|他撇弃 约瑟 的帐棚， 不拣选 以法莲 支派，
PS|78|68|却拣选 犹大 支派， 拣选他所喜爱的 锡安山 ；
PS|78|69|建造他的圣所如同高峰， 又像他所建立的永存之地。
PS|78|70|他拣选他的仆人 大卫 ， 从羊圈中将他召来，
PS|78|71|叫他不再牧放那些母羊， 为要牧养自己的百姓 雅各 和自己的产业 以色列 。
PS|78|72|于是，他以纯正的心牧养他们， 用巧妙的手引导他们。
PS|79|1|上帝啊，外邦人侵犯你的产业， 玷污你的圣殿，使 耶路撒冷 变成废墟，
PS|79|2|将你仆人的尸首交给天空的飞鸟为食， 把你圣民的肉交给地上的走兽，
PS|79|3|耶路撒冷 的周围流出他们的血如水， 无人埋葬。
PS|79|4|我们成为邻国羞辱的对象， 被四围的人嗤笑讥刺。
PS|79|5|耶和华啊，你发怒要到几时呢？ 要到永远吗？ 你的忌恨要如火焚烧吗？
PS|79|6|求你将你的愤怒倾倒在那不认识你的万邦 和那不求告你名的国度。
PS|79|7|因为他们吞了 雅各 ， 将他的住处变为废墟。
PS|79|8|求你不要记得我们先前世代的罪孽； 愿你的怜悯速速临到我们， 因为我们落到极卑微的地步。
PS|79|9|拯救我们的上帝啊，求你因你名的荣耀帮助我们！ 为你名的缘故搭救我们，赦免我们的罪。
PS|79|10|为何让列国说“他们的上帝在哪里”呢？ 求你让列国知道， 你在我们眼前伸你仆人流血的冤。
PS|79|11|愿被囚之人的叹息达到你面前， 求你以强大的膀臂存留那些将死的人。
PS|79|12|主啊，求你将我们邻邦所加给你的羞辱 七倍归到他们身上。
PS|79|13|这样，你的子民，你草场的羊， 要称谢你，直到永远； 要述说赞美你的话，直到万代。
PS|80|1|领 约瑟 如领羊群的 以色列 牧者啊，求你侧耳而听！ 在基路伯之上坐宝座的啊，求你发出光来！
PS|80|2|在 以法莲 、 便雅悯 、 玛拿西 面前 求你施展你的大能，拯救我们。
PS|80|3|上帝啊，求你使我们回转 ， 使你的脸发光，我们就会得救！
PS|80|4|耶和华─万军之上帝啊， 你因你百姓的祷告发怒，要到几时呢？
PS|80|5|你以眼泪当食物给他们吃， 量出满碗的眼泪给他们喝。
PS|80|6|你使邻邦因我们纷争， 我们的仇敌彼此戏笑。
PS|80|7|万军之上帝啊，求你使我们回转， 使你的脸发光，我们就会得救！
PS|80|8|你从 埃及 拔出一棵葡萄树， 赶出外邦人，把这树栽上。
PS|80|9|你在它面前清除杂物， 它就深深扎根，蔓延满地。
PS|80|10|它的影子遮蔽群山， 枝子好像高大的香柏树。
PS|80|11|它长出枝子，直到大海， 伸展嫩枝，延到 大河 。
PS|80|12|你为何拆毁这树的篱笆， 任凭路人摘取？
PS|80|13|林中的野猪践踏它， 田里的走兽吞吃它。
PS|80|14|万军之上帝啊，求你转回， 从天上垂看观察，眷顾这葡萄树；
PS|80|15|保护你右手所栽的根， 你为自己所坚固的幼苗。
PS|80|16|这树已经被火焚烧，被刀砍伐， 因你脸上的怒容就灭亡了。
PS|80|17|愿你的手扶持你右边的人， 你为自己所坚固的人子。
PS|80|18|这样，我们就不背离你； 求你救活我们，让我们得以求告你的名。
PS|80|19|耶和华─万军之上帝啊，求你使我们回转， 使你的脸发光，我们就会得救！
PS|81|1|你们当向上帝－我们的力量大声歌唱， 向 雅各 的上帝欢呼！
PS|81|2|高唱诗歌，击打手鼓， 弹奏悦耳的琴瑟。
PS|81|3|当在新月和满月－ 我们过节的日期吹角，
PS|81|4|因这是为 以色列 所定的律例， 是 雅各 上帝的典章。
PS|81|5|他攻击 埃及 地的时候， 曾立此为 约瑟 的法度。 我听见我所不明白的语言：
PS|81|6|“我使你 的肩头得脱重担， 使你的手放下筐子。
PS|81|7|你在急难中呼求，我就搭救你， 在雷的隐密处应允你， 在 米利巴 水那里考验你。（细拉）
PS|81|8|听啊，我的子民，我要劝戒你； 以色列 啊，我真愿你肯听从我。
PS|81|9|在你当中，不可有外族的神明； 外邦的神明，你也不可下拜。
PS|81|10|我是耶和华－你的上帝， 曾将你从 埃及 地领上来； 你要大大张口，我就使你满足。
PS|81|11|“无奈，我的子民不听我的声音， 以色列 不肯听从我。
PS|81|12|我就任凭他们心里顽梗， 随自己的计谋而行。
PS|81|13|我的子民若肯听从我， 以色列 肯行我的道，
PS|81|14|我就速速制伏他们的仇敌， 反手攻击他们的敌人。
PS|81|15|恨耶和华的人必来投降， 愿他们的厄运直到永远。
PS|81|16|他必拿上好的麦子给 以色列 吃， 又拿磐石出的蜂蜜使你饱足。 ”
PS|82|1|上帝站立在神圣的会中， 在诸神中施行审判。
PS|82|2|你们审判不秉公义， 抬举恶人的脸面，要到几时呢？（细拉）
PS|82|3|当为贫寒的人和孤儿伸冤， 为困苦和穷乏的人施行公义。
PS|82|4|当保护贫寒和贫穷的人， 救他们脱离恶人的手。
PS|82|5|他们愚昧，他们无知， 在黑暗中走来走去； 地的根基都摇动了。
PS|82|6|我曾说：“你们是诸神， 都是至高者的儿子。
PS|82|7|然而，你们要死去，与世人一样， 要仆倒，像任何一位王子一般。”
PS|82|8|上帝啊，求你起来审判全地， 因为你必得万国为业。
PS|83|1|上帝啊，求你不要静默！ 上帝啊，求你不要闭口，不要不作声！
PS|83|2|因为你的仇敌喧嚷， 恨你的抬起头来。
PS|83|3|他们同谋奸诈要害你的百姓， 彼此商议要害你所保护的人。
PS|83|4|他们说：“来吧，我们将他们除灭， 使他们不再成国！ 使 以色列 的名不再被人记念！”
PS|83|5|他们同心商议， 彼此结盟，要抵挡你；
PS|83|6|他们就是住帐棚的 以东 和 以实玛利 人， 摩押 和 夏甲 人，
PS|83|7|迦巴勒 、 亚扪 、 亚玛力 、 非利士 和 推罗 的居民。
PS|83|8|亚述 也与他们联合， 作 罗得 子孙的帮手。（细拉）
PS|83|9|求你待他们，如待 米甸 ， 如在 基顺河 待 西西拉 和 耶宾 一样。
PS|83|10|他们在 隐．多珥 灭亡， 成了地上的粪土。
PS|83|11|求你使他们的贵族像 俄立 和 西伊伯 ， 使他们的王子都像 西巴 和 撒慕拿 。
PS|83|12|因为他们说：“我们要得上帝的住处， 作自己的产业。”
PS|83|13|我的上帝啊，求你使他们像旋风中的尘土， 如风前的碎秸。
PS|83|14|火怎样焚烧树林， 火焰怎样烧着山岭，
PS|83|15|求你也照样用狂风追赶他们， 用暴雨恐吓他们。
PS|83|16|耶和华啊，求你使他们满面羞耻， 好叫他们寻求你的名！
PS|83|17|愿他们永远羞愧惊惶！ 愿他们惭愧灭亡！
PS|83|18|愿他们认识你的名是耶和华， 惟独你是掌管全地的至高者！
PS|84|1|万军之耶和华啊， 你的居所何等可爱！
PS|84|2|我羡慕渴想耶和华的院宇， 我的内心，我的肉体向永生上帝欢呼。
PS|84|3|万军之耶和华－我的王，我的上帝啊， 在你祭坛那里，麻雀为自己找到了家， 燕子为自己找着菢雏之窝。
PS|84|4|如此住在你殿中的有福了！ 他们不断地赞美你。（细拉）
PS|84|5|靠你有力量、心中向往 锡安 大道的， 这人有福了！
PS|84|6|他们经过“流泪谷” ，叫这谷变为泉源之地； 且有秋雨之福盖满了全谷。
PS|84|7|他们行走，力上加力， 各人到 锡安 朝见上帝。
PS|84|8|万军之耶和华上帝啊，求你听我的祷告！ 雅各 的上帝啊，求你侧耳而听！（细拉）
PS|84|9|上帝啊，我们的盾牌，求你观看， 求你垂顾你受膏者的面！
PS|84|10|在你的院宇一日， 胜似千日； 宁可在我上帝的殿中看门， 不愿住在恶人的帐棚里。
PS|84|11|因为耶和华上帝是太阳，是盾牌， 耶和华要赐下恩惠和荣耀。 他未尝留下福气不给那些行动正直的人。
PS|84|12|万军之耶和华啊， 倚靠你的人有福了！
PS|85|1|耶和华啊，你已经向你的地施恩， 救回被掳的 雅各 。
PS|85|2|你赦免了你百姓的罪孽， 遮盖了他们一切的过犯。（细拉）
PS|85|3|你收回所发的愤怒， 撤销你猛烈的怒气。
PS|85|4|拯救我们的上帝啊，求你使我们回转， 使你向我们所发的愤怒止息。
PS|85|5|你要向我们发怒到永远吗？ 要将你的怒气延留到万代吗？
PS|85|6|你不再将我们救活， 使你的百姓因你欢喜吗？
PS|85|7|耶和华啊，求你使我们得见你的慈爱， 又将你的救恩赐给我们。
PS|85|8|我要听上帝－耶和华所说的话， 因为他必应许赐平安给他的百姓，就是他的圣民； 他们却不可再转向愚昧 。
PS|85|9|他的救恩诚然与敬畏他的人相近， 使荣耀住在我们的地上。
PS|85|10|慈爱和诚实彼此相遇， 公义与和平彼此相亲。
PS|85|11|诚实从地而生， 公义从天而现。
PS|85|12|耶和华必赐福气给我们； 我们的地也要出土产。
PS|85|13|公义要行在他面前， 使他的脚踪有可走之路。
PS|86|1|耶和华啊，求你侧耳应允我， 因我是困苦贫穷的。
PS|86|2|求你保住我的性命，因我是虔诚的人。 我的上帝啊，求你拯救我这倚靠你的仆人！
PS|86|3|主啊，求你怜悯我， 因我终日求告你。
PS|86|4|主啊，求你使你的仆人心里欢喜， 因为我的心仰望你。
PS|86|5|主啊，你本为良善，乐于饶恕人， 以丰盛的慈爱对待凡求告你的人。
PS|86|6|耶和华啊，求你侧耳听我的祷告， 留心听我恳求的声音。
PS|86|7|我在患难之日要求告你， 因为你必应允我。
PS|86|8|主啊，诸神之中没有可与你相比的， 你的作为也无以为比。
PS|86|9|主啊，你所造的万民都要来敬拜你， 他们要荣耀你的名。
PS|86|10|因你本为大，且行奇妙的事， 惟独你是上帝。
PS|86|11|耶和华啊，求你将你的道指教我， 我要照你的真理而行； 求你使我专心敬畏你的名！
PS|86|12|主－我的上帝啊，我要一心称谢你； 我要荣耀你的名，直到永远。
PS|86|13|因为你的慈爱在我身上浩大， 你救了我的性命免入阴间的深处。
PS|86|14|上帝啊，骄傲的人起来攻击我， 又有一群强横的人寻索我的命； 他们没有将你放在眼里。
PS|86|15|主啊，你是有怜悯，有恩惠的上帝， 不轻易发怒，并有丰盛的慈爱和信实。
PS|86|16|求你转向我，怜悯我， 将你的力量赐给仆人，拯救你使女的儿子。
PS|86|17|求你向我显出恩待我的凭据， 使恨我的人看见就羞愧， 因为你－耶和华帮助我，安慰了我。
PS|87|1|耶和华所立的根基在圣山上。
PS|87|2|耶和华爱 锡安 的门， 胜于爱 雅各 一切的住处。
PS|87|3|上帝的城啊， 有荣耀的事是指着你说的。（细拉）
PS|87|4|我要提起 拉哈伯 和 巴比伦 人， 是在认识我之中的； 看哪， 非利士 、 推罗 和 古实 人， 个个生在那里。
PS|87|5|论到 锡安 ，必有话说： “这一个、那一个都生在其中”； 而且至高者必亲自坚立这城。
PS|87|6|当耶和华记录万民的时候， 他要写出人的出生地。（细拉）
PS|87|7|歌唱的、跳舞的，都要说： “我的泉源都在你里面。”
PS|88|1|耶和华－拯救我的上帝啊， 我昼夜在你面前呼求；
PS|88|2|愿我的祷告达到你面前， 求你侧耳听我的恳求！
PS|88|3|因为我心里满了患难， 我的性命临近阴间；
PS|88|4|我与下到地府的人同列， 如同无人帮助的人一样。
PS|88|5|我被丢在死人中， 好像被杀的人躺在坟墓里， 不再被你记得， 与你的手隔绝了。
PS|88|6|你把我放在极深的地府里， 在黑暗地，在深处。
PS|88|7|你的愤怒重压我身， 你用一切的波浪困住我。（细拉）
PS|88|8|你把我所认识的人隔在远处， 使我为他们所憎恶； 我被拘禁，不能出来。
PS|88|9|我的眼睛因困苦而昏花； 耶和华啊，我天天求告你，向你举手。
PS|88|10|你岂要行奇事给死人看吗？ 阴魂还能起来称谢你吗？（细拉）
PS|88|11|你的慈爱岂能在坟墓里被人述说吗？ 你的信实岂能在冥府 被人传扬吗？
PS|88|12|你的奇事岂能在幽暗里为人所知吗？ 你的公义岂能在遗忘之地为人所识吗？
PS|88|13|耶和华啊，至于我，我要呼求你； 每早晨，我的祷告要达到你面前。
PS|88|14|耶和华啊，你为何丢弃我？ 为何转脸不顾我？
PS|88|15|我自幼受苦，几乎死亡； 你使我惊恐，烦乱不安。
PS|88|16|你的烈怒漫过我身， 你用惊吓把我除灭。
PS|88|17|这些如水终日环绕我， 一起围困我。
PS|88|18|你把我的良朋密友隔在远处， 使我所认识的人都在黑暗里 。
PS|89|1|我要歌唱耶和华的慈爱，直到永远， 我要用口将你的信实传到万代。
PS|89|2|因我曾说：“你的慈爱必建立到永远， 你的信实必坚立在天上。”
PS|89|3|“我与我所拣选的人立了约， 向我的仆人 大卫 起了誓：
PS|89|4|‘我要坚立你的后裔，直到永远， 要建立你的宝座，直到万代。’”（细拉）
PS|89|5|耶和华啊，诸天要称谢你的奇事； 在圣者的会中，要称谢你的信实。
PS|89|6|因在天空谁能比耶和华呢？ 诸神之中，谁能像耶和华呢？
PS|89|7|在圣者的会中，他是大有威严的上帝， 比在他四围所有的更可畏惧。
PS|89|8|耶和华－万军之上帝啊， 哪一个大能者像耶和华？ 你的信实在你四围。
PS|89|9|你管辖海的狂傲； 波浪翻腾，你使它平静了。
PS|89|10|你打碎了 拉哈伯 ，使它如遭刺杀的人； 你用大能的膀臂打散了你的仇敌。
PS|89|11|天属你，地也属你； 世界和其中所充满的都为你所建立。
PS|89|12|南北为你所创造； 他泊 和 黑门 都因你的名欢呼。
PS|89|13|你有大能的膀臂， 你的手有力，你的右手也高举。
PS|89|14|公义和公平是你宝座的根基， 慈爱和信实行在你前面。
PS|89|15|知道向你欢呼的，那民有福了！ 耶和华啊，他们要行走在你脸的光中。
PS|89|16|他们因你的名终日欢乐， 因你的公义得以高举。
PS|89|17|你是他们力量的荣耀。 我们的角必被高举，因为你喜爱我们。
PS|89|18|我们的盾牌是耶和华， 我们的王是 以色列 的圣者。
PS|89|19|当时，你在异象中吩咐你的圣民，说： “我已把救助之力加在壮士身上， 高举了那从百姓中所拣选的人。
PS|89|20|我寻得我的仆人 大卫 ， 用我的圣膏膏他。
PS|89|21|我的手必使他坚立， 我的膀臂也必坚固他。
PS|89|22|仇敌必不勒索他， 凶恶之子也不苦害他。
PS|89|23|我要在他面前打碎他的敌人， 击杀那些恨他的人。
PS|89|24|我的信实和我的慈爱要与他同在； 因我的名，他的角必被高举。
PS|89|25|我要使他的手伸到海上， 右手伸到河上。
PS|89|26|他要称呼我说：‘你是我的父， 是我的上帝，是拯救我的磐石。’
PS|89|27|我也要立他为长子， 为世上最高的君王。
PS|89|28|我要为他存留我的慈爱，直到永远， 我与他所立的约必坚定不移。
PS|89|29|我也要使他的后裔存到永远， 使他的宝座如天之久。
PS|89|30|“倘若他的子孙离弃我的律法， 不照我的典章行，
PS|89|31|背弃我的律例， 不遵守我的诫命，
PS|89|32|我就要用杖责罚他们的过犯， 用鞭责罚他们的罪孽。
PS|89|33|只是我不将我的慈爱全然收回， 也不叫我的信实废除。
PS|89|34|我必不毁损我的约， 也不改变我口中所出的话。
PS|89|35|我仅此一次指着自己的神圣起誓， 我绝不向 大卫 说谎！
PS|89|36|他的后裔要存到永远， 他的宝座在我面前如太阳，
PS|89|37|又如月亮永远坚立； 天上的见证是确实的。”（细拉）
PS|89|38|但你恼怒你的受膏者， 拒绝他，离弃了他。
PS|89|39|你厌恶与你仆人所立的约， 将他的冠冕践踏于地。
PS|89|40|你拆毁了他一切的围墙， 使他的堡垒变为废墟。
PS|89|41|过路的人都抢夺他， 他成了邻邦羞辱的对象。
PS|89|42|你高举了他敌人的右手， 使他所有的仇敌欢喜。
PS|89|43|你叫他的刀剑卷刃， 使他在战争中站立不住。
PS|89|44|你使他的光辉止息， 将他的宝座推倒于地。
PS|89|45|你减少他年轻的日子， 又使他蒙羞。（细拉）
PS|89|46|耶和华啊，这要到几时呢？ 你要隐藏自己到永远吗？ 你的愤怒如火焚烧要到几时呢？
PS|89|47|求你想念我的生命是何等短暂。 你创造世人，要使他们归于何等的虚空呢？
PS|89|48|谁能常活不见死亡、 救自己脱离阴间的掌控呢？（细拉）
PS|89|49|主啊，你从前凭你的信实 向 大卫 起誓要施行的慈爱在哪里呢？
PS|89|50|主啊，求你记念仆人们所受的羞辱， 记念我怎样将万族所加的羞辱都放在我的胸怀。
PS|89|51|耶和华啊，这是你仇敌所加的羞辱， 羞辱了你受膏者的脚踪。
PS|89|52|耶和华是应当称颂的，直到永远。 阿们！阿们！ 神人摩西的祈祷。
PS|90|1|主啊，你世世代代作我们的居所。
PS|90|2|诸山未曾生出， 地与世界你未曾造成， 从亘古到永远，你是上帝。
PS|90|3|你使人归于尘土，说： “世人哪，你们要归回。”
PS|90|4|在你看来，千年如已过的昨日， 又如夜间的一更。
PS|90|5|你叫他们如水冲去， 他们如睡一觉。 早晨，他们如生长的草；
PS|90|6|早晨发芽生长， 晚上割下枯干。
PS|90|7|我们因你的怒气而消灭， 因你的愤怒而惊惶。
PS|90|8|你将我们的罪孽摆在你面前， 将我们的隐恶摆在你面光之中。
PS|90|9|我们经过的日子，都在你震怒之下， 我们度尽的年岁，好像一声叹息。
PS|90|10|我们一生的年日是七十岁， 若是强壮可到八十岁； 但其中所矜夸的不过是劳苦愁烦， 转眼即逝，我们便如飞而去。
PS|90|11|谁晓得你怒气的权势？ 谁因着敬畏你而晓得你的愤怒呢？
PS|90|12|求你指教我们怎样数算自己的日子， 好叫我们得着智慧的心。
PS|90|13|耶和华啊，我们要等到几时呢？ 求你转回，怜悯你的仆人们。
PS|90|14|求你使我们早早饱得你的慈爱， 好叫我们一生一世欢呼喜乐。
PS|90|15|求你照着你使我们受苦的日子， 和我们遭难的年岁，使我们喜乐。
PS|90|16|愿你的作为向你仆人们显现， 愿你的荣耀向他们子孙显明。
PS|90|17|愿主－我们上帝的恩宠归于我们身上。 愿你坚立我们手所做的工， 我们手所做的工，愿你坚立。
PS|91|1|住在至高者隐密处的， 必住在全能者的荫下。
PS|91|2|我要向耶和华说： “我的避难所、我的山寨、 我的上帝，你是我所倚靠的。”
PS|91|3|他必救你脱离捕鸟者的罗网 和毁灭人的瘟疫。
PS|91|4|他必用自己的翎毛遮蔽你； 你要投靠在他翅膀底下， 他的信实是大小的盾牌。
PS|91|5|你必不怕黑夜的惊骇， 或是白日飞的箭，
PS|91|6|也不怕黑夜流行的瘟疫， 或是午间灭人的灾害。
PS|91|7|虽有千人仆倒在你旁边， 万人仆倒在你右边， 这灾却不得临近你。
PS|91|8|你惟亲眼观看， 见恶人遭报。
PS|91|9|因为耶和华是我的避难所， 你以至高者为居所，
PS|91|10|祸患必不临到你， 灾害也不挨近你的帐棚。
PS|91|11|因他要为你命令他的使者， 在你所行的一切道路上保护你。
PS|91|12|他们要用手托住你， 免得你的脚碰在石头上。
PS|91|13|你要踹踏狮子和毒蛇， 践踏少壮狮子和大蛇。
PS|91|14|“因为他专心爱我，我要搭救他； 因为他认识我的名，我要把他安置在高处。
PS|91|15|他若求告我，我就应允他； 他在急难中，我与他同在； 我要搭救他，使他尊贵。
PS|91|16|我要使他享足长寿， 将我的救恩显明给他。”
PS|92|1|这是多么好啊！ 称谢耶和华， 歌颂你至高者的名，
PS|92|2|早晨传扬你的慈爱， 每夜传扬你的信实。
PS|92|3|用十弦的乐器和瑟， 用琴优雅的声音；
PS|92|4|因你－耶和华藉着你的作为使我高兴， 我要因你手的工作欢呼。
PS|92|5|耶和华啊，你的工作何其大！ 你的心思极其深！
PS|92|6|畜牲一般的人不晓得， 愚昧人也不明白。
PS|92|7|恶人虽茂盛如草， 作恶的人虽全都兴旺， 他们却要灭亡， 直到永远。
PS|92|8|耶和华啊，惟有你是至高， 直到永远。
PS|92|9|耶和华啊，看哪，你的仇敌， 看哪，你的仇敌都要灭亡； 作恶的全都要离散。
PS|92|10|你却高举了我的角，如野牛的角； 我是被新油膏抹的。
PS|92|11|我的眼睛看见我的仇敌遭报， 我的耳朵听见那些起来攻击我的恶人受罚。
PS|92|12|义人要兴旺如棕树， 生长如 黎巴嫩 的香柏树。
PS|92|13|他们栽于耶和华的殿中， 发旺在我们上帝的院里。
PS|92|14|他们发白的时候仍结果子， 而且鲜美多汁，
PS|92|15|好显明耶和华是正直的； 他是我的磐石，在他毫无不义。
PS|93|1|耶和华作王！ 他以威严为衣穿上； 耶和华以能力为衣，以能力束腰， 世界就坚定，不得动摇。
PS|93|2|你的宝座从太初立定， 你从亘古就有。
PS|93|3|耶和华啊，大水扬起， 大水发声，大水澎湃。
PS|93|4|耶和华在高处大有威力， 胜过诸水的响声，洋海的大浪。
PS|93|5|耶和华啊，你的法度最为确定； 你的殿宜称为圣，直到永远。
PS|94|1|耶和华啊，你是伸冤的上帝； 伸冤的上帝啊，求你发出光来！
PS|94|2|审判世界的主啊，求你挺身而立， 使骄傲的人受应得的报应！
PS|94|3|耶和华啊，恶人夸胜要到几时呢？ 要到几时呢？
PS|94|4|他们咆哮，说狂妄的话， 作恶的人全都夸耀自己。
PS|94|5|耶和华啊，他们强压你的百姓， 苦害你的产业。
PS|94|6|他们杀死寡妇和寄居的人， 又杀害孤儿。
PS|94|7|他们说：“耶和华必不看见， 雅各 的上帝必不留意。”
PS|94|8|百姓中像畜牲一般的人当思想， 你们愚昧人要到几时才有智慧呢？
PS|94|9|造耳朵的，难道自己听不见吗？ 造眼睛的，难道自己看不见吗？
PS|94|10|管教列国的，就是叫人得知识的， 难道自己不惩治人吗？
PS|94|11|耶和华知道人的意念是虚妄的。
PS|94|12|耶和华啊，你所管教、 用律法教导的人有福了！
PS|94|13|你使他在遭难的日子仍得平安， 直到为恶人挖好了坑。
PS|94|14|因为耶和华必不丢弃他的百姓， 也不离弃他的产业。
PS|94|15|审判要回复公义， 心里正直的，都必跟随它。
PS|94|16|谁肯为我起来攻击邪恶的？ 谁肯为我站起抵挡作恶的？
PS|94|17|若不是耶和华帮助我， 我早就住在寂静 之中了。
PS|94|18|我若说：“我失了脚！” 耶和华啊，你的慈爱必扶持我。
PS|94|19|我心里多忧多疑， 你的安慰使我欢乐。
PS|94|20|那藉着律例玩弄奸恶、 以权位肆行残害的，岂能与你交往呢？
PS|94|21|他们大家聚集攻击义人， 将无辜的人定了死罪。
PS|94|22|但耶和华向来作我的碉堡， 我的上帝作了我投靠的磐石。
PS|94|23|他叫他们的罪孽归到自己身上， 要因他们的邪恶剪除他们； 耶和华－我们的上帝要把他们剪除。
PS|95|1|来啊，我们要向耶和华歌唱， 向拯救我们的磐石欢呼！
PS|95|2|我们要以感谢来到他面前， 用诗歌向他欢呼！
PS|95|3|因耶和华是伟大的上帝， 是超越万神的大君王。
PS|95|4|地的深处在他手中； 山的高峰也属他。
PS|95|5|海洋属他，是他造的； 旱地也是他手造成的。
PS|95|6|来啊，我们要俯伏敬拜， 在造我们的耶和华面前跪拜。
PS|95|7|因为他是我们的上帝； 我们是他草场的百姓，是他手中的羊。 惟愿你们今天听他的话！
PS|95|8|你们不可硬着心，像在 米利巴 ， 就是在旷野 玛撒 的日子。
PS|95|9|那时，你们的祖宗试我，探我， 并且观看我的作为。
PS|95|10|四十年之久，我厌烦那世代，说： “这是心里迷糊的百姓， 竟不知道我的道路！”
PS|95|11|所以，我在怒中起誓： “他们断不可进入我的安息！”
PS|96|1|你们要向耶和华唱新歌！ 全地都要向耶和华歌唱！
PS|96|2|要向耶和华歌唱，称颂他的名！ 天天传扬他的救恩！
PS|96|3|在列国中述说他的荣耀！ 在万民中述说他的奇事！
PS|96|4|因耶和华本为大，当受极大的赞美； 他在万神之上，当受敬畏。
PS|96|5|因万民的神明都属虚无； 惟独耶和华创造诸天。
PS|96|6|有尊荣和威严在他面前， 有能力与华美在他圣所。
PS|96|7|民中的万族啊，要将荣耀、能力归给耶和华， 都归给耶和华！
PS|96|8|要将耶和华的名所当得的荣耀归给他， 拿供物来进入他的院宇。
PS|96|9|当敬拜神圣荣耀的耶和华 ， 全地都要在他面前战抖！
PS|96|10|要在列国中说：“耶和华作王了！ 世界坚定，不得动摇； 他要按公正审判万民。”
PS|96|11|愿天欢喜，愿地快乐！ 愿海和其中所充满的澎湃！
PS|96|12|愿田和其中所有的都欢乐！ 那时，林中的树木都要在耶和华面前欢呼。
PS|96|13|因为他来了，他来要审判全地。 他要按公义审判世界， 按信实审判万民。
PS|97|1|耶和华作王！愿地快乐！ 愿众海岛欢喜！
PS|97|2|密云和幽暗在他四围， 公义和公平是他宝座的根基。
PS|97|3|烈火在他前头行， 烧灭他四围的敌人。
PS|97|4|他的闪电光照世界， 大地看见就震动。
PS|97|5|诸山见耶和华的面， 就是全地之主的面，就如蜡熔化。
PS|97|6|诸天表明他的公义， 万民看见他的荣耀。
PS|97|7|愿所有事奉雕刻偶像、 靠虚无神明自夸的，都蒙羞愧。 万神哪，你们都当拜他。
PS|97|8|耶和华啊，因你的判断， 锡安 听见就欢喜； 犹大 的城镇 也都快乐。
PS|97|9|因为你－耶和华至高，超乎全地； 受尊崇，远超万神之上。
PS|97|10|你们爱耶和华的，都当恨恶罪恶； 他保护圣民的性命， 搭救他们脱离恶人的手。
PS|97|11|散播亮光是为义人 ， 喜乐归于心里正直的人。
PS|97|12|义人哪，你们当靠耶和华欢喜， 当颂扬他神圣的名字 。
PS|98|1|你们要向耶和华唱新歌！ 因为他行过奇妙的事， 他的右手和圣臂施行救恩。
PS|98|2|耶和华显明了他的救恩， 在列国眼前显出公义；
PS|98|3|记念他对 以色列 家的慈爱和信实。 地的四极都看见我们上帝的救恩。
PS|98|4|全地都要向耶和华欢呼， 要扬声，欢唱，歌颂！
PS|98|5|用琴歌颂耶和华， 用琴和诗歌的声音歌颂他！
PS|98|6|用号筒和角声， 在大君王耶和华面前欢呼！
PS|98|7|愿海和其中所充满的澎湃， 愿世界和住在其间的发声。
PS|98|8|愿大水拍掌， 愿诸山在耶和华面前一同欢呼；
PS|98|9|因为他来要审判全地。 他要按公义审判世界， 按公正审判万民。
PS|99|1|耶和华作王，万民当战抖！ 他坐在基路伯的宝座上，地当动摇。
PS|99|2|耶和华在 锡安 为大， 他超越万民之上。
PS|99|3|愿他们颂扬他大而可畏的名， 他本为圣！
PS|99|4|喜爱公平、大能的王啊，你坚立公正， 在 雅各 中施行公平和公义。
PS|99|5|当尊崇耶和华－我们的上帝， 在他脚凳前下拜。 他本为圣！
PS|99|6|在他的祭司中有 摩西 和 亚伦 ， 在求告他名的人中有 撒母耳 。 他们求告耶和华，他就应允他们。
PS|99|7|他在云柱中向他们说话， 他们遵守他的法度和他所赐给他们的律例。
PS|99|8|耶和华－我们的上帝啊，你应允了他们； 你是赦免他们的上帝， 却按他们所做的报应他们。
PS|99|9|当尊崇耶和华－我们的上帝， 在他的圣山下拜， 因为耶和华－我们的上帝本为圣！
PS|100|1|普天下当向耶和华欢呼！
PS|100|2|当乐意事奉耶和华， 当欢唱来到他面前！
PS|100|3|当认识耶和华是上帝！ 我们是他造的，也是属他的； 我们是他的民，是他草场的羊。
PS|100|4|当称谢进入他的门， 当赞美进入他的院。 当感谢他，称颂他的名！
PS|100|5|因为耶和华本为善； 他的慈爱存到永远， 他的信实直到万代。
PS|101|1|我要歌唱慈爱和公平， 耶和华啊，我要向你歌颂！
PS|101|2|我要用智慧行完全的道。 你几时到我这里来呢？ 我要以纯正的心行在我家中。
PS|101|3|邪僻的事，我都不摆在我眼前； 悖逆的人所做的事，我甚恨恶， 不容沾在我身上。
PS|101|4|歪曲的心思，我必远离； 邪恶的事情，我不知道。
PS|101|5|暗中谗害他邻居的，我必将他灭绝； 眼目高傲、心里骄纵的，我必不容忍。
PS|101|6|我眼要看顾地上诚实可靠的人，使他们与我同住； 行正直路的，他要侍候我。
PS|101|7|行诡诈的，必不得住在我家里； 说谎言的，必不得立在我眼前。
PS|101|8|我每日早晨要灭绝地上所有的恶人， 把作恶的从耶和华的城里全都剪除。
PS|102|1|耶和华啊，求你听我的祷告， 愿我的呼求达到你面前！
PS|102|2|我急难的日子，求你不要转脸不顾我！ 我呼求的日子，求你向我侧耳，快快应允我！
PS|102|3|因为我的年日在烟中消失 ， 我的骨头如火把烧着。
PS|102|4|我的心如草被踩碎而枯干， 甚至我忘记吃饭。
PS|102|5|因我叹息的声音， 我的肉紧贴骨头。
PS|102|6|我如同旷野的鹈鹕， 好像荒地的猫头鹰。
PS|102|7|我清醒难以入眠， 如同房顶上孤单的麻雀。
PS|102|8|我的仇敌整日辱骂我， 向我叫号的人指着我赌咒。
PS|102|9|我吃灰烬如同吃饭， 我喝的有眼泪搀杂。
PS|102|10|这都因你的恼恨和愤怒， 你把我举起，又把我摔下。
PS|102|11|我的年日如夕阳， 我也如草枯干。
PS|102|12|惟你－耶和华必永远坐在宝座上， 你的名 存到万代。
PS|102|13|你必起来怜悯 锡安 ； 因现在是可怜它的时候， 因所定的日期已经到了。
PS|102|14|你的仆人们喜爱 锡安 的石头， 怜悯它的尘土。
PS|102|15|列国要敬畏耶和华的名， 地上众王都要敬畏你的荣耀。
PS|102|16|因为耶和华建造了 锡安 ， 在他的荣耀里显现。
PS|102|17|他垂听穷乏人的祷告， 不藐视他们的祈求。
PS|102|18|这必为后代的人记下， 将来受造的百姓要赞美耶和华。
PS|102|19|因为他从至高的圣所垂看； 耶和华从天向地观看，
PS|102|20|要垂听被囚之人的叹息， 要释放将死的人，
PS|102|21|使人在 锡安 传扬耶和华的名， 在 耶路撒冷 传扬赞美他的话，
PS|102|22|就是在万民和列国 聚集事奉耶和华的时候。
PS|102|23|他使我的力量半途衰弱， 使我的年日短少。
PS|102|24|我说：“我的上帝啊， 不要使我中年去世。 你的年数世世无穷！”
PS|102|25|你起初立了地的根基， 天也是你手所造的。
PS|102|26|天地都会消灭，你却长存； 天地都会像外衣渐渐旧了。 你要将天地如内衣更换， 天地就都改变了。
PS|102|27|惟有你永不改变， 你的年数没有穷尽。
PS|102|28|你仆人的子孙要安然居住， 他们的后裔要坚立在你面前。
PS|103|1|我的心哪，你要称颂耶和华！ 凡在我里面的，都要称颂他的圣名！
PS|103|2|我的心哪，你要称颂耶和华！ 不可忘记他一切的恩惠！
PS|103|3|他赦免你一切的罪孽， 医治你一切的疾病。
PS|103|4|他救赎你的命脱离地府， 以仁爱和怜悯为你的冠冕。
PS|103|5|他用美物使你的生命 得以满足， 以致你如鹰返老还童。
PS|103|6|耶和华施行公义， 为所有受欺压的人伸冤。
PS|103|7|他使 摩西 知道他的法则， 使 以色列 人晓得他的作为。
PS|103|8|耶和华有怜悯，有恩惠， 不轻易发怒，且有丰盛的慈爱。
PS|103|9|他不长久责备， 也不永远怀怒。
PS|103|10|他没有按我们的罪待我们， 也没有照我们的罪孽报应我们。
PS|103|11|天离地何等的高， 他的慈爱向敬畏他的人也是何等的大！
PS|103|12|东离西有多远， 他叫我们的过犯离我们也有多远！
PS|103|13|父亲怎样怜悯他的儿女， 耶和华也怎样怜悯敬畏他的人！
PS|103|14|因为他知道我们的本体， 思念我们不过是尘土。
PS|103|15|至于世人，他的年日如草一样。 他兴旺如野地的花，
PS|103|16|经风一吹，就归无有， 它的原处也不再认识它。
PS|103|17|但耶和华的慈爱归于敬畏他的人， 从亘古到永远； 他的公义也归于子子孙孙，
PS|103|18|就是那些遵守他的约、 记念他的训词而遵行的人。
PS|103|19|耶和华在天上立定宝座， 他的国统管万有。
PS|103|20|听从他命令、成全他旨意、 有大能的天使啊，你们都要称颂耶和华！
PS|103|21|你们行他所喜悦的， 作他诸军，作他仆役的啊，都要称颂耶和华！
PS|103|22|你们一切被他造的， 在他所治理的各处， 都要称颂耶和华！ 我的心哪，你要称颂耶和华！
PS|104|1|我的心哪，你要称颂耶和华！ 耶和华－我的上帝啊，你为至大！ 你以尊荣威严为衣，
PS|104|2|披上亮光，如披外袍， 铺张穹苍，如铺幔子，
PS|104|3|在水中立楼阁的栋梁， 用云彩为车辇， 藉着风的翅膀而行，
PS|104|4|以风为使者， 以火焰为仆役，
PS|104|5|将地立在根基上， 使地永不动摇。
PS|104|6|你用深水遮盖地面，犹如衣裳； 诸水高过山岭。
PS|104|7|你的斥责一发，水就奔逃； 你的雷声一发，水就奔流。
PS|104|8|诸山上升，诸谷下沉， 归你为它所立定之地。
PS|104|9|你定了界限，使水不能超越， 不再转回淹没大地。
PS|104|10|耶和华使泉源涌在山谷， 流在山间，
PS|104|11|使野地的走兽有水喝， 野驴得解其渴。
PS|104|12|天上的飞鸟在水旁住宿， 在枝干间啼叫。
PS|104|13|他从楼阁中浇灌山岭； 因他作为的功效，地就丰足。
PS|104|14|他使草生长，给牲畜吃， 使菜蔬生长，供给人用 ， 使人从地里得食物，
PS|104|15|得酒能悦人心， 得油能润人面， 得粮能养人心。
PS|104|16|佳美的树木， 就是耶和华所栽种的 黎巴嫩 的香柏树， 都满了汁浆。
PS|104|17|雀鸟在其上搭窝， 鹳以松树 为家。
PS|104|18|高山为野山羊的居所， 岩石为石的藏身处。
PS|104|19|你安置月亮以定季节， 太阳自知沉落。
PS|104|20|你造黑暗为夜， 林中的百兽就都爬出来。
PS|104|21|少壮狮子吼叫觅食， 向上帝寻求食物。
PS|104|22|太阳一出，兽就躲避， 躺卧在洞里。
PS|104|23|人出去做工， 劳碌直到晚上。
PS|104|24|耶和华啊，你所造的何其多！ 都是你用智慧造成的， 全地遍满了你所造之物。
PS|104|25|那里有海，又大又广， 其中有无数的动物， 大小活物都有。
PS|104|26|那里有船行走， 有你所造的 力威亚探 悠游在其中。
PS|104|27|这些都仰望你按时给它们食物。
PS|104|28|你给它们，它们就拾起来； 你张手，它们就饱得美食。
PS|104|29|你转脸，它们就惊惶； 你收回它们的气，它们就死亡，归于尘土。
PS|104|30|你差遣你的灵，它们就受造； 你使地面更换为新。
PS|104|31|愿耶和华的荣耀存到永远！ 愿耶和华喜爱自己所造的！
PS|104|32|他看地，地便震动； 他摸山，山就冒烟。
PS|104|33|我一生要向耶和华唱诗！ 我还活的时候，要向我的上帝歌颂！
PS|104|34|愿他悦纳我的默念！ 我要因耶和华欢喜！
PS|104|35|愿罪人从世上消灭！ 愿恶人归于无有！ 我的心哪，你要称颂耶和华！ 哈利路亚 ！
PS|105|1|你们要称谢耶和华，求告他的名， 在万民中传扬他的作为！
PS|105|2|要向他唱诗，向他歌颂， 述说他一切奇妙的作为！
PS|105|3|要夸耀他的圣名！ 愿寻求耶和华的人心中欢喜！
PS|105|4|要寻求耶和华与他的能力， 时常寻求他的面。
PS|105|5|他仆人 亚伯拉罕 的后裔， 他所拣选 雅各 的子孙哪， 要记念他奇妙的作为和他的奇事， 并他口中的判语。
PS|105|6|
PS|105|7|他是耶和华－我们的上帝， 全地都有他的判断。
PS|105|8|他记念他的约，直到永远； 记念他吩咐的话，直到千代，
PS|105|9|就是与 亚伯拉罕 所立的约， 向 以撒 所起的誓。
PS|105|10|他将这约向 雅各 定为律例， 向 以色列 定为永远的约，
PS|105|11|说：“我必将 迦南 地赐给你， 作你们应得的产业。”
PS|105|12|当时，他们人丁有限， 数目稀少，在那地寄居。
PS|105|13|他们从这邦游到那邦， 从这国去到另一民族。
PS|105|14|他不容人欺负他们， 为他们的缘故责备君王：
PS|105|15|“不可伤害我的受膏者， 也不可恶待我的先知。”
PS|105|16|他命饥荒降在那地， 断绝日用的粮食 ，
PS|105|17|在他们以先差遣一个人前往， 约瑟 被卖为奴。
PS|105|18|人用脚镣伤他的脚， 他被铁的项链捆锁。
PS|105|19|耶和华的话试炼他， 直等所说的应验了。
PS|105|20|王差人将他解开， 治理万民的把他释放，
PS|105|21|立他为王家之主， 掌管他一切所有的，
PS|105|22|使他随意捆绑他的臣宰， 将智慧教导他的长老。
PS|105|23|以色列 也到了 埃及 ， 雅各 在 含 地寄居。
PS|105|24|耶和华使他的百姓生养众多， 使他们比敌人强盛，
PS|105|25|他使敌人的心转去恨他的百姓， 用诡计待他的仆人。
PS|105|26|他差遣他的仆人 摩西 和他所拣选的 亚伦 ，
PS|105|27|在敌人中间显他的神迹， 在 含 地显他的奇事。
PS|105|28|他差遣黑暗，就有黑暗； 他们没有违背他的话。
PS|105|29|他使 埃及 的水变为血， 令他们的鱼死了。
PS|105|30|在他们的地上，青蛙多多滋生， 王宫的内室也是如此。
PS|105|31|他一吩咐，苍蝇就成群飞来， 并有蚊子进入他们四境。
PS|105|32|他给他们降下冰雹为雨， 在他们的地上降下火焰。
PS|105|33|他击打他们的葡萄树和无花果树， 毁坏他们境内的树木。
PS|105|34|他一吩咐，就有蝗虫蝻子上来， 不计其数，
PS|105|35|吃光他们地上各样的菜蔬， 吞尽他们田地的出产。
PS|105|36|他又击杀他们国内 所有的长子， 就是他们强壮时头生的。
PS|105|37|他却带领自己的百姓带着金子银子出来， 他支派中没有一个走不动的。
PS|105|38|他们出来的时候， 埃及 人就欢喜； 因为 埃及 人惧怕他们。
PS|105|39|他铺张云彩当遮蔽， 夜间使火光照。
PS|105|40|他们祈求，他就使鹌鹑飞来， 并用天上的粮食使他们饱足。
PS|105|41|他敲开磐石，水就涌出； 在干旱之处，水流成河。
PS|105|42|这都因他记念他的圣言 和他的仆人 亚伯拉罕 。
PS|105|43|他带领自己的百姓欢乐而出， 带领自己的选民欢呼前往。
PS|105|44|他把列国的地赐给他们， 他们就承受万民劳碌得来的，
PS|105|45|好让他们遵他的律例， 守他的律法。 哈利路亚！
PS|106|1|哈利路亚！ 你们要称谢耶和华，因他本为善， 他的慈爱永远长存！
PS|106|2|谁能传扬耶和华的大能？ 谁能表明他一切的美德？
PS|106|3|凡遵守公平、常行公义的， 这人有福了！
PS|106|4|耶和华啊，你恩待你百姓的时候，求你记念我； 你拯救他们的时候，求你眷顾我，
PS|106|5|好使我经历你选民的福分， 享受你国民的喜乐， 与你的产业一同夸耀。
PS|106|6|我们与我们的祖宗一同犯罪， 偏邪行恶。
PS|106|7|我们的祖宗在 埃及 不明白你的奇事， 不记念你丰盛的慈爱， 反倒在 红海 行了悖逆。
PS|106|8|然而，他因自己的名拯救他们， 为要彰显他的大能。
PS|106|9|他斥责 红海 ，海就干了， 带领他们走过深海，如走旷野。
PS|106|10|他拯救他们脱离恨他们之人的手， 从仇敌手中救赎他们。
PS|106|11|水淹没他们的敌人， 没有一个存留。
PS|106|12|那时，他们才信他的话， 歌唱赞美他。
PS|106|13|很快地，他们就忘了他的作为， 不仰望他的指引，
PS|106|14|反倒在旷野起了贪婪之心， 在荒地试探上帝。
PS|106|15|他将他们所求的赐给他们， 却使他们心灵软弱。
PS|106|16|他们在营中嫉妒 摩西 和耶和华的圣者 亚伦 。
PS|106|17|地就裂开，吞下 大坍 ， 掩盖 亚比兰 一伙的人。
PS|106|18|有火在他们党中点燃， 有火焰烧毁了恶人。
PS|106|19|他们在 何烈山 造了牛犊， 叩拜铸成的像，
PS|106|20|将他们荣耀的主 换为吃草之牛的像，
PS|106|21|忘了上帝－他们的救主， 就是曾在 埃及 行大事，
PS|106|22|在 含 地行奇事， 在 红海 行可畏之事的那位。
PS|106|23|因此，他说要灭绝他们； 若非他所拣选的 摩西 在他面前站在破裂之处， 使他的愤怒转消， 恐怕他就灭绝他们了。
PS|106|24|他们又藐视那美地， 不信他的话，
PS|106|25|在自己帐棚内发怨言， 不听耶和华的声音。
PS|106|26|所以他向他们起誓， 必叫他们倒在旷野，
PS|106|27|叫他们的后裔倒在列国之中， 分散在各地。
PS|106|28|他们又与 巴力．毗珥 连合， 吃了祭死人的物。
PS|106|29|他们这样行，惹耶和华发怒， 就有瘟疫流行在他们中间。
PS|106|30|那时， 非尼哈 起而干预， 瘟疫这才止息。
PS|106|31|那就算他为义， 世世代代，直到永远。
PS|106|32|他们在 米利巴 水又惹耶和华发怒， 甚至 摩西 也因他们的缘故受亏损，
PS|106|33|是因他们触怒了他的灵， 摩西就用嘴说了急躁的话。
PS|106|34|他们不照耶和华所吩咐的 灭绝外邦人，
PS|106|35|反倒与列国相交， 学习他们的行为，
PS|106|36|事奉他们的偶像， 这就成了自己的圈套。
PS|106|37|他们把自己的儿女祭祀鬼魔，
PS|106|38|流无辜人的血， 就是自己儿女的血， 用他们祭祀 迦南 的偶像， 那地就被血玷污了。
PS|106|39|这样，他们被自己所做的玷污了， 在行为上犯了淫乱。
PS|106|40|耶和华的怒气向他的百姓发作， 他憎恶自己的产业，
PS|106|41|将他们交在外邦人手里， 恨他们的人就辖制他们。
PS|106|42|他们的仇敌欺压他们， 他们伏在敌人手下。
PS|106|43|他屡次搭救他们， 他们却图谋悖逆， 就因自己的罪孽降为卑下。
PS|106|44|然而，他听见他们哀告的时候， 就眷顾他们的急难，
PS|106|45|为了他们，他记念自己的约， 照他丰盛的慈爱改变心意，
PS|106|46|使他们在凡掳掠他们的人面前蒙怜悯。
PS|106|47|耶和华－我们的上帝啊，求你拯救我们， 从列国中召集我们， 我们好颂扬你的圣名， 以赞美你为夸胜。
PS|106|48|耶和华－ 以色列 的上帝是应当称颂的， 从亘古直到永远。 愿全体百姓都说：“阿们！” 哈利路亚！
PS|107|1|你们要称谢耶和华，因他本为善， 他的慈爱永远长存！
PS|107|2|愿耶和华救赎的百姓说这话， 就是他从敌人手中所救赎，
PS|107|3|从各地，从东从西， 从北从海那边召集来的。
PS|107|4|他们在旷野、在荒地飘流， 找不到可居住的城，
PS|107|5|又饥又渴， 心里发昏。
PS|107|6|于是他们在急难中哀求耶和华， 他就搭救他们脱离祸患，
PS|107|7|又领他们行走直路， 前往可居住的城。
PS|107|8|但愿人因耶和华的慈爱 和他向人所做的奇事都称谢他；
PS|107|9|因他使心里渴慕的人得以满足， 使饥饿的人得饱美食。
PS|107|10|那些坐在黑暗中、死荫里的人， 被困苦和铁链捆锁，
PS|107|11|是因他们违背上帝的言语， 藐视至高者的旨意。
PS|107|12|所以，他用劳苦制伏他们的心； 他们仆倒，无人扶助。
PS|107|13|于是他们在急难中哀求耶和华， 他就拯救他们脱离祸患。
PS|107|14|他从黑暗中、从死荫里领他们出来， 扯断他们的捆绑。
PS|107|15|但愿人因耶和华的慈爱 和他向人所做的奇事都称谢他；
PS|107|16|因为他打破了铜门， 砍断了铁闩。
PS|107|17|愚妄人因自己叛逆的行径 和自己的罪孽受苦楚。
PS|107|18|他们心里厌恶各样的食物， 就临近死亡之门。
PS|107|19|于是他们在急难中哀求耶和华， 他就拯救他们脱离祸患。
PS|107|20|他发出自己的话语医治他们， 救他们脱离阴府。
PS|107|21|但愿人因耶和华的慈爱 和他向人所做的奇事都称谢他。
PS|107|22|愿他们以感谢为祭献给他， 欢呼述说他的作为！
PS|107|23|那些搭船出海， 在大水中做生意的，
PS|107|24|他们看见耶和华的作为， 并他在深海中的奇事。
PS|107|25|他一出令，狂风卷起， 波浪翻腾。
PS|107|26|他们上到天空，下到海底， 他们的心因患难而消沉。
PS|107|27|他们摇摇晃晃，东倒西歪，好像醉酒的人， 他们的智慧无法可施。
PS|107|28|于是他们在急难中哀求耶和华， 他就领他们脱离祸患。
PS|107|29|他使狂风止息， 波浪平静，
PS|107|30|既平静了，他们就欢喜， 他就领他们到想要去的海港。
PS|107|31|但愿人因耶和华的慈爱 和他向人所做的奇事都称谢他。
PS|107|32|愿他们在百姓的会中尊崇他， 在长老的座位上赞美他！
PS|107|33|他使江河变为旷野， 叫水泉变为干涸之地，
PS|107|34|使肥沃之地变为荒芜的盐地， 都因当地居民的邪恶。
PS|107|35|他使旷野变为水潭， 叫旱地变为水泉，
PS|107|36|使饥饿的人住在那里， 建造可居住的城，
PS|107|37|又种田地，栽葡萄园， 得享所出产的果实。
PS|107|38|他赐福给他们，使他们生养众多， 也不叫他们的牲畜减少。
PS|107|39|但他们因欺压、患难、愁苦， 人口减少而且卑微。
PS|107|40|他使贵族蒙羞受辱， 使他们迷失在荒凉无路之地；
PS|107|41|却将穷乏人安置在高处，脱离苦难， 使他的家属多如羊群。
PS|107|42|正直的人看见就欢喜， 罪孽之辈却要哑口无言。
PS|107|43|凡有智慧的必在这些事上留心， 他必思想耶和华的慈爱。
PS|108|1|上帝啊，我心坚定； 我口 要唱诗歌颂！
PS|108|2|琴瑟啊，当醒起！ 我要唤起曙光！
PS|108|3|耶和华啊，我要在万民中称谢你， 在万族中歌颂你！
PS|108|4|因为你的慈爱大过诸天， 你的信实达到穹苍。
PS|108|5|上帝啊，愿你崇高过于诸天！ 愿你的荣耀高过全地！
PS|108|6|求你应允我，用右手施行拯救， 好让你所亲爱的人得救。
PS|108|7|上帝在他的圣所 说： “我要欢乐； 要划分 示剑 ， 丈量 疏割谷 。
PS|108|8|基列 是我的， 玛拿西 是我的， 以法莲 是护卫我头的， 犹大 是我的权杖。
PS|108|9|摩押 是我的沐浴盆， 我要向 以东 扔鞋， 我必因胜 非利士 而欢呼。”
PS|108|10|谁能领我进坚固城？ 谁能引我到 以东 地？
PS|108|11|上帝啊，你真的丢弃了我们吗？ 上帝啊，你不和我们的军队同去吗？
PS|108|12|求你帮助我们攻击敌人， 因为人的帮助是枉然的。
PS|108|13|我们倚靠上帝才得施展大能， 因为践踏我们敌人的就是他。
PS|109|1|我所赞美的上帝啊， 求你不要闭口不言。
PS|109|2|因为恶人的嘴和诡诈人的口张开攻击我， 他们用撒谎的舌头对我说话。
PS|109|3|他们围绕我，说怨恨的话， 又无故地攻打我。
PS|109|4|他们与我作对回报我的爱， 但我专心祈祷。
PS|109|5|他们向我以恶报善， 以恨报爱。
PS|109|6|求你派恶人辖制他， 派对头站在他右边！
PS|109|7|他受审判的时候， 愿他背负罪名而出！ 愿他的祈祷反成为罪！
PS|109|8|愿他的年岁短少！ 愿别人得他的职分！
PS|109|9|愿他的儿女成为孤儿， 他的妻子成为寡妇！
PS|109|10|愿他的儿女飘流讨饭， 从荒凉之处出来求乞 ！
PS|109|11|愿债主牢笼他一切所有的！ 愿陌生人抢走他劳碌得来的！
PS|109|12|愿无人向他布施恩惠， 无人恩待他的孤儿！
PS|109|13|愿他的后人断绝， 名字被涂去，不传于下代！
PS|109|14|愿耶和华记得他祖宗的罪孽， 不涂去他母亲的罪过！
PS|109|15|愿这些罪常在耶和华面前！ 愿他们的名字 从地上除灭！
PS|109|16|因为他从未想过要施恩， 却迫害困苦贫穷的和伤心的人， 把他们处死。
PS|109|17|他爱咒骂，咒骂就临到他； 他不喜爱祝福，祝福就远离他！
PS|109|18|他拿咒骂当衣服穿上； 这咒骂就如水进到他里面， 如油进入他骨头。
PS|109|19|愿这咒骂当他遮身的衣服， 作他经常束腰的带子！
PS|109|20|这就是那些与我作对、用恶言议论我的人 从耶和华所受的报应。
PS|109|21|但是你，主－耶和华啊， 求你因你的名采取行动； 因你的慈爱美好，求你搭救我！
PS|109|22|因为我困苦贫穷， 内心受伤。
PS|109|23|我如日影偏斜而去， 如蝗虫被抖出来。
PS|109|24|我因禁食，膝盖软弱； 我身体消瘦，不再丰润。
PS|109|25|我受他们的羞辱， 他们看见我就摇头。
PS|109|26|耶和华－我的上帝啊，求你帮助我， 照你的慈爱拯救我，
PS|109|27|好让他们知道这是你的手， 是你－耶和华所做的事。
PS|109|28|任凭他们咒骂，你却要赐福； 他们几时起来就必蒙羞， 你的仆人却要欢喜。
PS|109|29|愿与我作对的人披戴羞辱！ 愿他们以自己的羞愧作外袍遮身！
PS|109|30|我要用口极力称谢耶和华， 我要在众人中间赞美他；
PS|109|31|因为他必站在贫穷人的右边， 救他脱离定他死罪的人。
PS|110|1|耶和华对我主说： “你坐在我的右边， 等我使你仇敌作你的脚凳。”
PS|110|2|耶和华必使你从 锡安 伸出你能力的权杖； 你务要在仇敌中掌权。
PS|110|3|你在圣山上 掌权的日子， 你的子民必甘心跟随 ； 从晨曦初现， 你就有清晨 的甘露。
PS|110|4|耶和华起了誓，绝不改变： “你是照着 麦基洗德 的体系永远为祭司。”
PS|110|5|在你右边的主， 当他发怒的日子，必打伤列王。
PS|110|6|他要审判列国， 尸首就布满各处； 他要痛击遍地的领袖。
PS|110|7|他要喝路旁的河水， 因此必抬起头来。
PS|111|1|哈利路亚！ 我要在正直人的大会和会众中 一心称谢耶和华。
PS|111|2|耶和华的作为本为大， 被所有喜爱的人所探寻。
PS|111|3|他所做的是尊荣和威严， 他的公义存到永远。
PS|111|4|他行了奇事，使人记念； 耶和华有恩惠，有怜悯。
PS|111|5|他赐粮食给敬畏他的人， 他必永远记念他的约。
PS|111|6|他向百姓显出大能的作为， 将列国赐给他们为业。
PS|111|7|他手所做的信实公平， 他的训词全然可靠，
PS|111|8|是永永远远坚定的， 是按信实正直设立的。
PS|111|9|他向百姓施行救赎， 颁布他的约，直到永远； 他的名圣而可畏。
PS|111|10|敬畏耶和华是智慧的开端， 凡遵行他命令的有美好的见识。 耶和华是永远当赞美的！
PS|112|1|哈利路亚！ 敬畏耶和华，甚喜爱他命令的， 这人有福了！
PS|112|2|他的后裔在世必强盛， 正直人的后代必蒙福。
PS|112|3|他的家中有金银财宝， 他的义行存到永远。
PS|112|4|正直人在黑暗中有光向他照耀， 他有恩惠，有怜悯，有公义。
PS|112|5|施恩与人、借贷与人、秉公处事的人 必享美福，
PS|112|6|他永不动摇。 义人被记念，直到永远。
PS|112|7|他不惧怕凶恶的信息， 他的心坚定，倚靠耶和华。
PS|112|8|他的心确定，总不惧怕， 直到他看见敌人遭报。
PS|112|9|他施舍，赒济贫穷， 他的义行存到永远， 他的角必被高举，大有荣耀。
PS|112|10|恶人看见就愤怒，必咬牙而消亡， 恶人的心愿要归于幻灭。
PS|113|1|哈利路亚！ 耶和华的仆人哪，你们要赞美， 赞美耶和华的名！
PS|113|2|耶和华的名是应当称颂的， 从今时直到永远！
PS|113|3|从日出之地到日落之处， 耶和华的名是应当赞美的！
PS|113|4|耶和华超乎万国之上， 他的荣耀高过诸天。
PS|113|5|谁像耶和华－我们的上帝呢？ 他坐在至高之处，
PS|113|6|自己谦卑， 观看天上地下的事。
PS|113|7|他从灰尘里抬举贫寒的人， 从粪堆中提拔贫穷的人，
PS|113|8|使他们与贵族同坐， 与本国的贵族同坐。
PS|113|9|他使不孕的妇女安居家中， 成为快乐的母亲，儿女成群。 哈利路亚！
PS|114|1|以色列 出 埃及 ， 雅各 家离开说陌生语言之民时，
PS|114|2|犹大 作主的圣所， 以色列 为他所治理的国。
PS|114|3|沧海看见就奔逃， 约旦河 也倒流。
PS|114|4|大山踊跃如公羊， 小山跳舞如羔羊。
PS|114|5|沧海啊，你为何奔逃？ 约旦 哪，你为何倒流？
PS|114|6|大山哪，你为何踊跃如公羊？ 小山哪，你为何跳舞如羔羊？
PS|114|7|大地啊，在主的面前， 在 雅各 的上帝的面前，震动吧！
PS|114|8|他叫磐石变为水池， 使坚石变为泉源。
PS|115|1|耶和华啊，荣耀不要归与我们， 不要归与我们； 要因你的慈爱和信实归在你的名下！
PS|115|2|为何让列国说 “他们的上帝在哪里”呢？
PS|115|3|但是，我们的上帝在天上， 万事都随自己的旨意而行。
PS|115|4|他们的偶像是金的，是银的， 是人手所造的，
PS|115|5|有口却不能言， 有眼却不能看，
PS|115|6|有耳却不能听， 有鼻却不能闻，
PS|115|7|有手却不能摸， 有脚却不能走， 有喉却不能说话。
PS|115|8|造它们的要像它们一样， 凡靠它们的也必如此。
PS|115|9|以色列 啊，要倚靠耶和华！ 他是人的帮助和盾牌。
PS|115|10|亚伦 家啊，要倚靠耶和华！ 他是人的帮助和盾牌。
PS|115|11|敬畏耶和华的人哪，要倚靠耶和华！ 他是人的帮助和盾牌。
PS|115|12|耶和华向来眷念我们， 他还要赐福， 赐福给 以色列 家， 赐福给 亚伦 家。
PS|115|13|凡敬畏耶和华的，无论大小， 主必赐福给他。
PS|115|14|愿耶和华使你们 和你们的子孙日见增加。
PS|115|15|你们蒙了耶和华的福， 他是创造天地的主宰。
PS|115|16|天，是耶和华的天； 地，他却给了世人。
PS|115|17|死人不能赞美耶和华， 下到寂静 中的也都不能。
PS|115|18|但我们要称颂耶和华， 从今时直到永远。 哈利路亚！
PS|116|1|我爱耶和华， 因为他听了我的声音和我的恳求。
PS|116|2|他既向我侧耳， 我一生要求告他。
PS|116|3|死亡的绳索勒住我， 阴间的痛苦抓住我， 我遭遇患难愁苦。
PS|116|4|那时，我求告耶和华的名： “耶和华啊，求你救我！”
PS|116|5|耶和华有恩惠，有公义， 我们的上帝有怜悯。
PS|116|6|耶和华保护愚蒙的人； 我落到卑微的地步，他救了我。
PS|116|7|我的心哪！你要复归安宁， 因为耶和华用厚恩待你。
PS|116|8|主啊，你救我的命脱离死亡， 使我的眼不再流泪， 使我的脚不致跌倒。
PS|116|9|我行在耶和华面前， 走在活人之地。
PS|116|10|我信，尽管我说： “我受了极大的困苦。”
PS|116|11|我曾惊惶地说： “人都是说谎的！”
PS|116|12|耶和华向我赏赐一切厚恩， 我拿什么来报答他呢？
PS|116|13|我要举起救恩的杯， 称扬耶和华的名。
PS|116|14|我要在他的全体百姓面前 向耶和华还我所许的愿。
PS|116|15|在耶和华眼中， 圣民之死极为宝贵。
PS|116|16|耶和华啊，哦，我是你的仆人； 我是你的仆人，是你使女的儿子。 你已经解开我的捆索。
PS|116|17|我要以感谢为祭献给你， 又要求告耶和华的名。
PS|116|18|我要在 耶路撒冷 当中， 在耶和华殿的院内， 在他的全体百姓面前， 向耶和华还我所许的愿。 哈利路亚！
PS|116|19|
PS|117|1|万国啊，你们要赞美耶和华！ 万族啊，你们都要颂赞他！
PS|117|2|因为他向我们大施慈爱， 耶和华的信实存到永远。 哈利路亚！
PS|118|1|你们要称谢耶和华，因他本为善； 他的慈爱永远长存！
PS|118|2|愿 以色列 说： “他的慈爱永远长存！”
PS|118|3|愿 亚伦 家说： “他的慈爱永远长存！”
PS|118|4|愿敬畏耶和华的人说： “他的慈爱永远长存！”
PS|118|5|我在急难中求告耶和华， 耶和华就应允我，把我安置在宽阔之地。
PS|118|6|耶和华在我这边 ，我必不惧怕， 人能把我怎么样呢？
PS|118|7|在那帮助我的人中，有耶和华帮助我， 所以我要看见那些恨我的人遭报。
PS|118|8|投靠耶和华， 强似倚赖人；
PS|118|9|投靠耶和华， 强似倚赖权贵。
PS|118|10|列邦围绕我， 我靠耶和华的名必剿灭他们。
PS|118|11|他们围绕我，围困我， 我靠耶和华的名必剿灭他们。
PS|118|12|他们如同蜜蜂一般地围绕我， 他们熄灭，好像烧荆棘的火； 我靠耶和华的名，必剿灭他们。
PS|118|13|你用力推我，要叫我跌倒， 但耶和华帮助了我。
PS|118|14|耶和华是我的力量，是我的诗歌， 他也成了我的拯救。
PS|118|15|在义人的帐棚里，有欢呼拯救的声音， 耶和华的右手施展大能。
PS|118|16|耶和华的右手高举， 耶和华的右手施展大能。
PS|118|17|我不至于死，仍要存活， 并要传扬耶和华的作为。
PS|118|18|耶和华虽严严地惩治我， 却未曾将我交于死亡。
PS|118|19|给我敞开义门， 我要进去称谢耶和华！
PS|118|20|这是耶和华的门， 义人要进去！
PS|118|21|我要称谢你，因为你已经应允我， 又成了我的拯救！
PS|118|22|匠人所丢弃的石头 已成了房角的头块石头。
PS|118|23|这是耶和华所做的， 在我们眼中看为奇妙。
PS|118|24|这是耶和华所定的日子， 我们在其中要高兴欢喜！
PS|118|25|耶和华啊，求你拯救 ！ 耶和华啊，求你使我们顺利！
PS|118|26|奉耶和华的名来的是应当称颂的！ 我们从耶和华的殿中为你们祝福！
PS|118|27|耶和华是上帝， 他光照了我们。 你们要用绳索把祭牲拴住， 直牵到坛角。
PS|118|28|你是我的上帝，我要称谢你！ 我的上帝啊，我要尊崇你 ！
PS|118|29|你们要称谢耶和华，因他本为善； 他的慈爱永远长存！
PS|119|1|行为正直、遵行耶和华律法的， 这人有福了！
PS|119|2|遵守他的法度、一心寻求他的， 这人有福了！
PS|119|3|他们不做不义的事， 但遵行他的道。
PS|119|4|耶和华啊，你曾将你的训词吩咐我们， 为要我们切实遵守。
PS|119|5|但愿我行事坚定， 得以遵守你的律例。
PS|119|6|我看重你的一切命令， 就不致羞愧。
PS|119|7|我学习你公义的典章， 要以正直的心称谢你。
PS|119|8|我必遵守你的律例， 求你不要把我全然弃绝！
PS|119|9|青年要如何保持纯洁呢？ 是要遵行你的话！
PS|119|10|我曾一心寻求你， 求你不要使我偏离你的命令。
PS|119|11|我将你的话藏在心里， 免得我得罪你。
PS|119|12|耶和华啊，你是应当称颂的！ 求你将你的律例教导我！
PS|119|13|我用嘴唇传扬 你口中一切的典章。
PS|119|14|我喜爱你的法度， 如同喜爱一切的财物。
PS|119|15|我要默想你的训词， 看重你的道路。
PS|119|16|我要以你的律例为乐， 我不忘记你的话。
PS|119|17|求你用厚恩待你的仆人，使我存活， 我就遵守你的话。
PS|119|18|求你开我的眼睛， 使我看出你律法中的奇妙。
PS|119|19|我在地上是寄居的人， 求你不要向我隐藏你的命令！
PS|119|20|我时常切慕你的典章， 耗尽心力。
PS|119|21|受诅咒、偏离你命令的骄傲人， 你已经责备他们。
PS|119|22|求你除掉我所受的羞辱和藐视， 因我遵守你的法度。
PS|119|23|虽有掌权者坐着妄论我， 你仆人却思想你的律例。
PS|119|24|你的法度也是我的喜乐， 我的导师 。
PS|119|25|我的性命几乎归于尘土， 求你照你的话将我救活！
PS|119|26|我述说我所做的，你应允了我； 求你将你的律例教导我！
PS|119|27|求你使我明白你的训词， 我要默想你的奇事。
PS|119|28|我因愁苦身心耗尽， 求你照你的话使我坚立！
PS|119|29|求你使我离开奸诈的道路， 开恩将你的律法赐给我！
PS|119|30|我选择了忠信的道路， 将你的典章摆在我面前。
PS|119|31|我持守你的法度； 耶和华啊，求你不要叫我羞愧！
PS|119|32|你使我心胸开阔的时候， 我就往你命令的道路直奔。
PS|119|33|耶和华啊，求你将你的律例指教我， 我必遵守到底！
PS|119|34|求你赐我悟性，我就遵守你的律法， 且要一心遵守。
PS|119|35|求你叫我遵行你的命令， 因为这是我所喜爱的。
PS|119|36|求你使我的心趋向你的法度， 不趋向不义之财。
PS|119|37|求你叫我转眼不看虚假， 使我活在你的道路 中。
PS|119|38|求你向敬畏你的仆人 坚守你的话！
PS|119|39|求你使我所惧怕的羞辱远离我， 因你的典章本为美。
PS|119|40|看哪，我切慕你的训词， 求你因你的公义赐我生命 ！
PS|119|41|耶和华啊，求你使你的慈爱临到我， 照你的话使你的救恩临到我，
PS|119|42|我就有话回答那羞辱我的， 因我倚靠你的话。
PS|119|43|求你叫真理的话总不离开我的口， 因我仰望你的典章。
PS|119|44|我要常守你的律法， 直到永永远远。
PS|119|45|我要自由而行 ， 因我寻求了你的训词。
PS|119|46|我要在列王面前宣讲你的法度， 也不致羞愧。
PS|119|47|我以你的命令为乐， 这命令是我所喜爱的。
PS|119|48|我向我所爱的，就是你的命令高举双手 ， 我也要默想你的律例。
PS|119|49|求你记念你向仆人所说的话， 这话使我有盼望。
PS|119|50|你的话将我救活了； 这是我在患难中的安慰。
PS|119|51|骄傲的人极度地侮慢我， 我却未曾偏离你的律法。
PS|119|52|耶和华啊，我记念你从古以来的典章， 就得了安慰。
PS|119|53|我因恶人离弃你的律法， 怒火中烧。
PS|119|54|我在世寄居， 以你的律例为诗歌。
PS|119|55|耶和华啊，我夜间记念你的名， 我也要遵守你的律法。
PS|119|56|这临到我， 是因我谨守你的训词。
PS|119|57|耶和华是我的福分； 我曾说，我要遵守你的话。
PS|119|58|我一心恳求你的面， 求你照你的话怜悯我！
PS|119|59|我思想自己所行的道路， 我的脚步就转向你的法度。
PS|119|60|我速速遵守你的命令， 并不迟延。
PS|119|61|恶人的绳索缠绕我， 我却没有忘记你的律法。
PS|119|62|我因你公义的典章， 夜半起来称谢你。
PS|119|63|凡敬畏你、守你训词的人， 我都与他作伴。
PS|119|64|耶和华啊，遍地满了你的慈爱； 求你将你的律例教导我！
PS|119|65|耶和华啊，你照你的话， 善待你的仆人。
PS|119|66|求你教我明辨和知识， 因我信靠你的命令。
PS|119|67|我未受苦以先曾经迷失， 现在却遵守你的话。
PS|119|68|你本为善，所行的也善； 求你将你的律例教导我！
PS|119|69|骄傲的人编造谎言攻击我， 我却要一心遵守你的训词。
PS|119|70|他们的心蒙昧如蒙油脂， 我却喜爱你的律法。
PS|119|71|我受苦是与我有益， 为要使我学习你的律例。
PS|119|72|你口中的律法与我有益， 胜于千万金银。
PS|119|73|你的手造了我，塑造我； 求你赐我悟性学习你的命令！
PS|119|74|敬畏你的人看见我就欢喜， 因我仰望你的话。
PS|119|75|耶和华啊，我知道你的典章是公义的； 你使我受苦是以信实待我。
PS|119|76|求你照着你向仆人所说的话， 以慈爱安慰我。
PS|119|77|求你的怜悯临到我，使我存活， 因你的律法是我的喜乐。
PS|119|78|愿骄傲的人蒙羞，因为他们无理倾覆我； 但我要默想你的训词。
PS|119|79|愿敬畏你的人和知道你法度的人 都归向我。
PS|119|80|愿我的心在你的律例上完全， 使我不致蒙羞。
PS|119|81|我渴想你的救恩身心耗尽， 我仰望你的话。
PS|119|82|我因渴望你的话眼睛失明，说： “你何时安慰我呢？”
PS|119|83|我虽像烟薰的皮囊， 却不忘记你的律例。
PS|119|84|你仆人的年日有多少呢？ 你几时向迫害我的人施行审判呢？
PS|119|85|不顺从你律法的骄傲人 为我掘了坑。
PS|119|86|你的命令尽都信实； 他们无理迫害我，求你帮助我！
PS|119|87|他们几乎把我从世上除灭； 但我没有离弃你的训词。
PS|119|88|求你照你的慈爱将我救活， 我就遵守你口中的法度。
PS|119|89|耶和华啊，你的话安定在天， 直到永远。
PS|119|90|你的信实存到万代； 你坚立了地，地就长存。
PS|119|91|天地照你的典章存到今日； 万物都是你的仆役。
PS|119|92|我若不以你的律法为乐， 早就在苦难中灭绝了！
PS|119|93|我永不忘记你的训词， 因你用这训词将我救活。
PS|119|94|我是属你的，求你救我， 因我寻求了你的训词。
PS|119|95|恶人等着要灭绝我， 我却要揣摩你的法度。
PS|119|96|我看万事尽都有限， 惟有你的命令极其宽广。
PS|119|97|我何等爱慕你的律法， 终日不住地思想。
PS|119|98|你的命令常存在我心里， 使我比仇敌有智慧。
PS|119|99|我比我的教师更通达， 因我思想你的法度。
PS|119|100|我比年老的更明白， 因我谨守你的训词。
PS|119|101|我阻止我的脚走一切邪路， 为要遵守你的话。
PS|119|102|我没有偏离你的典章， 因为你教导了我。
PS|119|103|你的言语在我上膛何等甘美， 在我口中比蜜更甜！
PS|119|104|我藉着你的训词得以明白， 因此，我恨恶一切虚假的行径。
PS|119|105|你的话是我脚前的灯， 是我路上的光。
PS|119|106|你公义的典章，我曾起誓遵守， 我必按着誓言而行。
PS|119|107|我极其痛苦； 耶和华啊，求你照你的话将我救活！
PS|119|108|耶和华啊，求你悦纳我口中的赞美为甘心祭， 又将你的典章教导我！
PS|119|109|我的性命常在我手掌中 ， 我却不忘记你的律法。
PS|119|110|恶人为我设下罗网， 我却没有偏离你的训词。
PS|119|111|我以你的法度为永远的产业， 因这是我心中所喜爱的。
PS|119|112|我的心倾向你的律例， 谨守到底，直到永远。
PS|119|113|心怀二意的人为我所恨； 但你的律法为我所爱。
PS|119|114|你是我藏身之处，是我的盾牌； 我仰望你的话。
PS|119|115|作恶的人哪，你们离开我吧！ 我要遵守我上帝的命令。
PS|119|116|求你照你的话扶持我，使我存活， 不要叫我因失望而蒙羞。
PS|119|117|求你扶持我，使我得救， 时常看重你的律例。
PS|119|118|凡偏离你律例的人，你都轻看他们， 因为他们的诡诈必归虚空。
PS|119|119|你除掉地上所有的恶人，好像除掉渣滓 ； 因此我喜爱你的法度。
PS|119|120|我因惧怕你，肉体战栗； 我害怕你的典章。
PS|119|121|我行公平和公义， 求你不要撇下我，交给欺压我的人！
PS|119|122|求你保证你的仆人得福， 不容骄傲的人欺压我！
PS|119|123|我因盼望你的救恩 和你公义的言语眼睛失明。
PS|119|124|求你照你的慈爱待仆人， 将你的律例教导我。
PS|119|125|我是你的仆人，求你赐我悟性， 得以认识你的法度。
PS|119|126|这是耶和华采取行动的时候， 因人废弃了你的律法。
PS|119|127|所以，我喜爱你的命令胜于金子， 更胜于纯金。
PS|119|128|你的一切训词，在万事上我都以为正直； 我恨恶一切虚假的行径。
PS|119|129|你的法度奇妙， 所以我一心谨守。
PS|119|130|你的话一开启就发出亮光， 使愚蒙人通达。
PS|119|131|我大大张口，呼吸急促， 因我切慕你的命令。
PS|119|132|求你转向我，怜悯我， 就像你待那些喜爱你名的人。
PS|119|133|求你用你的言语使我脚步稳健， 不容罪孽辖制我。
PS|119|134|求你救我脱离人的欺压， 我要遵守你的训词。
PS|119|135|求你使你的脸向仆人发光， 又将你的律例教导我。
PS|119|136|我的眼睛流泪成河， 因为他们不守你的律法。
PS|119|137|耶和华啊，你是公义的； 你的典章正直！
PS|119|138|你所颁布的法度是公义的， 极其可靠。
PS|119|139|我的狂热把我烧灭， 因我敌人忘记你的话。
PS|119|140|你的言语极其精炼， 令你仆人喜爱。
PS|119|141|我渺小，被人藐视， 却不忘记你的训词。
PS|119|142|你的公义永远公义， 你的律法是确实的。
PS|119|143|我遭遇患难愁苦， 你的命令是我的喜乐。
PS|119|144|你的法度永远公义； 求你赐我悟性，使我存活。
PS|119|145|耶和华啊，我一心呼求你，求你应允我！ 我必谨守你的律例。
PS|119|146|我向你呼求，求你救我！ 我要遵守你的法度。
PS|119|147|天尚未亮我呼喊求救， 我仰望你的话。
PS|119|148|我终夜双眼睁开， 为要思想你的言语。
PS|119|149|求你按你的慈爱听我的声音， 耶和华啊，求你照你的典章将我救活！
PS|119|150|追逐奸恶的人 迫近了， 他们远离你的律法。
PS|119|151|耶和华啊，你就在我身边， 你一切的命令是确实的！
PS|119|152|我从你的法度早已知道， 这法度是你永远立定的。
PS|119|153|求你看顾我的苦难，搭救我， 因我不忘记你的律法。
PS|119|154|求你为我的冤屈辩护，救赎我， 照你的言语将我救活。
PS|119|155|救恩远离恶人， 因为他们不寻求你的律例。
PS|119|156|耶和华啊，你的怜悯本为大； 求你照你的典章将我救活。
PS|119|157|迫害我的、抵挡我的甚多， 我却没有偏离你的法度。
PS|119|158|我看见奸恶的人就憎恶， 因为他们不遵守你的言语。
PS|119|159|你看我何等喜爱你的训词！ 耶和华啊，求你按你的慈爱将我救活！
PS|119|160|你话语的精髓是真实的， 你一切公义的典章永远长存。
PS|119|161|掌权者无故迫害我， 然而我的心畏惧你的话。
PS|119|162|我喜爱你的言语， 好像人得到许多战利品。
PS|119|163|我恨恶，憎恶虚假； 惟喜爱你的律法。
PS|119|164|我因你公义的典章 一天七次赞美你。
PS|119|165|喜爱你律法的人大有平安， 任何事都不能使他们跌倒。
PS|119|166|耶和华啊，我仰望你的救恩， 遵行你的命令。
PS|119|167|我心谨守你的法度， 这法度我极其喜爱。
PS|119|168|我遵守你的训词和法度， 因我所行的道路都在你的面前。
PS|119|169|耶和华啊，愿我的呼求达到你面前， 求你照你的话赐我悟性。
PS|119|170|愿我的恳求达到你面前， 求你照你的言语搭救我。
PS|119|171|愿我的嘴唇发出赞美， 因为你将律例教导我。
PS|119|172|愿我的舌头歌唱你的言语， 因你一切的命令尽都公义。
PS|119|173|求你用你的手帮助我， 因我选择你的训词。
PS|119|174|耶和华啊，我切慕你的救恩！ 你的律法是我的喜乐。
PS|119|175|愿我的性命存活，得以赞美你！ 愿你的典章帮助我！
PS|119|176|我走迷了路如同失丧的羊，求你寻找你的仆人， 因我不忘记你的命令。
PS|120|1|我在急难中求告耶和华， 他就应允我。
PS|120|2|耶和华啊，求你救我脱离 说谎的嘴唇和诡诈的舌头！
PS|120|3|诡诈的舌头啊，他会给你什么呢？ 会加给你什么呢？
PS|120|4|就是勇士的利箭、 罗腾木 的炭火。
PS|120|5|祸哉！我寄居在 米设 ， 住在 基达 帐棚之中。
PS|120|6|我与那恨恶和平的人 许久同住。
PS|120|7|我愿和平， 当我发言，他们却要战争。
PS|121|1|我要向山举目， 我的帮助从何而来？
PS|121|2|我的帮助 从造天地的耶和华而来。
PS|121|3|他不叫你的脚摇动， 保护你的必不打盹！
PS|121|4|保护 以色列 的 必不打盹，也不睡觉。
PS|121|5|保护你的是耶和华， 耶和华在你右边荫庇你。
PS|121|6|白日，太阳必不伤你； 夜间，月亮也不害你。
PS|121|7|耶和华要保护你，免受一切的灾害， 他要保护你的性命。
PS|121|8|你出你入，耶和华要保护你， 从今时直到永远。
PS|122|1|我喜乐， 因人对我说：“我们到耶和华的殿去。”
PS|122|2|耶路撒冷 啊， 我们的脚站在你门内。
PS|122|3|耶路撒冷 被建造， 如同连结整齐的一座城。
PS|122|4|众支派就是耶和华的支派，上那里去， 按 以色列 的法度颂扬耶和华的名。
PS|122|5|他们在那里设立审判的宝座， 就是 大卫 家的宝座。
PS|122|6|你们要为 耶路撒冷 求平安： “愿爱你的人兴旺！
PS|122|7|愿你城中有平安！ 愿你宫内得平静！”
PS|122|8|为我弟兄和同伴的缘故，我要说： “愿你平安！”
PS|122|9|为耶和华－我们上帝殿的缘故， 我要为你求福！
PS|123|1|坐在天上的主啊， 我向你举目。
PS|123|2|看哪，仆人的眼睛怎样仰望主人的手， 婢女的眼睛怎样仰望女主人的手， 我们的眼睛也照样仰望耶和华－我们的上帝， 直到他怜悯我们。
PS|123|3|耶和华啊，求你怜悯我们，怜悯我们！ 因为我们受尽了藐视。
PS|123|4|我们受尽了安逸人的讥诮 和骄傲人的藐视。
PS|124|1|说吧， 以色列 ： “若不是耶和华帮助我们，
PS|124|2|若不是耶和华帮助我们， 当人起来攻击我们，
PS|124|3|那时，人向我们发怒， 就把我们活活吞了；
PS|124|4|那时，波涛必漫过我们， 河水必淹没我们；
PS|124|5|那时，狂傲的水 必淹没我们。”
PS|124|6|耶和华是应当称颂的！ 他没有把我们交给他们，作牙齿的猎物。
PS|124|7|我们好像雀鸟，从捕鸟人的罗网里逃脱， 罗网破裂，我们就逃脱了。
PS|124|8|我们得帮助， 是因造天地之耶和华的名。
PS|125|1|倚靠耶和华的人好像 锡安山 ， 安稳坐镇，永不动摇。
PS|125|2|众山怎样围绕 耶路撒冷 ， 耶和华也照样围绕他的百姓，从今时直到永远。
PS|125|3|恶人的杖必不在义人的土地上停留， 免得义人伸手作恶。
PS|125|4|耶和华啊，求你善待 行善和心里正直的人。
PS|125|5|至于那偏行弯曲道路的人， 耶和华必将他们和作恶的人一同驱逐出去。 愿平安归于 以色列 ！
PS|126|1|当耶和华使 锡安 被掳的人归回的时候， 我们好像做梦的人。
PS|126|2|那时，我们满口喜笑、 满舌欢呼； 那时，列国中就有人说： “耶和华为他们行了大事！”
PS|126|3|耶和华果然为我们行了大事， 我们就欢喜。
PS|126|4|耶和华啊，求你使我们这些被掳的人归回， 好像 尼革夫 的河水复流。
PS|126|5|流泪撒种的， 必欢呼收割！
PS|126|6|那带种流泪出去的， 必欢呼地带禾捆回来！
PS|127|1|若不是耶和华建造房屋， 建造的人就枉然劳力； 若不是耶和华看守城池， 看守的人就枉然警醒。
PS|127|2|你们清晨早起，夜晚安歇， 吃劳碌得来的饭，本是枉然； 惟有耶和华所亲爱的， 必叫他安然睡觉。
PS|127|3|看哪，儿女是耶和华所赐的产业， 所怀的胎是他所给的赏赐。
PS|127|4|人在年轻时生的儿女 好像勇士手中的箭。
PS|127|5|箭袋充满的人有福了！ 他们在城门口和仇敌争论时必不蒙羞。
PS|128|1|凡敬畏耶和华、 遵行他道的人有福了！
PS|128|2|你要吃劳碌得来的； 你要享福，凡事顺利。
PS|128|3|你妻子在你内室，好像多结果子的葡萄树； 你儿女围绕你的桌子，如同橄榄树苗。
PS|128|4|看哪，敬畏耶和华的人 必要这样蒙福！
PS|128|5|愿耶和华从 锡安 赐福给你！ 愿你一生一世看见 耶路撒冷 兴旺！
PS|128|6|愿你看见 你的子子孙孙！ 愿平安归于 以色列 ！
PS|129|1|说吧， 以色列 ： “从我幼年以来，人屡次苦害我；
PS|129|2|从我幼年以来，人屡次苦害我， 却没有胜过我。
PS|129|3|扶犁的人在我背上扶犁而耕， 耕的犁沟很长。”
PS|129|4|耶和华是公义的， 他砍断了恶人的绳索。
PS|129|5|愿恨恶 锡安 的 都蒙羞退后！
PS|129|6|愿他们像房顶上的草， 一发芽就枯干，
PS|129|7|收割的不够用手抓一把， 捆禾的也不够抱满怀。
PS|129|8|过路的也不说：“愿耶和华所赐的福归与你们！ 我们奉耶和华的名给你们祝福！”
PS|130|1|耶和华啊， 我从深处求告你！
PS|130|2|主啊，求你听我的声音！ 求你侧耳听我恳求的声音！
PS|130|3|耶和华啊，你若究察罪孽， 主啊，谁能站得住呢？
PS|130|4|但在你有赦免之恩， 要叫人敬畏你。
PS|130|5|我等候耶和华，我的心等候； 我也仰望他的话。
PS|130|6|我的心等候主，胜于守夜的等候天亮， 胜于守夜的等候天亮。
PS|130|7|以色列 啊，你当仰望耶和华， 因耶和华有慈爱，有丰盛的救恩。
PS|130|8|他必救赎 以色列 脱离一切的罪孽。
PS|131|1|耶和华啊，我的心不狂妄， 我的眼不高傲； 重大和测不透的事， 我也不敢行。
PS|131|2|我使我心安稳平静，好像母亲怀中断奶的孩子； 我的心在我里面如同断过奶的孩子。
PS|131|3|以色列 啊，你当仰望耶和华， 从今时直到永远！
PS|132|1|耶和华啊，求你记念 大卫 ， 记念他所受的一切苦难！
PS|132|2|他怎样向耶和华起誓， 向 雅各 的大能者许愿：
PS|132|3|“我必不进我的帐幕， 也不上我的床铺；
PS|132|4|我不容我的眼睛睡觉， 也不容我的眼皮打盹；
PS|132|5|直等到我为耶和华寻得所在， 为 雅各 的大能者寻得居所。”
PS|132|6|我们听说约柜在 以法他 ， 我们在 雅珥 的田野寻见它。
PS|132|7|“我们要进他的居所， 在他脚凳前下拜。”
PS|132|8|耶和华啊，求你兴起， 与你有能力的约柜同入安歇之所！
PS|132|9|愿你的祭司披上公义！ 愿你的圣民欢呼！
PS|132|10|求你因你仆人 大卫 的缘故， 不要厌弃你的受膏者！
PS|132|11|耶和华凭信实向 大卫 起了誓，绝不改变： “我要立你身所生的 坐在你的宝座上。
PS|132|12|你的众子若谨守我的约和我所教导他们的法度， 他们的子孙必永远坐在你的宝座上。”
PS|132|13|因为耶和华拣选了 锡安 ， 愿意当作自己的居所：
PS|132|14|“这是我永远安歇之所； 我要住在这地方，因为我愿意在这里。
PS|132|15|我要赐福使粮食丰足， 使其中的贫穷人饱享食物。
PS|132|16|我要使祭司披上救恩， 圣民就要大声欢呼！
PS|132|17|在那里我要使 大卫 的角茁壮， 为我的受膏者预备明灯。
PS|132|18|我要使他的仇敌披上羞耻； 但他的冠冕要在他头上发光。”
PS|133|1|看哪，弟兄和睦同住 是何等的善，何等的美！
PS|133|2|这好比那贵重的油浇在 亚伦 的头上， 流到胡须，又流到他的衣襟；
PS|133|3|又好比 黑门 的甘露降在 锡安山 ； 因为在那里有耶和华所命定的福，就是永远的生命。
PS|134|1|来，称颂耶和华！ 夜间侍立在耶和华殿中，耶和华的仆人，
PS|134|2|当向圣所举手， 称颂耶和华！
PS|134|3|愿造天地的耶和华 从 锡安 赐福给你们！
PS|135|1|哈利路亚！ 你们要赞美耶和华的名！ 侍立在耶和华殿中，耶和华的仆人， 侍立在我们上帝殿院中的，要赞美他！
PS|135|2|
PS|135|3|你们要赞美耶和华， 因耶和华本为善； 要歌颂他的名， 因为这是美好的。
PS|135|4|耶和华拣选 雅各 归自己， 拣选 以色列 作他宝贵的产业。
PS|135|5|我知道耶和华本为大， 也知道我们的主超乎万神之上。
PS|135|6|在天，在地，在海洋，在各深渊， 耶和华都随自己的旨意而行。
PS|135|7|他使云雾从地极上腾， 造电随雨而闪， 从仓库中吹出风来。
PS|135|8|他将 埃及 头生的， 连人带牲畜都击杀了。
PS|135|9|埃及 啊，他施行神迹奇事， 在你们中间，在法老和他所有臣仆身上。
PS|135|10|他击打许多国家， 杀戮大能的君王，
PS|135|11|就是 亚摩利 王 西宏 、 巴珊 王 噩 ， 和 迦南 一切的国度，
PS|135|12|他赏赐他们的地为业， 作为自己百姓 以色列 的产业。
PS|135|13|耶和华啊，你的名字存到永远！ 耶和华啊，你的称号 存到万代！
PS|135|14|耶和华要为自己的百姓伸冤， 为自己的仆人发怜悯。
PS|135|15|外邦的偶像是金的，是银的， 是人手所造的，
PS|135|16|有口却不能言， 有眼却不能看，
PS|135|17|有耳却不能听， 口中也没有气息。
PS|135|18|造它们的要像它们一样， 凡靠它们的也必如此。
PS|135|19|以色列 家啊，要称颂耶和华！ 亚伦 家啊，要称颂耶和华！
PS|135|20|利未 家啊，要称颂耶和华！ 你们敬畏耶和华的，要称颂耶和华！
PS|135|21|住在 耶路撒冷 的、 锡安 的耶和华， 是应当称颂的。 哈利路亚！
PS|136|1|你们要称谢耶和华，因他本为善； 他的慈爱永远长存。
PS|136|2|你们要称谢万神之神， 因他的慈爱永远长存。
PS|136|3|你们要称谢万主之主， 因他的慈爱永远长存。
PS|136|4|称谢那惟一能行大 奇事的， 因他的慈爱永远长存。
PS|136|5|称谢那用智慧造天的， 因他的慈爱永远长存。
PS|136|6|称谢那铺地在水以上的， 因他的慈爱永远长存。
PS|136|7|称谢那造成大光的， 因他的慈爱永远长存。
PS|136|8|他造太阳管白昼， 因他的慈爱永远长存。
PS|136|9|他造月亮星宿管黑夜， 因他的慈爱永远长存。
PS|136|10|称谢那击杀 埃及 凡是头生的， 因他的慈爱永远长存。
PS|136|11|他以大能的手和伸出来的膀臂， 因他的慈爱永远长存。 领 以色列 人从 埃及 人中出来， 因他的慈爱永远长存。
PS|136|12|
PS|136|13|称谢那分裂 红海 的， 因他的慈爱永远长存。
PS|136|14|他领 以色列 从其中经过， 因他的慈爱永远长存；
PS|136|15|却把法老和他的军队推落 红海 里， 因他的慈爱永远长存。
PS|136|16|称谢那引导自己子民行走旷野的， 因他的慈爱永远长存。
PS|136|17|称谢那击杀大君王的， 因他的慈爱永远长存。
PS|136|18|他杀戮威武的君王， 因他的慈爱永远长存；
PS|136|19|杀戮 亚摩利 王 西宏 ， 因他的慈爱永远长存；
PS|136|20|杀戮 巴珊 王 噩 ， 因他的慈爱永远长存。
PS|136|21|他赏赐他们的地为业， 因他的慈爱永远长存；
PS|136|22|作为他仆人 以色列 的产业， 因他的慈爱永远长存。
PS|136|23|我们身处卑微，他顾念我们， 因他的慈爱永远长存。
PS|136|24|他搭救我们脱离敌人， 因他的慈爱永远长存。
PS|136|25|凡有血有肉的，他赐粮食， 因他的慈爱永远长存。
PS|136|26|你们要称谢天上的上帝， 因他的慈爱永远长存。
PS|137|1|我们在 巴比伦 河边， 坐在那里，追想 锡安 ，就哭了。
PS|137|2|在一排柳树中， 我们挂上我们的竖琴。
PS|137|3|掳掠我们的在那里 要我们唱歌； 抢夺我们的要我们为他们作乐： “给我们唱一首 锡安 的歌吧！”
PS|137|4|我们怎能在外邦之土 唱耶和华的歌呢？
PS|137|5|耶路撒冷 啊，我若忘记你， 宁愿我的右手枯萎；
PS|137|6|我若不记得你，不看你过于我最喜乐的， 宁愿我的舌头贴于上膛！
PS|137|7|耶路撒冷 攻破的日子， 以东 人说：“拆毁！拆毁！ 直拆到根基！” 耶和华啊，求你记得！
PS|137|8|将要被灭的 巴比伦 哪， 用你待我们的恶行报复你的，那人有福了。
PS|137|9|抓起你的婴孩摔在磐石上的， 那人有福了。
PS|138|1|我要一心称谢你 ， 在诸神面前歌颂你。
PS|138|2|我要向你的圣殿下拜， 我要因你的慈爱和信实颂扬你的名； 因你使你的名和你的言语显为大， 超乎一切 。
PS|138|3|我呼求的日子，你应允我， 使我壮胆，心里有能力。
PS|138|4|耶和华啊，地上的君王都要称谢你， 因他们听见了你口中的言语。
PS|138|5|他们要歌颂耶和华的作为， 因耶和华大有荣耀。
PS|138|6|耶和华虽崇高，却看顾卑微的人； 骄傲的人，他从远处即能认出。
PS|138|7|我虽困在患难中，你必将我救活； 我的仇敌发怒，你必伸手抵挡他们， 你的右手也必拯救我。
PS|138|8|耶和华必成全他在我身上的旨意； 耶和华啊，你的慈爱永远长存！ 求你不要离弃你手所造的。
PS|139|1|耶和华啊，你已经鉴察我， 认识我。
PS|139|2|我坐下，我起来，你都晓得； 你从远处知道我的意念。
PS|139|3|我行路，我躺卧，你都细察； 你也深知我一切所行的。
PS|139|4|耶和华啊，我舌头上的话， 你没有一句不知道的。
PS|139|5|你前后环绕我， 按手在我身上。
PS|139|6|这样的知识奇妙，是我不能测的； 至高，是我不能及的。
PS|139|7|我往哪里去，躲避你的灵？ 我往哪里逃，躲避你的面？
PS|139|8|我若升到天上，你在那里； 我若躺在阴间，你也在那里。
PS|139|9|我若展开清晨的翅膀， 飞到海极居住，
PS|139|10|就是在那里，你的手必引导我， 你的右手也必扶持我。
PS|139|11|我若说“黑暗必定压碎我， 我周围的亮光必成为黑夜”，
PS|139|12|黑暗对你不再是黑暗， 黑夜却如白昼发亮。 黑暗和光明， 在你看来都是一样。
PS|139|13|我的肺腑是你所造的， 我在母腹中，你已编织 我。
PS|139|14|我要称谢你，因我受造奇妙可畏， 你的作为奇妙，这是我心深知道的。
PS|139|15|我在暗中受造，在地的深处被塑造； 那时，我的形体并不向你隐藏。
PS|139|16|我未成形的体质， 你的眼早已看见了； 你所定的日子，我尚未度一日， 都在你的册子写上了。
PS|139|17|上帝啊，你的意念向我何等宝贵！ 其数何等众多！
PS|139|18|我若数点，比海沙更多； 我睡醒的时候，仍和你同在。
PS|139|19|上帝啊，惟愿你杀戮恶人； 你们好流人血的，离开我去吧！
PS|139|20|他们说恶言顶撞你， 你的仇敌妄称你的名 。
PS|139|21|耶和华啊，恨恶你的，我岂不恨恶他们吗？ 攻击你的，我岂不憎恶他们吗？
PS|139|22|我恨恶他们到极点， 以他们为我的仇敌。
PS|139|23|上帝啊，求你鉴察我，知道我的心思， 试炼我，知道我的意念；
PS|139|24|看在我里面有什么恶行没有， 引导我走永生的道路。
PS|140|1|耶和华啊，求你救我脱离邪恶的人， 保护我脱离残暴的人！
PS|140|2|他们心中图谋奸恶， 日日不停挑起战争。
PS|140|3|他们的舌头锐利如蛇， 嘴唇里有毒蛇的毒液。（细拉）
PS|140|4|耶和华啊，求你庇护我脱离恶人的手， 保护我脱离残暴的人，他们想要推倒我。
PS|140|5|骄傲的人为我暗设罗网和绳索； 他们在路旁张开网，为我设下圈套。（细拉）
PS|140|6|我曾对耶和华说：“你是我的上帝。” 耶和华啊，求你侧耳听我恳求的声音！
PS|140|7|主－耶和华、我救恩的力量啊， 在战争的日子，你遮蔽了我的头。
PS|140|8|耶和华啊，求你不要遂恶人的心愿； 不要成就他们的计谋，免得他们自高。（细拉）
PS|140|9|至于那些昂首围困我的人， 愿他们嘴唇的奸恶陷害 自己！
PS|140|10|愿他们被丢在火中，火炭落在他们身上； 愿他们被抛在深坑里，不能再起来！
PS|140|11|愿说恶言的人在地上站立不住； 愿祸患猎取残暴的人，把他打倒。
PS|140|12|我知道耶和华必为困苦人伸冤， 为贫穷人辩护。
PS|140|13|义人必颂扬你的名， 正直人要在你面前居住。
PS|141|1|耶和华啊，我曾求告你， 求你快快临到我这里！ 我求告你的时候， 求你侧耳听我的声音！
PS|141|2|愿我的祷告如香呈到你面前！ 愿我的手举起 ，如献晚祭！
PS|141|3|耶和华啊，求你看守我的口， 把守我的嘴唇！
PS|141|4|不要使我的心偏向邪恶的事， 以致我和作恶的人一同行恶； 也不叫我吃他们的美食。
PS|141|5|任凭义人击打我，这算为仁慈； 任凭他责备我，这算为头上的膏油； 我的头不躲闪。 人正行恶的时候，我仍要祈祷。
PS|141|6|他们的审判官被扔在岩下， 他们就要听我的话，因为这话甘甜。
PS|141|7|我们的 骨头散落在阴间的口， 就像人耕田刨地 一样。
PS|141|8|主－耶和华啊，我的眼目仰望你； 我投靠你，求你不要使我的性命陷入危险！
PS|141|9|求你保护我脱离恶人为我设的罗网 和作恶之人的圈套！
PS|141|10|愿恶人落在自己的网中， 我却得以逃脱。
PS|142|1|我出声哀告耶和华， 出声恳求耶和华。
PS|142|2|我在他面前倾诉我的苦情， 在他面前陈说我的患难。
PS|142|3|我的灵在我里面发昏的时候， 你知道我的道路。 在我所行的路上， 人为我暗设罗网。
PS|142|4|求你留意向我右边观看， 无人认识我； 我无避难之处， 也无人眷顾我。
PS|142|5|耶和华啊，我曾向你哀求。 我说：“你是我的避难所， 在活人之地，你是我的福分。”
PS|142|6|求你留心听我的呼求， 因我落到极卑微之地； 求你救我脱离迫害我的人， 因为他们比我强盛。
PS|142|7|求你从被囚之地领我出来， 我好颂扬你的名。 义人必环绕我， 因为你用厚恩待我。
PS|143|1|耶和华啊，求你听我的祷告， 侧耳听我的恳求，凭你的信实和公义应允我。
PS|143|2|求你不要审问仆人， 因为在你面前，凡活着的人没有一个是义的。
PS|143|3|因为仇敌迫害我， 将我打倒在地， 使我住在幽暗之处， 像死了许久的人一样。
PS|143|4|我的灵在我里面发昏， 我的心在我里面颤栗。
PS|143|5|我追想古时之日，思想你的一切作为， 默念你手的工作。
PS|143|6|我向你举手， 我的心渴想你，如干旱之地盼雨一样。（细拉）
PS|143|7|耶和华啊，求你速速应允我！ 我的心神耗尽！ 求你不要转脸不顾我， 免得我像那些下入地府的人一样。
PS|143|8|求你使我清晨得听你慈爱的声音， 因我倚靠你； 求你使我知道当走的路， 因我的心仰望你。
PS|143|9|耶和华啊，求你救我脱离我的仇敌！ 我往你那里藏身。
PS|143|10|求你指教我遵行你的旨意， 因你是我的上帝； 愿你至善的灵 引我到平坦之地。
PS|143|11|耶和华啊，求你为你名的缘故将我救活， 凭你的公义，将我从患难中领出来，
PS|143|12|凭你的慈爱剪除我的仇敌， 灭绝所有苦待我的人，因我是你的仆人。
PS|144|1|耶和华─我的磐石是应当称颂的！ 他教导我的手争战， 教导我的指头打仗。
PS|144|2|他是我慈爱的主、我的山寨、 我的碉堡、我的救主、 我的盾牌，是我所投靠的。 他使我的百姓 服在我以下。
PS|144|3|耶和华啊，人算什么，你竟认识他！ 世人算什么，你竟顾念他！
PS|144|4|人不过像一口气， 他的年日如影消逝。
PS|144|5|耶和华啊，求你使天下垂，亲自降临； 求你摸山，使山冒烟。
PS|144|6|求你发出闪电，使仇敌四散， 射出你的箭，使他们混乱。
PS|144|7|求你从高处伸手救拔我， 救我脱离大水，脱离外邦人的手。
PS|144|8|他们的口说谎话， 他们的右手起假誓。
PS|144|9|上帝啊，我要向你唱新歌， 用十弦瑟向你歌颂。
PS|144|10|你是那拯救君王的， 你是那救仆人 大卫 脱离害命之刀的。
PS|144|11|求你救拔我， 救我脱离外邦人的手。 他们的口说谎话， 他们的右手起假誓。
PS|144|12|我们的儿子从幼年好像树苗长大， 我们的女儿如同房角石，按照建宫殿的样式凿成。
PS|144|13|我们的仓盈满，能供应各种粮食； 我们的羊在田野孳生千万。
PS|144|14|我们的牲口驮满货物， 没有人闯进来抢夺， 也没有人出去争战； 我们的街市上也没有哭号的声音。
PS|144|15|这样情况的百姓有福了！ 以耶和华为他们上帝的百姓有福了！
PS|145|1|我的上帝、我的王啊、我要尊崇你！ 我要永永远远称颂你的名！
PS|145|2|我要天天称颂你， 也要永永远远赞美你的名！
PS|145|3|耶和华本为大，该受大赞美， 其大无法测度。
PS|145|4|这一代要对那一代颂赞你的作为， 他们要传扬你的大能。
PS|145|5|他们要述说你威严荣耀的尊荣， 我要默念你奇妙的作为 。
PS|145|6|人要传讲你可畏的能力， 我也要传扬你的伟大。
PS|145|7|他们要将你可记念的大恩传开， 并要高唱你的公义。
PS|145|8|耶和华有恩惠，有怜悯， 不轻易发怒，大有慈爱。
PS|145|9|耶和华善待万有， 他的怜悯覆庇他一切所造的。
PS|145|10|耶和华啊，你一切所造的都要称谢你， 你的圣民也要称颂你。
PS|145|11|他们要传讲你国度的荣耀， 谈论你的大能，
PS|145|12|好让世人知道你大能的作为 和你国度威严的荣耀。
PS|145|13|你的国是永远的国！ 你执掌的权柄存到万代！ 耶和华一切的话信实可靠， 他一切的作为都有慈爱 。
PS|145|14|耶和华扶起所有跌倒的， 扶起所有被压下的。
PS|145|15|万有的眼目都仰望你， 你按时给他们食物。
PS|145|16|你张手， 使一切有生命的都随愿饱足。
PS|145|17|耶和华一切所行的，无不公义， 一切所做的，都有慈爱。
PS|145|18|耶和华临近凡求告他的， 临近所有诚心求告他的人。
PS|145|19|敬畏他的，他必成就他们的心愿， 也必听他们的呼求，拯救他们。
PS|145|20|耶和华保护凡爱他的人， 却要灭绝所有的恶人。
PS|145|21|我的口要述说赞美耶和华的话； 惟愿有血肉之躯的都永永远远称颂他的圣名。
PS|146|1|哈利路亚！ 我的心哪，你要赞美耶和华！
PS|146|2|我一生要赞美耶和华！ 我还活着的时候要歌颂我的上帝！
PS|146|3|你们不要倚靠君王，不要倚靠世人， 他一点也不能帮助。
PS|146|4|他的气一断，就归回尘土， 他所打算的，当日就消灭了。
PS|146|5|以 雅各 的上帝为帮助、 仰望耶和华－他上帝的，这人有福了！
PS|146|6|耶和华造天、地、海和其中的万物， 他守信实，直到永远。
PS|146|7|他为受欺压的伸冤， 赐食物给饥饿的人。 耶和华释放被囚的，
PS|146|8|耶和华开了盲人的眼睛， 耶和华扶起被压下的人， 耶和华喜爱义人。
PS|146|9|耶和华保护寄居的，扶持孤儿和寡妇， 却使恶人的道路弯曲。
PS|146|10|耶和华要作王，直到永远！ 锡安 哪，你的上帝要作王，直到万代！ 哈利路亚！
PS|147|1|哈利路亚！ 歌颂我们的上帝是美善的， 因为他是美好的，赞美他是合宜的。
PS|147|2|耶和华建造 耶路撒冷 ， 聚集 以色列 中被赶散的人。
PS|147|3|他医好伤心的人， 包扎他们的伤处。
PS|147|4|他数点星宿的数目， 一一称它们的名。
PS|147|5|我们的主本为大，大有能力， 他的智慧无法测度。
PS|147|6|耶和华扶持谦卑的人， 将恶人倾覆于地。
PS|147|7|你们要以感谢向耶和华歌唱， 用琴向我们的上帝歌颂。
PS|147|8|他用密云遮天，为地预备雨水， 使草生长在山上。
PS|147|9|他赐食物给走兽 和啼叫的小乌鸦。
PS|147|10|他不喜悦马的力大， 不喜爱人的腿快。
PS|147|11|耶和华喜爱敬畏他 和盼望他慈爱的人。
PS|147|12|耶路撒冷 啊，要颂赞耶和华！ 锡安 哪，要赞美你的上帝！
PS|147|13|因为他坚固了你的门闩， 赐福给你中间的儿女。
PS|147|14|他使你境内平安， 用上好的麦子使你满足。
PS|147|15|他向大地发出命令， 他的话速速颁行。
PS|147|16|他降雪如羊毛， 撒霜如灰烬。
PS|147|17|他掷下冰雹如碎渣， 他发出寒冷，谁能当得起呢？
PS|147|18|他一出令，这些就都融化， 他使风刮起，水便流动。
PS|147|19|他将他的道指示 雅各 ， 将他的律例典章指示 以色列 。
PS|147|20|他未曾这样对待别国， 至于他的典章，他们向来都不知道 。 哈利路亚！
PS|148|1|哈利路亚！ 你们要从天上赞美耶和华， 在高处赞美他！
PS|148|2|他的众使者啊，要赞美他！ 他的诸军啊，都要赞美他！
PS|148|3|太阳月亮啊，要赞美他！ 放光的星宿啊，都要赞美他！
PS|148|4|天上的天和天上的水啊， 你们都要赞美他！
PS|148|5|愿这些都赞美耶和华的名！ 因他一吩咐就都造成。
PS|148|6|他将这些设定，直到永永远远； 他订了律例，不能废去。
PS|148|7|你们哪，都当赞美耶和华： 地上一切所有的，大鱼和深洋，
PS|148|8|火和冰雹，雪和雾气， 成就他命令的狂风，
PS|148|9|大山和小山， 结果子的树木和一切香柏树，
PS|148|10|野兽和一切牲畜， 昆虫和飞鸟，
PS|148|11|世上的君王和万民， 领袖和世上所有的审判官，
PS|148|12|少年和少女， 老人和孩童，
PS|148|13|愿这些都赞美耶和华的名！ 因为独有他的名被尊崇，他的荣耀在天地之上。
PS|148|14|他高举自己百姓的角， 使他的圣民 以色列 人，就是与他相近的百姓得荣耀 。 哈利路亚！
PS|149|1|哈利路亚！ 你们要向耶和华唱新歌， 在圣民的会中赞美他！
PS|149|2|愿 以色列 因造他的主欢喜！ 愿 锡安 的民因他们的王快乐！
PS|149|3|愿他们跳舞赞美他的名， 击鼓弹琴歌颂他！
PS|149|4|因为耶和华喜爱自己的百姓， 他要用救恩当作谦卑人的妆饰。
PS|149|5|愿圣民因所得的荣耀欢乐！ 愿他们在床上也欢呼！
PS|149|6|愿他们口中称颂上帝为至高， 手里有两刃的剑，
PS|149|7|为要报复列国， 惩罚万民。
PS|149|8|要用链子捆他们的君王， 用铁镣锁他们的贵族，
PS|149|9|要在他们身上施行所记录的审判。 他的圣民都享荣耀。 哈利路亚！
PS|150|1|哈利路亚！ 你们要在上帝的圣所赞美他！ 在他显能力的穹苍赞美他！
PS|150|2|要因他大能的作为赞美他， 因他极其伟大赞美他！
PS|150|3|要用角声赞美他， 鼓瑟弹琴赞美他！
PS|150|4|击鼓跳舞赞美他！ 用丝弦的乐器和箫的声音赞美他！
PS|150|5|用大响的钹赞美他！ 用高声的钹赞美他！
PS|150|6|凡有生命的都要赞美耶和华！ 哈利路亚！
PROV|1|1|大卫 的儿子， 以色列 王 所罗门 的箴言：
PROV|1|2|要使人懂得智慧和训诲， 明白通达的言语，
PROV|1|3|使人领受明智的训诲， 就是公义、公平和正直，
PROV|1|4|使愚蒙人灵巧， 使年轻人有知识，有智谋。
PROV|1|5|智慧人听见，增长学问， 聪明人得着智谋，
PROV|1|6|明白箴言和譬喻， 懂得智慧人的言词和谜语。
PROV|1|7|敬畏耶和华是知识的开端； 愚妄人藐视智慧和训诲。
PROV|1|8|我儿啊，要听你父亲的训诲， 不可离弃你母亲的教诲；
PROV|1|9|因为这要作你头上恩惠的华冠， 作你颈上的项链。
PROV|1|10|我儿啊，罪人若引诱你， 你不可随从。
PROV|1|11|他们若说：“你与我们同去， 我们要埋伏杀人流血， 无故地潜藏，杀害无辜；
PROV|1|12|我们好像阴间，把他们活活吞下， 囫囵吞下，如吞下那下到地府的人；
PROV|1|13|我们必得各样宝物， 将所夺来的装满房屋；
PROV|1|14|你来与我们同伙， 共用一个钱囊。”
PROV|1|15|我儿啊，不要与他们走同一道路， 禁止你的脚走他们的路径。
PROV|1|16|因为他们的脚奔跑行恶， 他们急速杀人流血。
PROV|1|17|在飞鸟眼前张设网罗， 一定会徒劳无功；
PROV|1|18|同样，他们埋伏，是自流己血， 他们潜藏，是自害己命。
PROV|1|19|凡靠暴力敛财的，所行之路都是如此， 这种念头必夺去自己的生命。
PROV|1|20|智慧 在街市上呼喊， 在广场上高声呐喊，
PROV|1|21|在热闹街头呼叫， 在城门口，在城中，发出言语，说：
PROV|1|22|“你们无知的人喜爱无知， 傲慢人喜欢傲慢， 愚昧人恨恶知识， 要到几时呢？
PROV|1|23|你们当因我的责备回转， 我要将我的灵浇灌你们， 将我的话指示你们。
PROV|1|24|因为我呼唤，你们不听， 我招手，无人理会。
PROV|1|25|你们忽视我一切的劝戒， 拒听我的责备。
PROV|1|26|你们遭难，我就发笑； 惊恐临到你们， 惊恐如狂风来临， 灾难好像暴风来到， 急难痛苦临到你们身上， 我必嗤笑。
PROV|1|27|
PROV|1|28|那时，他们就会呼求我，我却不回答， 恳切寻求我，却寻不见。
PROV|1|29|因为他们恨恶知识， 选择不敬畏耶和华，
PROV|1|30|不听我的劝戒， 藐视我一切的责备，
PROV|1|31|所以他们要自食其果， 饱胀在自己的计谋中。
PROV|1|32|愚蒙人背道，害死自己， 愚昧人安逸，自取灭亡。
PROV|1|33|惟听从我的，必安然居住， 得享宁静，不怕灾祸。”
PROV|2|1|我儿啊，你若领受我的言语， 珍藏我的命令，
PROV|2|2|留心听智慧， 专心求聪明；
PROV|2|3|你若呼求明理， 扬声求聪明，
PROV|2|4|寻找她，如寻找银子， 搜寻她，如搜寻宝藏，
PROV|2|5|你就懂得敬畏耶和华， 得以认识上帝。
PROV|2|6|因为耶和华赏赐智慧， 知识和聪明都由他口而出。
PROV|2|7|他为正直人珍藏健全的知识， 给行为纯正的人作盾牌，
PROV|2|8|为要保护公正的路， 庇护虔诚人的道。
PROV|2|9|那时，你就明白公义、公平、 正直，和一切完善的道路。
PROV|2|10|因为智慧要进入你的心， 知识要使你内心欢愉。
PROV|2|11|智谋要庇护你， 聪明必保护你，
PROV|2|12|救你脱离恶人的道， 脱离言谈乖谬的人。
PROV|2|13|他们离弃正直的路， 行走黑暗的道，
PROV|2|14|喜欢作恶， 喜爱恶人的错谬。
PROV|2|15|他们的路歪曲， 他们偏离中道。
PROV|2|16|智慧要救你远离陌生女子， 远离那油嘴滑舌的外邦女子。
PROV|2|17|她离弃年轻时的配偶， 忘了自己神圣的盟约。
PROV|2|18|她的家陷入死亡， 她的路偏向阴魂。
PROV|2|19|凡到她那里去的，不得回转， 也得不到生命的路。
PROV|2|20|智慧使你行善人的道， 守义人的路。
PROV|2|21|正直人必在地上居住， 完全人必在其上存留；
PROV|2|22|惟恶人要从地上剪除， 奸诈人要被拔出。
PROV|3|1|我儿啊，不要忘记我的教诲， 你的心要谨守我的命令，
PROV|3|2|因为它们 必加给你长久的日子， 生命的年数与平安。
PROV|3|3|不可使慈爱和诚信离开你， 要系在你颈项上，刻在你心版上。
PROV|3|4|这样，你必在上帝和世人眼前 蒙恩惠，有美好的见识。
PROV|3|5|你要专心仰赖耶和华， 不可倚靠自己的聪明，
PROV|3|6|在你一切所行的路上都要认定他， 他必使你的道路平直。
PROV|3|7|不要自以为有智慧； 要敬畏耶和华，远离恶事。
PROV|3|8|这便医治你的肉体 ， 滋润你的百骨。
PROV|3|9|你要以财物 和一切初熟的土产尊崇耶和华，
PROV|3|10|这样，你的仓库必充满有余， 你的酒池有新酒盈溢。
PROV|3|11|我儿啊，不可轻看耶和华的管教， 也不可厌烦他的责备，
PROV|3|12|因为耶和华所爱的，他必责备， 正如父亲责备所喜爱的儿子。
PROV|3|13|得智慧，得聪明的， 这人有福了。
PROV|3|14|因为智慧的获利胜过银子， 所得的盈余强如金子，
PROV|3|15|比宝石 更宝贵， 你一切所喜爱的，都不足与其比较。
PROV|3|16|她的右手有长寿， 左手有富贵。
PROV|3|17|她的道是安乐， 她的路全是平安。
PROV|3|18|她给持守她的人作生命树， 谨守她的必定蒙福。
PROV|3|19|耶和华以智慧奠立地基， 以聪明铺设诸天，
PROV|3|20|以知识使深渊裂开， 使天空滴下甘露。
PROV|3|21|我儿啊，要谨守健全的知识和智谋， 不可使它们偏离你的眼目。
PROV|3|22|这样，它们必使你的生命有活力， 又作你颈项的美饰。
PROV|3|23|那时，你就坦然行路， 不致跌倒。
PROV|3|24|你躺下，必不惧怕； 你躺卧，睡得香甜。
PROV|3|25|忽然来的惊恐，你不要害怕； 恶人遭毁灭，也不要恐惧，
PROV|3|26|因为耶和华是你的倚靠， 他必保护你的脚不陷入罗网。
PROV|3|27|你的手若有行善的力量， 不可推辞，要施与那应得的人。
PROV|3|28|你若手头方便， 不可对邻舍说： “去吧，明天再来，我必给你。”
PROV|3|29|你的邻舍既在你附近安居， 不可设计害他。
PROV|3|30|人若未曾加害你， 不可无故与他相争。
PROV|3|31|不可嫉妒残暴的人， 不可选择他的任何道路。
PROV|3|32|因为走偏方向的人是耶和华所憎恶的； 正直人为他所亲密。
PROV|3|33|耶和华诅咒恶人的家； 义人的居所他却赐福。
PROV|3|34|他讥诮那爱讥诮的人； 但赐恩给谦卑的人。
PROV|3|35|智慧人必承受尊荣； 愚昧人高升却是羞辱。
PROV|4|1|孩子们，要听父亲的训诲， 留心明白道理。
PROV|4|2|因我给你们好的教导， 不可离弃我的教诲。
PROV|4|3|当我在父亲面前还是小孩， 是母亲独一娇儿的时候，
PROV|4|4|他教导我说：“你的心要持守我的话， 遵守我的命令，你就会存活。
PROV|4|5|要获得智慧，要获得聪明， 不可忘记， 也不可偏离我口中的言语。
PROV|4|6|不可离弃智慧，智慧就庇护你， 要爱她，她就保护你。
PROV|4|7|智慧为首，所以要获得智慧， 要用你一切所有的换取聪明。
PROV|4|8|高举智慧，她就使你升高， 拥抱智慧，她就使你尊荣。
PROV|4|9|她必将恩惠的华冠加在你头上， 把荣冕赐给你。”
PROV|4|10|我儿啊，要听，要领受我的言语， 你就必延年益寿。
PROV|4|11|我已指教你走智慧的道， 引导你行正直的路。
PROV|4|12|你行走，脚步没有阻碍； 你奔跑，也不致跌倒。
PROV|4|13|要持定训诲，不可放松； 要谨守它，因为它是你的生命。
PROV|4|14|不可行恶人的路， 不要走坏人的道；
PROV|4|15|要躲避，不可经过， 要转离而去。
PROV|4|16|他们若不行恶，难以成眠， 不使人跌倒，就睡卧不安；
PROV|4|17|因为他们以邪恶当饼吃， 以暴力当酒喝。
PROV|4|18|但义人的路好像黎明的光， 越照越明，直到正午。
PROV|4|19|恶人的道幽暗， 自己不知因何跌倒。
PROV|4|20|我儿啊，要留心听我的话， 侧耳听我的言语，
PROV|4|21|不可使它们偏离你的眼目， 要存记在你心中。
PROV|4|22|因为找到它们的，就找到生命， 得到全身的医治。
PROV|4|23|你要保守你心，胜过保守一切， 因为生命的泉源由心发出。
PROV|4|24|要离开歪曲的口， 转离偏邪的嘴唇。
PROV|4|25|你的两眼要向前看， 你的双目 直视前方。
PROV|4|26|要修平 你脚下的路， 你一切的道就必稳固。
PROV|4|27|不可偏左偏右， 你的脚要离开邪恶。
PROV|5|1|我儿啊，要留心听我的智慧， 侧耳听我的聪明，
PROV|5|2|为要使你谨守智谋， 嘴唇保护知识。
PROV|5|3|因为陌生女子的嘴唇滴下蜂蜜， 她的口比油更滑，
PROV|5|4|后来却苦似茵蔯， 锐利如两刃的剑。
PROV|5|5|她的脚坠落死亡， 她的脚步踏入阴间，
PROV|5|6|她无法找到生命的道路， 她的路变迁不定，自己却不知道。
PROV|5|7|孩子们，现在要听从我， 不可离弃我口中的言语。
PROV|5|8|你所行的道要远离她， 不可靠近她家的门口，
PROV|5|9|免得将你的尊荣给别人， 将你的岁月给残忍的人；
PROV|5|10|免得陌生人满得你的财富， 你劳苦所得的归入外邦人的家。
PROV|5|11|在你人生终结，你皮肉和身体衰残时， 你必唉声叹气，
PROV|5|12|说：“我为何恨恶管教， 心里轻看责备呢？
PROV|5|13|我不听从教师的话， 也没有侧耳听那教导我的。
PROV|5|14|在聚集的会众中， 我几乎坠入深渊。”
PROV|5|15|你要喝自己池中的水， 饮自己井里的活水。
PROV|5|16|你的泉源岂可溢流在外？ 你的河水岂可流到街上？
PROV|5|17|让它们惟独归你， 不可与陌生人同享。
PROV|5|18|要使你的泉源蒙福， 要喜爱你年轻时的妻子。
PROV|5|19|她如可爱的母鹿，如优美的母羊， 愿她的胸怀使你时时满足， 愿你常常迷恋她的爱情。
PROV|5|20|我儿啊，你为何迷恋陌生女子？ 为何拥抱外邦女子的胸怀？
PROV|5|21|因为人所行的道都在耶和华眼前， 他察验 人一切的路。
PROV|5|22|恶人被自己的罪孽抓住， 被自己罪恶的绳索缠绕。
PROV|5|23|他因不受管教而死亡， 因极度愚昧而走迷。
PROV|6|1|我儿啊，你若为朋友担保， 替陌生人击掌，
PROV|6|2|你就被口中的言语套住， 被嘴里的言语抓住。
PROV|6|3|我儿啊，你既落在朋友手中，当这样行才可救自己： 你要谦卑自己，去恳求你的朋友。
PROV|6|4|不要让你的眼睛睡觉， 不可容你的眼皮打盹。
PROV|6|5|要救自己，如羚羊脱离猎人的手， 如鸟脱离捕鸟人的手。
PROV|6|6|懒惰人哪， 你去察看蚂蚁的动作，就可得智慧。
PROV|6|7|蚂蚁没有领袖， 没有官长，没有君王，
PROV|6|8|尚且在夏天预备食物， 在收割时储存粮食。
PROV|6|9|懒惰人哪，你要睡到几时呢？ 你什么时候才睡醒呢？
PROV|6|10|再睡片时，打盹片时， 抱着双臂躺卧片时，
PROV|6|11|你的贫穷就如盗贼来到， 你的贫乏仿佛拿盾牌的人来临。
PROV|6|12|无赖的恶徒 行事全凭歪曲的口，
PROV|6|13|他眨眼传神， 以脚示意，用指点划，
PROV|6|14|存心乖谬， 常设恶谋，散播纷争。
PROV|6|15|所以，灾难必突然临到他， 他必顷刻被毁，无从医治。
PROV|6|16|耶和华所恨恶的有六样， 他心所憎恶的共有七样：
PROV|6|17|就是高傲的眼，撒谎的舌， 杀害无辜的手，
PROV|6|18|图谋恶计的心， 飞奔行恶的脚，
PROV|6|19|口吐谎言的假证人， 并在弟兄间散播纷争的人。
PROV|6|20|我儿啊，要遵守你父亲的命令， 不可离弃你母亲的教诲。
PROV|6|21|要常挂在你心上， 系在你颈项上。
PROV|6|22|你行走，她必引导你， 你躺卧，她必保护你， 你睡醒，她必与你谈论。
PROV|6|23|因为诫命是灯，教诲是光， 管教的责备是生命的道，
PROV|6|24|要保护你远离邪恶的妇女， 远离外邦女子谄媚的舌头。
PROV|6|25|你不要因她的美色而动心， 也不要被她的眼皮勾引。
PROV|6|26|因为连最后一块饼都会被妓女拿走 ； 有夫之妇会猎取宝贵的生命。
PROV|6|27|人若兜火在怀中， 他的衣服岂能不烧着呢？
PROV|6|28|人若走在火炭上， 他的脚岂能不烫伤呢？
PROV|6|29|与邻舍之妻同寝的，也是如此， 凡亲近她的，难免受罚。
PROV|6|30|贼因饥饿偷窃充饥， 人不藐视他，
PROV|6|31|但若被抓到，要赔偿七倍， 他必赔上家中一切财物。
PROV|6|32|与妇人行奸淫的，便是无知， 做这事的，必毁了自己。
PROV|6|33|他必受损伤和羞辱， 他的羞耻不得消除。
PROV|6|34|丈夫因嫉恨发怒， 报仇的时候绝不留情。
PROV|6|35|他不接受任何赔偿， 你送许多礼物，他也不肯和解。
PROV|7|1|我儿啊，要遵守我的言语， 存记我的命令。
PROV|7|2|遵守我的命令就得存活， 谨守我的教诲，好像保护眼中的瞳人。
PROV|7|3|要系在你指头上， 刻在你心版上。
PROV|7|4|对智慧说“你是我的姊妹”， 称呼聪明为亲人，
PROV|7|5|她就保护你远离陌生女子， 远离油嘴滑舌的外邦女子。
PROV|7|6|我曾在我房屋的窗户内， 透过窗格子往外观看，
PROV|7|7|看见在愚蒙人中， 注意到孩儿中有一个无知的青年，
PROV|7|8|从街上经过，靠近她的巷口， 直往她家的路去，
PROV|7|9|在黄昏，在傍晚， 在半夜，黑暗之中。
PROV|7|10|看哪，有一个女子来迎接他， 是妓女的打扮，有诡诈的心思。
PROV|7|11|她喧嚷，不守约束， 她的脚在家里留不住，
PROV|7|12|有时在街市，有时在广场， 或在各巷口等候。
PROV|7|13|她拉住那青年吻他， 厚着脸皮对他说：
PROV|7|14|“我已献了平安祭， 今日我还了所许的愿。
PROV|7|15|因此，我出来迎接你， 渴望见你的面，我总算找到你了！
PROV|7|16|我已在床上铺好被单， 是 埃及 麻织的花纹布，
PROV|7|17|又用没药、沉香、桂皮 薰了我的床。
PROV|7|18|你来，让我们饱享爱情，直到早晨， 让我们彼此亲爱欢乐。
PROV|7|19|因为我丈夫不在家， 出门远行，
PROV|7|20|他手带钱囊， 要到月圆才回家。”
PROV|7|21|这女子用许多巧言引诱他， 用谄媚的嘴唇催逼他。
PROV|7|22|青年立刻跟随她，好像牛去被宰杀， 又像愚妄人带着脚镣去受刑，
PROV|7|23|直到箭穿进他的肝，如同雀鸟急投罗网， 却不知会赔上自己的生命。
PROV|7|24|孩子们，现在要听从我， 要留心听我口中的言语。
PROV|7|25|你的心不可偏向她的道， 不要误入她的迷途。
PROV|7|26|因为她击倒许多人， 无数的人被她杀戮 。
PROV|7|27|她的家是在阴间之路， 下到死亡之宫。
PROV|8|1|智慧岂不呼唤？ 聪明岂不扬声？
PROV|8|2|她站立在十字路口， 在道路旁高处的顶上，
PROV|8|3|在城门旁，城门口， 入口处，她呼喊：
PROV|8|4|“人哪，我呼唤你们， 我向世人扬声。
PROV|8|5|愚蒙人哪，你们要学习灵巧， 愚昧人哪，你们的心要明辨。
PROV|8|6|你们当听，因我要说尊贵的事， 我要张开嘴唇讲正直的事。
PROV|8|7|我的口要发出真理， 我的嘴唇憎恶邪恶。
PROV|8|8|我口中的言语都是公义， 并无奸诈和歪曲。
PROV|8|9|聪明人看为正确， 有知识的，都以为正直。
PROV|8|10|你们当领受我的训诲，胜过领受银子， 宁得知识，强如得上选的金子。
PROV|8|11|“因为智慧比宝石更美， 一切可喜爱的都不足与其比较。
PROV|8|12|我－智慧以灵巧为居所， 又寻得知识和智谋。
PROV|8|13|敬畏耶和华就是恨恶邪恶； 我恨恶骄傲、狂妄、恶道，和乖谬的口。
PROV|8|14|我有策略和健全的知识， 我聪明，又有能力。
PROV|8|15|君王藉我治国， 王子藉我定公平，
PROV|8|16|王公贵族，所有公义的审判官， 都藉我掌权 。
PROV|8|17|爱我的，我也爱他， 恳切寻求我的，必寻见。
PROV|8|18|财富和尊荣在我， 恒久的财宝和繁荣 也在我。
PROV|8|19|我的果实胜过金子，强如纯金， 我的出产超乎上选的银子。
PROV|8|20|我在公义的道上走， 在公平的路中行，
PROV|8|21|使爱我的承受财产， 充满他们的库房。
PROV|8|22|“耶和华在造化的起头， 在太初创造万物之先，就有 了我。
PROV|8|23|从亘古，从太初， 未有大地以前，我已被立。
PROV|8|24|没有深渊， 没有大水的泉源，我已出生。
PROV|8|25|大山未曾奠定， 小山未有之先，我已出生。
PROV|8|26|那时，他还没有创造大地和田野， 并世上头一撮尘土。
PROV|8|27|他立高天，我在那里， 他在渊面的周围划出圆圈，
PROV|8|28|上使穹苍坚硬， 下使渊源稳固，
PROV|8|29|为沧海定出范围，使水不越过界限， 奠定大地的根基。
PROV|8|30|那时，我在他旁边为工程师， 天天充满喜乐，时时在他面前欢笑，
PROV|8|31|在他的全地欢笑， 喜爱住在人世间。
PROV|8|32|“孩子们，现在要听从我， 谨守我道的有福了。
PROV|8|33|要听训诲，得智慧， 不可弃绝。
PROV|8|34|听从我，天天在我门口守望， 在我门框旁等候的，那人有福了。
PROV|8|35|因为寻得我的，就寻得生命， 他必蒙耶和华的恩惠。
PROV|8|36|得罪我的，害了自己的生命， 凡恨恶我的，喜爱死亡。”
PROV|9|1|智慧建造房屋， 凿成七根柱子，
PROV|9|2|宰杀牲畜，调好美酒， 又摆设筵席，
PROV|9|3|派遣女仆出去， 自己在城中至高处呼唤：
PROV|9|4|“谁是愚蒙的人，让他转到这里来！” 又对那无知的人说：
PROV|9|5|“你们来，吃我的饼， 喝我调的酒。
PROV|9|6|你们要离弃愚蒙，就得存活， 并要走明智的道路。”
PROV|9|7|纠正傲慢人的，必招羞辱， 责备恶人的，必被侮辱。
PROV|9|8|不要责备傲慢人，免得他恨你； 要责备智慧人，他必爱你。
PROV|9|9|教导智慧人，他就越有智慧， 指示义人，他就增长学问。
PROV|9|10|敬畏耶和华是智慧的开端， 认识至圣者便是聪明。
PROV|9|11|藉着我，你的日子必增多， 你生命的年数也必加添。
PROV|9|12|你若有智慧，是自己有智慧； 你若傲慢，就自己承担。
PROV|9|13|愚昧的女子喧嚷， 她是愚蒙，一无所知。
PROV|9|14|她坐在自己家门口， 在城中高处的座位上，
PROV|9|15|呼唤过路的， 向那些在路上直走的人说：
PROV|9|16|“谁是愚蒙的人，让他转到这里来！” 又对那无知的人说：
PROV|9|17|“偷来的水是甜的， 暗藏的饼是美的。”
PROV|9|18|人却不知有阴魂在她那里， 她召唤的人是在阴间的深处。
PROV|10|1|所罗门的箴言： 智慧之子使父亲喜乐； 愚昧之子使母亲担忧。
PROV|10|2|不义之财毫无益处； 惟有公义能救人脱离死亡。
PROV|10|3|耶和华不使义人捱饿； 恶人所欲的，耶和华必拒绝。
PROV|10|4|手懒的，必致穷乏； 手勤的，却要富足。
PROV|10|5|夏天储存的，是智慧之子； 收割时沉睡的，是蒙羞之子。
PROV|10|6|福祉临到义人头上； 恶人的口藏匿残暴。
PROV|10|7|义人的称号带来祝福； 恶人的名字必然败坏。
PROV|10|8|智慧的心，领受诫命； 愚妄的嘴唇，必致倾倒。
PROV|10|9|行正直路的，步步安稳； 走弯曲道的，必致败露。
PROV|10|10|挤眉弄眼的，使人忧患； 愚妄的嘴唇，必致倾倒。
PROV|10|11|义人的口是生命的泉源； 恶人的口藏匿残暴。
PROV|10|12|恨能挑启争端； 爱能遮掩一切过错。
PROV|10|13|聪明人嘴里有智慧； 无知的人背上受刑杖。
PROV|10|14|智慧人积存知识； 愚妄人的口速致败坏。
PROV|10|15|有钱人的财物是他坚固的城； 贫寒人的贫乏使他败坏。
PROV|10|16|义人的报酬带来生命； 恶人的所得用来犯罪。
PROV|10|17|遵守训诲的，行在生命道上； 离弃责备的，走迷了路。
PROV|10|18|隐藏怨恨的，有说谎的嘴唇； 口出毁谤的，是愚昧人。
PROV|10|19|多言多语难免有过； 节制嘴唇是有智慧。
PROV|10|20|义人的舌如上选的银子； 恶人的心所值无几。
PROV|10|21|义人的嘴唇牧养多人； 愚妄人因无知而死亡。
PROV|10|22|耶和华所赐的福使人富足， 并不加上忧虑。
PROV|10|23|愚昧人以行恶为乐； 聪明人以智慧为乐。
PROV|10|24|恶人所怕的，必临到他； 义人的心愿，必蒙应允。
PROV|10|25|暴风一过，恶人归于无有； 义人却有永久的根基。
PROV|10|26|懒惰人使那差他的人， 如醋倒牙，如烟薰目。
PROV|10|27|敬畏耶和华使人长寿； 恶人的年岁必减少。
PROV|10|28|义人的盼望带来喜乐； 恶人的指望必致灭没。
PROV|10|29|耶和华的道是正直人的保障； 却成了作恶人的败坏。
PROV|10|30|义人永不动摇； 恶人不得住在地上。
PROV|10|31|义人的口结出智慧； 乖谬的舌必被割断。
PROV|10|32|义人的嘴唇懂得令人喜悦； 恶人的口只知乖谬。
PROV|11|1|诡诈的天平为耶和华所憎恶； 公平的法码为他所喜悦。
PROV|11|2|骄傲来，羞耻也来； 谦逊人却有智慧。
PROV|11|3|正直人的纯正必引导自己； 奸诈人的邪恶必毁灭自己。
PROV|11|4|遭怒的日子钱财无益； 惟有公义能救人脱离死亡。
PROV|11|5|完全人的义修平自己的路； 但恶人必因自己的恶跌倒。
PROV|11|6|正直人的义必拯救自己； 奸诈人必被自己的欲望缠住。
PROV|11|7|恶人一死，他的指望就灭绝； 罪人的盼望也必灭绝。
PROV|11|8|义人得脱离患难， 有恶人来代替他。
PROV|11|9|不虔敬的人用口败坏邻舍； 义人却因知识得救。
PROV|11|10|义人享福，全城喜乐； 恶人灭亡，人人欢呼。
PROV|11|11|因正直人的祝福，城必升高； 因邪恶人的口，它必倾覆。
PROV|11|12|藐视邻舍的，便是无知； 聪明人却静默不言。
PROV|11|13|到处传话的，泄漏机密； 内心老实的，保守秘密。
PROV|11|14|无智谋，民就败落； 谋士多，就必得胜。
PROV|11|15|为陌生人担保的，必受亏损； 恨恶击掌的，却得安稳。
PROV|11|16|恩慈的妇女得尊荣； 强壮的男子得财富。
PROV|11|17|仁慈的人善待自己； 残忍的人扰害己身。
PROV|11|18|恶人做事，得虚幻的报酬； 撒公义种子的，得实在的报偿。
PROV|11|19|真正行义的，必得生命； 追求邪恶的，必致死亡。
PROV|11|20|心中歪曲的，为耶和华所憎恶； 行为正直的，为他所喜悦。
PROV|11|21|击掌保证，恶人难免受罚； 义人的后裔必得拯救。
PROV|11|22|妇女美貌而无见识， 如同金环戴在猪鼻上。
PROV|11|23|义人的心愿尽是好的； 恶人的指望却带来愤怒。
PROV|11|24|有施舍的，钱财增添； 吝惜过度，反致穷乏。
PROV|11|25|慷慨待人，必然丰裕； 滋润人的，连自己也得滋润。
PROV|11|26|屯粮不卖的，百姓必诅咒他； 愿意出售的，祝福临到头上。
PROV|11|27|恳切求善的，就求得恩宠； 但那求恶的，恶必临到他。
PROV|11|28|倚靠财富的，自己必跌倒； 义人必兴旺如绿叶。
PROV|11|29|扰害己家的，必承受虚空 ； 愚妄人作心中有智慧者的仆人。
PROV|11|30|义人的果实是生命树； 智慧人必能得人。
PROV|11|31|看哪，义人在地上尚且受报， 何况恶人和罪人呢？
PROV|12|1|喜爱管教的，就是喜爱知识； 恨恶责备的，却像畜牲。
PROV|12|2|善人蒙耶和华的恩宠； 设诡计的，耶和华必定罪。
PROV|12|3|人靠恶行不能坚立； 义人的根必不动摇。
PROV|12|4|才德的妻子是丈夫的冠冕； 蒙羞的妇人使丈夫骨头朽烂。
PROV|12|5|义人的思念是公平； 恶人的计谋是诡诈。
PROV|12|6|恶人的言论埋伏流人的血； 正直人的口却拯救人。
PROV|12|7|恶人倾覆，归于无有； 义人的家却屹立不倒。
PROV|12|8|人按自己的智慧得称赞； 心中偏邪的，必被藐视。
PROV|12|9|被人藐视，但有自己仆人 的， 胜过妄自尊大，却缺乏食物。
PROV|12|10|义人顾惜他牲畜的命； 恶人的怜悯也是残忍。
PROV|12|11|耕种自己田地的，必得饱食； 追求虚浮的，却是无知。
PROV|12|12|恶人想得坏人的猎物； 义人的根结出果实。
PROV|12|13|嘴唇的过错是恶人的圈套； 但义人必脱离患难。
PROV|12|14|人因口所结的果实，必饱得美福； 人手所做的，必归到自己身上。
PROV|12|15|愚妄人所行的，在自己眼中看为正直； 惟智慧人从善如流。
PROV|12|16|愚妄人的恼怒立时显露； 通达人却能忍辱。
PROV|12|17|说出真话的，显明公义； 作假见证的，显出诡诈。
PROV|12|18|说话浮躁，犹如刺刀； 智慧人的舌头却能医治。
PROV|12|19|诚实的嘴唇永远坚立； 说谎的舌头只存片时。
PROV|12|20|图谋恶事的，心存诡诈； 劝人和睦的，便得喜乐。
PROV|12|21|义人不遭灾害； 恶人满受祸患。
PROV|12|22|说谎的嘴唇，为耶和华所憎恶； 行事诚实，为他所喜悦。
PROV|12|23|通达人隐藏知识； 愚昧人的心彰显愚昧。
PROV|12|24|殷勤人的手必掌权； 懒惰的人必服苦役。
PROV|12|25|人心忧虑，就必沉重； 一句良言，使心欢乐。
PROV|12|26|义人引导他的邻舍 ； 恶人的道叫人迷失。
PROV|12|27|懒惰的人不烤猎物； 殷勤的人却得宝贵的财物。
PROV|12|28|在公义的路上有生命； 在其道上并无死亡。
PROV|13|1|智慧之子听父亲的训诲； 傲慢人不听责备。
PROV|13|2|人因口所结的果实，必享美福； 奸诈人却意图残暴。
PROV|13|3|谨慎守口的，得保生命； 大张嘴唇的，必致败亡。
PROV|13|4|懒惰的人奢求，却无所得； 殷勤的人必然丰裕。
PROV|13|5|义人恨恶谎言； 恶人可憎可耻。
PROV|13|6|行为纯正的，有公义保护； 犯罪的，被罪恶倾覆。
PROV|13|7|假冒富足的，一无所有； 装作穷乏的，多有财物。
PROV|13|8|财富可作人的生命赎价； 穷乏人却听不见威吓的话。
PROV|13|9|义人的光使人欢喜 ； 恶人的灯要熄灭。
PROV|13|10|骄傲挑启纷争； 听劝言却有智慧。
PROV|13|11|不劳而获之财 必减少； 逐渐积蓄的必增多。
PROV|13|12|盼望迟延，令人心忧； 愿望实现，就是得到生命树。
PROV|13|13|藐视训言的，自取灭亡； 敬畏诫命的，必得善报。
PROV|13|14|智慧人的教诲是生命的泉源， 使人避开死亡的圈套。
PROV|13|15|美好的见识使人得宠； 奸诈人的道路恒久奸诈 。
PROV|13|16|通达人都凭知识行事； 愚昧人张扬自己的愚昧。
PROV|13|17|邪恶的使者必陷入祸患； 忠信的使臣带来医治。
PROV|13|18|弃绝管教的，必贫穷受辱； 领受责备的，必享尊荣。
PROV|13|19|愿望实现，心觉甘甜； 远离恶事，为愚昧人所憎恶。
PROV|13|20|与智慧人同行的，必得智慧； 和愚昧人作伴的，必受亏损。
PROV|13|21|祸患追赶罪人； 义人却得善报。
PROV|13|22|善人给子孙遗留产业； 罪人积财却归义人。
PROV|13|23|穷乏人开垦的地虽多产粮食， 却因不公而被夺走。
PROV|13|24|不忍用杖打儿子的，是恨恶他； 疼爱儿子的，勤加管教。
PROV|13|25|义人吃喝食欲满足； 恶人肚腹却是缺乏。
PROV|14|1|妇人的智慧建立家室； 愚昧却亲手拆毁它 。
PROV|14|2|行事正直的，敬畏耶和华； 偏离正路的，却藐视他。
PROV|14|3|在愚妄人的口中有骄傲的杖； 智慧人的嘴唇必保护自己。
PROV|14|4|没有牛，槽就空空； 土产丰盛却凭牛的力气。
PROV|14|5|诚实的证人不说谎； 虚假的证人口吐谎言。
PROV|14|6|傲慢人枉寻智慧； 聪明人易得知识。
PROV|14|7|不要到愚昧人面前， 你无法从他嘴唇里知道知识。
PROV|14|8|通达人的智慧使他认清自己的道路； 愚昧人的愚昧却是自欺。
PROV|14|9|愚妄人嘲笑赎愆祭 ； 但正直人蒙悦纳。
PROV|14|10|心中的苦楚，只有自己知道； 心里的喜乐，陌生人无法分享。
PROV|14|11|恶人的房屋必倒塌； 正直人的帐棚必兴旺。
PROV|14|12|有一条路，人以为正， 至终成为死亡之路。
PROV|14|13|人在喜笑中，心也会忧愁； 快乐的终点就是愁苦。
PROV|14|14|心中背道的，必满尝其果； 善人必从自己的行为得到回报。
PROV|14|15|无知的人什么话都信； 通达人谨慎自己的脚步。
PROV|14|16|智慧人有所惧怕，就远离恶事； 愚昧人却狂傲自恃。
PROV|14|17|轻易发怒的，行事愚昧； 擅长诡计的，被人恨恶。
PROV|14|18|愚蒙人承受愚昧为产业； 通达人得知识为冠冕。
PROV|14|19|坏人在善人面前俯伏； 恶人在义人门口也是如此。
PROV|14|20|穷乏人，连邻舍也恨他； 有钱人，爱他的人众多。
PROV|14|21|藐视邻舍的，这人有罪； 施恩给困苦人的，这人有福。
PROV|14|22|谋恶的，岂非走入迷途？ 谋善的，有慈爱和诚实。
PROV|14|23|任何勤劳总有收获； 仅耍嘴皮必致穷乏。
PROV|14|24|智慧人的冠冕是富有智慧； 愚昧人的愚昧终究是愚昧。
PROV|14|25|诚实作证，救人性命； 口吐谎言是诡诈。
PROV|14|26|敬畏耶和华的，大有倚靠； 他的儿女也有避难所。
PROV|14|27|敬畏耶和华是生命的泉源， 使人离开死亡的圈套。
PROV|14|28|君王的荣耀在乎民多； 没有百姓，王就衰败。
PROV|14|29|不轻易发怒的，大有聪明； 性情暴躁的，大显愚昧。
PROV|14|30|平静的心使肉体有生气； 嫉妒使骨头朽烂。
PROV|14|31|欺压贫寒人的，是蔑视造他的主； 怜悯贫穷人的，是尊敬主。
PROV|14|32|恶人因所行的恶必被推倒； 义人临死 ，有所投靠。
PROV|14|33|智慧安居在聪明人的心中， 在愚昧人的心中却不认识 。
PROV|14|34|公义使邦国高举； 罪恶是百姓的羞辱。
PROV|14|35|君王的恩宠临到智慧的臣仆； 但其愤怒临到蒙羞的臣仆。
PROV|15|1|回答柔和，使怒消退； 言语粗暴，触动怒气。
PROV|15|2|智慧人的舌善发知识； 愚昧人的口吐出愚昧。
PROV|15|3|耶和华的眼目无处不在， 恶人善人，他都鉴察。
PROV|15|4|温良的舌是生命树； 邪恶的舌使人心碎。
PROV|15|5|愚妄人藐视父亲的管教； 领受责备，使人精明。
PROV|15|6|义人家中多有财富； 恶人获利反受扰害。
PROV|15|7|智慧人的嘴传扬知识； 愚昧人的心并非如此。
PROV|15|8|恶人献祭，为耶和华所憎恶； 正直人祈祷，为他所喜悦。
PROV|15|9|恶人的道路，为耶和华所憎恶； 追求公义的，为他所喜爱。
PROV|15|10|背弃正路的，必受严刑； 恨恶责备的，必致死亡。
PROV|15|11|阴间和冥府 尚且在耶和华面前， 何况世人的心呢？
PROV|15|12|傲慢人不爱受责备， 也不去接近智慧人。
PROV|15|13|心中喜乐，面有喜色； 心里忧愁，灵就忧伤。
PROV|15|14|聪明人的心追求知识； 愚昧人的口吞吃愚昧。
PROV|15|15|困苦人的日子都是愁苦； 心中欢畅的，常享宴席。
PROV|15|16|财宝稀少，敬畏耶和华， 强如财宝众多，烦乱不安。
PROV|15|17|有爱，吃素菜， 强如相恨，吃肥牛。
PROV|15|18|暴怒的人挑启争端； 忍怒的人止息纷争。
PROV|15|19|懒惰人的道像荆棘的篱笆； 正直人的路是平坦大道。
PROV|15|20|智慧之子使父亲喜乐； 愚昧的人藐视母亲。
PROV|15|21|无知的人以愚昧为乐； 聪明的人按正直而行。
PROV|15|22|不先商议，所谋无效； 谋士众多，所谋得成。
PROV|15|23|口善应对，自觉喜乐； 话合其时，何等美好。
PROV|15|24|生命之道使智慧人上升， 使他远离底下的阴间。
PROV|15|25|耶和华必拆毁骄傲人的家， 却要立定寡妇的地界。
PROV|15|26|恶谋为耶和华所憎恶； 良言却是纯净的。
PROV|15|27|暴力敛财的，扰害己家； 恨恶贿赂的，必得存活。
PROV|15|28|义人的心思量应答； 恶人的口吐出恶言。
PROV|15|29|耶和华远离恶人， 却听义人的祈祷。
PROV|15|30|眼睛发光，使心喜乐； 好的信息，滋润骨头。
PROV|15|31|耳听使人得生命的责备， 必居住在智慧人之中。
PROV|15|32|弃绝管教的，轻看自己的生命； 领受责备的，却得智慧的心。
PROV|15|33|敬畏耶和华是智慧的训诲； 要得尊荣，先有谦卑。
PROV|16|1|心中的筹谋在乎人， 舌头的应对出于耶和华。
PROV|16|2|人一切所行的，在自己眼中看为纯洁， 惟有耶和华衡量人的内心。
PROV|16|3|你所做的，要交托耶和华， 你所谋的，就必坚立。
PROV|16|4|耶和华造万物各适其用， 就是恶人也为祸患的日子所造。
PROV|16|5|凡心里骄傲的，为耶和华所憎恶； 击掌保证，他难免受罚。
PROV|16|6|因慈爱和信实，罪孽得赎； 敬畏耶和华的，远离恶事。
PROV|16|7|人所行的若蒙耶和华喜悦， 耶和华也使仇敌与他和好。
PROV|16|8|少获利，行事公义， 强如多获利，行事不义。
PROV|16|9|人心筹算自己的道路； 惟耶和华指引他的脚步。
PROV|16|10|王的嘴唇有圣言， 审判之时，他的口必不差错。
PROV|16|11|公道的秤和天平属耶和华， 囊中一切的法码是他所定。
PROV|16|12|作恶，为王所憎恶， 因国位是靠公义坚立。
PROV|16|13|公义的嘴唇，王喜悦， 说正直话的，他喜爱。
PROV|16|14|王的震怒是死亡的使者， 但智慧人能平息王怒。
PROV|16|15|王脸上的光使人有生命， 他的恩惠好像云带来的春雨。
PROV|16|16|得智慧胜过得金子， 选聪明强如选银子。
PROV|16|17|正直人的道远离恶事， 谨守己路的，保全性命。
PROV|16|18|骄傲在败坏以先， 内心高傲在跌倒之前。
PROV|16|19|心里谦卑与困苦人来往， 强如与骄傲人同分战利品。
PROV|16|20|留心训言的 ，必得福乐； 倚靠耶和华的，这人有福。
PROV|16|21|心中有智慧的，必称为聪明人； 嘴唇的甜言，增长人的学问。
PROV|16|22|人有智慧就有生命的泉源； 愚妄人必受愚妄的惩戒。
PROV|16|23|智慧人的心使他的口谨慎， 又使他的嘴唇增长学问。
PROV|16|24|良言如同蜂巢， 使心甘甜，使骨得医治。
PROV|16|25|有一条路，人以为正， 至终却成为死亡之路。
PROV|16|26|劳力的人为自己劳力， 因为他的口腹催逼他。
PROV|16|27|匪徒图谋奸恶， 嘴唇上的言语仿佛烧焦的火。
PROV|16|28|乖谬的人散播纷争， 造谣的离间密友。
PROV|16|29|残暴的人引诱邻舍， 领他走不好的道路。
PROV|16|30|紧闭双目的，图谋乖谬； 紧咬嘴唇的，成就恶事。
PROV|16|31|白发是荣耀的冠冕， 行在公义道上的，必能得着。
PROV|16|32|不轻易发怒的，胜过勇士； 控制自己脾气的，强如取城。
PROV|16|33|人虽可掷签在膝上， 定事却由耶和华。
PROV|17|1|一块干饼，大家相安； 胜过宴席满屋，大家相争。
PROV|17|2|明智的仆人必管辖蒙羞的儿子， 并在兄弟中同分产业。
PROV|17|3|鼎为炼银，炉为炼金， 惟有耶和华熬炼人心。
PROV|17|4|行恶的，留心听恶毒的嘴唇； 说谎的，侧耳听邪恶的舌头。
PROV|17|5|讥笑穷乏人的，是蔑视造他的主； 幸灾乐祸的，难免受罚。
PROV|17|6|子孙为老人的冠冕； 父母是儿女的荣耀。
PROV|17|7|愚顽人说美言并不相宜， 君子说谎言也不合宜。
PROV|17|8|贿赂在馈赠者的眼中看为玉石， 随处运转都得顺利。
PROV|17|9|包容过错的，寻求友爱； 喋喋不休的，离间密友。
PROV|17|10|一句责备的话深入聪明人的心， 强如打愚昧人一百下。
PROV|17|11|恶人只寻求背叛， 残忍的使者必奉差攻击他。
PROV|17|12|宁可遇见失丧小熊的母熊， 也不愿遇见正行愚昧的愚昧人。
PROV|17|13|以恶报善的， 祸患必不离他的家。
PROV|17|14|纷争掀起，如同缺口的水； 因此，争端尚未爆发就当制止。
PROV|17|15|定恶人为义的，定义人为有罪的， 都为耶和华所憎恶。
PROV|17|16|愚昧人既无知， 为何手拿银钱去买智慧呢？
PROV|17|17|朋友时常亲爱， 弟兄为患难而生。
PROV|17|18|在邻舍面前击掌担保的， 是无知的人。
PROV|17|19|喜爱争吵的，是喜爱过犯； 门盖得高的，自取败坏。
PROV|17|20|心中歪曲的，得不着福乐； 舌头颠倒是非的，陷在祸患中。
PROV|17|21|生愚昧之子的，自己必愁苦； 愚顽人的父亲毫无喜乐。
PROV|17|22|喜乐的心能治好疾病； 忧伤的灵使骨头枯干。
PROV|17|23|恶人暗中受贿赂， 以致弯曲公正的路。
PROV|17|24|聪明人面前有智慧； 愚昧人眼望地的尽头。
PROV|17|25|愚昧的儿子使父亲愁烦， 使那生他的母亲忧苦。
PROV|17|26|刑罚义人实为不善， 责打正直的君子也不宜。
PROV|17|27|节制言语的，有见识； 性情温良的人，有聪明。
PROV|17|28|愚妄人若静默不言，可算为智慧， 闭上嘴唇也可算为聪明。
PROV|18|1|孤僻的人只顾自己的心愿 ， 他鄙视一切健全的知识。
PROV|18|2|愚昧人不喜爱聪明， 只喜爱表达自己的心意。
PROV|18|3|邪恶来，藐视跟着来； 羞耻到，辱骂同时到。
PROV|18|4|人的口所讲的话如同深水， 智慧之泉如涌流的河水。
PROV|18|5|偏袒恶人的情面，是不好的。 审判时使义人受屈，也是不善。
PROV|18|6|愚昧人的嘴唇挑起争端， 一开口就招鞭打。
PROV|18|7|愚昧人的口自取败坏， 他的嘴唇是自己生命的圈套。
PROV|18|8|造谣者的话如同美食， 深入人的肚腹。
PROV|18|9|做工懈怠的， 是破坏者的兄弟。
PROV|18|10|耶和华的名是坚固台， 义人奔入就得安稳。
PROV|18|11|有钱人的财物是他坚固的城， 在他幻想中，犹如高墙。
PROV|18|12|败坏之先，人心骄傲； 要得尊荣，先有谦卑。
PROV|18|13|未听完就回话的， 就是他的愚昧和羞辱。
PROV|18|14|人的心灵忍耐疾病； 心灵忧伤，谁能承当呢？
PROV|18|15|聪明人的心得知识； 智慧人的耳求知识。
PROV|18|16|人的礼物为他开路， 引他到高位的人面前。
PROV|18|17|先诉情由的，似乎有理； 另一人来到，就察出实情。
PROV|18|18|掣签能止息纷争， 也能化解双方激烈的争辩。
PROV|18|19|被冒犯的弟兄 强如难以攻下的坚城； 纷争如同城堡的门闩。
PROV|18|20|人的肚腹必因口所结的果实饱足； 他必因嘴唇所出的感到满足。
PROV|18|21|生死在舌头的掌握之下， 喜爱弄舌的，必吃它所结的果实。
PROV|18|22|得着妻子的，得着好处， 他是蒙了耶和华的恩惠。
PROV|18|23|穷乏人说哀求的话； 有钱人却用威吓的话回答。
PROV|18|24|朋友太多的人，必受损害 ； 但有一知己比兄弟更亲密。
PROV|19|1|行为纯正的穷乏人 胜过嘴唇歪曲的愚昧人。
PROV|19|2|热心而无见识，实为不善； 脚步急快的，易入歧途。
PROV|19|3|人因愚昧自毁前途， 他的心却埋怨耶和华。
PROV|19|4|财富使朋友增多； 贫寒人连仅有的朋友也离弃他。
PROV|19|5|作假见证的，难免受罚； 口吐谎言的，不能逃脱。
PROV|19|6|有权贵的，许多人求他赏脸； 爱送礼的，人都作他的朋友。
PROV|19|7|穷乏人连兄弟都恨他， 何况朋友，更是远离他！ 他用言语追随，他们却不在。
PROV|19|8|得着智慧的，爱惜生命； 持守聪明的，寻得好处。
PROV|19|9|作假见证的，难免受罚； 口吐谎言的，必定灭亡。
PROV|19|10|愚昧人奢华度日并不相宜， 仆人管辖王子，也不应该。
PROV|19|11|人有见识就不轻易发怒， 宽恕人的过失便是自己的荣耀。
PROV|19|12|王的愤怒好像狮子吼叫； 他的恩惠却如草上的甘露。
PROV|19|13|愚昧的儿子是父亲的祸患， 妻子的争吵如雨连连滴漏。
PROV|19|14|房屋钱财是祖宗所遗留的； 惟有贤慧的妻是耶和华所赐的。
PROV|19|15|懒惰使人沉睡， 懈怠的人必捱饿。
PROV|19|16|遵守诫命的，保全生命； 轻忽己路的，必致死亡。
PROV|19|17|怜悯贫寒人的，就是借给耶和华， 他的报偿，耶和华必归还他。
PROV|19|18|趁还有指望，管教你的儿子， 不可执意摧毁他。
PROV|19|19|暴怒的人必受惩罚， 你若救他，必须再救。
PROV|19|20|要听劝言，接受训诲， 使你终久有智慧。
PROV|19|21|人心多有计谋； 惟有耶和华的筹算才能成就。
PROV|19|22|仁慈的人令人喜爱 ， 穷乏人强如说谎言的。
PROV|19|23|敬畏耶和华的，得着生命， 他必饱足安居，不遭祸患。
PROV|19|24|懒惰人把手埋入盘里， 连缩回送进口中也不肯。
PROV|19|25|责打傲慢人，能使无知的人变精明； 责备聪明人，他就明白知识。
PROV|19|26|虐待父亲、驱逐母亲的， 是蒙羞致辱之子。
PROV|19|27|我儿啊，停止听 那叫你偏离知识言语的教导 。
PROV|19|28|卑劣的见证嘲笑公平， 恶人的口吞下罪孽。
PROV|19|29|刑罚是为傲慢人预备的， 鞭打则是为愚昧人的背预备的。
PROV|20|1|酒能使人傲慢，烈酒使人喧嚷， 凡沉溺其中的，都无智慧。
PROV|20|2|王的威吓如狮子吼叫， 激怒他的是自害己命。
PROV|20|3|止息纷争是人的尊荣， 愚妄人争闹不休。
PROV|20|4|懒惰人因冬寒不去耕种， 到收割时，他去寻找，一无所得。
PROV|20|5|人心中的筹算如同深水， 惟聪明人才能汲引出来。
PROV|20|6|很多人声称自己忠信， 但诚信的人谁能遇着呢？
PROV|20|7|义人行为纯正， 他后代的子孙有福了！
PROV|20|8|王坐在审判的位上， 以眼目驱散一切邪恶。
PROV|20|9|谁能说：“我已经洁净了我的心， 脱净了我的罪？”
PROV|20|10|两样的法码和两样的伊法 ， 都为耶和华所憎恶。
PROV|20|11|孩童的行动或纯洁，或正直， 都以行为显明自己。
PROV|20|12|能听的耳，能看的眼， 二者都为耶和华所造。
PROV|20|13|不要贪睡，免致贫穷； 眼要睁开，就可吃饱。
PROV|20|14|买东西的说：“不好，不好！” 及至离去，他却自夸。
PROV|20|15|有金子和许多宝石， 惟知识的嘴唇是贵重的珍宝。
PROV|20|16|谁为陌生人担保，就拿谁的衣服； 谁为外邦人作保，谁就要承当。
PROV|20|17|靠谎言而得的食物，令人愉悦； 到后来，他的口必充满碎石。
PROV|20|18|计谋凭筹算立定， 打仗要凭智谋。
PROV|20|19|到处传话的，泄漏机密； 口无遮拦的，不可与他结交。
PROV|20|20|咒骂父母的， 他的灯必熄灭，在漆黑中。
PROV|20|21|起初很快得来的产业， 终久却不是福。
PROV|20|22|你不要说：“我要以恶报恶”； 要等候耶和华，他必拯救你。
PROV|20|23|两样的法码为耶和华所憎恶， 诡诈的天平也为不善。
PROV|20|24|人的脚步为耶和华所定， 人岂能明白自己的道路呢？
PROV|20|25|人冒失地声称：“这是神圣的！” 许愿之后才细想，就是自陷圈套。
PROV|20|26|智慧的王驱散恶人， 用轮子滚过他们。
PROV|20|27|人的灵是耶和华的灯， 鉴察人的内心深处。
PROV|20|28|慈爱和诚实庇护君王， 他的王位因慈爱而立稳。
PROV|20|29|强壮是青年的荣耀； 白发为老人的尊荣。
PROV|20|30|鞭伤除净邪恶， 责打可洁净人心深处。
PROV|21|1|王的心在耶和华手中像河水， 他能使它随意流转。
PROV|21|2|人一切所行的，在自己眼中看为正直， 惟有耶和华衡量人心。
PROV|21|3|行公义和公平 比献祭更蒙耶和华悦纳。
PROV|21|4|眼高心傲，就是恶人的灯， 都是罪。
PROV|21|5|殷勤筹划的，足致丰裕； 行事急躁的，必致缺乏。
PROV|21|6|用诡诈之舌所得的财富 如被吹散的雾气，趋向灭亡 。
PROV|21|7|恶人的残暴必扫去自己， 因他们不肯按公平行事。
PROV|21|8|有罪的人其路弯曲； 纯洁的人行为正直。
PROV|21|9|宁可住在房顶的一角， 也不与好争吵的妇人同住。
PROV|21|10|恶人的心渴想邪恶， 他的眼并不怜悯邻舍。
PROV|21|11|傲慢人受惩罚，愚蒙人可得智慧； 智慧人受训诲，便得知识。
PROV|21|12|公义的上帝 鉴察恶人的家， 他倾覆恶人，以致灭亡。
PROV|21|13|塞耳不听贫寒人哀求的， 他自己呼求，也不蒙应允。
PROV|21|14|暗中送的礼物挽回怒气， 怀里的贿赂能止息暴怒。
PROV|21|15|秉公行义使义人喜乐， 却使作恶的人败坏。
PROV|21|16|人偏离智慧的路， 必与阴魂为伍 。
PROV|21|17|爱宴乐的，必致穷乏； 贪爱酒和油的，必不富足。
PROV|21|18|恶人作义人的赎价， 奸诈人代替正直人。
PROV|21|19|宁可住在旷野之地， 也不与争吵易怒的妇人同住。
PROV|21|20|智慧人的居所积蓄宝物与膏油 ； 愚昧人却挥霍一空。
PROV|21|21|追求公义慈爱的， 就寻得生命、公义 和尊荣。
PROV|21|22|智慧人爬上勇士的城墙， 摧毁他所倚靠的堡垒。
PROV|21|23|谨守口和舌的， 就保护自己免受灾难。
PROV|21|24|心骄气傲的人名叫傲慢， 他行事出于狂妄骄傲。
PROV|21|25|懒惰人的欲望害死自己， 因为他的手不肯做工；
PROV|21|26|有人终日贪得无餍， 义人却施舍而不吝惜。
PROV|21|27|恶人献的祭是可憎的， 何况他存恶意来献呢？
PROV|21|28|不实的见证必消灭； 惟聆听真情的，他的证词有力。
PROV|21|29|恶人脸无羞耻； 正直人行事坚定 。
PROV|21|30|没有人能以智慧、聪明、 谋略抵挡耶和华。
PROV|21|31|马是为打仗之日预备的； 得胜却在于耶和华。
PROV|22|1|美名胜过大财， 宏恩强如金银。
PROV|22|2|有钱人与穷乏人相遇 ， 他们都为耶和华所造。
PROV|22|3|通达人见祸就藏躲； 愚蒙人却前往受害。
PROV|22|4|敬畏耶和华心存谦卑， 就得财富、尊荣、生命为赏赐。
PROV|22|5|歪曲的人路上有荆棘和罗网， 保护自己生命的，必要远离。
PROV|22|6|教养孩童走当行的道， 就是到老他也不偏离。
PROV|22|7|有钱人管辖穷乏人， 欠债的是债主的仆人。
PROV|22|8|撒不义种子的必收割灾祸， 他逞怒的杖也必废掉。
PROV|22|9|眼目仁慈的必蒙福， 因他将食物分给贫寒人。
PROV|22|10|赶出傲慢人，争端就消除， 纷争和羞辱也必止息。
PROV|22|11|喜爱清心，嘴唇有恩言的， 王必与他为友。
PROV|22|12|耶和华的眼目保护知识， 却毁坏奸诈人的言语。
PROV|22|13|懒惰人说：“外面有狮子， 我在街上必被杀害。”
PROV|22|14|陌生女子的口是深坑， 耶和华所憎恶的，必陷在其中。
PROV|22|15|愚昧迷住孩童的心， 用管教的杖可以远远赶除。
PROV|22|16|欺压贫寒人为要利己的， 并送礼给有钱人的，都必缺乏。
PROV|22|17|你要侧耳听智慧人的言语 ， 留心领会我的知识。
PROV|22|18|你若心中存记， 嘴唇也准备就绪，这是美的。
PROV|22|19|我今日特地指教你， 为要使你倚靠耶和华。
PROV|22|20|谋略和知识的美事 ， 我岂没有写给你吗？
PROV|22|21|要使你明白真情实理， 好将实情回覆那差你来的人。
PROV|22|22|不可因人贫寒就抢夺他， 也不可在城门口欺压困苦人，
PROV|22|23|因耶和华必为他们辩护， 也必夺取那抢夺者的命。
PROV|22|24|不可结交好生气的人， 也不可与暴怒的人来往，
PROV|22|25|恐怕你效法他的行为， 自己就陷在圈套里。
PROV|22|26|不要为人击掌担保， 也不要为债务作保。
PROV|22|27|你若没有什么可偿还， 何必使人夺去你睡卧的床呢？
PROV|22|28|祖先所立的地界， 你不可挪移。
PROV|22|29|你看见办事殷勤的人吗？ 他必侍立在君王面前， 不在平庸的人面前。
PROV|23|1|你若与长官坐席， 要留意在你面前的是谁。
PROV|23|2|你若是胃口大的人， 就当拿刀放在喉咙上。
PROV|23|3|不可贪恋长官的美食， 因为那是欺哄人的食物。
PROV|23|4|不要劳碌求富， 要有聪明来节制。
PROV|23|5|你定睛在财富，它就消失， 因为它必长翅膀，如鹰向天飞去。
PROV|23|6|守财奴 的饭，你不要吃， 也不要贪恋他的美味；
PROV|23|7|因为他的心怎样算计 ， 他为人就是这样。 他虽对你说：请吃，请喝， 他的心却与你相背。
PROV|23|8|你所吃的那点食物必吐出来， 你恭维的话语也必落空。
PROV|23|9|不要说话给愚昧人听， 因他必藐视你智慧的言语。
PROV|23|10|不可挪移古时的地界， 也不可侵占孤儿的田地，
PROV|23|11|因他们的救赎者 大有能力， 他必向你为他们辩护。
PROV|23|12|你要留心领受训诲， 侧耳听从知识的言语。
PROV|23|13|不可不管教孩童， 因为你用杖打他，他不会死。
PROV|23|14|你用杖打他， 就可以救他的性命免下阴间。
PROV|23|15|我儿啊，你若心存智慧， 我的心就甚欢喜。
PROV|23|16|你的嘴唇若说正直话， 我的心肠也必快乐。
PROV|23|17|你的心不要羡慕罪人， 却要羡慕常常敬畏耶和华的人，
PROV|23|18|因为你必有前途， 你的指望也不致断绝。
PROV|23|19|我儿啊，你当听，当存智慧， 好在正道上引导你的心。
PROV|23|20|不可与好饮酒的人在一起， 也不要跟贪吃肉的人来往，
PROV|23|21|因为贪食好酒的，必致贫穷， 爱睡觉的，必穿破烂衣服。
PROV|23|22|你要听从生你的父亲； 不可因母亲年老而轻看她。
PROV|23|23|你当获得真理，不可出卖， 智慧、训诲和聪明也是一样。
PROV|23|24|义人的父亲必大大快乐， 生智慧儿子的，必因他欢喜。
PROV|23|25|愿你的父母欢喜， 愿那生你的母亲快乐。
PROV|23|26|我儿啊，要将你的心归我， 你的眼目也要喜爱 我的道路。
PROV|23|27|妓女是深坑， 外邦女子是窄井。
PROV|23|28|她像强盗埋伏， 她使奸诈的人增多。
PROV|23|29|谁有祸患？谁有灾难？ 谁有纷争？谁有焦虑？ 谁无故受伤？谁的眼目红赤？
PROV|23|30|就是那流连饮酒的人， 常去寻找调和的酒。
PROV|23|31|酒发红，在杯中闪烁时， 你不可观看； 虽下咽舒畅， 终究它必咬你如蛇，刺你如毒蛇。
PROV|23|32|
PROV|23|33|你的眼睛必看见怪异的事， 你的心必发出乖谬的话。
PROV|23|34|你必像躺在深海中， 或卧在桅杆顶上，
PROV|23|35|说：“人击打我，但我未受伤， 重击我，我不觉得。 我几时清醒， 还要再去寻酒。”
PROV|24|1|你不要嫉妒恶人， 也不要渴望与他们相处，
PROV|24|2|因为他们的心图谋暴行， 他们的嘴唇谈论奸恶。
PROV|24|3|房屋因智慧建造， 因聪明立稳；
PROV|24|4|又因知识， 屋内充满各样美好宝贵的财物。
PROV|24|5|有智慧的勇士大有能力， 有知识的人力上加力。
PROV|24|6|你去打仗，要凭智谋； 谋士众多，就必得胜。
PROV|24|7|对愚妄人，智慧高不可及， 所以他在城门不敢开口。
PROV|24|8|图谋行恶的， 必称为奸诈人。
PROV|24|9|愚妄人的筹划尽是罪恶， 傲慢者为人所憎恶。
PROV|24|10|在患难时你若灰心， 你的力量就微小。
PROV|24|11|人被拉到死亡，你要解救； 人将被杀，你须拦阻。
PROV|24|12|你若说：“看哪，这事我们不知道”， 那衡量人心的岂不明白吗？ 保护你性命的岂不知道吗？ 他岂不按各人所做的报应各人吗？
PROV|24|13|我儿啊，你要吃蜜，因为它是美好的， 要让甘甜的蜜滴入你的口。
PROV|24|14|你要知道，智慧对你的生命正像如此。 你若找着，必有前途， 你的指望也不致断绝。
PROV|24|15|你这恶人，不可埋伏攻击义人的家， 也不可毁坏他安居之所。
PROV|24|16|因为义人虽七次跌倒，仍必兴起； 恶人却被祸患倾倒。
PROV|24|17|你的仇敌跌倒，你不要欢喜， 他倾倒，你的心不要快乐；
PROV|24|18|恐怕耶和华看见就不喜悦， 将怒气从仇敌身上转过来。
PROV|24|19|不要为作恶的心怀不平， 也不要嫉妒恶人，
PROV|24|20|因为坏人没有前途， 恶人的灯也必熄灭。
PROV|24|21|我儿啊，你要敬畏耶和华与君王， 不可结交反覆无常的人，
PROV|24|22|因为他们的灾难必忽然兴起。 谁能知道耶和华与君王所施行的毁灭呢？
PROV|24|23|以下也是智慧人的箴言： 审判时看人情面是不好的。
PROV|24|24|对恶人说“你是义人”的， 万民必诅咒，万族必恼恨。
PROV|24|25|责备恶人的，必得喜悦， 美好的福分也必临到他。
PROV|24|26|应对合宜的， 犹如与人亲吻。
PROV|24|27|你要在外面预备材料， 在田间为自己准备齐全， 然后才建造你的房屋。
PROV|24|28|不可无故作证反对邻舍， 也不可用嘴唇欺骗人。
PROV|24|29|不可说：“人怎样待我，我也怎样待他， 我必照他所做的报复他。”
PROV|24|30|我经过懒惰人的田地， 走过无知人的葡萄园，
PROV|24|31|看哪，它长满了荆棘， 荨麻盖地面， 石墙也坍塌了。
PROV|24|32|我看见就留心思想， 我看着就领受训诲。
PROV|24|33|再睡片时，打盹片时， 抱着双臂躺卧片时，
PROV|24|34|你的贫穷就如盗贼来到， 你的贫乏仿佛拿盾牌的人来临。
PROV|25|1|以下也是 所罗门 的箴言，是 犹大 王 希西家 的人所誊录的。
PROV|25|2|隐藏事情是上帝的荣耀； 查明事情乃君王的荣耀。
PROV|25|3|天之高，地之深， 君王之心测不透。
PROV|25|4|除去银子的渣滓， 银匠就做出器皿来。
PROV|25|5|除去王面前的恶人， 国位就靠公义坚立。
PROV|25|6|不可在君王面前妄自尊大， 也不要站在大人的位上。
PROV|25|7|宁可让人家说“请你上到这里来”， 强如在你觐见的贵人面前令你退下。
PROV|25|8|不要冒失出去与人争讼 ， 免得你的邻舍羞辱你， 最后你就不知怎么做。
PROV|25|9|要与邻舍争辩你的案情， 不可泄漏他人的隐密，
PROV|25|10|恐怕听见的人责骂你， 你就难以摆脱臭名。
PROV|25|11|一句话说得合宜， 就如金苹果在银网子里
PROV|25|12|智慧人的劝戒在顺从的人耳中， 好像金环和金首饰。
PROV|25|13|忠信的使者对那差他的人， 就如收割时有冰雪的凉气， 使主人的心舒畅。
PROV|25|14|人空夸礼物而不肯赠送， 就好像有风有云却无雨。
PROV|25|15|恒常的忍耐可以劝服君王， 柔和的舌头能折断骨头。
PROV|25|16|你得了蜜，吃够就好， 免得过饱就吐出来。
PROV|25|17|你的脚要少进邻舍的家， 免得他厌烦你，恨恶你。
PROV|25|18|作假见证陷害邻舍的， 就是大锤，是利刀，是快箭。
PROV|25|19|患难时倚靠奸诈的人， 好像牙齿断裂，又如脚脱臼。
PROV|25|20|对伤心的人唱歌， 就如冷天脱他的衣服， 又如在碱上倒醋 。
PROV|25|21|你的仇敌若饿了，就给他饭吃， 若渴了，就给他水喝；
PROV|25|22|因为你这样做，就是把炭火堆在他的头上， 耶和华必回报你。
PROV|25|23|正如北风生雨， 毁谤的舌头也生怒容。
PROV|25|24|宁可住在房顶的一角， 也不与好争吵的妇人同住。
PROV|25|25|有好消息从遥远的地方来， 就如凉水滋润口渴的人。
PROV|25|26|义人在恶人面前退缩， 好像搅浑之泉，污染之井。
PROV|25|27|吃蜜过多是不好的， 自求荣耀也是一样。
PROV|25|28|人不克制自己的心， 就像毁坏的城没有墙。
PROV|26|1|愚昧人得尊荣不相宜， 正如夏天落雪，收割时下雨。
PROV|26|2|诅咒不会无故临到 ， 正如麻雀掠过，燕子翻飞。
PROV|26|3|鞭子是为打马，辔头是为勒驴， 刑杖正是为打愚昧人的背。
PROV|26|4|不要照愚昧人的愚昧话回答他， 免得你与他一样。
PROV|26|5|要照愚昧人的愚昧话回答他， 免得他自以为有智慧。
PROV|26|6|藉愚昧人的手寄信的， 就像砍断双脚，喝下残暴。
PROV|26|7|箴言在愚昧人的口中， 正如瘸子的脚悬空无用。
PROV|26|8|将尊荣给愚昧人的， 就像石头绑在弹弓上。
PROV|26|9|箴言在愚昧人的口中， 好像荆棘刺入醉汉的手。
PROV|26|10|雇愚昧人的，与雇过路人的， 就像弓箭手射伤任何人。
PROV|26|11|愚昧人重复做愚昧之事， 就如狗转过来吃自己所吐的。
PROV|26|12|你看见自以为有智慧的人吗？ 愚昧人比他更有指望。
PROV|26|13|懒惰人说：“道路有猛狮， 街上有壮狮。”
PROV|26|14|懒惰人在床上， 就像门在轴心上转动一样。
PROV|26|15|懒惰人把手埋入盘里， 就是送进口中也觉得累。
PROV|26|16|懒惰人眼看自己 比七个善于应对的人更有智慧。
PROV|26|17|过路时卷入与己无关的纷争， 好像人揪住狗耳一般。
PROV|26|18|人欺骗邻舍，却说 “我只是开玩笑而已”， 他就像疯狂的人抛掷致死的火把和利箭。
PROV|26|19|
PROV|26|20|火缺了柴就必熄灭； 无人造谣，纷争就止息。
PROV|26|21|好争吵的人煽动争端， 就如余火加炭，火上加柴一样。
PROV|26|22|造谣者的话如同美食， 深入人的肚腹。
PROV|26|23|火热的 嘴唇，邪恶的心， 好像银渣包在瓦器上。
PROV|26|24|仇敌用嘴唇掩饰， 心里却藏着诡诈；
PROV|26|25|他用甜言蜜语，你不能相信他， 因为他心中有七样可憎恶的事。
PROV|26|26|他虽用诡诈掩饰怨恨， 他的邪恶必在集会中显露。
PROV|26|27|挖陷坑的，自己必陷在其中； 滚石头的，石头反滚在他身上。
PROV|26|28|虚谎的舌憎恨他所压伤的人； 谄媚的口败坏人的事。
PROV|27|1|不要为明天自夸， 因为你不知道每天会发生何事。
PROV|27|2|要让陌生人夸奖你，不可用口自夸； 让外邦人称赞你，不可用嘴唇称赞自己。
PROV|27|3|石头沉，沙土重， 愚妄人的恼怒比这两样更沉重。
PROV|27|4|愤怒为残忍，怒气像狂澜， 惟有嫉妒，谁能挡得住呢？
PROV|27|5|当面的责备 胜过隐藏的爱情。
PROV|27|6|朋友加的伤痕出于忠诚； 敌人的亲吻却是多余。
PROV|27|7|人吃饱了，厌恶蜂房的蜜； 人饥饿了，一切苦物都觉甘甜。
PROV|27|8|人离故乡漂泊， 就像雀鸟离窝四处飞翔。
PROV|27|9|膏油与香料使人心喜悦， 朋友诚心的劝勉也是如此甘美。
PROV|27|10|你的朋友和父亲的朋友， 你都不可离弃。 你遭难时，不要上兄弟的家去； 相近的邻舍强如远方的兄弟。
PROV|27|11|我儿啊，你要做智慧人，好叫我的心欢喜， 使我可以回答那辱骂我的人。
PROV|27|12|通达人见祸就藏躲； 愚蒙人却前往受害。
PROV|27|13|谁为陌生人担保，就拿谁的衣服； 谁为外邦女子作保，谁就要承当。
PROV|27|14|清晨起来大声给朋友祝福的， 就算是诅咒他。
PROV|27|15|下雨天连连滴漏， 好争吵的妇人就像这样；
PROV|27|16|拦阻她的，就是拦阻风， 又像用右手抓油。
PROV|27|17|以铁磨铁，越磨越利， 朋友当面琢磨，也是如此。
PROV|27|18|看守无花果树的，必吃树上的果子； 敬奉主人的，必得尊荣。
PROV|27|19|水中照脸，彼此相符； 人心相映，也是如此。
PROV|27|20|阴间和冥府 永不满足， 人的眼目也是如此。
PROV|27|21|鼎为炼银，炉为炼金， 口中的称赞也试炼人。
PROV|27|22|用杵把愚妄人与谷粒一同捣在臼中， 他的愚昧还是离不了他。
PROV|27|23|你要详细知道你羊群的景况， 留心照顾你的牛群，
PROV|27|24|因为财富不能永留， 冠冕岂能存到万代？
PROV|27|25|青草除去，嫩草长出， 山上的菜蔬也被采收。
PROV|27|26|绵羊可以做衣服， 公山羊可作田地的价值，
PROV|27|27|并有母山羊奶够你吃， 够你养家和女仆的生活。
PROV|28|1|恶人虽无人追赶也逃跑； 义人却胆壮像狮子。
PROV|28|2|地上因有罪过，君王就多更换； 因聪明和有见识的人，国必长存。
PROV|28|3|穷乏人欺压贫寒人， 好像暴雨扫过，不留粮食。
PROV|28|4|离弃律法的，夸奖恶人； 遵守律法的，却与恶人相争。
PROV|28|5|恶人不明白公义； 惟有寻求耶和华的，无不明白。
PROV|28|6|行为纯正的穷乏人 胜过行事歪曲的有钱人。
PROV|28|7|谨守教诲的，是聪明之子； 与贪食者为伍的，却羞辱其父。
PROV|28|8|人以厚利增加财富， 是给那怜悯贫寒人的积财。
PROV|28|9|转耳不听教诲的， 他的祈祷也可憎。
PROV|28|10|诱惑正直人行恶道的，必掉在自己的坑里； 惟有完全人必承受福分。
PROV|28|11|有钱人自以为有智慧， 但聪明的贫寒人能看穿他。
PROV|28|12|义人高升，有大荣耀； 恶人兴起，人就躲藏。
PROV|28|13|遮掩自己过犯的，必不顺利； 承认且离弃过犯的，必蒙怜悯。
PROV|28|14|常存敬畏的，这人有福了； 心里刚硬的，必陷在祸患里。
PROV|28|15|邪恶的君王压制贫民， 好像吼叫的狮子，又如觅食的熊。
PROV|28|16|无知的君王多行暴虐； 恨恶非分之财的，必年长日久。
PROV|28|17|背负流人血之罪的，必逃跑直到地府； 愿无人帮助他！
PROV|28|18|行为正直的，必蒙拯救； 行事弯曲的，立时跌倒。
PROV|28|19|耕种自己田地的，粮食充足； 追求虚浮的，穷困潦倒。
PROV|28|20|诚实人必多得福； 想要急速发财的，难免受罚。
PROV|28|21|看人情面是不好的； 却有人因一块饼而犯法。
PROV|28|22|守财奴 想要急速发财， 却不知穷乏必临到他身上。
PROV|28|23|责备人的，后来蒙人喜悦， 多于那用舌头谄媚人的。
PROV|28|24|抢夺父母竟说“这不是罪过”， 此人与毁灭者同类。
PROV|28|25|心中贪婪的，挑起争端； 倚靠耶和华的，必得丰裕。
PROV|28|26|心中自以为是的，就是愚昧人； 凭智慧行事的，必蒙拯救。
PROV|28|27|赒济穷乏人的，不致缺乏； 遮眼不看的，多受诅咒。
PROV|28|28|恶人兴起，人就躲藏； 恶人败亡，义人必增多。
PROV|29|1|人屡次受责罚，仍然硬着颈项， 他必顷刻被毁，无从医治。
PROV|29|2|义人增多，民就喜乐； 恶人掌权，民就叹息。
PROV|29|3|爱慕智慧的，使父亲喜乐； 结交妓女的，却浪费钱财。
PROV|29|4|王藉公平，使国坚定； 强索贡物的，使它毁坏。
PROV|29|5|谄媚邻舍的， 就是设网罗绊他的脚。
PROV|29|6|恶人犯罪，自陷圈套； 惟独义人欢呼喜乐。
PROV|29|7|义人关注贫寒人的案情； 恶人不明了这种知识。
PROV|29|8|傲慢人煽动全城； 智慧人止息众怒。
PROV|29|9|智慧人与愚妄人有争讼， 或怒或笑，总不得安宁。
PROV|29|10|好流人血的，恨恶完全人， 正直人却顾惜 他的性命。
PROV|29|11|愚昧人怒气全发； 智慧人自我平息。
PROV|29|12|君王若听谎言， 他一切臣仆都是奸恶。
PROV|29|13|穷乏人和欺压者相遇 ， 耶和华使他们的眼目明亮。
PROV|29|14|君王凭诚信判断贫寒人， 他的国位必永远坚立。
PROV|29|15|杖打和责备能增加智慧； 任性的少年使母亲羞愧。
PROV|29|16|恶人多，过犯也加多， 义人必看见他们败亡。
PROV|29|17|管教你的儿子，他就使你得安宁， 也使你心里喜乐。
PROV|29|18|没有异象 ，民就放肆； 惟遵守律法的，便为有福。
PROV|29|19|仆人不能靠言语受教； 他即使明白，也不回应。
PROV|29|20|你见过言语急躁的人吗？ 愚昧人比他更有指望。
PROV|29|21|人将仆人从小娇养， 至终必带来忧伤 。
PROV|29|22|好生气的人挑起争端， 暴怒的人多多犯错。
PROV|29|23|人的高傲使自己蒙羞； 心里谦逊的，必得尊荣。
PROV|29|24|与盗贼分赃的，是恨恶自己的性命； 他虽听见发誓的声音，也不告诉人。
PROV|29|25|惧怕人的，陷入圈套； 惟有倚靠耶和华的，必得安稳。
PROV|29|26|求王恩的人多； 人获公正来自耶和华。
PROV|29|27|不义之人，义人憎恶； 行事正直的，恶人憎恶。
PROV|30|1|雅基 的儿子、 玛撒 人 亚古珥 的言语 ，是这人对 以铁 和 乌甲 说的。
PROV|30|2|我比众人更像畜牲， 也没有人的聪明。
PROV|30|3|我没有学好智慧， 也不认识至圣者。
PROV|30|4|谁升天又降下来？ 谁聚风在手掌中？ 谁包水在衣服里？ 谁立定地的四极？ 他名叫什么？ 他儿子名叫什么？ 你知道吗？
PROV|30|5|上帝的言语句句都是炼净的， 投靠他的，他便作他们的盾牌。
PROV|30|6|你不可加添他的言语， 恐怕他责备你，你就显为说谎的。
PROV|30|7|我求你两件事， 在我未死之先，不要拒绝我：
PROV|30|8|求你使虚假和谎言远离我， 使我不贫穷也不富足， 赐给我需用的饮食。
PROV|30|9|免得我饱足了，就不认你，说： “耶和华是谁呢？” 又恐怕我贫穷就偷窃， 以致亵渎我上帝的名。
PROV|30|10|不要向主人谗害他的仆人， 恐怕他诅咒你，你便算为有罪。
PROV|30|11|有一类人，诅咒父亲， 不给母亲祝福。
PROV|30|12|有一类人，自以为纯洁， 却没有洗净自己的污秽。
PROV|30|13|有一类人，眼目何其高傲， 眼皮也是高举。
PROV|30|14|有一类人，牙如剑，齿如刀， 要吞灭地上的困苦人和世间的贫穷人。
PROV|30|15|水蛭有两个女儿： “给呀，给呀。” 有三样不知足的， 不说“够了”的有四样：
PROV|30|16|阴间和不生育的子宫， 吸水不足的地，还有不说“够了”的火。
PROV|30|17|嘲笑父亲、藐视而不听从母亲的， 谷中的乌鸦必啄他的眼睛，小鹰也必吃它。
PROV|30|18|我所测不透的奇妙有三样， 我所不知道的有四样：
PROV|30|19|就是鹰在空中飞的道， 蛇在磐石上爬的道， 船在海中行的道， 男与女交合的道。
PROV|30|20|淫妇的道是这样， 她吃了，把嘴一擦就说： “我没有行恶。”
PROV|30|21|使地震动的有三样， 地承担不起的有四样：
PROV|30|22|就是仆人作王， 愚顽人吃得饱足，
PROV|30|23|令人憎恶的女子出嫁， 婢女取代她的女主人。
PROV|30|24|地上有四样东西虽小，却甚聪明：
PROV|30|25|蚂蚁是无力之类， 却在夏天预备粮食。
PROV|30|26|石獾并非强壮之类， 却在岩石中造房子。
PROV|30|27|蝗虫没有君王， 却分队而出。
PROV|30|28|壁虎你用手就可抓住， 它却住在王宫。
PROV|30|29|脚步威武的有三样， 行走威武的有四样：
PROV|30|30|狮子－百兽中最勇猛的、 无论遇见什么绝不退缩，
PROV|30|31|猎狗，公山羊， 和有整排士兵的君王。
PROV|30|32|你若行事愚顽，自高自傲， 或是设计恶谋，就当用手捂口。
PROV|30|33|搅动牛奶必成乳酪， 扭鼻子必出血， 照样，激发烈怒必挑起争端。
PROV|31|1|玛撒 王 利慕伊勒 的言语，就是他母亲教导他的 。
PROV|31|2|我儿，怎么了？ 我腹中生的儿，怎么了？ 我许愿而得的儿，怎么了？
PROV|31|3|不要将你的精力给妇女， 也不要有败坏君王的行为。
PROV|31|4|利慕伊勒 啊，君王不宜，君王不宜喝酒， 王子寻找烈酒也不相宜；
PROV|31|5|恐怕喝了就忘记所颁的法令， 颠倒所有困苦人的是非。
PROV|31|6|可以把烈酒给将亡的人喝， 把酒给心里愁苦的人喝，
PROV|31|7|让他喝了，就忘记他的贫穷， 不再记得他的苦楚。
PROV|31|8|你当为不能自辩的人 开口， 为所有孤独无助者伸冤。
PROV|31|9|你当开口按公义判断， 当为困苦和贫穷的人辩护。
PROV|31|10|才德的妇人谁能得着呢？ 她的价值远胜过宝石。
PROV|31|11|她丈夫心里信赖她， 必不缺少利益；
PROV|31|12|她终其一生， 使丈夫有益无损。
PROV|31|13|她寻找羊毛和麻， 欢喜用手做工。
PROV|31|14|她好像商船， 从远方运来粮食，
PROV|31|15|未到黎明她就起来， 把食物分给家中的人， 将当做的工分派女仆。
PROV|31|16|她想得田地，就去买来， 用手中的成果栽葡萄园。
PROV|31|17|她以能力束腰， 使膀臂有力。
PROV|31|18|她觉得自己获利不错， 她的灯终夜不灭。
PROV|31|19|她伸手拿卷线杆， 她的手掌把住纺车。
PROV|31|20|她张手赒济困苦人， 伸手帮助贫穷人。
PROV|31|21|她不因下雪为家里的人担心， 因为全家都穿上朱红衣服。
PROV|31|22|她为自己制作被单， 她的衣服是细麻和紫色布做的。
PROV|31|23|她丈夫在城门口与本地的长老同坐， 为人所认识。
PROV|31|24|她做细麻布衣裳来卖， 又将腰带卖给商家。
PROV|31|25|能力和威仪是她的衣服， 她想到日后的景况就喜笑。
PROV|31|26|她开口就发智慧， 她舌上有仁慈的教诲。
PROV|31|27|她管理家务， 并不吃闲饭。
PROV|31|28|她的儿女起来称她有福， 她的丈夫也称赞她：
PROV|31|29|“才德的女子很多， 惟独你超过一切。”
PROV|31|30|魅力是虚假的，美貌是虚浮的； 惟敬畏耶和华的妇女必得称赞。
PROV|31|31|她手中的成果你们要赏给她， 愿她的工作在城门口荣耀她。
ECCL|1|1|在 耶路撒冷 作王、 大卫 的儿子、传道者的言语。
ECCL|1|2|传道者说：虚空的虚空， 虚空的虚空，全是虚空。
ECCL|1|3|人一切的劳碌， 就是他在日光之下的劳碌，有什么益处呢？
ECCL|1|4|一代过去，一代又来， 地却永远长存。
ECCL|1|5|太阳上升，太阳下落， 急归所出之地。
ECCL|1|6|风往南刮，又向北转， 不停旋转，绕回原路。
ECCL|1|7|江河都往海里流，海却不满； 江河从何处流，仍归回原处。
ECCL|1|8|万事令人厌倦， 人不能说尽。 眼看，看不饱； 耳听，听不足。
ECCL|1|9|已有的事，后必再有； 已行的事，后必再行。 日光之下并无新事。
ECCL|1|10|有一件事人指着说：“看，这是新的！” 它在我们以前的世代早已有了。
ECCL|1|11|已过的事，无人记念； 将来的事，后来的人也不记念。
ECCL|1|12|我传道者在 耶路撒冷 作过 以色列 的王。
ECCL|1|13|我用智慧专心探寻、考察天下所发生的一切事：上帝给世人何等沉重的担子，使他们在其中劳苦！
ECCL|1|14|我见日光之下所发生的一切事，看哪，全是虚空，全是捕风。
ECCL|1|15|弯曲的，不能变直； 缺乏的，不计其数。
ECCL|1|16|我心里说：“看哪，我大有智慧，胜过在我以前所有统治 耶路撒冷 的人；我的心也多经历智慧和知识的事。”
ECCL|1|17|我专心想要明白智慧，想要明白狂妄与愚昧，方知这也是捕风。
ECCL|1|18|因为多有智慧，就多有愁烦； 增加知识，就增加忧伤。
ECCL|2|1|我心里说：“来吧，让我用喜乐试试你，使你享福！”看哪，这也是虚空。
ECCL|2|2|论嬉笑，我说：“这是狂妄。”论享乐，“这有什么用呢？”
ECCL|2|3|我心以智慧引导我，我心里探究，如何用酒使身体舒畅，如何抓住愚昧，直等我看明世人在天下短暂一生中，当行何事为美。
ECCL|2|4|我大兴土木，为自己建造房屋，栽葡萄园，
ECCL|2|5|修造庭园和公园，在其中栽种各样果树，
ECCL|2|6|挖造水池，用以灌溉林中的幼树。
ECCL|2|7|我买了仆婢，也有生在家中的仆婢；又有许多牛群羊群，胜过我以前所有在 耶路撒冷 的人。
ECCL|2|8|我为自己积蓄金银，搜集各君王、各省份的财宝；又为自己得男女歌手和世人所喜爱的物，以及一个又一个的妃嫔。
ECCL|2|9|这样，我就日渐昌盛，胜过我以前所有在 耶路撒冷 的人。我的智慧仍然存留。
ECCL|2|10|凡我眼所求的，我没有克制它；我心所乐的，我没有不享受。因我的心要为一切的劳碌快乐，这是我从一切劳碌中所得的报偿 。
ECCL|2|11|后来，我回顾我手所经营的一切和我劳碌所做的工。看哪，全是虚空，全是捕风；在日光之下毫无益处。
ECCL|2|12|我转而回顾智慧、狂妄和愚昧。在王以后来的人又如何呢？不过做先前所做的就是了。
ECCL|2|13|于是我看出智慧胜过愚昧，如同光明胜过黑暗。
ECCL|2|14|智慧人的眼目光明 ，愚昧人却在黑暗里行。但我知道他们都有相同的遭遇。
ECCL|2|15|我心里就说：“愚昧人所遇见的，我也一样遇见，那么我何必更有智慧呢？”我心里说：“这也是虚空。”
ECCL|2|16|智慧人和愚昧人一样，不会长久被人记念，因为日后都被遗忘。可叹！智慧人和愚昧人都一样会死亡。
ECCL|2|17|于是我恨恶生命，因为在日光之下所发生的事我都以为烦恼，全是虚空，全是捕风。
ECCL|2|18|我恨恶一切的劳碌，就是我在日光之下所劳碌的，因为我所得的必须留给我以后的人。
ECCL|2|19|那人是智慧是愚昧，谁能知道呢？他竟要掌管我在日光之下用智慧劳碌所得的。这也是虚空。
ECCL|2|20|我转想我在日光之下所劳碌的一切工作，心就绝望。
ECCL|2|21|因为有人用智慧、知识、灵巧劳碌工作，所得来的却要遗留给未曾劳碌的人作产业。这也是虚空，大大不幸。
ECCL|2|22|人一切的劳碌操心，就是他在日光之下所劳碌的，又得着了什么呢？
ECCL|2|23|他日日忧虑，他的劳苦成为愁烦，连夜间心也不得休息。这也是虚空。
ECCL|2|24|难道一个人有吃有喝，且在劳碌中享福，不是福气吗？我看这也是出于上帝的手。
ECCL|2|25|论到吃用、享福，谁能胜过我呢？
ECCL|2|26|上帝喜爱谁，就给谁智慧、知识和喜乐；惟有罪人，上帝使他劳苦，将他所储藏、所堆积的归给上帝所喜爱的人。这也是虚空，也是捕风。
ECCL|3|1|凡事都有定期， 天下每一事务都有定时。
ECCL|3|2|生有时，死有时； 栽种有时，拔出 有时；
ECCL|3|3|杀戮有时，医治有时； 拆毁有时，建造有时；
ECCL|3|4|哭有时，笑有时； 哀恸有时，跳舞有时；
ECCL|3|5|丢石头有时，捡石头有时； 怀抱有时，不抱有时；
ECCL|3|6|寻找有时，失落有时； 保存有时，抛弃有时；
ECCL|3|7|撕裂有时，缝补有时； 沉默有时，说话有时；
ECCL|3|8|喜爱有时，恨恶有时； 战争有时，和平有时。
ECCL|3|9|这样，做事的人在他所劳碌的事上得到什么益处呢？
ECCL|3|10|我观看上帝给世人的担子，使他们在其中劳苦：
ECCL|3|11|上帝造万物，各按其时成为美好，又将永恒安放在世人心里；然而上帝从始至终的作为，人不能测透。
ECCL|3|12|我知道，人除了终身喜乐纳福，没有一件幸福的事。
ECCL|3|13|并且人人吃喝，在他的一切劳碌中享福，这也是上帝的赏赐。
ECCL|3|14|我知道上帝所做的都必存到永远；无所增添，无所减少。上帝这样做，是要人在他面前存敬畏的心。
ECCL|3|15|现今的事以前就有了，将来的事也早已有了，并且上帝使已过的事重新再来 。
ECCL|3|16|我又见日光之下，应有公平之处有奸恶，应有公义之处也有奸恶。
ECCL|3|17|我心里说：“上帝必审判义人和恶人，因为在那里，各样事务，一切工作，都有定时。”
ECCL|3|18|我心里说：“为世人的缘故，上帝考验他们，让他们看见自己不过像走兽一样。”
ECCL|3|19|因为世人遭遇的，走兽也遭遇，所遭遇的都一样：这个怎样死，那个也怎样死，他们都有一样的气息。人不能强于走兽，全是虚空；
ECCL|3|20|都归一处，都是出于尘土，也都归于尘土。
ECCL|3|21|谁知道人的气息是往上升，走兽的气息是下入地呢？
ECCL|3|22|总而言之，人能够在他经营的事上喜乐，是最好不过了，因为这是他应得的报偿。他身后的事谁能领他回来看呢？
ECCL|4|1|我转而观看日光之下所发生的一切欺压之事。看哪，受欺压的流泪，无人安慰；欺压他们的有权势，也无人安慰。
ECCL|4|2|因此，我赞叹那已死的死人，胜过那还活着的活人。
ECCL|4|3|但那尚未出生，就是未曾见过日光之下所发生之恶事的，比这两种人更幸福。
ECCL|4|4|我见人因彼此嫉妒而有一切的劳碌和各样工作的成就，这也是虚空，也是捕风。
ECCL|4|5|愚昧人抱着双臂， 自食其肉。
ECCL|4|6|一掌满满而得享安静， 胜过两掌满满而劳碌捕风。
ECCL|4|7|我转而观看日光之下有一件虚空的事：
ECCL|4|8|有人孤单无双，无子无兄弟，竟劳碌不息，眼目也不以财富为满足。他说：“我劳碌，自己却不享福，到底是为了谁呢？”这也是虚空，是极沉重的担子。
ECCL|4|9|两个人总比一个人好，他们劳碌同得美好的报偿。
ECCL|4|10|若是跌倒，这人可以扶起他的同伴；倘若孤身跌倒，没有别人扶起他来，这人就有祸了。
ECCL|4|11|再者，二人同睡就都暖和，一人独睡怎能暖和呢？
ECCL|4|12|若遇敌攻击，孤身难挡，二人就能抵挡他；三股合成的绳子不易折断。
ECCL|4|13|贫穷而有智慧的年轻人，胜过年老不再纳谏的愚昧王，
ECCL|4|14|那人从监牢里出来作王，在国中原是出身贫寒。
ECCL|4|15|我见日光之下所有行走的活人，都跟随那年轻人，就是接续作王的那位。
ECCL|4|16|他的百姓，就是他所治理的众人，多得无数；但后来的人还是不喜欢他。这也是虚空，也是捕风。
ECCL|5|1|你到上帝的殿要谨慎你的脚步；近前听，胜过愚昧人献祭，他们不知道自己在作恶。
ECCL|5|2|在上帝面前你不可冒失开口，也不可心急发言；因为上帝在天上，你在地上，所以你的话语要少。
ECCL|5|3|事务多，令人做梦；话语多，显出愚昧。
ECCL|5|4|你向上帝许愿，还愿不可迟延，因他不喜欢愚昧人，你许的愿应当偿还。
ECCL|5|5|你许愿不还，不如不许。
ECCL|5|6|不可放任你的口使肉体犯罪，也不可在使者 面前说是错许了。为何使上帝因你的声音发怒，败坏你手所做的呢？
ECCL|5|7|多梦多言，其中多有虚空，你只要敬畏上帝。
ECCL|5|8|你若在一个地区看见穷人受欺压，公义公平被掠夺，不要因此惊奇；有一位高过居高位的在鉴察，在他们之上还有更高的。
ECCL|5|9|况且地的益处归众人，就是君王也受田地的供应。
ECCL|5|10|喜爱银子的，不因得银子满足；喜爱财富的，也不因得利益知足。这也是虚空。
ECCL|5|11|货物增添，吃的人也增添，物主得什么益处呢？不过眼看而已！
ECCL|5|12|劳碌的人不拘吃多吃少，睡得香甜；富人的丰足却不容他睡觉。
ECCL|5|13|我见日光之下有一件令人忧伤的祸患，就是财主积存财富，反害自己。
ECCL|5|14|他因遭遇不幸 ，财产尽失；他生了儿子，手里却一无所有。
ECCL|5|15|他怎样从母胎赤身而来，也必照样赤身而去；他所劳碌得来的，手中分毫不能带去。
ECCL|5|16|这是一件令人忧伤的祸患。他来的时候怎样，去的时候也必怎样。他为风劳碌有什么益处呢？
ECCL|5|17|并且他终身在黑暗中吃喝 ，多有烦恼、病痛和怒气。
ECCL|5|18|看哪，我所见为善为美的，就是人在上帝赐他一生的日子吃喝，享受日光之下劳碌得来的好处，因为这是他应得的报偿。
ECCL|5|19|而且，一个人蒙上帝赏赐财富与资产，又使他能享用，能获取自己当有的报偿 ，在他的劳碌中喜乐，这是上帝的赏赐。
ECCL|5|20|他不多思念自己一生的日子，因为上帝使他的心充满喜乐。
ECCL|6|1|我见日光之下有一件祸患重压在人身上，
ECCL|6|2|就是人蒙上帝赐他财富、资产和尊荣，以致他心里所愿的一样都不缺，只是上帝使他不能享用，反被外人享用。这是虚空，也是祸患。
ECCL|6|3|人若生一百个儿子，活许多岁数；他即使寿命很长，心里却不因福乐而满足，又不得埋葬；我说，那流掉的胎比他倒好。
ECCL|6|4|因为这胎虚虚而来，暗暗而去，名字被黑暗遮蔽，
ECCL|6|5|而且没有见过天日，什么都不知道，这胎比那人倒享安息。
ECCL|6|6|那人虽然活千年，再活千年，却不能享福；众人岂不都归同一个地方去吗？
ECCL|6|7|人的劳碌都为口腹，心里却不知足。
ECCL|6|8|智慧人比愚昧人有什么益处呢？困苦人在众人面前知道如何行，有什么益处呢？
ECCL|6|9|眼睛所看的比心里妄想的倒好。这也是虚空，也是捕风。
ECCL|6|10|先前所有的，早已起了名，人早知道人是如何的，不能与比自己强壮的相争。
ECCL|6|11|话语多，虚空也增多，这对人有什么益处呢？
ECCL|6|12|人一生虚度的日子，如影儿经过，谁知道什么才是对他有益呢？谁能告诉他身后在日光之下会发生什么事呢？
ECCL|7|1|名誉强如美好的膏油， 人死去的日子胜过他出生的日子。
ECCL|7|2|往丧家去， 强如往宴乐的家， 因为死是众人的结局， 活人必将这事放在心上。
ECCL|7|3|忧愁强如喜笑， 因为面带愁容，终必使心喜乐。
ECCL|7|4|智慧人的心在遭丧之家； 愚昧人的心在快乐之家。
ECCL|7|5|听智慧人的责备， 强如听愚昧人歌唱；
ECCL|7|6|因为愚昧人的笑声， 好像锅子下面烧荆棘的爆声， 这也是虚空。
ECCL|7|7|勒索使智慧人变为愚妄， 贿赂能败坏人的心。
ECCL|7|8|事情的终局强如它的起头； 存心忍耐的，胜过居心骄傲的。
ECCL|7|9|你的心不要急躁恼怒， 因为恼怒存在愚昧人的怀中。
ECCL|7|10|不要说： 为什么先前的日子强过现今的日子呢？ 你这样问不是出于智慧。
ECCL|7|11|智慧加上产业是美好的， 对见天日的人都有益处。
ECCL|7|12|因为智慧庇护人， 好像金钱庇护人一样； 智慧能保全智慧者的生命， 这就是知识的益处。
ECCL|7|13|你要观看上帝的作为， 谁能使他所弯曲的变直呢？
ECCL|7|14|顺利时要喜乐；患难时当思考。上帝使这两样都发生，因此，人不知将会发生什么事。
ECCL|7|15|在虚度的日子里，我见过各样的事情，义人在他的义中灭亡，恶人在他的恶中倒享长寿。
ECCL|7|16|不要行义过分，也不要过于自逞智慧，何必自取败亡呢？
ECCL|7|17|不要行恶过分，也不要为人愚昧，何必未到期而死呢？
ECCL|7|18|你持守这个，那个也不要松手才好。敬畏上帝的人，这一切都能兼得。
ECCL|7|19|智慧使拥有智慧的人比城中十个官长更有能力。
ECCL|7|20|其实世上没有行善而不犯罪的义人。
ECCL|7|21|人所说的话，你不要都放在心上，免得听见你的仆人诅咒你。
ECCL|7|22|因为你心里知道，自己也曾屡次诅咒别人。
ECCL|7|23|我曾用智慧试验这一切事，我说：“要得智慧。”智慧却离我远。
ECCL|7|24|万事之理遥不可及，太深奥，谁能测透呢？
ECCL|7|25|我转念，一心要知道，要考察，要寻求智慧和万事的来由，要知道邪恶为愚昧，愚昧为狂妄。
ECCL|7|26|我发现有一种妇人比死还苦毒：她本身是陷阱，她的心是罗网，手是锁链。凡蒙上帝喜爱的人必能躲开她；有罪的人却被她缠住了。
ECCL|7|27|传道者说：“你看，我考察一件又一件，为要寻求万事的来由，这是我所寻得的：
ECCL|7|28|我继续寻找，却未找到；一千当中，我找到一个男的，但在这一切当中，却找不到一个女的。
ECCL|7|29|你看，我所找到的只有一件，就是上帝造的人是正直的，但他们却寻出许多诡计。”
ECCL|8|1|谁如 智慧人呢？ 谁知道事情的解释呢？ 人的智慧使他的脸发光， 改变他脸上的暴戾之气 。
ECCL|8|2|我劝你 因上帝誓言的缘故，当遵守王的命令。
ECCL|8|3|不要急躁离开王的面前，不要固执行恶，因为他凡事都随自己心意而行。
ECCL|8|4|王的话本有权力，谁能对他说：“你在做什么？”
ECCL|8|5|凡遵守命令的，必不经历祸患；智慧人的心知道适当的时机和必经的过程。
ECCL|8|6|各样事务都有时机和过程，但人有苦难重压在身。
ECCL|8|7|他不知道将来的事，其实将来如何，谁能告诉他呢？
ECCL|8|8|没有人能掌握生命，将生命留住；也没有人有权力掌管死期。这场争战无人能免；邪恶也不能救那行邪恶的人。
ECCL|8|9|这一切我都见过，我专心考察日光之下所发生的一切事，有时这人管辖那人，令他受害。
ECCL|8|10|我见恶人埋葬；从前他们进出圣地，他们在城中的作为被人忘记。这也是虚空。
ECCL|8|11|判罪之后不立刻执行，所以世人满怀作恶的心思。
ECCL|8|12|罪人虽然作恶百次，倒享长寿；然而我也知道，福乐必临到敬畏上帝的人，就是在他面前心存敬畏的人。
ECCL|8|13|恶人却不得福乐，他的日子好像影儿不得长久，因为他不敬畏上帝。
ECCL|8|14|世上有一件虚空的事，就是义人所遭遇的，反而照恶人所做的；恶人所遭遇的，反而照义人所做的。我说，这也是虚空。
ECCL|8|15|我就称赞快乐，原来人在日光之下，最大的福气莫过于吃喝快乐；他在日光之下，上帝赐他一生的日子，要从劳碌中享受所得。
ECCL|8|16|我专心想要明白智慧，要观看世上所发生的事。有人昼夜不得阖眼睡觉。
ECCL|8|17|我观看上帝一切的作为，知道人不能探求日光之下所发生的事；任凭他费多少力探索，都找不出来，智慧人虽说他明白，仍不能找出来。
ECCL|9|1|我将这一切事放在心上，详细研究这些，就知道义人和智慧人，并他们的作为都在上帝手中；或是爱，或是恨，都在他们面前，但人不能知道。
ECCL|9|2|凡临到众人的际遇都一样：义人和恶人，好人 ，洁净的人和不洁净的人，献祭的和不献祭的，都一样。好人如何，罪人也如何；起誓的如何，怕起誓的也如何。
ECCL|9|3|在日光之下发生的一切事中有一件祸患，就是众人的际遇都一样，并且世人的心充满了恶；活着的时候心里狂妄，后来就归死人那里去了。
ECCL|9|4|与一切活人相连的，那人还有指望，因为活着的狗胜过死了的狮子。
ECCL|9|5|活着的人知道必死；死了的人毫无所知，也不再得赏赐，因为他们的名 已被遗忘。
ECCL|9|6|他们的爱，他们的恨，他们的嫉妒，早就消灭了。在日光之下所发生的一切事，他们永不再有份了。
ECCL|9|7|你只管欢欢喜喜吃你的饭，心中快乐喝你的酒，因为上帝已经悦纳你的作为。
ECCL|9|8|你的衣服要时时洁白，你头上也不要缺少膏油。
ECCL|9|9|在你一生虚空的日子，就是上帝赐你在日光之下虚空 的日子，当与你所爱的妻快活度日，因为那是你一生中在日光之下劳碌所得的报偿。
ECCL|9|10|凡你手所当做的事，要尽力去做；因为在你所必须去的阴间没有工作，没有谋算，没有知识，也没有智慧。
ECCL|9|11|我转而回顾日光之下，快跑的未必能赢，强壮的未必战胜，智慧的未必得粮食，聪明的未必得财富，有学问的未必得人喜悦，全在乎各人遇上的时候和机会。
ECCL|9|12|人不知道自己的定期。鱼被险恶的网圈住，鸟被罗网捉住，祸患的时刻忽然临到，世人陷在其中也是如此。
ECCL|9|13|我见日光之下有一样智慧，在我看来是伟大的，
ECCL|9|14|就是有一人口稀少的小城，遇大君王前来攻击，修筑营垒，将城围困。
ECCL|9|15|城中有一个贫穷的智慧人，他用智慧救了那城，却没有人记念那穷人。
ECCL|9|16|我就说，智慧胜过勇力；然而那贫穷人的智慧被人藐视，他的话也无人听从。
ECCL|9|17|宁可听智慧人安静的话语，不听掌权者在愚昧人中的喊声。
ECCL|9|18|智慧胜过打仗的兵器；但一个罪人能败坏许多善事。
ECCL|10|1|死苍蝇使做香的膏油散发臭气； 同样，一点愚昧也能压倒智慧和尊荣。
ECCL|10|2|智慧人的心居右； 愚昧人的心居左。
ECCL|10|3|愚昧人的行径显出无知， 对众人说，他是愚昧人。
ECCL|10|4|掌权者的怒气若向你发作， 不要离开你的本位， 因为镇定能平息大过。
ECCL|10|5|我见日光之下有一件祸患， 似乎出于统治者的错误，
ECCL|10|6|就是愚昧人立在高位； 有钱人却坐在低位。
ECCL|10|7|我见仆人骑马， 王子像仆人在地上步行。
ECCL|10|8|挖陷坑的，自己必陷在其中； 拆城墙的，自己必被蛇咬。
ECCL|10|9|开凿石头的，会受损伤； 劈开木头的，必遭危险。
ECCL|10|10|铁器钝了，若不将刃磨快，就必多费力气； 但智慧的益处在于使人成功。
ECCL|10|11|尚未行法术，蛇若咬人， 行法术的人就得不到什么好处了。
ECCL|10|12|智慧人的口说出恩言； 愚昧人的嘴吞灭自己，
ECCL|10|13|他口中的话语起头是愚昧， 终局是邪恶的狂妄。
ECCL|10|14|愚昧人多有话语。 人不知将来会发生什么事， 他身后的事谁能告诉他呢？
ECCL|10|15|愚昧人的劳碌使自己困乏， 连进城的路他也不知道。
ECCL|10|16|邦国啊，你的君王若年少， 你的群臣早晨宴乐， 你就有祸了！
ECCL|10|17|邦国啊，你的君王若是贵族之子， 你的群臣按时吃喝， 是为强身，不为酒醉， 你就有福了！
ECCL|10|18|因人懒惰，房顶塌下； 因人手懒，房屋滴漏。
ECCL|10|19|摆设宴席是为欢乐。 酒能使人快活， 钱能叫万事应心。
ECCL|10|20|不可诅咒君王， 连起意也不可， 在卧室里也不可诅咒富人； 因为空中的飞鸟必传扬这声音， 有翅膀的必述说这事。
ECCL|11|1|当将你的粮食撒在水面上， 因为日子久了，你必能得着它。
ECCL|11|2|将你所拥有的分给七人，或八人， 因为你不知道会有什么灾祸临到地上。
ECCL|11|3|云若满了雨，就必倾倒在地上。 树向南倒，或向北倒， 树倒在何处，就留在何处。
ECCL|11|4|看风的，必不撒种； 望云的，必不收割。
ECCL|11|5|你不知道气息如何进入孕妇的骨头里 ；照样，造万物之上帝的作为，你也无从得知。
ECCL|11|6|早晨要撒种，晚上也不要歇手，因为你不知道哪一样发旺；前者或后者，或两者都一样好。
ECCL|11|7|光是甜美的，眼见日光是多么好啊！
ECCL|11|8|人活多少年，就当快乐多少年，然而也当想到黑暗的日子；因为这样的日子必多，所要来临的全是虚空。
ECCL|11|9|年轻人哪，你在年少时当快乐；在年轻时使你的心欢畅，做你心所愿做的，看你眼所爱看的；却要知道，为这一切，上帝必审问你。
ECCL|11|10|所以，当从心中除掉愁烦，从肉体除去痛苦；因为年少和年轻之时，全是虚空。
ECCL|12|1|你趁着年轻、衰老的日子尚未来到，就是你所说，我毫无喜悦的那些岁月来临之前，当记念造你的主。
ECCL|12|2|不要等到太阳、光明、月亮、星宿变为黑暗，雨后云又返回；
ECCL|12|3|看守房屋的发颤，强壮的屈身，推磨的妇女因人少而停工，从窗户往外看的眼光变为昏暗；
ECCL|12|4|街门关闭，推磨的声音微小，鸟一叫，就惊醒，唱歌女子的声音也都微弱；
ECCL|12|5|人怕高处，路上有惊慌；杏树开花，蚱蜢成为重担，欲望不再挑起；因为人归他永远的家，吊丧的在街上往来。
ECCL|12|6|不要等到银链折断 ，金罐破裂，瓶子在泉旁损坏，水轮在井口断裂，
ECCL|12|7|尘土仍归于地，像原来一样，气息仍归于赐气息的上帝。
ECCL|12|8|传道者说：“虚空的虚空，全是虚空。”
ECCL|12|9|再者，传道者因有智慧，将知识教导众人；他思量，考察，并列举出许多箴言。
ECCL|12|10|传道者专心寻求可喜悦的言语，是凭正直写的诚实话。
ECCL|12|11|智慧人的话语如同刺棒；这些嘉言好像钉稳的钉子，都是一个牧者所赐的。
ECCL|12|12|我儿，还有一点，你当受劝戒：著书多，没有穷尽；读书多，身体疲倦。
ECCL|12|13|这些事都已听见了，结论就是：敬畏上帝，谨守他的诫命，这是人当尽的本分。
ECCL|12|14|因为人所做的事，连一切隐藏的事，无论是善是恶，上帝都必审问。
SONG|1|1|所罗门 的雅歌 。
SONG|1|2|愿他用口与我亲吻。 你的爱情比酒更美，
SONG|1|3|你的膏油馨香， 你的名如倾泻而出的香膏， 所以童女都爱你。
SONG|1|4|愿你吸引我跟随你；让我们快跑吧！ 王领我进入他的内室。 我们必因你欢喜快乐， 我们要思念你的爱情， 胜似思念美酒。 她们爱你是理所当然的。
SONG|1|5|耶路撒冷 的女子啊， 我虽然黑，却是秀美， 如同 基达 的帐棚， 好像 所罗门 的幔子，
SONG|1|6|不要因太阳把我晒黑了就瞪着我。 我母亲的儿子向我发怒， 他们使我看守葡萄园； 我自己的葡萄园我却没有看守。
SONG|1|7|我心所爱的啊，请告诉我， 你在何处牧羊？ 正午在何处使羊歇卧？ 我何必像蒙着脸的女子 在你同伴的羊群旁边呢？
SONG|1|8|你这女子中最美丽的， 你若不知道， 只管跟随羊群的脚踪行， 在牧人的帐棚边，牧放你的小山羊。
SONG|1|9|我的佳偶， 你好比法老战车上的骏马。
SONG|1|10|你的两颊因发辫而秀美， 你的颈项因珠串而华丽。
SONG|1|11|我们要为你编上金链，镶上银饰。
SONG|1|12|王正坐席的时候， 我的哪哒香膏散发香味。
SONG|1|13|我的良人好像一袋没药， 在我胸怀中。
SONG|1|14|我的良人好像一束凤仙花， 在 隐．基底 的葡萄园中。
SONG|1|15|看哪，我的佳偶，你真美丽！ 看哪，你真美丽！你的眼睛是鸽子。
SONG|1|16|看哪，我的良人，你多英俊可爱！ 让我们以青草为床榻，
SONG|1|17|以香柏树为房子的栋梁， 以松树作屋顶的椽木。
SONG|2|1|我是 沙仑 的玫瑰花， 是谷中的百合花。
SONG|2|2|我的佳偶在女子中， 好像荆棘里的百合花。
SONG|2|3|我的良人在男子中， 如同苹果树在树林里。 我欢欢喜喜坐在他的荫下， 尝他果子的滋味，觉得甘甜。
SONG|2|4|他领我进入宴会厅， 为我插上爱的旗帜。
SONG|2|5|请你们用葡萄饼增补我力， 以苹果畅快我的心， 因我为爱而生病。
SONG|2|6|他的左手在我头下， 他的右手将我环抱。
SONG|2|7|耶路撒冷 的女子啊， 我指着羚羊或田野的母鹿嘱咐你们， 不要唤醒，不要挑动爱情，等它自发。
SONG|2|8|听啊！我良人的声音， 看哪！他穿山越岭而来。
SONG|2|9|我的良人像羚羊，像小鹿。 看哪，他站在我们的墙壁边， 从窗户往里观看， 从窗格子往里窥探。
SONG|2|10|我的良人对我说： “我的佳偶，起来！ 我的美人，与我同去！
SONG|2|11|看哪，因为冬天已逝， 雨水止住，已经过去了。
SONG|2|12|地上百花开放， 歌唱的时候到了， 斑鸠的声音在我们境内也听见了。
SONG|2|13|无花果树的果子渐渐成熟， 葡萄树开花，散发香气。 我的佳偶，起来！ 我的美人，与我同去！
SONG|2|14|我的鸽子啊，你在磐石穴中， 在陡岩的隐密处。 求你容我得见你的面貌， 求你容我得听你的声音； 因你的声音悦耳， 你的容貌秀美。
SONG|2|15|请为我们擒拿狐狸， 就是毁坏葡萄园的小狐狸， 我们的葡萄正在开花。”
SONG|2|16|我的良人属我，我也属他， 他在百合花中放牧。
SONG|2|17|我的良人哪， 等到天起凉风、 日影飞去的时候， 愿你归回，像羚羊， 像小鹿，在崎岖的山 上。
SONG|3|1|我夜间躺卧在床上， 寻找我心所爱的； 我寻找他，却寻不着。
SONG|3|2|“我要起来，绕行城中， 在街市上，在广场上， 寻找我心所爱的。” 我寻找他，却寻不着。
SONG|3|3|城中巡逻的守卫遇见我， “你们看见我心所爱的没有？”
SONG|3|4|我刚离开他们，就遇见我心所爱的。 我拉住他，不放他走， 领他进入我母亲的家， 到怀我者的内室。
SONG|3|5|耶路撒冷 的女子啊， 我指着羚羊或田野的母鹿嘱咐你们， 不要唤醒，不要挑动爱情，等它自发。
SONG|3|6|那如烟柱从旷野上来， 薰了没药、乳香，扑上商人各样香粉的是谁呢？
SONG|3|7|看哪，是 所罗门 的轿， 周围有六十个勇士， 都是 以色列 中的勇士。
SONG|3|8|他们的手都持刀，善于争战， 各人腰间佩刀，防备夜间恐怖的攻击。
SONG|3|9|所罗门 王用 黎巴嫩 木 为自己制作轿子。
SONG|3|10|轿柱是用银做的， 轿底是用金做的， 坐垫是紫色的， 其中所铺的是 耶路撒冷 女子的爱情。
SONG|3|11|锡安的女子啊， 你们要出去观看 所罗门 王！ 他头戴冠冕，就是在他结婚当天 心中喜乐的时候，他母亲给他戴上的。
SONG|4|1|看哪，我的佳偶，你真美丽！看哪，你真美丽！ 你的眼睛在面纱后好像鸽子。 你的头发如同一群山羊，从 基列山 下来。
SONG|4|2|你的牙齿如新剪毛的一群母羊，洗净之后走上来， 它们成对，没有一颗是单独的。
SONG|4|3|你的唇好像一条朱红线， 你的嘴秀美。 你的鬓角在面纱后， 如同迸开的石榴。
SONG|4|4|你的颈项犹如 大卫 为收藏军器而造的高塔， 其上悬挂一千个盾牌， 都是勇士的盾牌。
SONG|4|5|你的两乳好像百合花中吃草的一对小鹿， 是母鹿双生的。
SONG|4|6|我要往没药山和乳香冈去， 直到天起凉风、 日影飞去的时候。
SONG|4|7|我的佳偶，你全然美丽， 毫无瑕疵！
SONG|4|8|我的新娘，请你与我一同离开 黎巴嫩 ， 与我一同离开 黎巴嫩 。 从 亚玛拿 山巅， 从 示尼珥 ，就是 黑门山 顶， 从狮子的洞， 从豹子的山往下观看。
SONG|4|9|我的妹子，我的新娘， 你夺了我的心。 你明眸一瞥， 你颈项的链子， 夺了我的心！
SONG|4|10|我的妹子，我的新娘， 你的爱情 何其美！ 你的爱情比酒甜美！ 你膏油的馨香胜过一切香料！
SONG|4|11|我的新娘，你的唇滴下蜂蜜， 你的舌下有蜜，有奶。 你衣服的香气宛如 黎巴嫩 的芬芳。
SONG|4|12|我的妹子，我的新娘 是上锁的园子， 是禁闭的园子 ， 是封闭的泉源。
SONG|4|13|你园内所种的结了石榴， 有佳美的果子， 并凤仙花与哪哒树。
SONG|4|14|有哪哒和番红花， 香菖蒲和桂树， 并各样乳香木、没药、沉香， 与一切上等的香料。
SONG|4|15|你是园中的泉，活水的井， 是从 黎巴嫩 涌流而下的溪水。
SONG|4|16|北风啊，兴起！ 南风啊，吹来！ 吹在我的园内， 使其中的香气散发出来。 愿我的良人进入自己园里， 吃他佳美的果子。
SONG|5|1|我的妹子，我的新娘， 我进入我的园中， 采了我的没药和香料， 吃了我的蜂房和蜂蜜， 喝了我的酒和奶。 我的朋友，请吃！ 我亲爱的，请喝，多多地喝！
SONG|5|2|我身躺卧，我心却醒。 这是我良人的声音； 他敲门： “我的妹子，我的佳偶， 我的鸽子，我完美的人儿， 请你为我开门； 因我的头沾满露水， 我的发被夜露滴湿。”
SONG|5|3|我脱了衣裳，怎能再穿上呢？ 我洗了脚，怎可再弄脏呢？
SONG|5|4|我的良人从门缝里伸进他的手， 我便因他动了心。
SONG|5|5|我起来，要为我的良人开门。 我的两手滴下没药， 我的指头有没药汁滴在门闩上。
SONG|5|6|我为我的良人开了门， 我的良人却已转身走了。 他说话的时候，我魂不守舍。 我寻找他，竟寻不着， 我呼叫他，他却不回答。
SONG|5|7|城中巡逻的守卫遇见我， 打了我，伤了我， 看守城墙的人夺去我的披肩。
SONG|5|8|耶路撒冷 的女子啊，我嘱咐你们： 若遇见我的良人， 要告诉他，我为爱而生病。
SONG|5|9|你这女子中最美丽的， 你的良人有什么胜过别的良人呢？ 你的良人有什么胜过别的良人， 使你这样嘱咐我们？
SONG|5|10|我的良人红润发亮， 超乎万人之上。
SONG|5|11|他的头像千足的纯金， 他的发绺卷曲，黑如乌鸦。
SONG|5|12|他的眼如溪水旁的鸽子， 沐浴在奶中，安得合式 。
SONG|5|13|他的两颊如香花园， 如香草台 ； 他的嘴唇像百合花， 滴下没药汁。
SONG|5|14|他的双手宛如金条， 镶嵌水苍玉； 他的身体如同雕刻的象牙， 周围镶嵌蓝宝石。
SONG|5|15|他的腿好比白玉石柱， 安在精金座上； 他的容貌如 黎巴嫩 ， 佳美如香柏树。
SONG|5|16|他的口甘甜， 他全然可爱。 耶路撒冷 的女子啊， 这是我的良人， 这是我的朋友。
SONG|6|1|你这女子中最美丽的， 你的良人往何处去？ 你的良人转向何处去了？ 我们好与你同去寻找他。
SONG|6|2|我的良人进入自己园中， 到香花园， 在园内放牧， 采百合花。
SONG|6|3|我属我的良人， 我的良人属我； 他在百合花中放牧。
SONG|6|4|我的佳偶啊，你美丽如 得撒 ， 秀美如 耶路撒冷 ， 威武如展开旌旗的军队。
SONG|6|5|求你转开眼睛不要看我， 因你的眼睛使我慌乱。 你的头发如同一群山羊，从 基列山 下来。
SONG|6|6|你的牙齿如一群母羊，洗净之后走上来， 它们成对，没有一颗是单独的。
SONG|6|7|你的鬓角在面纱后， 如同迸开的石榴。
SONG|6|8|虽有六十王后、八十妃嫔， 并有无数的童女。
SONG|6|9|她是我独一的鸽子、我完美的人儿， 是她母亲独生的， 是生养她的所宠爱的。 女子见了都称她有福， 王后妃嫔见了也赞美她。
SONG|6|10|那俯视如晨曦、 美丽如月亮、皎洁如太阳、 威武如展开旌旗军队的是谁呢？
SONG|6|11|我下到坚果园， 要看谷中青翠的植物， 要看葡萄可曾发芽， 石榴可曾放蕊；
SONG|6|12|不知不觉， 我仿佛坐在我百姓高官 的战车中。
SONG|6|13|回来，回来， 书拉密 的女子； 回来，回来，我们要看你。 你们为何要观看 书拉密 的女子， 像观看两队人马在跳舞 呢？
SONG|7|1|尊贵的女子啊，你的脚在鞋中何等秀美！ 你的大腿圆润，好像美玉， 是巧匠的手做成的。
SONG|7|2|你的肚脐如圆杯， 不缺调和的酒。 你的肚子如一堆麦子， 周围有百合花。
SONG|7|3|你的两乳好像一对小鹿， 是母鹿双生的。
SONG|7|4|你的颈项如象牙塔， 你的眼睛像 希实本 、 巴特．拉并 门旁的水池， 你的鼻子仿佛朝向 大马士革 的 黎巴嫩 塔。
SONG|7|5|你的头在你身上好像 迦密山 ， 你头上的发呈紫色， 王被这发绺系住了。
SONG|7|6|我亲爱的，喜乐的女子啊， 你何等美丽！何等令人喜悦！
SONG|7|7|你的身材好像棕树， 你的两乳如同累累的果实。
SONG|7|8|我说：我要爬上棕树，抓住枝子。 愿你的两乳好像葡萄累累， 愿你鼻子的香气如苹果；
SONG|7|9|你的上颚如美酒， 直流入我良人的口里， 流入沉睡者的口中 。
SONG|7|10|我属我的良人， 他也恋慕我。
SONG|7|11|来吧！我的良人， 让我们往田间去， 在村庄住宿。
SONG|7|12|早晨让我们起来往葡萄园去， 看葡萄树发芽没有， 花开了没有， 石榴放蕊没有， 在那里我要将我的爱情给你。
SONG|7|13|曼陀罗草 散发香味， 在我们的门内有各样新陈佳美的果子； 我的良人，这都是我为你保存的。
SONG|8|1|惟愿你像我的兄弟， 像吃我母亲奶的兄弟。 我在外头遇见你就与你亲吻， 谁也不轻看我。
SONG|8|2|我必引导你， 领你进入我母亲的家， 她必教导我， 我必使你喝石榴汁酿的香酒。
SONG|8|3|他的左手在我头下， 他的右手将我环抱。
SONG|8|4|耶路撒冷 的女子啊， 我嘱咐你们， 不要唤醒、不要挑动爱情，等它自发。
SONG|8|5|那靠着良人从旷野上来的是谁呢？ 在苹果树下，我叫醒了你； 在那里，你母亲曾为了生你而阵痛， 在那里，生你的为你阵痛。
SONG|8|6|求你将我放在你心上如印记， 带在你臂上如戳记。 因为爱情如死之坚强， 热恋如阴间之牢固， 所发的光是火焰的光， 是极其猛烈的火焰 。
SONG|8|7|爱情，众水不能熄灭， 江河也不能淹没。 若有人拿家中所有的财宝要换爱情， 就全被藐视。
SONG|8|8|我们有一小妹， 她还没有乳房， 人来提亲的日子， 我们当为她怎么办呢？
SONG|8|9|她若是墙， 我们要在其上建造银塔； 她若是门， 我们要用香柏木板围护她。
SONG|8|10|我是墙， 我的两乳像塔。 那时，我在他眼中是找到平安的人。
SONG|8|11|所罗门 在 巴力．哈们 有一葡萄园， 他将这葡萄园租给看守的人， 每人为其中的果子要交一千银子。
SONG|8|12|我有属自己的葡萄园。 所罗门 哪，一千归你， 两百归看守果子的人。
SONG|8|13|你这住在园中的， 同伴都要听你的声音， 求你使我也得以听见。
SONG|8|14|我的良人哪，求你快来！ 像羚羊，像小鹿，在香草山上。
ISA|1|1|当 乌西雅 、 约坦 、 亚哈斯 、 希西家 作 犹大 王的时候， 亚摩斯 的儿子 以赛亚 见异象，论到 犹大 和 耶路撒冷 。
ISA|1|2|天哪，要听！地啊，侧耳而听！ 因为耶和华说： “我养育儿女，将他们养大， 他们竟悖逆我。
ISA|1|3|牛认识主人， 驴认识主人的槽； 以色列 却不认识， 我的民却不明白。”
ISA|1|4|祸哉！犯罪的国民， 担着罪孽的百姓， 行恶的族类， 败坏的儿女！ 他们离弃耶和华， 藐视 以色列 的圣者， 背向他，与他疏远。
ISA|1|5|你们为什么屡次悖逆，继续受责打呢？ 你们已经满头疼痛， 全心发昏；
ISA|1|6|从脚掌到头顶， 没有一处是完好的， 尽是创伤、瘀青，与流血的伤口， 未曾挤净，未曾包扎， 也没有用膏滋润。
ISA|1|7|你们的土地荒芜， 城镇被火烧毁； 你们的田地在你们眼前被陌生人侵吞， 既被陌生人倾覆，就成为荒芜 。
ISA|1|8|仅存的 锡安 ， 好似葡萄园的草棚， 如瓜田中的茅屋， 又如被围困的城。
ISA|1|9|若不是万军之耶和华为我们留下一些幸存者， 我们早已变成 所多玛 ，像 蛾摩拉 一样了。
ISA|1|10|所多玛 的官长啊， 你们要听耶和华的言语！ 蛾摩拉 的百姓啊， 要侧耳听我们上帝的教诲！
ISA|1|11|耶和华说： “你们许多的祭物于我何益呢？ 公绵羊的燔祭和肥畜的油脂， 我已经腻烦了； 公牛、羔羊、公山羊的血， 我都不喜悦。
ISA|1|12|“你们来朝见我， 谁向你们的手要求这些， 使你们践踏我的院宇呢？
ISA|1|13|不要再献无谓的供物了， 香是我所憎恶的。 我不能容忍行恶又守严肃会： 初一、安息日和召集的大会。
ISA|1|14|你们的初一和节期，我心里恨恶， 它们成了我的重担， 担当这些，令我厌烦。
ISA|1|15|你们举手祷告，我必遮眼不看， 就算你们多多祈祷，我也不听； 你们的手沾满了血。
ISA|1|16|你们要洗涤、自洁， 从我眼前除掉恶行； 要停止作恶，
ISA|1|17|学习行善， 寻求公平， 帮助受欺压的 ， 替孤儿伸冤， 为寡妇辩护。”
ISA|1|18|耶和华说： “来吧，我们彼此辩论。 你们的罪虽像朱红，必变成雪白； 虽红如丹颜，必白如羊毛。
ISA|1|19|你们若甘心听从， 必吃地上的美物；
ISA|1|20|若不听从，反倒悖逆， 必被刀剑吞灭； 这是耶和华亲口说的。”
ISA|1|21|忠信的城竟然变为妓女！ 从前充满了公平， 公义居在其中， 现今却有凶手居住。
ISA|1|22|你的银子变为渣滓， 你的酒用水冲淡。
ISA|1|23|你的官长悖逆， 与盗贼为伍， 全都喜爱贿赂， 追求赃物； 他们不为孤儿伸冤， 寡妇的案件也呈不到他们面前。
ISA|1|24|因此，主－万军之耶和华、 以色列 的大能者说： “唉！我要向我的对头雪恨， 向我的敌人报仇。
ISA|1|25|我必反手对付你， 如碱炼净你的渣滓， 除尽你的杂质。
ISA|1|26|我必回复你的审判官，像起初一样， 回复你的谋士，如起先一般。 然后，你必称为公义之城， 忠信之邑。”
ISA|1|27|锡安 必因公平得蒙救赎， 其中归正的人必因公义得蒙救赎。
ISA|1|28|但悖逆的和犯罪的必一同败亡， 离弃耶和华的必致消灭。
ISA|1|29|那等人必因所喜爱的圣树抱愧； 你们必因所选择的园子 蒙羞，
ISA|1|30|因为你们必如叶子枯干的橡树， 如无水的园子。
ISA|1|31|有权势的必如麻线， 他的作为好像火花， 都要一同焚烧，无人扑灭。
ISA|2|1|亚摩斯 的儿子 以赛亚 所见，有关 犹大 和 耶路撒冷 的事。
ISA|2|2|末后的日子，耶和华殿的山必坚立， 超乎诸山，高举过于万岭； 万国都要流归这山。
ISA|2|3|必有许多民族前往，说： “来吧，我们登耶和华的山， 到 雅各 上帝的殿。 他必将他的道教导我们， 我们也要行他的路。” 因为教诲必出于 锡安 ， 耶和华的言语必出于 耶路撒冷 。
ISA|2|4|他必在万国中施行审判， 为许多民族断定是非。 他们要将刀打成犁头， 把枪打成镰刀； 这国不举刀攻击那国， 他们也不再学习战事。
ISA|2|5|雅各 家啊， 来吧！让我们在耶和华的光明中行走。
ISA|2|6|你离弃了你的百姓 雅各 家， 因为他们充满了东方的习俗 ， 又像 非利士 人一样观星象， 并与外邦人击掌。
ISA|2|7|他们的国满了金银， 财宝也无穷； 他们的地满了马匹， 战车也无数。
ISA|2|8|他们的地满了偶像； 他们跪拜自己手所造的， 就是自己手指所做的。
ISA|2|9|有人屈膝， 有人下跪； 所以，不要饶恕他们。
ISA|2|10|当进入磐石，藏在土中， 躲避耶和华的惊吓和他威严的荣光。
ISA|2|11|到那日，眼目高傲的必降卑， 狂妄的人必屈膝； 惟独耶和华被尊崇。
ISA|2|12|因万军之耶和华的一个日子 要临到所有骄傲狂妄的， 临到一切自高的， 使他们降为卑；
ISA|2|13|临到 黎巴嫩 高大的香柏树、 巴珊 的橡树，
ISA|2|14|临到一切高山、 一切峻岭，
ISA|2|15|临到一切碉堡、 一切坚固的城墙，
ISA|2|16|临到 他施 一切的船只、 一切华丽的船艇。
ISA|2|17|人的骄傲必屈膝， 人的狂妄必降卑； 在那日，惟独耶和华被尊崇，
ISA|2|18|偶像必全然废弃。
ISA|2|19|耶和华兴起使地大震动的时候， 人就进入石洞和土穴里， 躲避耶和华的惊吓和他威严的荣光。
ISA|2|20|到那日，人必将造来敬拜的金偶像、银偶像 抛给田鼠和蝙蝠。
ISA|2|21|耶和华兴起使地大震动的时候， 人就进入磐缝和岩隙里， 躲避耶和华的惊吓和他威严的荣光。
ISA|2|22|你们不要倚靠世人， 他只不过鼻孔里有气息， 算得了什么呢？
ISA|3|1|看哪，主－万军之耶和华要从 耶路撒冷 和 犹大 除掉众人所倚靠的，所仰赖的， 就是所倚靠的粮，所仰赖的水；
ISA|3|2|除掉勇士和战士， 审判官和先知， 占卜的和长老，
ISA|3|3|除掉五十夫长和显要、 谋士和巧匠， 以及擅长法术的人。
ISA|3|4|我必使孩童作他们的领袖， 幼儿管辖他们。
ISA|3|5|百姓要彼此欺压， 各人欺压邻舍； 青年要侮慢老人， 卑贱的要侮慢尊贵的。
ISA|3|6|人在父家拉住自己的兄弟： “你有外衣，来作我们的官长， 让这些败坏的事归于你的手下吧！”
ISA|3|7|那时，他必扬声说： “我不作医治你们的人； 我家里没有粮食，也没有衣服， 你们不可立我作百姓的官长。”
ISA|3|8|耶路撒冷 败落， 犹大 倾倒； 因为他们的舌头和行为与耶和华相悖， 无视于他荣光的眼目。
ISA|3|9|他们的脸色证明自己不正， 他们述说自己像 所多玛 一样的罪恶，毫不隐瞒。 他们有祸了！因为作恶自害。
ISA|3|10|你们要对义人说，他是有福的， 因为他必吃自己行为所结的果实。
ISA|3|11|恶人有祸了！他必遭灾难！ 因为他要按自己手所做的受报应。
ISA|3|12|至于我的百姓， 统治者剥削你们， 放高利贷的人管辖你们 。 我的百姓啊，引导你的使你走错， 并毁坏你所行的道路。
ISA|3|13|耶和华兴起诉讼， 站着审判万民。
ISA|3|14|耶和华必审问他国中的长老和领袖： “你们，你们摧毁葡萄园， 抢夺困苦人，囤积在你们家中。
ISA|3|15|你们为何压碎我的百姓， 碾磨困苦人的脸呢？” 这是万军之主耶和华说的。
ISA|3|16|耶和华说： 因为 锡安 狂傲， 行走挺项，卖弄眼目， 俏步徐行，脚下玎珰，
ISA|3|17|主必使 锡安 头顶长疮， 耶和华又暴露其下体。
ISA|3|18|到那日，主必除掉华美的足饰、额带、月牙圈、
ISA|3|19|耳环、手镯、面纱、
ISA|3|20|头巾、足链、华带、香盒、符囊、
ISA|3|21|戒指、鼻环、
ISA|3|22|礼服、外套、披肩、皮包、
ISA|3|23|手镜、细麻衣、头饰、纱巾。
ISA|3|24|必有腐烂代替馨香， 绳子代替腰带， 光秃代替美发， 麻衣系腰代替华服， 烙痕代替美貌。
ISA|3|25|你的男丁必倒在刀下， 你的勇士必死在阵上。
ISA|3|26|锡安 的城门必悲伤、哀号； 它必荒凉，坐在地上。
ISA|4|1|在那日，七个女人必拉住一个男人，说：“我们吃自己的食物，穿自己的衣服，但求你允许我们归你名下，除掉我们的羞耻。”
ISA|4|2|在那日，耶和华的苗必华美尊荣，地的出产必成为幸存的 以色列 民的骄傲和光荣。
ISA|4|3|主以公平的灵和焚烧的灵洗净 锡安 居民 的污秽，又除净在 耶路撒冷 流人血的罪。那时，剩在 锡安 、留在 耶路撒冷 的，就是一切住 耶路撒冷 、在生命册上记名的，必称为圣。
ISA|4|4|
ISA|4|5|耶和华必在整座 锡安山 ，在会众之上，白天造云，黑夜发出烟和火焰的光，因为在一切荣耀之上必有华盖；
ISA|4|6|这要作为棚子，白天可以遮荫避暑，暴风雨侵袭时，可作藏身处和避难所。
ISA|5|1|我要为我亲爱的唱歌， 我所爱的、他的葡萄园之歌。 我亲爱的有葡萄园 在肥沃的山冈上。
ISA|5|2|他刨挖园子，清除石头， 栽种上等的葡萄树， 在园中盖了一座楼， 又凿出酒池； 指望它结葡萄， 反倒结了野葡萄。
ISA|5|3|耶路撒冷 的居民和 犹大 人哪， 现在，请你们在我与我的葡萄园之间断定是非。
ISA|5|4|我为我葡萄园所做的之外， 还有什么可做的呢？ 我指望它结葡萄， 怎么倒结了野葡萄呢？
ISA|5|5|现在我告诉你们， 我要向我的葡萄园怎么做。 我必撤去篱笆，使它被烧毁； 拆毁围墙，使它被践踏。
ISA|5|6|我必使它荒废，不再修剪， 不再锄草，任荆棘蒺藜生长； 我也必吩咐密云， 不再降雨在其上。
ISA|5|7|万军之耶和华的葡萄园就是 以色列 家； 他所喜爱的树就是 犹大 人。 他指望公平， 看哪，却有流血； 指望公义， 看哪，却有冤声。
ISA|5|8|祸哉！你们以房接房， 以地连地， 以致不留余地， 只顾自己独居境内。
ISA|5|9|我耳闻万军之耶和华说： “许多房屋必然荒废； 宏伟华丽，无人居住。
ISA|5|10|十亩 的葡萄园只酿出一罢特的酒， 一贺梅珥的谷种只结一伊法粮食。”
ISA|5|11|祸哉！那些清晨早起，追寻烈酒， 因酒狂热，流连到深夜的人，
ISA|5|12|他们在宴席上 弹琴，鼓瑟，击鼓，吹笛，饮酒， 却不留意耶和华的作为， 也不留心他手所做的。
ISA|5|13|所以，我的百姓因无知就被掳去； 尊贵的人甚是饥饿， 平民也极其干渴。
ISA|5|14|因此，阴间胃口 大开， 张开无限量的口； 令 耶路撒冷 的贵族与平民、狂欢的与作乐的人 都掉落其中。
ISA|5|15|人为之屈膝， 人就降为卑； 高傲的眼目也降为卑。
ISA|5|16|惟有万军之耶和华因公平显为崇高， 神圣的上帝因公义显为圣。
ISA|5|17|羔羊必来吃草，如同在自己的草场； 在富有人的废墟，流浪的牲畜也来吃 。
ISA|5|18|祸哉！那些以虚假的绳子牵引罪孽， 以套车的绳索紧拉罪恶的人。
ISA|5|19|他们说： “任 以色列 的圣者急速前行，快快成就他的作为， 好让我们看看； 任他的筹算临近成就， 好使我们知道。”
ISA|5|20|祸哉！那些称恶为善，称善为恶， 以暗为光，以光为暗， 以苦为甜，以甜为苦的人。
ISA|5|21|祸哉！那些在自己眼中有智慧， 在自己面前有通达的人。
ISA|5|22|祸哉！那些以饮酒称雄， 以调烈酒称霸的人。
ISA|5|23|他们因受贿赂，就称恶人为义， 将义人的义夺去。
ISA|5|24|火苗怎样吞灭碎秸， 干草怎样落在火焰之中， 照样，他们的根必然腐朽， 他们的花像灰尘扬起； 因为他们厌弃万军之耶和华的教诲， 藐视 以色列 圣者的言语。
ISA|5|25|因此，耶和华的怒气向他的百姓发作。 他伸手攻击他们，山岭就震动； 他们的尸首在街市上好像粪土。 虽然如此，他的怒气并未转消， 他的手依然伸出。
ISA|5|26|他必竖立大旗，召集远方的国民， 把他们从地极叫来。 看哪，他们必急速奔来，
ISA|5|27|其中没有疲倦的，绊跌的； 没有打盹的，睡觉的； 腰带并不放松， 鞋带也不拉断。
ISA|5|28|他们的箭锐利， 弓也上了弦； 马蹄如坚石， 车轮像旋风。
ISA|5|29|他们要吼叫，像母狮， 咆哮，像少壮狮子； 他们要咆哮，抓取猎物， 稳稳叼走，无人能救回。
ISA|5|30|那日，他们要向 以色列 人咆哮， 像海浪澎湃； 人若望地，看哪，只有黑暗与祸患， 光明因密云而变黑暗。
ISA|6|1|当 乌西雅 王崩的那年，我看见主坐在高高的宝座上。他的衣裳下摆遮满圣殿。
ISA|6|2|上有撒拉弗侍立，各有六个翅膀：两个翅膀遮脸，两个翅膀遮脚，两个翅膀飞翔，
ISA|6|3|彼此呼喊说： “圣哉！圣哉！圣哉！万军之耶和华； 他的荣光遍满全地！”
ISA|6|4|因呼喊者的声音，门槛的根基震动，殿里充满了烟云。
ISA|6|5|那时我说：“祸哉！我灭亡了！因为我是嘴唇不洁的人，住在嘴唇不洁的民中，又因我亲眼看见大君王－万军之耶和华。”
ISA|6|6|有一撒拉弗向我飞来，手里拿着烧红的炭，是用火钳从坛上取下来的，
ISA|6|7|用炭沾我的口，说：“看哪，这炭沾了你的嘴唇，你的罪孽便除掉，你的罪恶就赦免了。”
ISA|6|8|我听见主的声音说：“我可以差遣谁呢？谁肯为我们去呢？”我说：“我在这里，请差遣我！”
ISA|6|9|他说：“你去告诉这百姓说： ‘你们听了又听，却不明白； 看了又看，却不晓得。’
ISA|6|10|要使这百姓心蒙油脂， 耳朵发沉， 眼睛昏花； 恐怕他们眼睛看见， 耳朵听见， 心里明白， 回转过来，就得医治。”
ISA|6|11|我就说：“主啊，这到几时为止呢？”他说： “直到城镇荒凉，无人居住， 房屋空无一人，土地极其荒芜；
ISA|6|12|耶和华将人迁到远方， 国内被撇弃的土地很多。
ISA|6|13|国内剩下的人若还有十分之一， 也必被吞灭。 然而如同大树与橡树，虽被砍伐， 残干却仍存留， 圣洁的苗裔是它的残干。”
ISA|7|1|乌西雅 的孙子， 约坦 的儿子， 犹大 王 亚哈斯 在位的时候， 亚兰 王 利汛 和 利玛利 的儿子 以色列 王 比加 上来攻打 耶路撒冷 ，却不能攻取。
ISA|7|2|有人告诉 大卫 家说：“ 亚兰 与 以法莲 已经结盟。”王的心和百姓的心就都颤动，好像林中的树被风吹动一样。
ISA|7|3|耶和华对 以赛亚 说：“你和你的儿子 施亚．雅述 要出去，到 上池 的水沟尽头，往漂布地的大路上，迎见 亚哈斯 ，
ISA|7|4|对他说：‘你要谨慎，要镇定，不要害怕，不要因 利汛 和 亚兰 ，以及 利玛利 的儿子这两个冒烟火把的头所发的烈怒而心里胆怯。
ISA|7|5|因为 亚兰 、 以法莲 ，和 利玛利 的儿子设恶谋要害你，说：
ISA|7|6|我们要上去攻击 犹大 ，扰乱它，攻破它来归我们，在其中立 他比勒 的儿子为王。
ISA|7|7|主耶和华如此说： 这事必站立不住， 也不得成就。
ISA|7|8|因为 亚兰 的首都是 大马士革 ， 大马士革 的领袖是 利汛 ； 六十五年之内， 以法莲 必然国破族亡，
ISA|7|9|以法莲 的首都是 撒玛利亚 ； 撒玛利亚 的领袖是 利玛利 的儿子。 你们若是不信， 必站立不稳。’”
ISA|7|10|耶和华又吩咐 亚哈斯 ：
ISA|7|11|“你向耶和华－你的上帝求一个预兆：在阴间的深渊，或往上的高处。”
ISA|7|12|但 亚哈斯 说：“我不求；我不试探耶和华。”
ISA|7|13|以赛亚 说：“听啊， 大卫 家！你们使人厌烦岂算小事，还要使我的上帝厌烦吗？
ISA|7|14|因此，主自己要给你们一个预兆，看哪，必有童女怀孕生子，给他起名叫 以马内利 。
ISA|7|15|到他晓得弃恶择善的时候，他必吃乳酪与蜂蜜。
ISA|7|16|因为在这孩子还不晓得弃恶择善之先，你所憎恶的那两个王的土地必被撇弃。
ISA|7|17|耶和华必使 亚述 王临到你和你的百姓，并你的父家，自从 以法莲 脱离 犹大 的时候，未曾有过这样的日子。
ISA|7|18|“那时，耶和华要呼叫，召来 埃及 江河源头的苍蝇和 亚述 地的蜂；
ISA|7|19|它们都必飞来，停在陡峭的谷中、岩石缝里、一切荆棘丛中和片片草场上。
ISA|7|20|“那时，主必用 大河 外雇来的剃刀，就是 亚述 王，剃去你的头发和脚毛，并要剃净你的胡须。
ISA|7|21|“那时，每一个人要养活一头母牛犊和两只母羊；
ISA|7|22|因为奶量充足，他就有乳酪可吃，国内剩余的人也都能吃乳酪与蜂蜜。
ISA|7|23|“那时，凡种一千棵葡萄树、价值一千银子的地方，必长出荆棘和蒺藜。
ISA|7|24|人到那里去，必带弓箭，因为遍地长满了荆棘和蒺藜。
ISA|7|25|所有锄头刨过的山地，你因惧怕荆棘和蒺藜，不敢到那里去；只能作放牛之处，羊群践踏之地。”
ISA|8|1|耶和华对我说：“你取一块大板子，拿人的笔 ，写上‘玛黑珥．沙拉勒．哈施．罢斯’ 。
ISA|8|2|我 要用可靠的证人， 乌利亚 祭司和 耶比利家 的儿子 撒迦利亚 为我作证。”
ISA|8|3|我亲近女先知 ；她就怀孕生子，耶和华对我说：“给他起名叫 玛黑珥．沙拉勒．哈施．罢斯 ；
ISA|8|4|因为在这孩子还不晓得叫爸爸妈妈以前， 大马士革 的财宝和 撒玛利亚 的掳物必被 亚述 王掠夺一空。”
ISA|8|5|耶和华又吩咐我：
ISA|8|6|“这百姓既厌弃 西罗亚 缓流的水，喜欢 利汛 以及 利玛利 的儿子，
ISA|8|7|因此，看哪，主必使 亚述 王和他的威势如 大河 翻腾汹涌的水上涨，盖过他们，必上涨超过一切水道，涨过两岸，
ISA|8|8|必冲入 犹大 ，涨溢泛滥，直到颈项。他展开翅膀，遮蔽你的全地。 以马内利 啊！”
ISA|8|9|万民哪，任凭你们行恶 ，终必毁灭； 远方的众人哪，当侧耳而听！ 任凭你们束腰，终必毁灭； 你们束起腰来，终必毁灭。
ISA|8|10|任凭你们筹算什么，终必无效； 不管你们讲定什么，总不成立； 因为上帝与我们同在。
ISA|8|11|耶和华以大能的手训诫我不可行 这百姓所行的道，对我这样说：
ISA|8|12|“这百姓说同谋背叛的，你们不要说同谋背叛。他们所怕的，你们不要怕，也不要畏惧；
ISA|8|13|但要尊万军之耶和华为圣，他才是你们所当怕的，所当畏惧的。
ISA|8|14|他必作为圣所，却向 以色列 的两家成为绊脚的石头，使人跌倒的磐石；作 耶路撒冷 居民的罗网和圈套。
ISA|8|15|许多人在其上绊倒，他们跌倒，甚至跌伤，并且落入陷阱，被抓住了。”
ISA|8|16|你要卷起律法书，在我门徒中间封住教诲。
ISA|8|17|我要等候那转脸不顾 雅各 家的耶和华，也要仰望他。
ISA|8|18|看哪，我与耶和华所赐给我的儿女成了 以色列 的预兆和奇迹，这是从住在 锡安山 万军之耶和华来的。
ISA|8|19|有人对你们说：“当求问招魂的与行巫术的，他们唧唧喳喳，念念有词。”然而，百姓不当求问自己的上帝吗？岂可为活人求问死人呢？
ISA|8|20|当以教诲和律法书为准；人所说的若不与此相符，必没有黎明。
ISA|8|21|他必经过这地，遇艰难，受饥饿；饥饿的时候，心中焦躁，咒骂自己的君王和上帝。他仰观上天，
ISA|8|22|俯察下地，看哪，尽是艰难、黑暗和骇人的昏暗。他必被赶入幽暗中去。
ISA|9|1|但那受过痛苦的必不再见幽暗。 从前上帝使 西布伦 地和 拿弗他利 地被藐视，末后却使这沿海的路， 约旦河 东，外邦人居住的 加利利 地得荣耀。
ISA|9|2|在黑暗中行走的百姓看见了大光； 住在死荫之地的人有光照耀他们。
ISA|9|3|你使这国民众多 ， 使他们喜乐大增； 他们在你面前欢喜， 好像收割时的欢喜， 又像人分战利品那样的快乐。
ISA|9|4|因为他们所负的重轭 和肩头上的杖， 并欺压者的棍， 你都已经折断， 如同在 米甸 的日子一般。
ISA|9|5|战士在战乱中所穿的靴子， 以及那滚在血中的衣服， 都必当作柴火燃烧。
ISA|9|6|因有一婴孩为我们而生； 有一子赐给我们。 政权必担在他的肩头上； 他名称为“奇妙策士、全能的上帝、永在的父、和平的君”。
ISA|9|7|他的政权与平安必加增无穷。 他必在 大卫 的宝座上治理他的国， 以公平公义使国坚定稳固， 从今直到永远。 万军之耶和华的热心必成就这事。
ISA|9|8|主向 雅各 家发出言语， 主的话临到 以色列 家。
ISA|9|9|众百姓，就是 以法莲 和 撒玛利亚 的居民， 都将知道； 他们凭骄傲自大的心说：
ISA|9|10|“砖块掉落了，我们要凿石头重建； 桑树砍了，我们要改种香柏树。”
ISA|9|11|因此，耶和华兴起 利汛 的敌人 前来攻击 以色列 ， 要激起它的仇敌，
ISA|9|12|东有 亚兰 人，西有 非利士 人； 他们张口吞吃 以色列 。 虽然如此，耶和华的怒气并未转消； 他的手依然伸出。
ISA|9|13|这百姓还没有归向击打他们的主， 也没有寻求万军之耶和华。
ISA|9|14|耶和华在一日之间 从 以色列 中剪除了头与尾－ 棕树枝与芦苇－
ISA|9|15|长老和显要就是头， 以谎言教人的先知就是尾。
ISA|9|16|因为引导这百姓的使他们走入迷途， 被引导的都必被吞灭。
ISA|9|17|所以，主不喜爱 他们的青年， 也不怜悯他们的孤儿和寡妇； 因为他们都是亵渎的，行恶的， 并且各人的口都说愚妄的话。 虽然如此，耶和华的怒气并未转消； 他的手依然伸出。
ISA|9|18|邪恶如火焚烧， 吞灭荆棘和蒺藜， 在稠密的树林中点燃， 成为烟柱，旋转上腾。
ISA|9|19|因万军之耶和华的烈怒，地都烧遍了； 百姓成为柴火， 无人怜惜弟兄。
ISA|9|20|有人右边抢夺，犹受饥饿； 左边吞吃，仍不饱足， 各人吃自己膀臂上的肉。
ISA|9|21|玛拿西 吞吃 以法莲 ， 以法莲 吞吃 玛拿西 ， 他们又一同攻击 犹大 。 虽然如此，耶和华的怒气并未转消； 他的手依然伸出。
ISA|10|1|祸哉！那些设立不义之律例的， 和记录奸诈之判词的，
ISA|10|2|为要扭曲贫寒人的案件， 夺去我民中困苦人的理， 以寡妇当作掳物， 以孤儿当作掠物。
ISA|10|3|到降罚的日子，灾祸从远方临到， 那时，你们要怎么办呢？ 你们要向谁逃奔求救呢？ 你们的财宝要存放何处呢？
ISA|10|4|他们只得屈身在被掳的人之下， 仆倒在被杀的人中间 。 虽然如此，耶和华的怒气并未转消； 他的手依然伸出。
ISA|10|5|祸哉！ 亚述 ，我怒气的棍！ 他们手中的杖是我的恼恨。
ISA|10|6|我要差遣他攻击亵渎的国， 吩咐他对付我所恼怒的民， 抢走掳物，夺取掠物， 将他们践踏，如同街上的泥土一般。
ISA|10|7|然而，这并非他的意念， 他的心不是这样打算； 他的心要摧毁， 要剪除不少的国家。
ISA|10|8|他说：“我的官长岂不都是君王吗？
ISA|10|9|迦勒挪 岂不像 迦基米施 吗？ 哈马 岂不像 亚珥拔 吗？ 撒玛利亚 岂不像 大马士革 吗？
ISA|10|10|既然我的手已伸到了这些有偶像的国， 他们所雕刻的偶像 过于 耶路撒冷 和 撒玛利亚 的偶像，
ISA|10|11|我岂不照样待 耶路撒冷 和其中的偶像， 如同我待 撒玛利亚 和其中的偶像吗？”
ISA|10|12|主在 锡安山 和 耶路撒冷 成就他一切工作的时候，说：“我必惩罚 亚述 王自大的心和他高傲尊贵的眼目。”
ISA|10|13|因为他说： “我所成就的事是靠我手的能力 和我的智慧， 因为我本有聪明。 我挪移列国的地界， 抢夺他们所积蓄的财宝， 并且像勇士，使坐宝座的降为卑。
ISA|10|14|我的手夺取列国的财宝， 好像人夺取鸟窝； 我得了全地， 好像人拾起被弃的鸟蛋； 没有振动翅膀的， 没有张嘴的，也没有鸣叫的。”
ISA|10|15|斧岂可向用斧砍伐的自夸呢？ 锯岂可向拉锯的自大呢？ 这好比棍挥动那举棍的， 好比杖举起那不是木头的人。
ISA|10|16|因此，主－万军之耶和华 必使 亚述 王的壮士变为瘦弱， 在他的荣华之下必有火点燃， 如同火在燃烧一般。
ISA|10|17|以色列 的光必变成火， 它的圣者必成为火焰； 一日之间，将 亚述 王的荆棘和蒺藜焚烧净尽，
ISA|10|18|又毁灭树林和田园的荣华， 连魂带体，好像病重的人消逝 一样。
ISA|10|19|他林中只剩下稀少的树木， 连孩童也能写其数目。
ISA|10|20|到那日， 以色列 所剩下的和 雅各 家所逃脱的，必不再倚靠那击打他们的，却要诚心仰赖耶和华－ 以色列 的圣者。
ISA|10|21|所剩下的，就是 雅各 家的余民，必归回全能的上帝。
ISA|10|22|以色列 啊，你的百姓虽多如海沙，惟有剩下的归回。灭绝之事已成定局，公义必如水涨溢。
ISA|10|23|因为万军之主耶和华在全地必成就所定的灭绝之事。
ISA|10|24|所以，万军之主耶和华如此说：“住 锡安 我的百姓啊， 亚述 王虽然用棍击打你，又如 埃及 举杖攻击你，你不要怕他。
ISA|10|25|因为还有一点点时候，我向你们发的愤怒就要结束，我的怒气要使他们灭亡。
ISA|10|26|万军之耶和华要举起鞭子来攻击他，好像在 俄立 磐石那里击打 米甸 人一样。他的杖向海伸出，他必把杖举起，如在 埃及 一般。
ISA|10|27|到那日， 亚述 王的重担必离开你的肩头，他的轭必离开你的颈项；那轭必因肥壮而撑断 。”
ISA|10|28|亚述 王来到 亚叶 ， 经过 米矶仑 ， 在 密抹 安放辎重。
ISA|10|29|他们过了隘口， 要在 迦巴 住宿。 拉玛 战兢， 扫罗 的 基比亚 逃命。
ISA|10|30|迦琳 哪，要高声呼喊！ 注意听， 莱煞 啊！ 困苦的 亚拿突 啊 ！
ISA|10|31|玛得米那 躲避， 基柄 的居民逃遁。
ISA|10|32|当那日， 亚述 王要在 挪伯 停留， 挥手攻击 锡安 的山， 就是 耶路撒冷 的山。
ISA|10|33|看哪，主－万军之耶和华 以猛撞削断树枝； 巨木必被砍下， 高大的树必降为低。
ISA|10|34|稠密的树林，他要用铁器砍下， 黎巴嫩 必被大能者伐倒 。
ISA|11|1|从 耶西 的残干必长出嫩枝， 他的根所抽的枝子必结果实。
ISA|11|2|耶和华的灵必住在他身上， 就是智慧和聪明的灵， 谋略和能力的灵， 知识和敬畏耶和华的灵。
ISA|11|3|他必以敬畏耶和华为乐； 行审判不凭眼见， 断是非也不凭耳闻；
ISA|11|4|却要以公义审判贫寒人， 以正直判断地上的困苦人， 以口中的棍击打全地， 以嘴里的气杀戮恶人。
ISA|11|5|公义必当他的腰带， 信实必作他胁下的带子。
ISA|11|6|野狼必与小绵羊同住， 豹子与小山羊同卧； 少壮狮子、牛犊和肥畜同群 ； 孩童要牵引它们。
ISA|11|7|牛必与熊同食， 牛犊与小熊同卧； 狮子与牛一样吃草。
ISA|11|8|吃奶的婴孩在虺蛇的洞口玩耍， 断奶的幼儿必按手在毒蛇的穴上。
ISA|11|9|在我圣山各处， 它们都不伤人，不害物； 因为认识耶和华的知识要遍满全地， 好像水充满海洋一般。
ISA|11|10|到那日， 耶西 的根立作万民的大旗；列国的人必寻求他，他安歇之所大有荣耀。
ISA|11|11|当那日，主必再度伸手救回自己百姓中所剩余的，就是在 亚述 、 埃及 、 巴特罗 、 古实 、 以拦 、 示拿 、 哈马 ，并众海岛所剩下的。
ISA|11|12|他要向列国竖立大旗， 召集 以色列 被赶散的人， 又从地极四方聚集分散的 犹大 人。
ISA|11|13|以法莲 的嫉妒必消散， 苦待 犹大 的也被剪除； 以法莲 必不嫉妒 犹大 ， 犹大 也不苦待 以法莲 。
ISA|11|14|他们要飞向西方， 扑在 非利士 人的肩头上， 他们要一同掳掠东方人， 他们的手伸到 以东 和 摩押 ； 亚扪 人也必顺服他们。
ISA|11|15|耶和华必使 埃及 的海湾全然毁坏 ， 他举手在 大河 之上刮起了暴热的风， 击打它，使它分成七条溪流， 人穿鞋便可渡过。
ISA|11|16|必有一条大道， 为百姓中从 亚述 逃脱生还的余民而开， 如当日为 以色列 从 埃及 上来一样。
ISA|12|1|在那日，你要说： “耶和华啊，我要称谢你！ 因为你虽然向我发怒， 你的怒气却已转消； 你又安慰了我。
ISA|12|2|“看哪！上帝是我的拯救； 我要倚靠他，并不惧怕。 因为主耶和华是我的力量， 是我的诗歌， 他也成了我的拯救。”
ISA|12|3|你们必从救恩的泉源欢然取水。
ISA|12|4|在那日，你们要说： “当称谢耶和华，求告他的名； 在万民中传扬他的作为， 宣告他的名已被尊崇。
ISA|12|5|“你们要向耶和华唱歌， 因他所做的十分宏伟； 但愿这事遍传全地。
ISA|12|6|锡安 的居民哪，当扬声欢呼， 因为在你们当中的 以色列 圣者最为伟大。”
ISA|13|1|亚摩斯 的儿子 以赛亚 所见，有关 巴比伦 的默示。
ISA|13|2|你们要在荒凉的山上竖立大旗， 向他们扬声， 挥手招呼他们进入贵族之门。
ISA|13|3|我吩咐我所分别为圣的人， 召唤我的勇士， 就是我那狂喜高傲的人， 为要执行我的怒气。
ISA|13|4|听啊，山间有喧闹的声音， 好像有许多百姓聚集， 听啊，多国之民聚集闹哄的声音； 这是万军之耶和华召集作战的军队。
ISA|13|5|他们从远方来， 从天边来， 耶和华和他恼恨的兵器 要毁灭全地。
ISA|13|6|你们要哀号， 因为耶和华的日子临近了！ 这日来到，好像毁灭从全能者来到。
ISA|13|7|因此，人的手都变软弱， 人的心都必惶惶。
ISA|13|8|他们必惊恐， 悲痛和愁苦将他们抓住。 他们阵痛，好像临产的妇人一样， 彼此惊奇对看，脸如火焰。
ISA|13|9|看哪！耶和华的日子临到， 必有残忍、愤恨、烈怒， 使这地荒芜， 除灭其中的罪人。
ISA|13|10|天上的星宿都不发光， 太阳一升起就变黑暗， 月亮也不放光。
ISA|13|11|我必因邪恶惩罚世界， 因罪孽惩罚恶人， 我要止息骄傲人的狂妄， 制伏残暴者的傲慢。
ISA|13|12|我要使人比纯金更少， 比 俄斐 的赤金还少。
ISA|13|13|我，万军之耶和华狂怒，就是发烈怒的日子， 要令天震动， 地必摇撼，离其本位。
ISA|13|14|人如被追赶的羚羊， 像无人聚集的羊群， 各自归回本族， 逃到本地。
ISA|13|15|凡被追上的必被刺死， 凡被捉拿的必倒在刀下。
ISA|13|16|他们的婴孩必在他们眼前被摔死， 他们的房屋被抢劫， 他们的妻子被污辱。
ISA|13|17|看哪，我必激起 玛代 人攻击他们， 玛代 人并不看重银子， 也不喜爱金子。
ISA|13|18|他们必用弓击溃青年， 不怜悯妇人所生的； 眼也不顾惜孩子。
ISA|13|19|巴比伦 为列国的荣耀， 为 迦勒底 人所夸耀的华美， 必像上帝所倾覆的 所多玛 、 蛾摩拉 一样；
ISA|13|20|国中必永无人烟， 世世代代无人居住； 阿拉伯 人不在那里支搭帐棚， 牧羊的人也不使羊群躺卧在那里。
ISA|13|21|旷野的走兽躺卧在那里， 咆哮的动物挤满栖身之所； 鸵鸟住在那里， 山羊鬼魔也在那里跳舞。
ISA|13|22|土狼必在它的宫殿 呼号， 野狗在华美的殿里吼叫。 巴比伦 的时辰临近了， 它的日子必不长久。
ISA|14|1|耶和华要怜悯 雅各 ，再度拣选 以色列 ，将他们安顿在本地。寄居的必与他们联合，加入 雅各 家。
ISA|14|2|外邦人要将他们带回本地。 以色列 家必在耶和华的地上得外邦人为仆婢，也要掳掠先前掳掠他们的，辖制先前欺压他们的。
ISA|14|3|当耶和华使你得享安息，脱离愁苦、烦恼，和被迫做苦工的日子，
ISA|14|4|你必唱这诗歌嘲讽 巴比伦 王说： “欺压人的竟然灭亡！ 他的凶暴 竟然止息！
ISA|14|5|耶和华折断恶人的杖， 打断统治者的权杖；
ISA|14|6|他们在愤怒中连连攻击万民， 在怒气中辖制列国， 逼迫他们，毫不留情。
ISA|14|7|现在全地得安息，享平静， 人都出声欢呼。
ISA|14|8|松树和 黎巴嫩 的香柏树 都因你欢乐： 自从你仆倒， 再也无人上来砍伐我们。
ISA|14|9|下面的阴间因你震动， 迎接你的到来； 在世曾为领袖的阴魂为你惊动， 那曾为列国君王的，都从宝座起立。
ISA|14|10|他们都要发言，对你说： ‘你也变为软弱，像我们一样吗？ 你也成了我们的样子吗？’
ISA|14|11|你的威严和琴瑟的声音都下到阴间。 你下面铺的是虫，上面盖的是蛆。
ISA|14|12|“明亮之星，早晨之子啊， 你竟然从天坠落！ 你这攻败列国的，竟然被砍倒在地上！
ISA|14|13|你心里曾说： ‘我要升到天上， 我要高举我的宝座在上帝的众星之上， 我要坐在会众聚集的山上，在极北的地方。
ISA|14|14|我要升到高云之上， 我要与至高者同等。’
ISA|14|15|然而，你必坠落阴间， 到地府极深之处。
ISA|14|16|凡看见你的都要定睛望你， 留意看你，说： ‘就是这个人吗？ 他使大地颤抖， 使列国震动，
ISA|14|17|使世界如同荒野， 使城镇倾覆； 是他，不释放被掳的人归家。’
ISA|14|18|列国的君王各自在自己的坟墓中， 在尊荣里长眠。
ISA|14|19|惟独你被抛弃在你的坟墓之外， 有如被厌恶的枝子 ， 被许多用刀刺透杀死的人覆盖着， 一同坠落地府的石头那里， 像被践踏的尸首。
ISA|14|20|你不得与君王同葬， 因为你毁坏你的国，杀戮你的民。 “恶人的后裔永不留名。
ISA|14|21|为了祖先的罪孽， 要预备他子孙的屠宰场， 免得他们兴起，夺得全地， 使城市遍满地面。”
ISA|14|22|万军之耶和华说： “我必起来攻击他们， 将 巴比伦 的名号和剩余的人， 连子带孙一并剪除； 这是耶和华说的。
ISA|14|23|“我必使 巴比伦 为豪猪占据， 成为泥沼之地； 我要用灭命的扫帚扫净它； 这是万军之耶和华说的。”
ISA|14|24|万军之耶和华起誓说： “我怎样思想，必照样成就； 我怎样定意，必照样坚立，
ISA|14|25|要在我的地上击破 亚述 ， 在我的山上将它践踏。 它的轭必离开受压制的人， 它的重担必离开他们的肩头。”
ISA|14|26|这是向全地所定的旨意， 向万国所伸出的手。
ISA|14|27|万军之耶和华既然定意，谁能阻挠呢？ 他的手已经伸出，谁能使它缩回呢？
ISA|14|28|亚哈斯 王崩的那年，有默示如下：
ISA|14|29|“全 非利士 啊， 不要因击打你的杖折断就喜乐。 因为蛇必生出毒蛇， 它所生的是会飞的火蛇。
ISA|14|30|贫寒人的长子必有得吃； 贫穷人必安然躺卧。 我必以饥荒灭绝你的根， 它 必杀尽你所剩余的人。
ISA|14|31|门哪，哀号吧！ 城啊，呼喊吧！ 全 非利士 都熔化了！ 因为有烟从北方而来， 在它的行伍中没有掉队的。”
ISA|14|32|当如何回答外邦的使者呢？ “耶和华建立了 锡安 ， 在其中他困苦的百姓必有倚靠。”
ISA|15|1|论 摩押 的默示。 一夜之间， 摩押 的 亚珥 变为荒废， 归于无有； 一夜之间， 摩押 的 基珥 变为荒废， 归于无有。
ISA|15|2|摩押 上到神庙和 底本 的丘坛去哭泣； 它因 尼波 和 米底巴 哀号， 各人头上光秃，胡须剃净。
ISA|15|3|他们在街市上腰束麻布， 都在房顶和广场上哀号， 泪流不停。
ISA|15|4|希实本 和 以利亚利 呼喊， 他们的声音达到 雅杂 ， 所以 摩押 的士兵高声喊叫， 他们的心战兢。
ISA|15|5|我的心 为 摩押 哀号； 它的难民逃到 琐珥 ， 逃到 伊基拉．施利施亚 。 他们上 鲁希坡 ，随走随哭， 在 何罗念 的路上，因毁灭发出哀声。
ISA|15|6|宁林 的水干涸， 青草枯干，嫩草死光， 青绿之物，一无所有。
ISA|15|7|因此， 摩押 人所得的财物和积蓄 都要运过 柳树河 。
ISA|15|8|哀声遍传 摩押 四境， 哀号的声音达到 以基莲 ， 哀号的声音远及 比珥．以琳 。
ISA|15|9|底们 的水充满了血， 然而我还要加添 底们 的灾难， 让狮子追上 摩押 的难民 和那地 剩余的人。
ISA|16|1|你们当将 羔羊奉送给那地的掌权者， 从 西拉 往旷野，送到 锡安 的山。
ISA|16|2|摩押 的居民 来到 亚嫩 渡口， 如逃遁的飞鸟，被赶离鸟巢 。
ISA|16|3|求你赐谋略，行公平， 使你的影子在正午如黑夜， 掩护逃亡的人，不泄露逃难者的行踪。
ISA|16|4|愿我 摩押 逃亡的人 寄居在你那里， 你作他们的避难所，躲避灭命者的面。 勒索的人消失， 毁灭的事止息， 欺压者从国中除灭，
ISA|16|5|在 大卫 帐幕中必有宝座因慈爱坚立， 必有一位君王凭信实坐在其上， 施行审判，寻求公平，迅速行公义。
ISA|16|6|我们听闻 摩押 的骄傲， 极其骄傲； 它狂妄、骄傲、自大， 它夸大的言词都是空的。
ISA|16|7|因此， 摩押 人必为 摩押 哀号， 人人都要哀号。 你们要为 吉珥．哈列设 的葡萄饼哀叹， 极其忧伤。
ISA|16|8|因为 希实本 的田地 和 西比玛 的葡萄树都衰残了， 列国的君主折断它的枝干， 这枝子曾长到 雅谢 ，延伸到旷野， 嫩枝向外伸出，直伸过海；
ISA|16|9|所以，我要为 西比玛 的葡萄树哀哭， 像 雅谢 人一样哀哭。 希实本 、 以利亚利 啊， 我要以眼泪浇灌你， 你因夏天果子和收割的庄稼， 欢呼声已经止息了。
ISA|16|10|田园中不再有欢喜快乐， 葡萄园里必无人歌唱，无人欢呼， 在压酒池中踹酒的不再踹酒了， 我使欢呼的声音止息了 。
ISA|16|11|因此，我的心肠为 摩押 哀鸣如琴， 我的内心为 吉珥．哈列设 哀哭。
ISA|16|12|当 摩押 人出现在丘坛，筋疲力尽时，虽然到自己的圣所祈祷，却仍无济于事。
ISA|16|13|这是耶和华曾论到 摩押 的话。
ISA|16|14|但现在，耶和华说：“三年之内，按照雇工年数的算法， 摩押 的荣华必变为羞辱，人口虽曾众多，剩余的又少又弱。”
ISA|17|1|论 大马士革 的默示。 看哪， 大马士革 不再为城市， 变为废墟。
ISA|17|2|亚罗珥 的城镇被撇弃 ， 将成为牧羊之处， 羊群在那里躺卧， 无人使它们惊吓。
ISA|17|3|以法莲 不再有堡垒， 大马士革 失去其王国， 亚兰 的百姓所剩无几， 如 以色列 人的荣美消失一般； 这是万军之耶和华说的。
ISA|17|4|到那日， 雅各 的荣美必失色， 它肥胖的身躯渐渐消瘦；
ISA|17|5|像人收割成熟的禾稼， 用手臂割取麦穗， 又像人在 利乏音谷 拾取穗子；
ISA|17|6|其间所剩不多，好像人打橄榄树， 在最高的树梢上只剩两、三颗橄榄， 在多结果子的旁枝上只剩四、五颗； 这是耶和华－ 以色列 的上帝说的。
ISA|17|7|当那日，人必仰望造他们的主，眼目看着 以色列 的圣者。
ISA|17|8|他们必不仰望自己手所筑的祭坛，也不理会自己指头所造的 亚舍拉 和香坛。
ISA|17|9|当那日，他们坚固的城必因 以色列 人的缘故，如同树林中和山顶上所撇弃的地方 。这样，地就荒芜了。
ISA|17|10|因你忘记拯救你的上帝， 忘记那保护你的磐石； 所以，你虽栽上佳美的树苗， 插上别样的枝子，
ISA|17|11|栽种的日子，你使它生长， 栽种的早晨，你使它开花， 但在愁苦、极其伤痛的日子， 所收割的都归无有。
ISA|17|12|唉！万民闹哄，好像海浪澎湃， 列邦喧闹，如同洪水滔滔，
ISA|17|13|列邦喧闹，如同大水滔滔； 但上帝一斥责，他们就远远躲避， 他们被追赶，如同山上风前的糠秕， 又如暴风前的碎秸；
ISA|17|14|看哪，晚上有惊吓，未到早晨它就消失无踪。 这是掳掠我们之人的厄运，是抢夺我们之人的报应。
ISA|18|1|祸哉！ 古实河 的那一边、翅膀刷刷作响之地，
ISA|18|2|差遣使者在水面上， 坐蒲草船过海。 你们这些疾行的使者， 要到高大光滑的民那里去； 那民远近都畏惧， 是强大好征服的国， 土地有河流穿过。
ISA|18|3|世上所有的居民，住在地上的人哪， 山上大旗竖起时，你们要看， 号角吹响时，你们要听。
ISA|18|4|耶和华对我如此说： “我要安静，从我的居所观看， 如同日光下闪烁的热气， 又如收割时 露水蒸发的云雾。”
ISA|18|5|收割之前，花蕾先谢， 花成了将熟的葡萄； 他必用刀削去嫩枝， 砍掉蔓延的枝条，
ISA|18|6|一起丢给山间的鸷鸟和地上的野兽； 鸷鸟要在其上避暑， 地上一切的野兽都在那里过冬。
ISA|18|7|到那时，这高大光滑的民， 远近都畏惧的民、 强大好征服之国、 土地有河流穿过； 他们必被当作 礼物献给万军之耶和华， 献到 锡安山 － 万军之耶和华立他名的地方。
ISA|19|1|论 埃及 的默示。 看哪，耶和华乘驾快云， 临到 埃及 ； 埃及 的偶像在他面前战兢， 埃及 人的心在里面消溶。
ISA|19|2|我要激起 埃及 人攻击 埃及 人， 弟兄攻击弟兄， 邻舍攻击邻舍， 这城攻击那城， 这国攻击那国。
ISA|19|3|埃及 人的心神在里面耗尽， 我要破坏他们的计谋。 他们必求问偶像和念咒的， 求问招魂的与行巫术的人。
ISA|19|4|我要将 埃及 人交在严厉的主人手中， 残暴的君王必管辖他们； 这是主－万军之耶和华说的。
ISA|19|5|海水枯竭， 河流干涸，
ISA|19|6|江河发臭， 埃及 的河水必然减少而枯干。 芦苇和芦荻枯萎，
ISA|19|7|尼罗河 旁的植物 ，在 尼罗河 的沿岸， 并 尼罗河 旁所种的一切 全都枯焦，被风吹去，归于无有。
ISA|19|8|打鱼的哀哭， 所有在 尼罗河 钓鱼的都必悲伤， 在水上撒网的也都衰残。
ISA|19|9|以细致的麻编织的必羞愧， 织布的必变苍白 ；
ISA|19|10|织布的心情沮丧 ， 所有的佣工心都愁烦。
ISA|19|11|琐安 的官长极其愚昧， 法老智慧的谋士筹划愚谋； 你们怎敢对法老说： “我是智慧人的子孙， 是古代国王的后裔？”
ISA|19|12|你的智慧人在哪里？ 万军之耶和华向 埃及 所定的旨意， 他们既然知道，就让他们告诉你吧！
ISA|19|13|琐安 的官长愚昧， 挪弗 的官长受蒙蔽； 作 埃及 支派栋梁的， 带领 埃及 走错了路。
ISA|19|14|耶和华使歪曲的灵渗入 埃及 中间， 让他们使 埃及 一切所做的都出差错， 好像醉酒之人呕吐时东倒西歪一样。
ISA|19|15|在 埃及 ，无论是头是尾， 棕树枝与芦苇，所做的事都不得成就。
ISA|19|16|到那日， 埃及 必像妇人一样，因万军之耶和华挥手攻击而战兢惧怕。
ISA|19|17|犹大 地必使 埃及 惊恐，不论向谁提起，他都惧怕。这是因万军之耶和华向 埃及 所定的旨意。
ISA|19|18|当那日， 埃及 地必有五个城市的人说 迦南 的语言，又指着万军之耶和华起誓。有一城必称为“太阳城” 。
ISA|19|19|在那日，在 埃及 地将有献给耶和华的一座坛，边界上必有为耶和华立的一根柱子。
ISA|19|20|这都要在 埃及 地为万军之耶和华作记号和证据。 埃及 人因受欺压哀求耶和华，他就差遣一位救主作护卫者，拯救他们，
ISA|19|21|耶和华就被 埃及 所认识。在那日， 埃及 人要认识耶和华，献牲祭和素祭敬拜他，并向耶和华许愿还愿。
ISA|19|22|耶和华必击打 埃及 ，又击打又医治， 埃及 人就归向耶和华。他必应允他们的祷告，医治他们。
ISA|19|23|在那日，必有从 埃及 通往 亚述 的大道。 亚述 人要进入 埃及 ， 埃及 人也要进入 亚述 ； 埃及 人要与 亚述 人一同敬拜。
ISA|19|24|在那日， 以色列 将与 埃及 、 亚述 三国一起，使地上的人得福。
ISA|19|25|万军之耶和华必赐福给他们，说：“ 埃及 －我的百姓， 亚述 －我手的工作， 以色列 －我的产业，都有福了！”
ISA|20|1|亚述 元帅 受 亚述 王 撒珥根 派遣往 亚实突 的那年，他攻打 亚实突 ，将城攻取。
ISA|20|2|那时，耶和华吩咐 亚摩斯 的儿子 以赛亚 说：“你去解掉你腰间的麻布，脱下你脚上的鞋。” 以赛亚 就这样做，赤身赤脚行走。
ISA|20|3|耶和华说：“我仆人 以赛亚 怎样赤身赤脚行走三年，作为关于 埃及 和 古实 的预兆奇迹，
ISA|20|4|照样， 亚述 王必掳去 埃及 人，掠去 古实 人，无论老少，都赤身赤脚，露出下体，使 埃及 蒙羞。
ISA|20|5|以色列 人必惊惶羞愧，因为他们仰望 古实 ，以 埃及 为荣。
ISA|20|6|“那时，沿海一带的居民必说：‘看哪，我们素来所仰望的，就是为躲避 亚述 王所逃往 求救的，不过如此！我们怎能逃脱呢？’”
ISA|21|1|论海边旷野的默示。 它像 尼革夫 的旋风扫过， 从旷野，从可怕之地而来。
ISA|21|2|有凄惨的异象向我揭示： “诡诈的在行诡诈，毁灭的在行毁灭。 以拦 哪，前进吧！ 玛代 啊，围攻吧！ 我使它一切的叹息停止了。”
ISA|21|3|为此，我腰部满是疼痛， 痛苦将我抓住， 好像临产的妇人一样的痛。 我疼痛甚至不能听， 我惊惶甚至不能看 。
ISA|21|4|我心慌乱，惊恐威吓我。 我所渴望的黄昏，反成为我的恐惧。
ISA|21|5|有人摆设筵席， 铺上地毯，又吃又喝。 “官长啊，起来， 抹亮盾牌。”
ISA|21|6|主对我如此说： “你去设立守望者， 让他报告他所看见的。
ISA|21|7|他会看见一对一对骑着马的军队， 又看见驴队，骆驼队， 他要留心听，仔细地听。”
ISA|21|8|他如狮子般吼叫 ： “主啊，我白天常站在暸望楼， 彻夜立在我的暸望台。”
ISA|21|9|看哪，有一对一对骑着马的军队前来。 他就回应说：“ 巴比伦 倾倒了！倾倒了！ 他把 巴比伦 神明的一切雕刻偶像都打碎在地上了。”
ISA|21|10|我被打的禾稼，我禾场上的谷物啊， 我从万军之耶和华－ 以色列 的上帝那里所听见的，都告诉你们了。
ISA|21|11|论 度玛 的默示。 有人声从 西珥 呼喊： “守望的啊，夜里如何？ 守望的啊，夜里如何？”
ISA|21|12|守望者说： “早晨来到，黑夜将临。 你们若要问，问吧， 也可以回头再来。”
ISA|21|13|论 阿拉伯 的默示。 底但 的旅行商队啊， 你们在 阿拉伯 的树林中住宿。
ISA|21|14|提玛 地的居民哪， 提水来迎接口渴的人， 带饼来迎接难民。
ISA|21|15|他们躲避刀剑和出了鞘的刀， 躲避上了弦的弓与战争的重灾。
ISA|21|16|主对我这样说：“一年之内，按照雇工年数的算法， 基达 一切的繁华必归无有。
ISA|21|17|基达 人中强壮弓箭手剩下的数目甚为稀少，这是耶和华－ 以色列 的上帝说的。”
ISA|22|1|论异象谷的默示。 什么事使你们上去， 全都上到屋顶呢？
ISA|22|2|你这四处呐喊、大声喧哗的城、 欢乐的邑啊， 你被杀的并非被刀所杀， 也不是因打仗阵亡。
ISA|22|3|你所有的官长一同奔逃， 不用弓箭就被捆绑 ； 你们即使逃往远方， 也要被找到，一同被捆绑。
ISA|22|4|因此我说： “不要看我， 让我痛哭吧！ 不要因我百姓 的毁灭竭力安慰我。”
ISA|22|5|因为这是万军之主耶和华使异象谷 混乱、践踏、烦扰的日子； 城墙被攻破， 哀声达到山上。
ISA|22|6|以拦 提着箭袋， 有战车、士兵、骑兵； 吉珥 亮出盾牌，
ISA|22|7|你佳美的山谷遍布战车， 骑兵排列在城门前。
ISA|22|8|他除掉 犹大 的防御。 那时，你指望森林库里的兵器。
ISA|22|9|你们看见 大卫城 缺口很多，就汇集 下池 的水；
ISA|22|10|你们数点 耶路撒冷 的房屋，拆毁房屋，用以修补城墙，
ISA|22|11|又在两道城墙中间挖水池，用以盛旧池的水，却不仰望成就这事的主，也不顾念从古时定这事的主。
ISA|22|12|当那日，万军之主耶和华使人哭泣哀号， 头上光秃，身披麻布。
ISA|22|13|看哪，人却欢喜快乐， 宰牛杀羊，吃肉喝酒： “让我们吃吃喝喝吧！因为明天要死了。”
ISA|22|14|万军之耶和华开启我的耳朵： “这罪孽直到你们死，断不得赦免！” 这是万军之主耶和华说的。
ISA|22|15|万军之主耶和华如此说：“你到 舍伯那 宫廷总管那里去，说：
ISA|22|16|‘你在这里凭什么？你在这里靠谁？竟敢在这里为自己凿坟墓，在高处为自己凿坟墓，在岩石中为自己挖安身之所！
ISA|22|17|你这伟大的人，看哪，耶和华必将你用力抛出，将你紧紧缠裹。
ISA|22|18|他必将你卷成一团，好像抛球一样抛向宽阔之地。你这主人家的羞辱啊，你必死在那里，你引以为荣的战车也毁在那里。
ISA|22|19|我要革除你的官职，你必从原位被逐 。’
ISA|22|20|“到那日，我要召 希勒家 的儿子─我的仆人 以利亚敬 来，
ISA|22|21|将你的外袍给他穿上，将你的腰带给他系紧，将你的政权交在他手中。他必作 耶路撒冷 居民和 犹大 家的父。
ISA|22|22|我要将 大卫 家的钥匙放在他肩头上。他开了，无人能关；他关了，无人能开。
ISA|22|23|我要使他立稳，像钉子钉在坚固的地方；他必成为他父家荣耀的宝座。
ISA|22|24|他父家所有的荣耀，连儿女带子孙，有如杯碗、瓶罐的小器皿，都挂在他身上。
ISA|22|25|当那日，万军之耶和华说，钉在坚固处的钉子必挪移，被砍断落地，挂在上面的各样重担都被切断。这是耶和华说的。”
ISA|23|1|论 推罗 的默示。 哀号吧， 他施 的船只！ 因为 推罗 已成废墟，没有房屋存留， 他们从 基提 地来的时候，得到这个消息 。
ISA|23|2|沿海的居民， 西顿 的商家啊， 当静默无声。 你差人航海 ，
ISA|23|3|在大水之上， 西曷河 的粮食、 尼罗河 的庄稼是 推罗 的进项， 它就成为列国的商埠。
ISA|23|4|西顿 ，你这海洋中的堡垒啊，应当羞愧， 因为大海说 ： “我未经历产痛，也没有生产， 未曾养育男孩，也没有抚养女孩。”
ISA|23|5|推罗 的风声传到 埃及 时， 他们为这风声极其疼痛。
ISA|23|6|你们当渡到 他施 去， 哀号吧，沿海的居民！
ISA|23|7|这就是你们那古老欢乐的城市吗？ 它的脚曾带人到远方居住。
ISA|23|8|谁定意 推罗 有这样的遭遇呢？ 它本是赐冠冕的， 它的商家是王子， 生意人是世上尊贵的人。
ISA|23|9|这是万军之耶和华所定的， 为要贬抑一切荣耀的狂傲， 使地上一切尊贵的人被藐视。
ISA|23|10|他施 啊， 你要像 尼罗河 一样在你的地泛滥， 不再有腰带的束缚了。
ISA|23|11|耶和华已经向海伸手， 震动列国； 他出令对付 迦南 ， 要拆毁其中的堡垒。
ISA|23|12|他说：“受欺压的少女 西顿 哪， 你必不再欢乐。 起来！渡到 基提 去， 就是在那里也不得安歇。
ISA|23|13|看哪， 迦勒底 人之地，这国民如今已不复存在。 亚述 人使它 成为住旷野者的居所。他们建筑自己的了望楼，拆毁它的宫殿，使它成为荒凉。
ISA|23|14|哀号吧， 他施 的船只！ 因你们的堡垒已成废墟。
ISA|23|15|到那时， 推罗 必被忘记七十年，就是一位君王的年数。七十年后， 推罗 的景况必如妓女之歌：
ISA|23|16|“你这被遗忘的妓女啊， 带着琴周游城内， 弹得美妙，唱许多歌， 好让人记得你。”
ISA|23|17|七十年后，耶和华必巡视 推罗 ，使它再度获利 ，与地面上的世界各国贸易 。
ISA|23|18|它的收益和获利都要归耶和华为圣，不再私自屯积存留；因为它的收益必归给住在耶和华面前的人，使他们吃饱，穿华丽的衣服。
ISA|24|1|看哪，耶和华使地空虚，变为荒芜， 地面扭曲，居民四散。
ISA|24|2|那时，百姓如何，祭司也如何； 仆人如何，主人也如何； 婢女如何，主母也如何； 买主如何，卖主也如何； 放债的如何，借贷的也如何； 债主如何，欠债的也如何。
ISA|24|3|地必全然空虚，尽都荒芜， 因为这话是耶和华说的。
ISA|24|4|大地悲哀凋零， 世界败落衰残， 地上居高位的人也没落了。
ISA|24|5|地被其上的居民所污秽， 因为他们犯了律法， 废了律例，背了永约。
ISA|24|6|所以，诅咒吞灭大地， 住在其上的都有罪； 地上的居民被火焚烧， 剩下的人稀少。
ISA|24|7|新酒悲哀，葡萄树凋残， 心中欢乐的都叹息。
ISA|24|8|击鼓之乐停止， 狂欢者的喧哗止住， 弹琴之乐也停止了。
ISA|24|9|人不再饮酒唱歌， 喝烈酒的，必以为苦。
ISA|24|10|荒凉的城拆毁了， 各家关闭，无法进入。
ISA|24|11|有人在街上嚷着要酒喝， 一切的喜乐变为昏暗， 地上的欢乐全都消失。
ISA|24|12|城里尽是荒凉， 城门全都摧毁。
ISA|24|13|地上的万民正像打过的橄榄树， 又如葡萄酿酒以后再去摘取，所剩无几。
ISA|24|14|他们要高声欢呼， 从海那边扬声赞美耶和华的威严。
ISA|24|15|因此，你们要在日出之地荣耀耶和华， 在众海岛荣耀耶和华－ 以色列 上帝的名。
ISA|24|16|我们听见从地极有人歌唱： “荣耀归于公义的那一位！” 我却说：“我灭亡了！ 我灭亡了，我有祸了！ 诡诈的还在行诡诈， 诡诈的还在大行诡诈。”
ISA|24|17|地上的居民哪， 惊吓、陷阱、罗网都临到你；
ISA|24|18|躲过惊吓之声的坠入陷阱， 逃离陷阱的又被罗网缠住， 因为天上的窗户都打开， 地的根基也震动。
ISA|24|19|地必全然破坏，尽都崩裂， 剧烈震动。
ISA|24|20|地要摇摇晃晃，好像醉酒的人， 又如小屋子摇来摇去； 罪过重压其上， 它就塌陷，不能复起。
ISA|24|21|到那日，耶和华在天上必惩罚天上的军队， 在地上必惩罚地上的列王。
ISA|24|22|他们必被聚集， 像囚犯困在牢里， 他们被关在监狱， 多日之后便受惩罚。
ISA|24|23|那时，月亮要蒙羞，太阳要惭愧， 因为万军之耶和华必在 锡安山 ， 在 耶路撒冷 作王， 在他众长老面前彰显荣耀。
ISA|25|1|耶和华啊，你是我的上帝， 我要尊崇你，称颂你的名。 因为你以信实忠信 行远古所定奇妙的事。
ISA|25|2|你使城市变为废墟， 使坚固的城荒凉， 使外邦人的城堡不再为城， 永远不再重建。
ISA|25|3|所以，强大的民必尊敬你， 残暴之国的城必敬畏你。
ISA|25|4|因为你是贫寒人的保障， 贫穷人急难中的保障， 暴风雨之避难所， 炎热地之阴凉处。 当残暴者盛气凌人的时候， 如暴风直吹墙壁，
ISA|25|5|如干旱地的热气， 你要制止外邦人的喧嚷， 残暴者的歌要停止， 好像热气因云的阴影而消失。
ISA|25|6|在这山上，万军之耶和华必为万民摆设宴席，有肥甘与美酒，就是满有骨髓的肥甘与精酿的美酒。
ISA|25|7|在这山上，他必吞灭缠裹万民的面纱和那遮盖列国的遮蔽物。
ISA|25|8|他已吞灭死亡直到永远。主耶和华必擦干各人脸上的眼泪，在全地除去他百姓的羞辱；这是耶和华说的。
ISA|25|9|到那日，人必说：“看哪，这是我们的上帝，我们向来等候他，他必拯救我们。这是耶和华，我们向来等候他，我们必因他的救恩欢喜快乐。”
ISA|25|10|耶和华的手必按住这山， 摩押 人要被践踏在他底下，好像干草被践踏在粪池 里。
ISA|25|11|他们要在其中伸展双手，好像游泳的人伸手游泳。他们的手虽灵巧，耶和华却使他们的骄傲降为卑下。
ISA|25|12|他使你城墙上坚固的碉堡倾倒，夷为平地，化为尘土。
ISA|26|1|当那日，在 犹大 地，人必唱这歌： “我们有坚固的城， 耶和华赐救恩为城墙，为城郭。
ISA|26|2|你们要敞开城门， 使守信的公义之民得以进入。
ISA|26|3|坚心倚赖你的，你必保守他十分平安， 因为他倚靠你。
ISA|26|4|你们当倚靠耶和华，直到永远， 因为耶和华，耶和华是永远的磐石。
ISA|26|5|他使居住高处的与高处的城市一同降为卑下， 将城拆毁，夷为平地，化为尘土，
ISA|26|6|使它被脚践踏， 就是被困苦人和贫寒人的脚践踏。”
ISA|26|7|义人的道是正直的， 正直的主啊，你修平义人的路。
ISA|26|8|耶和华啊，我们在你行审判的路上等候你 ， 我们心里所渴慕的，就是你的名和你的称号 。
ISA|26|9|夜间，我的心渴想你， 我里面的灵切切寻求你。 因为你在地上行审判的时候， 世上的居民就学习公义。
ISA|26|10|恶人虽然领受恩惠， 仍未学到公义。 在正直之地，他行不义， 也不看耶和华的威严。
ISA|26|11|耶和华啊，你的手高举，他们不观看； 愿他们观看你为百姓发的热心而羞愧， 愿火吞灭你的敌人。
ISA|26|12|耶和华啊，你必赏赐我们平安， 因为我们所做的一切，都是你为我们成就的。
ISA|26|13|耶和华－我们的上帝啊， 在你以外曾有别的主管辖我们， 但我们惟独称扬你的名。
ISA|26|14|死去的不能再复活， 阴魂不能再兴起； 你惩罚他们，使他们毁灭， 他们的名号 就全然消灭。
ISA|26|15|耶和华啊，你增添国民， 你增添国民，得了荣耀， 又拓展国土的疆界。
ISA|26|16|耶和华啊，他们在急难中寻求你。 你的管教临到他们身上时， 他们倾吐低声的祷告。
ISA|26|17|妇人怀孕，临产疼痛， 在痛苦之中喊叫； 耶和华啊，我们在你面前也是如此。
ISA|26|18|我们曾怀孕，曾疼痛， 所生产的竟像风一样， 并未带给地上任何拯救； 世上也未曾有居民生下来 。
ISA|26|19|你的死人要复活， 我的尸首要起来。 睡在尘土里的啊，要醒起歌唱！ 你的甘露好像晨曦 的甘露， 地要交出阴魂。
ISA|26|20|我的百姓啊，要进入内室， 关上你的门，躲避片刻， 等到愤怒过去。
ISA|26|21|因为，看哪，耶和华从他的居所出来， 要惩罚地上居民的罪孽。 地必露出其中的血， 不再掩盖被杀的人。
ISA|27|1|到那日，耶和华必用他坚硬锐利的大刀惩罚 力威亚探 ，就是那爬得快的蛇，惩罚 力威亚探 ，就是那弯弯曲曲的蛇，并杀死海里的大鱼。
ISA|27|2|当那日，你们要唱这美好 葡萄园的歌：
ISA|27|3|“我－耶和华看守葡萄园，按时灌溉， 昼夜看守，免得有人损害。
ISA|27|4|我心中不存愤怒。 惟愿在战争中我有荆棘和蒺藜， 我就起步攻击他， 把他一同焚烧；
ISA|27|5|或者让他紧靠我，以我为避难所， 与我和好， 与我和好。”
ISA|27|6|将来 雅各 要扎根， 以色列 要发芽开花， 果实遍满地面。
ISA|27|7|耶和华击打 以色列 ， 岂像击打那些击打他们的人吗？ 以色列 被杀戮， 岂像其他人所遭遇的杀戮吗？
ISA|27|8|你驱赶他们，放逐他们， 与他们相争。 在刮东风的日子， 他以暴风赶逐他们。
ISA|27|9|所以， 雅各 的罪孽藉此得赦免， 除罪的效果尽在乎此； 他使祭坛的石头变为粉碎的石灰， 使 亚舍拉 和香坛不再立起。
ISA|27|10|因为坚固的城变为荒凉， 成了被撇弃的居所，像旷野一样； 牛犊在那里吃草， 在那里躺卧，吃尽其中的树枝。
ISA|27|11|它的枝条一枯干，就被折断， 妇女用以点火燃烧。 因为这百姓蒙昧无知， 所以，造他们的必不怜悯他们， 造成他们的也不施恩给他们。
ISA|27|12|到那日， 以色列 人哪，耶和华必像人打树拾果一般，从 大河 的支流，直到 埃及 的溪谷，将你们一一收集。
ISA|27|13|当那日，号角大响；在 亚述 地将亡的，与被赶散至 埃及 地的，都要前来，在 耶路撒冷 圣山上敬拜耶和华。
ISA|28|1|祸哉！ 以法莲 酒徒高傲的冠冕， 其荣美竟如花凋残； 他们在肥沃的山谷顶上， 被酒击败。
ISA|28|2|看哪，主有一位大能大力者， 如强烈的冰雹， 如毁灭的暴风雨， 如涨溢的洪水， 他必亲手将他们摔落在地。
ISA|28|3|以法莲 酒徒高傲的冠冕， 必被脚践踏；
ISA|28|4|那如凋残之花的荣美， 在肥沃的山谷顶上， 必如夏令前初熟的无花果， 让看见的人注意， 摘到手里，随即吞吃。
ISA|28|5|到那日，万军之耶和华 必成为他余民的荣冠华冕，
ISA|28|6|成为在位审判者的公平之灵， 和城门口制敌的力量。
ISA|28|7|这些人也因酒摇晃， 因烈酒东倒西歪。 祭司和先知因烈酒摇晃， 被酒所困， 因烈酒东倒西歪。 他们错解默示， 审判时不分是非。
ISA|28|8|筵席上都满了呕吐的污秽， 没有一处干净。
ISA|28|9|“他要将知识指教谁呢？ 要向谁阐明信息呢？ 是向那些刚断奶的， 离开母亲胸怀的吗？
ISA|28|10|因为他咕哝咕哝，咕哝咕哝， 唠唠叨叨，唠唠叨叨， 这里一点，那里一点。”
ISA|28|11|耶和华要藉嘲弄的嘴唇和外邦人的舌头， 向这百姓说话。
ISA|28|12|他曾对他们说： “这是安歇之所， 你们要使疲乏的人得安歇， 这是歇息之处。” 他们却不肯听。
ISA|28|13|耶和华的话对他们而言是 “咕哝咕哝，咕哝咕哝， 唠唠叨叨， 唠唠叨叨， 这里一点，那里一点”； 以致他们往前行， 却后仰跌倒，甚至跌伤， 落入陷阱，被抓住了。
ISA|28|14|因此，你们这些傲慢的人， 就是管辖住 耶路撒冷 这百姓的， 要听耶和华的话。
ISA|28|15|你们曾说： “我们已与死亡立约， 与阴间结盟， 不可挡的鞭子挥过时， 必不临到我们； 因我们以谎言为避难所， 靠虚假来藏身”；
ISA|28|16|所以，主耶和华如此说： “看哪，我在 锡安 放一块石头作为根基， 是衡量的石头， 是宝贵的房角石，稳固的根基； 信靠他的人必不致惊恐。
ISA|28|17|我以公平为准绳， 以公义为铅垂线； 冰雹必冲去谎言的避难所， 大水必漫过藏身之处。
ISA|28|18|你们与死亡所立的约必废除， 与阴间所结的盟不得坚立； 不可挡的鞭子挥过时， 你们必被践踏。
ISA|28|19|每逢它挥来，必将你们掳去； 每早晨它必挥过， 白昼黑夜都是如此。 明白这信息的都必惊恐。”
ISA|28|20|床榻短，人不能伸展； 被子窄，人无从裹身。
ISA|28|21|耶和华必兴起，像在 毗拉心山 ， 他必发怒，如在 基遍谷 ； 为要做成他的工，就是非常的工， 成就他的事，就是奇异的事。
ISA|28|22|现在你们不可傲慢， 免得捆绑你们的绳索更结实， 因为我从万军之主耶和华那里听见， 在全地施行灭绝的事已定。
ISA|28|23|你们当侧耳听我的声音， 留心听我的言语。
ISA|28|24|那为撒种而耕地的 会不停地耕地，松土，耙地吗？
ISA|28|25|他铲平了地面， 岂不就种小茴香， 播种大茴香， 按行列种小麦， 在定处种大麦， 在田边种粗麦吗？
ISA|28|26|他的上帝教导他， 指导他合宜的方法。
ISA|28|27|原来打小茴香，不用尖利的器具， 轧大茴香，也不是用车轮； 却要用杖打小茴香， 用棍打大茴香。
ISA|28|28|谷要打， 但不能持续地捣， 用车轮和马轧， 却不轧碎它。
ISA|28|29|这也是出于万军之耶和华， 他的谋略奇妙， 他的智慧广大。
ISA|29|1|祸哉！ 亚利伊勒 ， 亚利伊勒 ， 大卫 安营的城， 任凭你年复一年， 节期照常循环，
ISA|29|2|我却要使 亚利伊勒 遭难； 它必悲伤哀号， 它对我是 亚利伊勒 。
ISA|29|3|我必四围安营攻击你， 筑台围困你， 堆垒攻击你。
ISA|29|4|你必败落，从地里说话， 你的言语细微出于尘埃。 你的声音必像那招魂者的声音出于地， 你的言语呢喃出于尘埃。
ISA|29|5|你那成群的陌生人 要像细尘， 暴民要像吹起的糠秕； 这事必顷刻之间忽然临到。
ISA|29|6|万军之耶和华必使雷轰、地震、巨响、旋风、暴风， 并吞灭的火焰临到它。
ISA|29|7|那时，攻击 亚利伊勒 列国的军队， 与一切攻击 亚利伊勒 和它城堡， 并带给它患难的， 必如梦，如夜间的异象；
ISA|29|8|又像饥饿的人在梦中吃饭， 醒了仍觉饥肠辘辘； 或像口渴的人在梦中喝水， 醒了仍觉发昏，心里想喝。 攻击 锡安山 列国的军队也必如此。
ISA|29|9|你们等候惊奇吧！ 你们沉迷宴乐吧！ 他们醉了，却非因酒； 东倒西歪，却非因烈酒。
ISA|29|10|因为耶和华将沉睡的灵浇灌你们， 遮住你们的眼， 眼就是先知， 覆盖你们的头， 头就是先见。
ISA|29|11|所有的默示，在你们看来都如封住的书卷，人将这书卷交给识字的人，说：“请念吧！”他说：“我不能念，因为它封住了。”
ISA|29|12|又将这书卷交给不识字的人，说：“请念吧！”他说：“我不识字。”
ISA|29|13|主说：“因这百姓以口亲近我， 用嘴唇尊敬我， 心却远离我； 他们敬畏我， 不过是领受前人的命令。
ISA|29|14|所以，看哪，我要在这百姓中行奇妙的事， 就是奇妙又奇妙的事。 他们智慧人的智慧必然消灭， 聪明人的聪明必然消失。”
ISA|29|15|祸哉！那些向耶和华深藏谋略的， 他们在暗中行事，说： “有谁看见我们呢？ 谁会注意我们呢？”
ISA|29|16|你们把事情颠倒了， 岂可看陶匠如陶土呢？ 受造物岂可论创造者说， “他并没有造我”？ 制成物岂可论制作者说， “他根本不懂”？
ISA|29|17|黎巴嫩 变为田园， 田园看似森林， 不是只需要一些时间吗？
ISA|29|18|那时，聋子必听见这书上的话； 盲人的眼必从迷蒙黑暗中看见。
ISA|29|19|困苦的人必因耶和华增添欢喜， 人间贫穷的必因 以色列 的圣者快乐。
ISA|29|20|因为残暴的人归于无有， 傲慢的人已经灭绝， 一切存心作恶的都被剪除。
ISA|29|21|他们凭一句话定一个人有罪， 为在城门口断是非的设下罗网， 又用虚无的事屈枉义人。
ISA|29|22|所以，救赎 亚伯拉罕 的耶和华 论到 雅各 家时如此说： “ 雅各 必不再羞愧， 面容也不再变色。
ISA|29|23|当他的儿女看见 我的手在他们当中所成就的事情 ， 他们就必尊我的名为圣， 尊 雅各 的圣者为圣， 他们必敬畏 以色列 的上帝。
ISA|29|24|心中迷糊的必明白， 发怨言的必领受训诲。”
ISA|30|1|耶和华说： “祸哉！这悖逆的儿女。 他们同谋，却不出于我， 结盟，却不出于我的灵， 以致罪上加罪。
ISA|30|2|他们没有寻求我的指示，就起身下 埃及 去， 要倚靠法老的庇护坚固自己， 并投在 埃及 的荫下。
ISA|30|3|但法老的庇护反成为你们的羞辱； 你们投在 埃及 荫下，反使你们惭愧。
ISA|30|4|他们的领袖已在 琐安 ， 他们的使臣到了 哈内斯 。
ISA|30|5|他们必因那无益于他们的民蒙羞； 那民并非帮助，也非有益， 只带来羞耻和凌辱。”
ISA|30|6|论 尼革夫 牲畜的默示。 他们将财物驮在驴背上， 将宝物驮在骆驼的背脊， 经过艰难困苦之地， 就是母狮、公狮、毒蛇、飞蛇之地， 往那无益于他们的民那里去。
ISA|30|7|埃及 的帮助是徒然的， 因此，我称它为“毫不中用的 拉哈伯 ” 。
ISA|30|8|现在你要去， 在他们面前将这话刻在版上， 写在书上， 以便流传后世，直到永永远远 。
ISA|30|9|因为他们是悖逆的百姓、说谎的儿女， 是不肯听从耶和华训诲的儿女。
ISA|30|10|他们对先见说：“不要再看了”； 对先知说：“不要向我们预言正直的事； 要对我们说好听的话， 预言虚幻的事。
ISA|30|11|要离开这道，偏离这路， 不要在我们面前再提说 以色列 的圣者。”
ISA|30|12|所以， 以色列 的圣者如此说： “因你们藐视这话， 倚赖欺压和诡诈，以此为可靠，
ISA|30|13|因此，这罪孽在你们身上， 好像高墙里有凸起的裂缝， 顷刻之间忽然坍下来了；
ISA|30|14|它被砸碎，好像把陶匠的瓦器摔碎， 毫不顾惜， 甚至在碎块中找不到一片 可用以从炉内取火，或从池中舀水。
ISA|30|15|主耶和华－ 以色列 的圣者如此说： “你们得救在乎归回安息， 得力在乎平静安稳。” 你们却是不肯，
ISA|30|16|你们说：“不然，我们要骑马奔走”， 所以你们必然奔走。 你们又说：“我们要骑快马”， 所以追赶你们的，也必飞快。
ISA|30|17|一人叱喝，令千人逃跑， 五人叱喝，你们都逃跑； 以致剩下的如山顶的旗杆， 如山冈上的大旗。
ISA|30|18|耶和华必然等候，要施恩给你们； 必然兴起，好怜悯你们。 因为耶和华是公平的上帝； 凡等候他的都是有福的！
ISA|30|19|住在 锡安 、居于 耶路撒冷 的百姓啊，你必不再哭泣。主必因你哀求的声音施恩给你，他听见的时候就必应允你。
ISA|30|20|主虽然以艰难给你当饼，以困苦给你当水，你的教师却不再隐藏，你的眼睛必看见你的教师。
ISA|30|21|你或向左或向右，必听见后边有声音说：“这是正路，要行在其间。”
ISA|30|22|你要玷污那雕刻偶像所包的银子和铸造偶像所镀的金子。你要抛弃它们，如抛弃污秽之物；对偶像说：“去吧！”
ISA|30|23|你撒种在地里，主必降雨在其上，使地所出的粮食肥美丰盛。那时，你的牲畜必在辽阔的草场吃草。
ISA|30|24|耕地的牛和驴必吃加盐的饲料，是用铲子和杈子扬净的。
ISA|30|25|在大行杀戮的日子，城楼倒塌的时候，高山峻岭必有川河涌流。
ISA|30|26|当耶和华包扎他百姓的伤口，医治他所击打伤痕的日子，月光必像日光，日光必加七倍，像七日的光一样。
ISA|30|27|看哪，耶和华的名从远方来， 他的怒气烧起，浓烟上腾。 他的嘴唇满有愤恨， 他的舌头像吞灭的火。
ISA|30|28|他的气息如涨溢的河水，直涨到颈项， 要用毁灭的筛网筛净列国， 并在众民口中安放导错方向的嚼环。
ISA|30|29|你们必唱歌，像守圣节的夜间一样；并且心中喜乐，像人吹笛，来到耶和华的山，到 以色列 的磐石那里。
ISA|30|30|耶和华必使人听见他威严的声音，又以极大的愤怒、吞灭的火焰、雷雨、暴风和像石块的冰雹，使人看见他降罚的膀臂。
ISA|30|31|亚述 必因耶和华的声音惊惶，耶和华必用杖击打它。
ISA|30|32|耶和华必将定规要打 的杖加在它身上；每打一下，都必配合击鼓弹琴的节奏。打仗时，耶和华必振臂与它交战。
ISA|30|33|原来 陀斐特 早已预备好了，是为君王预备的；又深又宽，堆满了火和木柴；耶和华的气息犹如一股硫磺使它燃起。
ISA|31|1|祸哉！那些下 埃及 求帮助的， 他们仰赖马匹，倚靠甚多的战车， 并倚靠强壮的骑兵， 却不仰望 以色列 的圣者， 也不求问耶和华。
ISA|31|2|其实，耶和华有智慧， 他降灾祸， 并不撤回自己的话， 却要兴起攻击作恶之家， 攻击那帮助人作恶的。
ISA|31|3|埃及 人不过是人，并非上帝， 他们的马不过是血肉，并不是灵。 耶和华一伸手， 那帮助人的必绊跌，受帮助的也必跌倒， 都一同灭亡。
ISA|31|4|耶和华对我如此说， 狮子和少壮狮子为猎物而咆哮， 许多牧人被召来攻击它， 它总不因他们的声音惊惶， 也不因他们的喧嚷退缩； 万军之耶和华也必如此 降临在 锡安 的大小山冈上争战。
ISA|31|5|雀鸟盘旋护卫， 万军之耶和华也必照样保护 耶路撒冷 ； 他必保护拯救， 必逾越而搭救。
ISA|31|6|以色列 人哪，要归向你们严重悖逆的那一位！
ISA|31|7|到那日，你们各人要抛弃亲手所造、陷自己于罪中的金偶像和银偶像。
ISA|31|8|亚述 必倒在刀下，并非人的刀； 有刀要将它吞灭，并非人的刀。 它要逃避这刀， 它的年轻人必做苦工。
ISA|31|9|它的磐石必因惊吓而消失， 它的领袖必因大旗惊惶； 这是那有火在 锡安 、 有炉在 耶路撒冷 的耶和华说的。
ISA|32|1|看哪，必有一位君王凭公义执政， 必有王子藉公平掌权。
ISA|32|2|必有一人如避风港， 如暴风雨的藏身处； 如干旱地的溪流， 又如干燥地巨石的阴影。
ISA|32|3|看的人眼睛不再昏花， 听的人耳朵必留心听。
ISA|32|4|性急的人懂得分辨， 口吃的人说话流畅。
ISA|32|5|愚顽人不再称为君子， 流氓不再称为绅士。
ISA|32|6|因为愚顽人必说愚妄的话， 他的心作恶 ， 行亵渎的事， 传播恶言攻击耶和华， 使饥饿的人仍然饥饿， 口渴的人无水可喝。
ISA|32|7|流氓的手段邪恶， 他图谋恶计， 用谎言毁灭困苦人； 贫穷人讲求公理时， 他也是如此行。
ISA|32|8|君子却图谋高尚的事， 他必因高尚的事站立得稳。
ISA|32|9|安逸的妇女啊，起来听我的声音！ 无虑的女子啊，侧耳听我的言语！
ISA|32|10|无虑的女子啊，再过一年，你们必颤栗， 因为无葡萄可摘， 也无果实可收。
ISA|32|11|安逸的妇女啊，要战兢； 无虑的女子啊，要颤栗， 要脱去衣服，赤着身体， 腰束麻布。
ISA|32|12|你们要为美好的田地 和多结果子的葡萄树捶胸哀哭。
ISA|32|13|刺草和荆棘要长在我百姓的田地上， 长在欢乐城中一切快乐家园上。
ISA|32|14|宫殿必被撇下， 繁华的城必被抛弃， 堡垒和了望楼永为洞穴， 成为野驴的乐土， 羊群的草场。
ISA|32|15|等到圣灵从高处浇灌我们， 旷野将变为田园， 田园看似森林。
ISA|32|16|公平要居住在旷野， 公义要安歇在田园。
ISA|32|17|公义的果实是平安， 公义的效果是平静和安稳，直到永远。
ISA|32|18|我的百姓要住在平安的居所， 安稳的住处，宁静的安歇之地。
ISA|32|19|虽有冰雹击倒树林， 城也夷为平地；
ISA|32|20|然而你们在水边撒种， 牧放牛驴的有福了！
ISA|33|1|祸哉！你这未遭毁灭而毁灭人的人， 人未以诡诈待你而你以诡诈待人的人！ 等你行完了毁灭， 自己必被毁灭； 你行完了诡诈， 人必以诡诈待你。
ISA|33|2|耶和华啊，求你施恩给我们， 我们等候你。 求你每早晨作我们的膀臂， 遭难时作我们的拯救。
ISA|33|3|轰然之声一发出，万民就奔逃； 你一兴起 ，列国就四散。
ISA|33|4|你们的掳物必被敛尽， 有如蚂蚱敛尽禾稼； 人为掳物奔走，宛如蝗虫蹦跳。
ISA|33|5|耶和华受尊崇，居高处， 使公平和公义充满 锡安 。
ISA|33|6|他是你这世代安定的力量， 丰盛的救恩、 智慧和知识； 敬畏耶和华是 锡安 的至宝。
ISA|33|7|看哪，他们的英雄在外面哀号 ， 求和的使臣在痛哭。
ISA|33|8|大路荒凉，行人止息； 盟约撕毁，见证 被弃， 人也不受尊重。
ISA|33|9|大地悲哀衰残， 黎巴嫩 羞愧且枯干， 沙仑 好像旷野， 巴珊 和 迦密 必凋残。
ISA|33|10|耶和华说： “现在我要兴起， 要高升， 要受尊崇。
ISA|33|11|你们怀的是糠秕，生的是碎秸； 你们的气息如火吞灭自己。
ISA|33|12|万民必像烧着的石灰， 又如斩断的荆棘，在火里燃烧。”
ISA|33|13|你们远方的人，当听我所做的事； 你们近处的人，当承认我的大能。
ISA|33|14|锡安 的罪人都惧怕， 战兢抓住不敬虔的人。 我们中间有谁能与吞噬的火同住？ 我们中间有谁能与不灭的火共存呢？
ISA|33|15|那行事公义、说话正直、 憎恶欺压所得之财、 摇手不受贿赂、 掩耳不听流血的计谋、 闭眼不看邪恶之事的，
ISA|33|16|这人必居高处， 他的保障是磐石的堡垒， 必有粮食赐给他， 饮水也不致断绝。
ISA|33|17|你必亲眼看见君王的荣美， 看见辽阔之地。
ISA|33|18|你的心必回想那些恐怖的事： “那数算的人在哪里？ 秤重的人在哪里？ 数点城楼的又在哪里呢？”
ISA|33|19|你必不再看见那凶暴的民， 他们嘴唇说艰涩的言语，难以理解； 舌头结巴，说无意义的话。
ISA|33|20|你要注视 锡安 ，我们守圣节的城！ 你必亲眼看见 耶路撒冷 成为安静的居所， 成为不挪移的帐幕， 橛子永不拔出， 绳索一根也不折断。
ISA|33|21|在那里，威严的耶和华对我们是宽阔的江河， 其中必没有摇桨的小船来往， 也没有巨大的船舶经过。
ISA|33|22|耶和华是审判我们的， 耶和华为我们设立律法； 耶和华是我们的君王， 他必拯救我们。
ISA|33|23|船上的绳索松开， 不能稳住桅杆， 也无法扬起船帆。 那时许多掳物被瓜分， 连瘸腿的也能夺走掠物。
ISA|33|24|城内的居民无人说：“我病了”； 城里居住的百姓，罪孽都蒙赦免。
ISA|34|1|列国啊，要近前来听！ 万民哪，要侧耳而听！ 全地和其上所充满的， 世界和其中所出的，都应当听！
ISA|34|2|因为耶和华向列国发怒， 向他们的全军发烈怒， 要将他们灭尽，任人杀戮。
ISA|34|3|被杀的人必被抛弃， 尸首臭气上腾， 诸山为他们的血所融化。
ISA|34|4|天上万象都要朽坏， 天被卷起，有如书卷， 其上的万象尽都衰残； 如葡萄树的叶子凋落， 又如无花果树枯萎一样。
ISA|34|5|因为我的刀在天上将要显现 ； 看哪，这刀临到 以东 和我所诅咒的民， 要施行审判。
ISA|34|6|耶和华的刀沾满了血， 是用油脂和羔羊、公山羊的血， 并公绵羊肾上的油脂滋润的； 因为在 波斯拉 有祭物献给耶和华， 在 以东 地有大屠杀。
ISA|34|7|野牛与他们一起倒下， 牛犊和壮牛也一同倒下。 他们的地被血染遍， 他们的尘土因油脂肥润。
ISA|34|8|这是耶和华报仇之日， 为 锡安 伸冤的报应之年。
ISA|34|9|它的河水要变为柏油， 尘埃变为硫磺， 大地成为燃烧的柏油，
ISA|34|10|昼夜总不熄灭， 它的烟永远上腾， 必世世代代成为荒废， 永永远远无人经过。
ISA|34|11|鹈鹕、豪猪要得它为业， 猫头鹰、乌鸦要住在其间。 耶和华必将空虚的准绳、 混沌的石垂线，拉在 以东 之上。
ISA|34|12|人必宣称那里没有王国， 它的贵族和所有领袖都归于无有。
ISA|34|13|以东 的宫殿要长出荆棘， 城堡要生长蒺藜和刺草； 成为野狗的住处， 鸵鸟的居所。
ISA|34|14|野兽要和土狼相遇， 山羊鬼魔要与同伴对唱， 莉莉丝 必在那里栖身， 为自己寻找安歇之处。
ISA|34|15|箭头蛇要在那里做窝， 下蛋，孵蛋，并招聚幼蛇在其保护之下； 鹞鹰也与伴侣聚集在那里。
ISA|34|16|你们要查考并诵读耶和华的书； 这些现象必然存在， 没有一样动物缺少伴侣。 因为是他，藉着我的口 吩咐， 他的灵将它们聚集。
ISA|34|17|他为它们抽签， 亲手用准绳为它们分地； 直到它们永远得地为业， 世世代代住在其间。
ISA|35|1|旷野和干旱之地必然欢喜， 沙漠也必快乐； 又如玫瑰绽放，
ISA|35|2|朵朵繁茂， 其乐融融，而且欢呼。 黎巴嫩 的荣耀， 并 迦密 与 沙仑 的华美，必赐给它。 人要看见耶和华的荣耀， 看见我们上帝的荣美。
ISA|35|3|你们要使软弱的手强壮， 使无力的膝盖稳固；
ISA|35|4|对心里焦急的人说： “要刚强，不要惧怕。 看哪，你们的上帝要来施报， 要施行极大的报应， 他必来拯救你们。”
ISA|35|5|那时，盲人的眼必睁开， 聋子的耳必开通。
ISA|35|6|那时，瘸子必跳跃如鹿， 哑巴的舌头必欢呼。 在旷野有水喷出， 在沙漠有江河涌流。
ISA|35|7|火热之地要变为水池， 干渴之地要变为泉源。 野狗躺卧休息之处 必长出青草、芦苇和蒲草。
ISA|35|8|在那里必有一条大道， 就是一条路 ，称为圣路。 污秽的人不得经过， 是专为走路的人 预备的， 愚昧的人也不会迷路。
ISA|35|9|在那里没有狮子， 猛兽也不经过； 在那里它们未现踪迹， 只有救赎的民在那里行走。
ISA|35|10|耶和华救赎的民必归回， 歌唱来到 锡安 ； 永远的快乐必归到他们头上， 他们必得着欢喜快乐， 忧伤叹息尽都逃避。
ISA|36|1|希西家 王十四年， 亚述 王 西拿基立 上来攻击 犹大 的一切坚固的城，将城攻取。
ISA|36|2|亚述 王从 拉吉 差遣将军 率领大军前往 耶路撒冷 ，到 希西家 王那里去。将军站在 上池 的水沟旁，在往漂布地的大路上。
ISA|36|3|希勒家 的儿子 以利亚敬 宫廷总管、 舍伯那 书记和 亚萨 的儿子 约亚 史官，出来见他。
ISA|36|4|将军对他们说：“你们去告诉 希西家 ，大王 亚述 王如此说：‘你倚靠什么，让你如此自信满满？
ISA|36|5|我说 ，你有打仗的计谋和能力，我看不过是空话。你到底倚靠谁，竟敢背叛我呢？
ISA|36|6|看哪，你所倚靠的 埃及 是那断裂的苇杖，人若倚靠这杖，它就刺进他的手，穿透它。 埃及 王法老向所有倚靠他的人都是这样。
ISA|36|7|你若对我说：我们倚靠耶和华－我们的上帝， 希西家 岂不是将上帝的丘坛和祭坛废去，并且吩咐 犹大 和 耶路撒冷 的人说：你们只当在这一个坛前敬拜吗？
ISA|36|8|现在你与我主 亚述 王打赌，我给你两千匹马，看你能否派得出骑士来骑它们。
ISA|36|9|若不然，怎能使我主臣仆中最小的一个军官转脸而逃呢？你难道要倚靠 埃及 的战车和骑兵吗？
ISA|36|10|现在我上来攻击毁灭这地，岂不是出于耶和华吗？耶和华吩咐我说，你上去攻击这地，毁灭它吧！’”
ISA|36|11|以利亚敬 、 舍伯那 、 约亚 对将军说：“求你用 亚兰 话对仆人说，因为我们听得懂；不要用 犹大 话对我们说，免得传到城墙上百姓的耳中。”
ISA|36|12|将军说：“我主差遣我来，岂是单对你和你的主人说这些话吗？不也是对这些坐在城墙上，要与你们一同吃自己粪、喝自己尿的人说的吗？”
ISA|36|13|于是 亚述 将军站着，用 犹大 话大声喊着说：“你们当听大王 亚述 王的话，
ISA|36|14|王如此说：‘你们不要被 希西家 欺哄了，因他不能拯救你们。
ISA|36|15|不要听凭 希西家 说服你们倚靠耶和华，他说，耶和华必要拯救我们，这城必不交在 亚述 王的手中。’
ISA|36|16|你们不要听 希西家 的话！因 亚述 王如此说：‘你们要与我讲和，出来投降，各人就可以吃自己葡萄树和无花果树的果子，喝自己井里的水，
ISA|36|17|等我来领你们到一个地方，与你们本地一样，就是有五谷和新酒之地，有粮食和葡萄园之地。
ISA|36|18|恐怕 希西家 误导你们说，耶和华必拯救我们。列国的神明有哪一个曾救它本国脱离 亚述 王的手呢？
ISA|36|19|哈马 和 亚珥拔 的神明在哪里呢？ 西法瓦音 的神明在哪里呢？它们曾救 撒玛利亚 脱离我的手吗？
ISA|36|20|这些国的神明有谁曾救自己的国家脱离我的手呢？难道耶和华能救 耶路撒冷 脱离我的手吗？’”
ISA|36|21|百姓静默不言，一句不答，因为 希西家 王曾吩咐说：“不要回答他。”
ISA|36|22|当下 希勒家 的儿子 以利亚敬 宫廷总管、 舍伯那 书记，和 亚萨 的儿子 约亚 史官都撕裂衣服，来到 希西家 那里，将 亚述 将军的话告诉他。
ISA|37|1|希西家 王听见了，就撕裂衣服，披上麻布，进了耶和华的殿。
ISA|37|2|他差遣 以利亚敬 宫廷总管和 舍伯那 书记，并祭司中年长的，都披上麻布，到 亚摩斯 的儿子 以赛亚 先知那里去。
ISA|37|3|他们对他说：“ 希西家 如此说：‘今日是急难、惩罚、凌辱的日子，就如婴孩快要出生，却没有力气生产。
ISA|37|4|或许耶和华－你的上帝听见 亚述 将军的话，就是他主人 亚述 王差他来辱骂永生上帝的话，耶和华－你的上帝就斥责所听见的这些话。求你为幸存的余民扬声祷告。’”
ISA|37|5|希西家 王的臣仆就来到 以赛亚 那里。
ISA|37|6|以赛亚 对他们说：“要对你们的主人这样说，耶和华如此说：‘你听见 亚述 王的仆人亵渎我的话，不要惧怕。
ISA|37|7|看哪，因为我必惊动他的心 ，他要听见风声就归回本地，在那里我必使他倒在刀下。’”
ISA|37|8|亚述 将军听见 亚述 王已拔营离开 拉吉 ，就启程返回，正遇见 亚述 王去攻打 立拿 。
ISA|37|9|亚述 王听见有人谈论 古实 王 特哈加 说：“他出来要与你争战。” 亚述 王一听见，就差使者去见 希西家 ，说：
ISA|37|10|“你们要对 犹大 王 希西家 如此说：‘不要听你所倚靠的上帝欺哄你说： 耶路撒冷 必不交在 亚述 王的手中。
ISA|37|11|看哪，你总听说 亚述 诸王向列国所行的是尽行灭绝，难道你能幸免吗？
ISA|37|12|我祖先所毁灭的，就是 歌散 、 哈兰 、 利色 和 提．拉撒 的 伊甸 人；这些国的神明何曾拯救他们呢？
ISA|37|13|哈马 的王， 亚珥拔 的王， 西法瓦音城 的王， 希拿 和 以瓦 的王，都在哪里呢？’”
ISA|37|14|希西家 从使者手里接过书信，看完了，就上耶和华的殿，在耶和华面前展开书信。
ISA|37|15|希西家 向耶和华祷告说：
ISA|37|16|“坐在基路伯之上万军之耶和华－ 以色列 的上帝啊，你，惟有你是地上万国的上帝，你创造了天和地。
ISA|37|17|耶和华啊，求你侧耳而听；耶和华啊，求你睁眼而看，听 西拿基立 差遣使者辱骂永生上帝的一切话。
ISA|37|18|耶和华啊， 亚述 诸王果然使列国和列国之地变为荒芜，
ISA|37|19|将列国的神明扔在火里，因为它们不是神明，是人手所造的，是木头、石头，所以被灭绝了。
ISA|37|20|耶和华－我们的上帝啊，现在求你救我们脱离 亚述 王的手，使地上万国都知道惟有你是耶和华。”
ISA|37|21|亚摩斯 的儿子 以赛亚 就差人去见 希西家 ，说：“耶和华－ 以色列 的上帝如此说，你因 亚述 王 西拿基立 的事向我祈求，
ISA|37|22|所以耶和华论他这样说： ‘少女 锡安 藐视你，嘲笑你； 耶路撒冷 向你摇头。
ISA|37|23|“‘你辱骂谁，亵渎谁， 扬起声来，高举眼目攻击谁呢？ 你攻击的是 以色列 的圣者。
ISA|37|24|你藉臣仆辱骂主说： 我率领许多战车登上高山， 到 黎巴嫩 的顶端； 我要砍伐其中高大的香柏树 和上好的松树。 我必上到极高之处， 进入茂盛的森林里。
ISA|37|25|我已经挖井喝水 我必用脚掌踏干 埃及 一切的河流。
ISA|37|26|“‘你岂没有听见 我早先所定、古时所立、现今实现的事吗？ 就是让你去毁坏坚固的城镇，使它们变为废墟；
ISA|37|27|城里居民的力量甚小， 他们惊惶羞愧； 像野草，像青菜， 如房顶上的草， 被东风刮散 。
ISA|37|28|“‘你站起，你坐下，你出去，你进来， 你向我发烈怒，我都知道。
ISA|37|29|因你向我发烈怒， 你的狂傲上达我耳中， 我要用钩子钩住你的鼻子， 将嚼环放在你口里， 使你从原路转回去。’
ISA|37|30|“我赐给你的预兆：你们今年要吃野生的，明年也要吃自长的；后年，你们就要耕种收割，栽葡萄园，吃其中的果子。
ISA|37|31|犹大 家所逃脱剩余的，仍要往下扎根，向上结果。
ISA|37|32|必有剩余的民从 耶路撒冷 而出；有逃脱的人从 锡安山 而来。万军之耶和华的热心必成就这事。
ISA|37|33|“所以耶和华论 亚述 王如此说：他必不得来到这城，也不在这里射箭，不得拿盾牌到城前，也不能建土堆攻城。
ISA|37|34|他从哪条路来，必从那条路回去，必不得来到这城。这是耶和华说的。
ISA|37|35|因我为自己的缘故，又为我仆人 大卫 的缘故，必保护拯救这城。”
ISA|37|36|耶和华的使者出去，在 亚述 营中杀了十八万五千人。清早有人起来，看哪，都是死尸。
ISA|37|37|亚述 王 西拿基立 就拔营回去，住在 尼尼微 。
ISA|37|38|一日，他在他的神明 尼斯洛 庙里叩拜，他儿子 亚得米勒 和 沙利色 用刀杀了他，然后逃到 亚拉腊 地；他儿子 以撒．哈顿 接续他作王。
ISA|38|1|那些日子， 希西家 病得要死， 亚摩斯 的儿子 以赛亚 先知来见他，对他说：“耶和华如此说：‘你当留遗嘱给你的家，因为你必死，不能活了。’”
ISA|38|2|希西家 就转脸朝墙，向耶和华祷告，
ISA|38|3|说：“耶和华啊，求你记念我在你面前怎样存完全的心，按诚实行事，又做你眼中看为善的事。” 希西家 就痛哭。
ISA|38|4|耶和华的话临到 以赛亚 说：
ISA|38|5|“你去告诉 希西家 说，耶和华－你祖先 大卫 的上帝如此说：‘我听见了你的祷告，看见了你的眼泪。看哪，我必加添你十五年的寿数；
ISA|38|6|我要救你和这城脱离 亚述 王的手，也要保护这城。’
ISA|38|7|“耶和华必成就他所说的这话。这是耶和华给你的预兆：
ISA|38|8|看哪，我要使 亚哈斯 日晷上随太阳前进的影子，往后退十度。”于是，在日晷上照下来的日影果然往后退了十度。
ISA|38|9|犹大 王 希西家 患病痊愈后的诗：
ISA|38|10|我说，在如日中天的时候我就走了， 将剩余的年岁交给阴间的门。
ISA|38|11|我说，我必不得见耶和华，不得在活人之地见耶和华， 也不再看见世人，就是短暂世界 中的居民。
ISA|38|12|我的住处好像牧人的帐棚， 遭人掀起，离我而去； 我将性命卷起， 像织布的卷布一样。 他从织布机头那里将我剪断， 你使我命丧于旦夕。
ISA|38|13|我令自己安静 直到天亮； 他像狮子折断我所有的骨头， 你使我命丧于旦夕。
ISA|38|14|我像燕子呢喃， 像白鹤鸣叫， 又如鸽子哀鸣； 我因仰望，眼睛困倦。 主啊，我受欺压， 求你为我作保。
ISA|38|15|我还有什么可说的呢？ 他应许我的 ，他已成就了。 我因心里的苦楚， 在一生的年日必谦卑而行 。
ISA|38|16|主啊，人得存活是在乎此， 我的灵存活也全在乎此 ； 求你使我痊愈，仍然存活。
ISA|38|17|看哪，我受大苦是为使我得平安； 你爱我，救我的性命脱离败坏的地府， 将我一切的罪扔在你背后。
ISA|38|18|原来，阴间不能称谢你， 死亡不能颂扬你， 下到地府的人也不能盼望你的信实。
ISA|38|19|只有活人，活人必称谢你， 像我今日称谢你一样。 为父的，必使儿女知道你的信实。
ISA|38|20|耶和华肯救我， 所以，我们要一生一世 在耶和华殿中 弹奏我弦乐的歌。
ISA|38|21|以赛亚 说：“拿一块无花果饼来，贴在疮上，王必痊愈。”
ISA|38|22|希西家 说：“我能上耶和华的殿，有什么预兆呢？”
ISA|39|1|那时， 巴拉但 的儿子， 巴比伦 王 米罗达．巴拉但 听见 希西家 病得痊愈，就送书信和礼物给他。
ISA|39|2|希西家 欢喜见使者，就将自己宝库里的金子、银子、香料、贵重的膏油和他军械库里一切的兵器，以及他所有的财宝，都给他们看；在他家中和全国之内， 希西家 没有一样不给他们看的。
ISA|39|3|于是 以赛亚 先知到 希西家 王那里去，对他说：“这些人说了些什么？他们从哪里来见你？” 希西家 说：“他们从远方的 巴比伦 来见我。”
ISA|39|4|以赛亚 说：“他们在你家里看见了什么？” 希西家 说：“凡我家中所有的，他们都看见了；我财宝中没有一样东西不给他们看的。”
ISA|39|5|以赛亚 对 希西家 说：“你要听万军之耶和华的话，
ISA|39|6|耶和华说：‘看哪，日子将到，凡你家里所有的，并你祖先积蓄到如今的一切，都要被掳到 巴比伦 去，不留下一样；
ISA|39|7|从你本身所生的孩子，其中必有被掳到 巴比伦 王宫当太监的。’”
ISA|39|8|希西家 对 以赛亚 说：“你所说耶和华的话甚好。”因为他想：“在我有生之年必有太平和安稳。”
ISA|40|1|你们的上帝说： “要安慰，安慰我的百姓。
ISA|40|2|要对 耶路撒冷 说安慰的话， 向它宣告， 它的战争已结束， 它的罪孽已赦免； 它为自己一切的罪， 已从耶和华手中加倍受罚。”
ISA|40|3|有声音呼喊着： “要在旷野为耶和华预备道路， 在沙漠为我们的上帝修直大道。
ISA|40|4|一切山洼都要填满， 大小山冈都要削平； 陡峭的要变为平坦， 崎岖的必成为平原。
ISA|40|5|耶和华的荣耀必然显现， 凡有血肉之躯的都一同看见， 因为这是耶和华亲口说的。”
ISA|40|6|有声音说：“你喊叫吧！” 我 说：“我喊叫什么呢？” 凡有血肉之躯的尽都如草， 他的一切荣美像野地的花。
ISA|40|7|耶和华吹一口气， 草就枯干，花也凋谢。 百姓诚然是草；
ISA|40|8|草必枯干，花必凋谢， 惟有我们上帝的话永远立定。
ISA|40|9|报好信息的 锡安 哪， 要登高山； 报好信息的 耶路撒冷 啊， 要极力扬声。 扬声不要惧怕， 对 犹大 的城镇说： “看哪，你们的上帝！”
ISA|40|10|看哪，主耶和华必以大能临到， 他的膀臂必为他掌权； 看哪，他的赏赐在他那里， 他的报应在他面前。
ISA|40|11|他要像牧人牧养自己的羊群， 用膀臂聚集羔羊，抱在胸怀， 慢慢引导那乳养小羊的。
ISA|40|12|谁曾用手心量诸水， 用手虎口量苍天， 用升斗盛大地的尘土， 用秤称山岭， 用天平称冈陵呢？
ISA|40|13|谁曾测度耶和华的灵， 或作他的谋士指教他呢？
ISA|40|14|他与谁商议， 谁教导他， 以公平的路指示他， 将知识传授与他， 又将通达的道指教他呢？
ISA|40|15|看哪，列国都像水桶里的一滴， 又如天平上的微尘； 看哪，他举起众海岛，好像举起极微小之物。
ISA|40|16|黎巴嫩 不够当柴烧， 其中的走兽也不够作燔祭。
ISA|40|17|列国在他面前如同不存在， 在他看来微不足道，只是虚空。
ISA|40|18|你们究竟将谁比上帝， 用什么形像与他相较呢？
ISA|40|19|至于偶像，匠人铸造它， 银匠用金子包裹它， 又为它铸造银链。
ISA|40|20|没有能力捐献的人， 就挑选不易朽坏的木头， 为自己寻找巧匠， 竖立不会倒的偶像。
ISA|40|21|你们岂不知道吗？ 岂未曾听见吗？ 难道没有人从起头就告诉你们吗？ 自从地的根基立定， 你们岂不明白吗？
ISA|40|22|上帝坐在地的穹窿之上， 地上的居民有如蚱蜢。 他铺张穹苍如幔子， 展开诸天如可住的帐棚。
ISA|40|23|他使君王归于虚无， 使地上的审判官成为虚空。
ISA|40|24|他们刚栽上， 刚种好， 根也刚扎在地里， 经他一吹，就都枯干； 旋风将他们吹去，像碎秸一样。
ISA|40|25|那圣者说：“你们将谁与我相比， 与我相等呢？”
ISA|40|26|你们要向上举目， 看是谁创造这万象， 按数目领出它们， 一一称其名， 以他的权能 和他的大能大力， 使它们一个都不缺。
ISA|40|27|雅各 啊，你为何说， 以色列 啊，你为何言， “我的道路向耶和华隐藏， 我的冤屈上帝并不查问”？
ISA|40|28|你岂不曾知道吗？ 你岂未曾听见吗？ 永在的上帝耶和华，创造地极的主， 他不疲乏，也不困倦； 他的智慧无法测度。
ISA|40|29|疲乏的，他赐能力； 软弱的，他加力量。
ISA|40|30|就是年轻人也要疲乏困倦， 强壮的也必全然跌倒。
ISA|40|31|但那等候耶和华的必重新得力。 他们必如鹰展翅上腾； 他们奔跑却不困倦， 行走却不疲乏。
ISA|41|1|众海岛啊，在我面前静默； 万民要重新得力， 让他们近前来陈述， 我们可以彼此辩论。
ISA|41|2|谁从东方兴起一人， 凭公义召他来到脚前？ 谁将列国交给他， 使他管辖列王， 把他们如灰尘交与他的刀， 如风吹的碎秸交与他的弓？
ISA|41|3|他追赶君王， 安然走过， 快速地脚不落地 。
ISA|41|4|谁做成这事， 从起初宣召历代呢？ 就是我－耶和华！ 我是首先的， 也与末后的同在。
ISA|41|5|众海岛看见就都害怕， 地极也都战兢， 他们近前来；
ISA|41|6|各人互相帮助， 对弟兄说：“壮胆吧！”
ISA|41|7|木匠鼓励银匠， 用锤子打光的鼓励打砧的， 对焊工说：“焊得好！” 又用钉子钉稳，免得它倒下。
ISA|41|8|惟你 以色列 ，我的仆人， 雅各 ，我所拣选的， 我朋友 亚伯拉罕 的后裔，
ISA|41|9|你是我从地极领来， 从地角召来的， 我对你说：“你是我的仆人； 我拣选你，并不弃绝你。”
ISA|41|10|你不要害怕，因为我与你同在； 不要惊惶，因为我是你的上帝。 我必坚固你，帮助你， 用我公义的右手扶持你。
ISA|41|11|看哪，凡向你发怒的都抱愧蒙羞， 与你相争的必如无有，并要灭亡。
ISA|41|12|与你争斗的，你要寻找他们，却遍寻不着； 与你争战的必如无有，成为虚无。
ISA|41|13|因为我耶和华－你的上帝 必搀扶你的右手， 对你说：“不要害怕！ 我必帮助你。”
ISA|41|14|虫子 雅各 ， 以色列 人哪， 不要害怕！ 我必帮助你； 救赎你的是 以色列 的圣者。 这是耶和华说的。
ISA|41|15|看哪，我使你成为 全新的打谷机，齿轮锐利； 你要把山岭打得粉碎， 使冈陵如同糠秕。
ISA|41|16|你要簸扬它们，风要将它们吹去； 旋风要刮散它们。 你却要以耶和华为喜乐， 因 以色列 的圣者夸耀。
ISA|41|17|困苦贫穷人寻找水，却寻不着； 他们因口渴，舌头干燥。 我－耶和华必应允他们， 我─ 以色列 的上帝必不离弃他们。
ISA|41|18|我要在光秃的高地开江河， 在谷中开泉源； 我要使沙漠变为水池， 使干地变为涌泉。
ISA|41|19|我要在旷野栽植香柏树、 皂荚树、番石榴树，和野橄榄树。 在沙漠一同栽上松树、杉树， 和黄杨树，
ISA|41|20|好叫人看见，知道， 思想，明白； 这是耶和华亲手做的， 是 以色列 的圣者所造的。
ISA|41|21|耶和华说： “你们要呈上你们的案件。” 雅各 的君王说： “你们要提出你们的理由。”
ISA|41|22|让它们近前来，告诉我们将来要发生什么事！ 你们要说明先前发生的事，好让我们思索； 或者告诉我们将来的事，使我们得知事情的结局。
ISA|41|23|你们要指明未来的事， 使我们知道你们是神明！ 你们或降福，或降祸， 好使我们惊奇，一同观看。
ISA|41|24|看哪，你们属乎虚无， 你们的作为也属虚空； 那选择你们的是可憎恶的。
ISA|41|25|我从北方兴起一人， 他从日出之地而来， 是求告我名的； 他必踩踏 掌权者，如踩踏泥土， 又如陶匠踹泥一般。
ISA|41|26|有谁从起初宣布这事，使我们知道呢？ 有谁从先前指明，使我们说“他是对的”呢？ 没有人宣布， 没有人指明， 也没有人听见你们的话。
ISA|41|27|我首先对 锡安 说，看哪，他们在此！ 我要将一位报好信息的赐给 耶路撒冷 。
ISA|41|28|然而我观看，并无一人； 我询问的时候， 他们中间也没有谋士可回答。
ISA|41|29|看哪，他们尽是麻烦 ， 所做的工都属虚无； 所铸的偶像是风，是虚空。
ISA|42|1|看哪，我的仆人， 我所扶持、所拣选、心所喜悦的！ 我已将我的灵赐给他， 他必将公理传给万邦。
ISA|42|2|他不喧嚷，不扬声， 也不使街上听见他的声音。
ISA|42|3|压伤的芦苇，他不折断； 将残的灯火，他不吹灭。 他凭信实将公理传开。
ISA|42|4|他不灰心，也不丧胆， 直到他在地上设立公理； 众海岛都等候他的训诲。
ISA|42|5|那创造诸天，铺张穹苍， 铺开地与地的出产， 赐气息给地上众人， 赐生命给行走其上之人的 上帝耶和华如此说：
ISA|42|6|“我－耶和华凭公义召你， 要搀扶你的手，保护你， 要藉着你与百姓立约， 使你成为万邦之光，
ISA|42|7|开盲人的眼， 领囚犯出监狱， 领坐在黑暗中的出地牢。
ISA|42|8|我是耶和华，这是我的名； 我必不将我的荣耀归给别神 ， 也不将我所得的颂赞归给雕刻的偶像。
ISA|42|9|看哪，先前的事已经成就， 现在我要指明新事， 告诉你们尚未发生的事。
ISA|42|10|航海的人和海中一切所有的， 众海岛和其中的居民， 都当向耶和华唱新歌， 从地极赞美他。
ISA|42|11|旷野和其中的城镇， 并 基达 人居住的村庄都当扬声 ； 西拉 的居民当欢呼， 在山顶上大声呼喊。
ISA|42|12|愿他们将荣耀归给耶和华， 在海岛中传扬颂赞他的话。
ISA|42|13|耶和华必如勇士出征， 如战士激起愤恨， 他要喊叫，大声呐喊， 击败他的敌人。
ISA|42|14|我许久闭口不言，沉默不语； 现在我要像临产的妇人，大声喊叫， 呼吸急促而喘气。
ISA|42|15|我要使大小山冈变为荒芜， 使其上的花草都枯干； 我要使江河变为沙洲， 使水池尽都干涸。
ISA|42|16|我要引导盲人行他们所不认识的道， 引领他们走他们未曾走过的路； 我在他们面前使黑暗变为光明， 使弯曲变为平直。 这些事我都要做， 并不离弃他们。
ISA|42|17|但那倚靠雕刻的偶像， 对铸造的偶像说： “你是我们的神明”； 这种人要退后，大大蒙羞。
ISA|42|18|你们这耳聋的，听吧！ 你们这眼瞎的，看吧， 使你们得以看见！
ISA|42|19|谁比我的仆人眼瞎呢？ 谁比我所差遣的使者耳聋呢？ 谁瞎眼像那献身给我的人？ 谁瞎眼 像耶和华的仆人呢？
ISA|42|20|看见许多事却不领会， 耳朵开通却听不见。
ISA|42|21|耶和华因自己的公义， 乐意使律法为大为尊。
ISA|42|22|但这百姓是被抢被夺的， 全都陷在洞穴中，关在监牢里； 他们成了掠物，无人拯救， 成了掳物，无人索还。
ISA|42|23|你们中间谁肯侧耳听这话， 谁肯留心听，以防将来呢？
ISA|42|24|谁将 雅各 交出作为掳物， 将 以色列 交给抢夺者呢？ 岂不是耶和华 ─我们所得罪的那位吗？ 他们不肯遵行他的道， 也不听从他的训诲。
ISA|42|25|所以，他将猛烈的怒气和战争的威力 倾倒在 以色列 身上； 在他周围如火燃起，他竟然不知， 烧着了，他也不在意。
ISA|43|1|雅各 啊，创造你的耶和华， 以色列 啊，造成你的那位， 现在如此说： “你不要害怕，因为我救赎了你； 我曾提你的名召你，你是属我的。
ISA|43|2|你从水中经过，我必与你同在， 你渡过江河，水必不漫过你； 你在火中行走，也不被烧伤， 火焰必不烧着你身。
ISA|43|3|因为我是耶和华－你的上帝， 是 以色列 的圣者－你的救主； 我使 埃及 作你的赎价， 使 古实 和 西巴 代替你。
ISA|43|4|因我看你为宝贝为尊贵； 又因我爱你， 所以使人代替你， 使万民替换你的生命。
ISA|43|5|你不要害怕，因我与你同在； 我必领你的后裔从东方来， 又从西方召集你。
ISA|43|6|我要对北方说，交出来！ 对南方说，不可扣留！ 要将我的儿子从远方带来， 将我的女儿从地极领回，
ISA|43|7|就是凡称为我名下的人， 是我为自己的荣耀创造的， 是我所塑造，所做成的。”
ISA|43|8|你要将有眼却瞎、 有耳却聋的民都带出来！
ISA|43|9|任凭万国聚集， 任凭万民会合。 他们当中谁能说明， 并将先前的事指示我们呢？ 让他们带来见证，显明他们有理， 看是否听见的人会说：“果然是真的。”
ISA|43|10|你们是我的见证， 是我所拣选的仆人， 为了要使你们知道，且信服我， 又明白我就是耶和华。 在我以前没有任何被造的真神， 在我以后也必没有。 这是耶和华说的。
ISA|43|11|我，惟有我是耶和华； 除我以外没有救主。
ISA|43|12|我曾指示，我曾拯救，我曾说明， 并没有外族的神明 在你们中间。 你们是我的见证， 我是上帝。 这是耶和华说的。
ISA|43|13|自有日子以来，我就是上帝， 谁也不能救人脱离我的手。 我要行事，谁能逆转呢？
ISA|43|14|耶和华─你们的救赎主、 以色列 的圣者如此说： “因你们的缘故， 我已派遣人到 巴比伦 去； 要使 迦勒底 人都如难民， 坐自己素来宴乐的船下来。
ISA|43|15|我是耶和华－你们的圣者， 是创造 以色列 的，是你们的君王。”
ISA|43|16|那在沧海中开道， 在大水中开路， 使战车、马匹、军兵、勇士一同出来， 使他们仆倒，不再起来， 使他们灭没，好像熄灭之灯火的耶和华如此说：
ISA|43|17|
ISA|43|18|“你们不要追念从前的事， 也不要思想古时的事。
ISA|43|19|看哪，我要行一件新事， 如今就要显明，你们岂不知道吗？ 我必在旷野开道路， 在沙漠开江河 。
ISA|43|20|野地的走兽要尊敬我， 野狗和鸵鸟也必尊敬我。 因我使旷野有水， 使沙漠有河， 好赐给我的百姓、我的选民喝。
ISA|43|21|这百姓是我为自己造的， 为要述说我的美德。”
ISA|43|22|“ 雅各 啊，你并没有求告我； 以色列 啊，你倒厌烦我。
ISA|43|23|你并没有将你的羊带来献给我做燔祭， 也没有用牲祭尊敬我； 我未曾因素祭使你操劳， 也没有因乳香使你厌烦。
ISA|43|24|你没有用银子为我买香菖蒲， 也没有用祭物的油脂使我饱足； 倒使我因你的罪恶操劳， 使我因你的罪孽厌烦。
ISA|43|25|我，惟有我为自己的缘故涂去你的过犯， 我也不再记得你的罪恶。
ISA|43|26|你尽管提醒我，让我们来辩论； 尽管陈述，自显为义。
ISA|43|27|你的始祖犯罪， 你的师傅违背我；
ISA|43|28|因此，我要凌辱圣所的领袖 ， 使 雅各 遭毁灭， 使 以色列 受辱骂。”
ISA|44|1|“我的仆人 雅各 ， 我所拣选的 以色列 啊， 现在你当听。
ISA|44|2|那位造你，使你在母腹中成形， 并要帮助你的耶和华如此说： 我的仆人 雅各 ， 我所拣选的 耶书仑 哪， 不要害怕！
ISA|44|3|因为我要把水浇灌干渴的地方， 使水涌流在干旱之地。 我要将我的灵浇灌你的后裔， 使我的福临到你的子孙。
ISA|44|4|他们要在草丛中生长 ， 如溪水旁的柳树。
ISA|44|5|这个要说：‘我是属耶和华的’， 那个要以 雅各 的名自称， 又有一个在手上写着：‘归耶和华’， 并自称为 以色列 。”
ISA|44|6|耶和华－ 以色列 的君王， 以色列 的救赎主－万军之耶和华如此说： “我是首先的，也是末后的； 除我以外再没有上帝。
ISA|44|7|自从古时我设立了人， 谁能像我宣告，指明，又为自己陈说呢？ 让他指明未来的事和必成的事吧！
ISA|44|8|你们不要恐惧，也不要害怕。 我岂不是从上古就告诉并指示你们了吗？ 你们是我的见证人！ 除我以外，岂有上帝呢？ 诚然没有磐石，就我所知，一个也没有！”
ISA|44|9|制造偶像的人尽都虚空，他们所喜悦的全无益处；偶像的见证人毫无所见，毫无所知，以致他们羞愧。
ISA|44|10|谁制造神像，铸造偶像？这些都是无益的。
ISA|44|11|看哪，他的同伙都必羞愧。工匠不过是人，任他们聚集，任他们站立吧！他们都必惧怕，一同羞愧。
ISA|44|12|铁匠用工具在火炭上工作 ，用锤打出形状，用他有力的膀臂来锤。他因饥饿而无力气；因未喝水而疲倦。
ISA|44|13|木匠拉线，用笔划出样子，用刨子刨成形状，又用圆规划了模样。他仿照人的体态，做出美妙的人形，放在庙里。
ISA|44|14|他砍伐香柏树，又取杉树和橡树，在树林中让它茁壮；或栽种松树，得雨水滋润长大。
ISA|44|15|这树，人可用以生火；他拿一些来取暖，又搧火烤饼，而且做神像供跪拜，做雕刻的偶像向它叩拜。
ISA|44|16|他将一半的木头烧在火中，用它烤肉来吃；吃饱了，就自己取暖说：“啊哈，我暖和了，我看到火了！”
ISA|44|17|然后又用剩下的一半做了一个神明，就是雕刻的偶像，向这偶像俯伏叩拜，向它祷告说：“求你拯救我，因你是我的神明。”
ISA|44|18|他们既无知，又不思想；因为耶和华蒙蔽他们的眼，使他们看不见，塞住他们的心，使他们不明白。
ISA|44|19|没有一个心里醒悟，有知识，有聪明，能说：“我曾拿一部分用火燃烧，在炭火上烤饼，也烤肉来吃。这剩下的，我岂要做可憎之像吗？我岂可向木头叩拜呢？”
ISA|44|20|他以灰尘为食，心里迷糊，以致偏邪，不能自救，也不能说：“我右手中岂不是有虚谎吗？”
ISA|44|21|雅各 啊，要思念这些事； 以色列 啊，你是我的仆人。 我造了你，你是我的仆人， 以色列 啊，我必不忘记你 。
ISA|44|22|我涂去你的过犯，像厚云消散； 涂去你的罪恶，如薄雾消失。 你当归向我，因我救赎了你。
ISA|44|23|诸天哪，应当歌唱， 因为耶和华成就这事。 地的深处啊，应当欢呼； 众山哪，要出声歌唱； 树林和其中所有的树木啊，你们都当歌唱！ 因为耶和华救赎了 雅各 ， 并要因 以色列 荣耀自己。
ISA|44|24|从你在母腹中就造了你，你的救赎主－耶和华如此说： “我－耶和华创造万物， 独自铺张诸天，亲自展开大地 ；
ISA|44|25|我使虚谎的预兆失效， 愚弄占卜的人， 使智慧人退后， 使他的知识变为愚拙；
ISA|44|26|却使我仆人的话站得住， 成就我使者的筹算。 我论 耶路撒冷 说：‘必有人居住’； 论 犹大 的城镇说：‘必被建造， 我必重建其中的废墟。’
ISA|44|27|我对深渊说：‘干了吧！ 我要使你的江河干涸’；
ISA|44|28|论 居鲁士 说：‘他是我的牧人， 他要成就我所喜悦的， 下令建造 耶路撒冷 ， 发命令立稳圣殿的根基。’”
ISA|45|1|耶和华对所膏的 居鲁士 如此说， 他的右手我曾搀扶， 使列国降服在他面前， 列王的腰带我曾松开， 使城门在他面前敞开， 不得关闭：
ISA|45|2|“我要在你前面行， 修平崎岖之地。 我必打破铜门， 砍断铁闩。
ISA|45|3|我要将暗中的宝物和隐藏的财富赐给你， 使你知道提名召你的 就是我－耶和华， 以色列 的上帝。
ISA|45|4|因我的仆人 雅各 ， 我所拣选的 以色列 ， 我提名召你； 你虽不认识我， 我也加给你名号。
ISA|45|5|我是耶和华，再没有别的了； 除了我以外再没有上帝。 你虽不认识我， 我必给你束腰。
ISA|45|6|从日出之地到日落之处使人都知道 除我以外，没有别的。 我是耶和华，再没有别的了。
ISA|45|7|我造光，又造暗； 施平安，又降灾祸； 做成这一切的是我－耶和华。
ISA|45|8|“诸天哪，要如雨倾盆而降， 云要降下公义， 地要裂开，救恩涌出 ， 使公义也一同滋长； 这都是我－耶和华造的。”
ISA|45|9|“那与造他的主争论的人有祸了！ 他不过是地上瓦块中的一片 。 泥土岂可对塑造它的说：‘你做的是什么？ 你所做的物怎么没有把手呢？ ’
ISA|45|10|有人对父亲说， ‘你生的是什么’， 对母亲 说， ‘你生产的是什么’； 这人有祸了！”
ISA|45|11|耶和华－ 以色列 的圣者， 就是造 以色列 的如此说： “难道我孩子的未来，你们能质问我， 我手的工作，你们可以吩咐我吗？
ISA|45|12|我造大地，又创造人在地上。 我亲手铺张诸天， 天上万象也是我所任命的。
ISA|45|13|我凭公义兴起 居鲁士 ， 又要修直他一切的道路。 他必建造我的城， 释放我被掳的民， 不为工价，也不为奖赏。” 这是万军之耶和华说的。
ISA|45|14|耶和华如此说： “ 埃及 的出产和 古实 的货物必归你； 身量高大的 西巴 人，他们必过来归你，为你所有。 他们必带着锁链过来跟随你， 向你下拜，祈求你说： ‘上帝真是在你中间，再没有别的， 没有别的上帝。’”
ISA|45|15|救主－ 以色列 的上帝啊， 你诚然是隐藏自己的上帝。
ISA|45|16|制造偶像的都要抱愧蒙羞， 他们要一同归于惭愧。
ISA|45|17|惟有 以色列 必蒙耶和华拯救， 得永远的救恩。 你们必不蒙羞，也不抱愧， 直到永世无尽。
ISA|45|18|耶和华如此说， 他创造诸天，他是上帝； 他造了地，形成它，坚固它， 并非创造它为荒凉， 而是要给人居住： “我是耶和华，再没有别的。
ISA|45|19|我不在隐密黑暗之地说话， 也没有对 雅各 的后裔说， ‘你们寻求我是徒然的’， 我－耶和华所讲的是公义， 所说的是正直。”
ISA|45|20|“你们从列国逃脱的人， 要一同聚集前来。 那些抬着雕刻的木偶、 祈求不能救人之神明的， 毫无知识。
ISA|45|21|你们要近前来说明， 让他们彼此商议。 谁从古时指明这事？ 谁从上古述说它？ 不是我－耶和华吗？ 除了我以外，再没有上帝； 我是公义的上帝，又是救主； 除了我以外，再没有别的了。
ISA|45|22|“地的四极都当转向我， 就必得救； 因为我是上帝，再没有别的。
ISA|45|23|我指着自己起誓， 公义从我的口发出，这话并不返回： ‘万膝必向我跪拜， 万口必凭我起誓。’
ISA|45|24|人论我说 ， “公义、能力，惟独在乎耶和华。 人必归向他， 凡向他发怒的都必蒙羞。
ISA|45|25|以色列 的后裔必因耶和华得称为义， 并要彼此夸耀。”
ISA|46|1|彼勒 叩拜， 尼波 屈身； 巴比伦 的偶像驮在走兽和牲畜背上。 你们所抬的成了重驮， 使牲畜疲乏。
ISA|46|2|这些神明一同屈身叩拜， 不能救自己 ， 反倒遭人掳去。
ISA|46|3|雅各 家， 以色列 家所有的余民哪， 你们自从生下就蒙我抱， 自出母胎便由我来背， 你们都要听从我。
ISA|46|4|直到你们年老，我不改变； 直到你们发白，我仍扶持。 我已造你，就必背你； 我必抱你，也必拯救。
ISA|46|5|你们将谁与我相比，与我相等， 将谁与我相较，使我们相似呢？
ISA|46|6|他们从钱囊中倒出金子， 用天平秤出银子， 雇银匠造成神像， 他们又俯伏，又叩拜。
ISA|46|7|他们抬起神像，扛在肩上， 安置在定处，使它站立， 不离本位； 人呼求它，它却不回答， 也无法救人脱离灾难。
ISA|46|8|你们当记得这事，立定心意 。 叛逆的人哪，要留心思想。
ISA|46|9|要追念上古的事， 因为我是上帝，并无别的； 我是上帝，没有能与我相比的。
ISA|46|10|我从起初就指明末后的事， 从古时便言明未成的事， 说：“我的筹算必立定； 凡我所喜悦的，我必成就。”
ISA|46|11|我召鸷鸟从东方来， 召那成就我筹算的人从远方来。 我已说出，就必成就； 我已谋定，也必做成。
ISA|46|12|你们这些心中顽固、 远离公义的人，要听从我。
ISA|46|13|我使我的公义临近，它已不远。 我的救恩必不迟延。 我要为 以色列 －我的荣耀 在 锡安 施行救恩。
ISA|47|1|少女 巴比伦 哪， 下来坐在尘埃； 迦勒底 啊， 没有宝座，要坐在地上； 你不再称为柔弱娇嫩。
ISA|47|2|要用磨磨面， 揭去面纱， 脱去长裙， 露腿渡河。
ISA|47|3|你的下体必被露出； 你的羞辱必被看见。 我要报复， 谁也不宽容 。
ISA|47|4|我们的救赎主是 以色列 的圣者， 他的名为万军之耶和华。
ISA|47|5|迦勒底 啊， 你要静坐，进入黑暗中， 因你不再称为万国之后。
ISA|47|6|我向我的百姓发怒， 使我的产业受凌辱， 将他们交在你手中； 然而你毫不怜悯他们， 连老年人你也加极重的轭。
ISA|47|7|你说：“我必永远为后。” 你不将这事放在心上， 也不思想事情的结局。
ISA|47|8|你这专好宴乐、以为地位稳固的， 现在当听这话。 你心中说： “惟有我，除我以外再没有别的。 我必不致寡居， 也不经历丧子之痛。”
ISA|47|9|哪知，丧子、寡居这两件事 一日之间忽然临到你； 你虽多行邪术、广施魔咒， 这两件事必全然临到你身上。
ISA|47|10|你倚靠自己的恶行，说： “无人看见我。” 你的智慧聪明使你走偏， 你心里说： “惟有我，除我以外再没有别的了。”
ISA|47|11|但灾祸临到你， 你不知如何驱除； 灾害落在你身上， 你也无法除掉， 你所不知道的毁灭必忽然临到你身上。
ISA|47|12|尽管使用从幼年就施行的魔符和众多的邪术吧！ 或许有些帮助， 或许可以致胜。
ISA|47|13|你筹划太多，以致疲倦。 让那些观天象，看星宿， 在初一说预言的都起来， 救你脱离所要临到你的事！
ISA|47|14|看哪，他们要像碎秸被火焚烧， 无法救自己脱离火焰的魔掌； 没有炭火可以取暖 ， 你也不能坐在火旁。
ISA|47|15|你所操劳的事都像这样； 从你幼年以来与你交易的都各奔己路， 没有一人来救你。
ISA|48|1|雅各 家，称为 以色列 名下， 从 犹大 的源头而出的啊， 你们指着耶和华的名起誓， 提说 以色列 的上帝， 却不凭诚信，也不凭公义； 你们自称为圣城之民， 倚靠名为万军之耶和华－ 以色列 的上帝； 现在，当听我言：
ISA|48|2|
ISA|48|3|“先前的事，我自古已说明， 已从我口而出， 是我所指示的； 我瞬间行事，事便成就。
ISA|48|4|因为我知道你是顽梗的； 你的颈项是铁的， 你的额头是铜的。
ISA|48|5|所以，我自古就给你说明， 在事未成以先指示你， 免得你说：‘这些事是我的偶像所行的， 是我雕刻的偶像和铸造的神像所命定的。’
ISA|48|6|“你既已听见，现在要察看这一切； 你们不是要说明吗？ 从今以后，我要指示你新事， 就是你所不知道的隐密事。
ISA|48|7|这事是现今造的，并非自古就有， 在今日以先，你未曾听见； 免得你说：‘看哪，这事我早已知道了。’
ISA|48|8|诚然你未曾听见，也未曾知道； 你的耳朵从来未曾开通。 我原知道你行事极其诡诈， 你自从出母胎以来， 就称为悖逆的。
ISA|48|9|“我为我的名暂且忍怒， 为了我的荣耀向你容忍， 不将你剪除。
ISA|48|10|看哪，我熬炼你，却不像熬炼银子； 你在苦难的火炉中，我试炼 你。
ISA|48|11|我为自己的缘故必做这事， 我岂能被亵渎？ 我必不将我的荣耀归给别神 。
ISA|48|12|雅各 －我所选召的 以色列 啊， 当听从我： 我是耶和华， “我是首先的，也是末后的。
ISA|48|13|我亲手立了地的根基， 以右手铺张诸天； 我一召唤，天地就都立定。
ISA|48|14|你们都当聚集而听， 偶像 之中谁曾说明这些事？ 耶和华爱他，他必向 巴比伦 成就耶和华的旨意， 耶和华的膀臂也要加在 迦勒底 人身上 。
ISA|48|15|我，惟有我曾说过， 我选召他，领他来， 他的道路必亨通。
ISA|48|16|你们要接近我来听这话， 我从起初就未曾在隐密之处说话， 万事之始，我就在那里。” 现在，主耶和华差遣了我， 带着他的灵而来 。
ISA|48|17|耶和华－你的救赎主， 以色列 的圣者如此说： “我是耶和华－你的上帝， 我教导你，使你得益处， 指引你当走的路。
ISA|48|18|甚愿你听从我的命令， 你的平安就会如河水， 你的公义如海浪，
ISA|48|19|你的后裔必多如海沙， 你腹中所生的必多如沙粒。 他的名绝不从我面前剪除， 也不灭绝。”
ISA|48|20|你们要从 巴比伦 出来， 从 迦勒底 人中逃脱， 以欢呼的声音宣告， 将这事传扬到地极，说： 耶和华救赎了他的仆人 雅各 ！
ISA|48|21|他引导他们经过沙漠， 他们却未尝干渴； 他为他们使水从磐石流出， 磐石裂开，水就涌出。
ISA|48|22|耶和华说： “恶人必不得平安！”
ISA|49|1|众海岛啊，当听从我！ 远方的众民哪，要留心听！ 自出母胎，耶和华就选召我； 自出母腹，他就称呼我的名。
ISA|49|2|他使我的口如快刀， 把我藏在他手荫之下； 又使我成为磨利的箭， 把我藏在他箭袋之中；
ISA|49|3|对我说：“你是我的仆人 以色列 ； 我必因你得荣耀。”
ISA|49|4|我却说：“我劳碌是徒然， 我尽力是虚无虚空。 耶和华诚然以公平待我， 我的赏赐在我的上帝那里。”
ISA|49|5|现在耶和华说话，他从我出母胎，就造我作他的仆人， 要使 雅各 归向他， 使 以色列 聚集在他那里。 耶和华看我为尊贵， 我的上帝是我的力量。
ISA|49|6|他说：“你作我的仆人， 使 雅各 众支派复兴， 使 以色列 中蒙保存的人归回； 然而此事尚小， 我还要使你作万邦之光， 使你施行我的救恩，直到地极。”
ISA|49|7|救赎主－ 以色列 的圣者耶和华 对那被人藐视、本国憎恶、 统治者奴役的如此说： “君王看见就站起来， 领袖也要下拜； 这都是因信实的耶和华， 因拣选你的 以色列 的圣者。”
ISA|49|8|耶和华如此说： “在悦纳的时候，我应允了你； 在拯救的日子，我帮助了你。 我要保护你， 要藉着你与百姓立约， 为了复兴遍地， 使人承受荒芜之地为业；
ISA|49|9|对那被捆绑的人说：‘出来吧！’ 对在黑暗里的人说：‘显现吧！’ 他们在路上必得饮食， 在光秃的高地必有食物。
ISA|49|10|他们不饥不渴， 炎热和烈日必不伤害他们； 因为怜悯他们的必引导他们， 领他们到水泉旁边。
ISA|49|11|我必在众山开辟路径， 大道也要填高。
ISA|49|12|看哪，他们从远方来； 有些从北方来，有些从西方来， 有些从 色弗尼 地来。”
ISA|49|13|诸天哪，应当欢呼！ 大地啊，应当快乐！ 众山哪，应当扬声歌唱！ 因为耶和华已经安慰他的百姓， 他要怜悯他的困苦之民。
ISA|49|14|锡安 说：“耶和华离弃了我， 主忘记了我。”
ISA|49|15|妇人焉能忘记她吃奶的婴孩， 不怜悯她所生的儿子？ 即或有忘记的， 我却不忘记你。
ISA|49|16|看哪，我将你铭刻在我掌上， 你的城墙常在我眼前。
ISA|49|17|建立你的胜过毁坏你的， 使你荒废的必都离你而去。
ISA|49|18|你举目向四围观看， 他们都聚集来到你这里。 我指着我的永生起誓， 你定要以他们为妆饰佩戴， 带着他们，像新娘一样。 这是耶和华说的。
ISA|49|19|至于你荒废凄凉之处， 并你被毁坏之地， 如今居民必嫌太窄， 吞灭你的必离你遥远。
ISA|49|20|你要再听见丧失子女后所生的儿女说： “这地方我居住太窄， 请你给我地方居住。”
ISA|49|21|那时你心里必说：“我既丧子不育， 被掳，飘流在外 ， 谁给我生了这些？ 谁将他们养大呢？ 看哪，我被撇下独自一人时， 他们都在哪里呢？”
ISA|49|22|主耶和华如此说： “看哪，我必向列国举手， 向万民竖立大旗； 他们必将你的儿子抱在怀中带来， 将你的女儿背在肩上扛来。
ISA|49|23|列王必作你的养父， 王后必作你的乳母。 他们必以脸伏地，向你下拜， 并舔你脚上的尘土。 你就知道我是耶和华， 等候我的必不致羞愧。”
ISA|49|24|勇士抢去的岂能夺回？ 被残暴者掳掠的岂能得解救呢？
ISA|49|25|但耶和华如此说： “就是勇士所掳掠的，也可以夺回； 残暴者所抢的，也可以得解救。 与你相争的，我必与他相争， 我也要拯救你的儿女。
ISA|49|26|我必使那欺压你的吃自己的肉， 饮自己的血，如喝甜酒喝醉一样。 凡有血肉之躯的都必知道我－耶和华是你的救主， 是你的救赎主，是 雅各 的大能者。”
ISA|50|1|耶和华如此说： “我休了你们的母亲， 她的休书在哪里呢？ 我将你们卖给了我哪一个债主呢？ 看哪，你们被卖是因你们的罪孽； 你们的母亲被休，是因你们的过犯。
ISA|50|2|我来的时候，为何没有人呢？ 我呼唤的时候，为何无人回应呢？ 我的膀臂岂是过短、不能救赎吗？ 我岂无拯救之力吗？ 看哪，我一斥责，海就干了； 我使江河变为旷野， 其中的鱼因无水腥臭，干渴而死。
ISA|50|3|我使诸天以黑暗为衣， 以麻布为遮盖。”
ISA|50|4|主耶和华赐我受教者的舌头， 使我知道怎样用言语扶助疲乏的人。 主每天早晨唤醒，唤醒我的耳朵， 使我能听，像受教者一样。
ISA|50|5|主耶和华开启我的耳朵， 我并未违背，也未退后。
ISA|50|6|人打我的背，我任他打； 人拔我两颊的胡须，我由他拔； 人侮辱我，向我吐唾沫，我并不掩面。
ISA|50|7|主耶和华必帮助我， 所以我不抱愧。 我硬着脸面好像坚石， 也知道我必不致蒙羞。
ISA|50|8|称我为义的与我相近； 谁与我争论， 让我们来对质； 谁与我作对， 让他近前来吧！
ISA|50|9|看哪，主耶和华必帮助我， 谁能定我有罪呢？ 看哪，他们都要像衣服渐渐破旧， 被蛀虫蛀光。
ISA|50|10|你们当中有谁是敬畏耶和华， 听从他仆人的话语， 却行在黑暗中，没有亮光的， 当倚靠耶和华的名， 仰赖自己的上帝。
ISA|50|11|看哪，你们当中所有点火、以火把围绕自己的人， 当行走在你们的火焰 里， 并你们所点的火把中。 这是我亲手为你们定的： 你们必躺卧在悲惨之中。
ISA|51|1|追求公义、 寻求耶和华的人哪， 当听从我！ 你们要追想自己是从哪块磐石凿出， 从哪个岩穴挖掘而来；
ISA|51|2|要追想你们的祖宗 亚伯拉罕 和生你们的 撒拉 ； 因为我选召 亚伯拉罕 时，他只有一个人， 但我赐福给他， 使他增多。
ISA|51|3|耶和华已经安慰 锡安 ， 安慰了 锡安 一切的废墟， 使旷野如 伊甸 ， 使沙漠像耶和华的园子； 其中必有欢喜、快乐、感谢， 和歌唱的声音。
ISA|51|4|我的民哪，要留心听我， 我的国啊，要向我侧耳； 因为训诲必从我而出， 我必使我的公理成为万民之光。
ISA|51|5|我的公义临近， 我的救恩发出。 我的膀臂要审判万民， 众海岛都要等候我，倚赖我的膀臂。
ISA|51|6|你们要向天举目， 观看下面的地； 天必像烟云消散， 地必如衣服渐渐破旧； 其上的居民也要如此 死亡。 惟有我的救恩永远长存， 我的公义也不废掉。
ISA|51|7|知道公义、将我的训诲存在心中的人哪， 当听从我！ 不要怕人的辱骂， 也不要因人的毁谤惊惶。
ISA|51|8|因为他们必像衣服被蛀虫蛀； 像羊毛被虫子咬。 惟有我的公义永远长存， 我的救恩直到万代。
ISA|51|9|耶和华的膀臂啊，兴起，兴起！ 以能力为衣穿上， 像古时的年日，像上古的世代一样兴起！ 从前砍碎 拉哈伯 、 刺透大鱼的，不是你吗？
ISA|51|10|使海与深渊的水干涸， 在海的深处开路， 使救赎的民走过的，不是你吗？
ISA|51|11|耶和华救赎的民必归回， 歌唱来到 锡安 ； 永恒的喜乐必归到他们头上。 他们必得着欢喜快乐， 忧伤叹息尽都逃避。
ISA|51|12|我，惟有我是安慰你们的。 你是谁，竟怕那必死的人， 怕那生命如草的世人，
ISA|51|13|却忘记铺张诸天、立定地基、 造你的耶和华？ 你因欺压者图谋毁灭所发的暴怒， 终日害怕， 其实那欺压者的暴怒在哪里呢？
ISA|51|14|被掳的即将得释放， 不至于死而下入地府， 也不致缺乏食物。
ISA|51|15|我是耶和华－你的上帝， 我搅动大海，使海中的波浪澎湃， 万军之耶和华是我的名。
ISA|51|16|我已将我的话放在你口中， 用我的手影遮蔽你， 为要安定诸天，立定地基， 并对 锡安 说：“你是我的百姓。”
ISA|51|17|耶路撒冷 啊，兴起，兴起！ 站起来！ 你从耶和华手中喝了他愤怒的杯， 那使人东倒西歪的杯，直到喝尽。
ISA|51|18|她所生育的孩子中，没有一个搀她的； 她所抚养的孩子中，没有一个扶她的。
ISA|51|19|这双重的灾难临到你， 有谁怜悯你呢？ 破坏和毁灭，饥荒和战争临到， 我如何能安慰你呢 ？
ISA|51|20|你的孩子发昏， 在各街头躺卧， 如同网罗里的羚羊， 满了耶和华的愤怒， 满了你上帝的斥责。
ISA|51|21|因此，你这困苦却非因酒而醉的， 当听这话，
ISA|51|22|你的主，耶和华， 就是为他百姓辩护的上帝如此说： “看哪，我已从你手中接过 那使人东倒西歪的杯， 就是我愤怒的杯， 你必不再喝。
ISA|51|23|我必将这杯递在苦待你的人 手中。 他们曾对你说：‘你屈身， 任我们践踏过去吧！’ 你就以背为地， 又如街道，任人走过。
ISA|52|1|锡安 哪，兴起！兴起！ 穿上你的能力！ 圣城 耶路撒冷 啊，穿上你华美的衣服！ 因为从今以后， 未受割礼、不洁净的必不再进入你中间。
ISA|52|2|耶路撒冷 啊，抖去尘埃， 起来坐在王位上！ 被掳的 锡安 哪， 解开你颈上的锁链！
ISA|52|3|耶和华如此说：“你们白白地被卖，也必不用银子赎回。”
ISA|52|4|主耶和华如此说：“先前我的百姓下到 埃及 ，在那里寄居，末后又有 亚述 人欺压他们。”
ISA|52|5|我的百姓既是白白地被掳，如今我在这里做什么呢？这是耶和华说的。辖制他们的人欢呼 ，我的名终日不断受亵渎，这是耶和华说的。
ISA|52|6|因此，我的百姓必认识我的名；在那日，他们必知道说这话的就是我。看哪，是我！”
ISA|52|7|在山上报佳音，传平安， 报好信息，传扬救恩， 那人的脚踪何等佳美啊！ 他对 锡安 说：“你的上帝作王了！”
ISA|52|8|听啊，你守望之人的声音， 他们扬声一同欢唱； 因为他们必亲眼看见耶和华返回 锡安 。
ISA|52|9|耶路撒冷 的废墟啊， 要出声一同欢唱； 因为耶和华安慰了他的百姓， 救赎了 耶路撒冷 。
ISA|52|10|耶和华在万国眼前露出圣臂， 地的四极都要看见我们上帝的救恩。
ISA|52|11|离开吧！离开吧！ 你们要从 巴比伦 出来。 你们扛抬耶和华器皿的人哪， 不要沾不洁净的东西， 离去时务要保持洁净。
ISA|52|12|你们出来必不致匆忙， 也不致奔逃； 因为耶和华要在你们前头行， 以色列 的上帝必作你们的后盾。
ISA|52|13|看哪，我的仆人行事必有智慧， 他必被高升，高举， 升到至高之处。
ISA|52|14|许多人因他 惊奇 ─他的面貌比别人憔悴， 他的外表比世人枯槁─
ISA|52|15|同样，他也必使许多国家惊奇 ， 君王要向他闭口。 未曾传给他们的，他们必看见； 未曾听见过的事，他们要明白。
ISA|53|1|我们所传的有谁信呢？ 耶和华的膀臂向谁显露呢？
ISA|53|2|他在耶和华面前生长如嫩芽， 像根出于干地。 他无佳形美容使我们注视他， 也无美貌使我们仰慕他。
ISA|53|3|他被藐视，被人厌弃； 多受痛苦，常经忧患。 他被藐视， 好像被人掩面不看的一样， 我们也不尊重他。
ISA|53|4|他诚然担当我们的忧患， 背负我们的痛苦； 我们却以为他受责罚， 是被上帝击打苦待。
ISA|53|5|他为我们的过犯受害， 为我们的罪孽被压伤。 因他受的惩罚，我们得平安； 因他受的鞭伤，我们得医治。
ISA|53|6|我们都如羊走迷， 各人偏行己路； 耶和华使我们众人的罪孽都归在他身上。
ISA|53|7|他被欺压受苦， 却不开口； 他像羔羊被牵去宰杀， 又像羊在剪毛的人手下无声， 他也是这样不开口。
ISA|53|8|因受欺压和审判，他被夺去， 谁能想到他的世代呢？ 因为他从活人之地被剪除， 为我百姓 的罪过他被带到死里 。
ISA|53|9|他虽然未行残暴， 口中也没有诡诈， 人还使他与恶人同穴， 与财主同墓 。
ISA|53|10|耶和华的旨意要压伤他， 使他受苦。 当他的生命作为赎罪祭时 ， 他必看见后裔，他的年日必然长久。 耶和华所喜悦的事，必在他手中亨通。
ISA|53|11|因自己的劳苦，他必看见光 就心满意足。 因自己的认识，我的义仆使许多人得称为义， 他要担当他们的罪孽。
ISA|53|12|因此，我要使他与位大的同份， 与强盛的均分掳物。 因为他倾倒自己的生命，以致于死， 也列在罪犯之中。 他却担当多人的罪， 为他们的过犯代求 。
ISA|54|1|你这不怀孕、不生育的，要欢呼； 你这未曾经过产难的，要欢呼，扬声呼喊； 因为被遗弃的妇人， 比有丈夫的人儿女更多； 这是耶和华说的。
ISA|54|2|要扩张你帐幕之地， 伸展你居所的幔子，不要缩回； 要放长你的绳子， 坚固你的橛子。
ISA|54|3|因为你要向左向右开展， 你的后裔必得列国为业， 又使荒废的城镇有人居住。
ISA|54|4|不要惧怕，因你必不致蒙羞； 不要抱愧，因你必不致受辱。 你必忘记年轻时的羞愧， 不再记得守寡的耻辱。
ISA|54|5|因为造你的是你的丈夫， 万军之耶和华是他的名； 救赎你的是 以色列 的圣者， 他必称为全地之上帝。
ISA|54|6|耶和华召你， 如同召回心中忧伤遭遗弃的妇人， 就是年轻时所娶被遗弃的妻子； 这是你的上帝说的。
ISA|54|7|我离弃你不过片时， 却要大施怜悯将你寻回。
ISA|54|8|我因涨溢的怒气， 一时向你转脸， 但我要以永远的慈爱怜悯你； 这是耶和华－你的救赎主说的。
ISA|54|9|这事于我有如 挪亚 的洪水； 我怎样起誓不再使 挪亚 的洪水淹没全地， 也照样起誓不再向你发怒， 且不斥责你。
ISA|54|10|大山可以挪开， 小山可以迁移， 但我的慈爱必不离开你， 我平安的约也不迁移； 这是怜悯你的耶和华说的。
ISA|54|11|你这受困苦、被暴风卷走、不得怜悯的城， 看哪，我必以灰泥来做你的石头， 以蓝宝石立你的根基，
ISA|54|12|又以红宝石造你的女墙， 以晶莹的珠玉造你的城门， 以珍贵的宝石造你四围的边界。
ISA|54|13|你的儿女都要领受耶和华的教导， 你的儿女必大享平安。
ISA|54|14|你必因公义得坚立， 必远离欺压，毫不惧怕； 你必远离惊吓，惊吓必不临近你。
ISA|54|15|若有人攻击你，这非出于我； 凡攻击你的，必因你仆倒。
ISA|54|16|看哪，我造了那吹炭火、打造合用兵器的铁匠； 我也造了那残害人、行毁灭的人。
ISA|54|17|凡为攻击你而造的兵器必无效用； 在审判时兴起用口舌攻击你的， 你必驳倒他。 这是耶和华仆人的产业， 是他们从我所得的义； 这是耶和华说的。
ISA|55|1|来！你们所有干渴的，都当来到水边； 没有银钱的也可以来。 你们都来，买了吃； 不用银钱，不付代价， 就可买酒和奶。
ISA|55|2|你们为何花钱买那不是食物的东西， 用劳碌得来的买那无法使人饱足的呢？ 你们要留意听从我的话，就能吃那美物， 得享肥甘，心中喜乐。
ISA|55|3|当侧耳而听，来到我这里； 要听，就必存活。 我要与你们立永约， 就是应许给 大卫 那可靠的慈爱。
ISA|55|4|看哪，我已立他作万民的见证， 立他作万民的君王和发令者。
ISA|55|5|看哪，你要召集素不认识的国民， 素不认识的国民要奔向你； 这都因耶和华─你的上帝， 因 以色列 的圣者已经荣耀了你。
ISA|55|6|当趁耶和华可寻找的时候寻找他， 在他接近的时候求告他。
ISA|55|7|恶人当离弃自己的道路， 不义的人应除掉自己的意念。 归向耶和华，耶和华就必怜悯他； 当归向我们的上帝，因为他必广行赦免。
ISA|55|8|我的意念非同你们的意念， 我的道路非同你们的道路。 这是耶和华说的。
ISA|55|9|天怎样高过地， 照样，我的道路高过你们的道路， 我的意念高过你们的意念。
ISA|55|10|雨雪从天而降，并不返回， 却要滋润土地，使地面发芽结实， 使撒种的有种，使要吃的有粮。
ISA|55|11|我口所出的话也必如此， 绝不徒然返回， 却要成就我的旨意， 达成我差它的目的。
ISA|55|12|你们必欢欢喜喜出来， 平平安安蒙引导。 大山小山必在你们面前欢呼， 田野的树木也都拍掌。
ISA|55|13|松树长出，代替荆棘； 番石榴长出，代替蒺藜。 这要为耶和华留名， 作为永不磨灭的证据。
ISA|56|1|耶和华如此说： “你们当守公平，行公义； 因我的救恩临近， 我的公义将要显现。
ISA|56|2|谨守安息日不予干犯， 禁止己手不作恶， 如此行、如此持守的人有福了！”
ISA|56|3|与耶和华联合的外邦人不要说： “耶和华将我和他的子民分别出来。” 太监也不要说：“看哪，我是枯树。”
ISA|56|4|因为耶和华如此说： “那些谨守我的安息日， 选择我旨意， 持守我约的太监，
ISA|56|5|我必使他们在我殿中，在我墙内， 有纪念碑，有名号， 胜过有儿有女； 我必赐他们永远的名，不能剪除。
ISA|56|6|“那些与耶和华联合， 事奉他，爱他名， 作他仆人的外邦人， 凡谨守安息日不予干犯， 又持守我约的人，
ISA|56|7|我必领他们到我的圣山， 使他们在我的祷告的殿中喜乐。 他们的燔祭和祭物， 在我坛上必蒙悦纳， 因我的殿必称为万民祷告的殿。
ISA|56|8|我还要召集更多的人 归并到这些被召集的人中。 这是召集被赶散的 以色列 人的 主耶和华说的。”
ISA|56|9|野地的走兽，你们都来吞吃吧！ 林中的野兽，你们也来吞吃！
ISA|56|10|以色列 的守望者都瞎了眼， 没有知识； 都是哑狗，不会吠叫， 只知做梦，躺卧，贪睡，
ISA|56|11|这些狗贪食，不知饱足。 这些牧人不知明辨， 他们都偏行己路， 人人追求自己的利益。
ISA|56|12|他们说：“来吧！我去拿酒， 让我们畅饮烈酒吧！ 明天必和今天一样， 甚至更好！”
ISA|57|1|义人死亡， 无人放在心上； 虔诚的人被接去， 无人理解； 义人被接去，以免祸患。
ISA|57|2|行为正直的人进入平安， 得以在床上安歇 。
ISA|57|3|到这里来吧！ 你们这些巫婆的儿子， 奸夫和妓女的后代；
ISA|57|4|你们向谁戏笑？ 向谁张口吐舌呢？ 你们岂不是叛逆所生的儿女， 虚谎所生的后代吗？
ISA|57|5|你们在橡树 中间，在各青翠的树下欲火攻心； 在山谷间，在岩隙下杀了儿女；
ISA|57|6|去拜谷中光滑的石头有你们的份， 这些就是你们的命运。 你向它们献浇酒祭，献供物， 这事我岂能容忍吗？
ISA|57|7|你在高而又高的山上安设床铺， 上那里去献祭。
ISA|57|8|你在门后，在门框后， 立起你的牌来； 你离弃了我，赤露己身， 又爬上自己所铺宽阔的床铺， 与它们立约； 你喜爱它们的床，看着它们的赤体 。
ISA|57|9|你带了油到 摩洛 那里， 加上许多香水。 你派遣使者往远方去， 甚至降到阴间，
ISA|57|10|因路途遥远，你就疲倦， 却不说，这是枉然， 以为能找到复兴之力， 所以不觉疲惫。
ISA|57|11|你怕谁，因谁恐惧， 竟说谎，不记得我， 不将这事放在心上。 是否因我许久闭口不言， 你就不怕我了呢？
ISA|57|12|我可以宣告你的公义和你的作为， 但它们与你无益。
ISA|57|13|你哀求的时候， 让你所搜集的神像 拯救你吧！ 风要把它们全都刮散， 吹一口气就都吹走。 但那投靠我的必得地产， 承受我的圣山为业。
ISA|57|14|耶和华说： “你们要修筑，修筑，要预备道路， 除掉我百姓路中的绊脚石。”
ISA|57|15|那至高无上、永远长存、 名为圣者的如此说： “我住在至高至圣的所在， 却与心灵痛悔的谦卑人同住； 要使谦卑的人心灵苏醒， 使痛悔的人内心复苏。
ISA|57|16|我必不长久控诉，也不永远怀怒， 因为我虽使灵性发昏，我也造了人的气息。
ISA|57|17|我因人贪婪的罪孽，发怒击打他； 我转脸向他发怒， 他却仍随意背道而行。
ISA|57|18|我看见他的行为， 要医治他，引导他 ， 使他和与他一同哀伤的人都得安慰。
ISA|57|19|我要医治他， 他要结出嘴唇的果实。 平安，平安，归给远处和近处的人！ 这是耶和华说的。”
ISA|57|20|但是恶人好像翻腾的海， 不得平静； 其中的水常涌出污秽和淤泥。
ISA|57|21|我的上帝说：“恶人必不得平安！”
ISA|58|1|你要大声喊叫，不要停止； 要扬声，好像吹角； 向我的百姓宣告他们的过犯， 向 雅各 家陈述他们的罪恶。
ISA|58|2|他们天天寻求我， 乐意明白我的道， 好像行义的国家， 未离弃它的上帝的典章； 他们向我求问公义的判词， 喜悦亲近上帝。
ISA|58|3|“我们禁食，你为何不看呢？ 我们刻苦己心，你为何不理会呢？” 看哪，你们禁食的时候仍追求私利， 剥削为你们做苦工的人。
ISA|58|4|看哪，你们禁食，却起纷争兴讼， 以凶恶的拳头打人。 你们今日这种禁食 无法使你们的声音听闻于高处。
ISA|58|5|这岂是我所要的禁食， 为人所用以刻苦己心的日子吗？ 我难道只是叫人如芦苇般低头， 铺上麻布和灰烬吗？ 你能称此为禁食， 为耶和华所悦纳的日子吗？
ISA|58|6|我所要的禁食，岂不是要你松开凶恶的绳， 解开轭上的索， 使被欺压的得自由， 折断一切的轭吗？
ISA|58|7|岂不是要你把食物分给饥饿的人， 将流浪的穷人接到家中， 见赤身的给他衣服遮体， 而不隐藏自己避开你的骨肉吗？
ISA|58|8|这样，必有光如晨光破晓照耀你， 你也要快快得到医治； 你的公义在你前面行， 耶和华的荣光必作你的后盾。
ISA|58|9|那时你求告，耶和华必应允； 你呼求，他必说：“我在这里。” 你若从你中间除掉重轭 和指摘人的指头，并发恶言的事，
ISA|58|10|向饥饿的人施怜悯， 使困苦的人得满足； 你在黑暗中就必得着光明， 你的幽暗必变如正午。
ISA|58|11|耶和华必时常引导你， 在干旱之地使你心满意足， 又使你骨头强壮。 你必如有水浇灌的园子， 又像水流不绝的泉源。
ISA|58|12|你们中间必有人起来修造久已荒废之处， 立起代代相承的根基。 你必称为修补裂痕的， 和重修路径给人居住的。
ISA|58|13|你若禁止自己的脚践踏安息日， 不在我的圣日做自己高兴的事， 称安息日为“可喜乐的”， 称耶和华的圣日为“可尊重的”， 尊敬这日， 不走自己的道路， 不求自己的喜悦， 也不随意说话；
ISA|58|14|那么，你就会以耶和华为乐。 耶和华要使你乘驾于地的高处， 又要以你祖先 雅各 的产业养育你； 这是耶和华亲口说的。
ISA|59|1|看哪，耶和华的膀臂并非过短，不能拯救， 耳朵并非发沉，不能听见，
ISA|59|2|但你们的罪孽使你们与上帝隔绝， 你们的罪恶使他转脸不听你们。
ISA|59|3|因你们的手掌被血沾染， 你们的指头被罪玷污， 你们的嘴唇说谎言， 你们的舌头出恶语。
ISA|59|4|无人按公义控诉， 也无人凭诚实辩白； 却倚靠虚妄，口说谎言， 怀毒害，生罪孽。
ISA|59|5|他们孵毒蛇蛋， 结蜘蛛网。 凡吃这蛋的必死， 蛋一打破，就孵出蛇来。
ISA|59|6|所结的网不能当衣服， 无法掩盖自己所作所为。 他们的行为全是邪恶， 手所做的尽都残暴。
ISA|59|7|他们的脚奔跑行恶， 急速流无辜者的血； 他们的思想全是恶念， 走过的路尽是破坏与毁灭。
ISA|59|8|平安的路，他们不知道， 所行的事无一公平。 他们为自己修筑弯曲的路， 凡走这路的都不得平安。
ISA|59|9|因此，公平离我们甚远， 公义追不上我们。 我们指望光亮，看哪，却只有黑暗， 指望光明，却行在幽暗中。
ISA|59|10|我们用手摸墙，好像盲人， 四处摸索，如同失明的人； 中午时我们绊倒，如在黄昏一样， 在强壮的人中，我们好像死人一般。
ISA|59|11|我们全都咆哮如熊， 哀鸣如鸽子； 指望公平，却得不着； 指望救恩，它却远离。
ISA|59|12|我们的过犯在你面前增加， 罪恶作证控告我们； 过犯与我们同在。 至于我们的罪孽，我们都知道：
ISA|59|13|就是悖逆，否认耶和华， 转去不跟从我们的上帝， 口说欺压和叛逆的话， 心怀谎言，随即说出；
ISA|59|14|公平转而退后， 公义站在远处， 诚实仆倒在广场上， 正直不得进入；
ISA|59|15|诚实少见， 离弃邪恶的人反成掠物。 那时，耶和华见没有公平， 就不喜悦。
ISA|59|16|他见无人， 竟无一人代求，甚为诧异， 就用自己的膀臂拯救他， 以公义扶持他。
ISA|59|17|他穿上公义为铠甲， 戴上救恩为头盔， 穿上报复为衣服， 披戴热心为外袍。
ISA|59|18|他必按人的行为报应， 恼怒他的敌人， 报复他的仇敌， 向众海岛施行报应。
ISA|59|19|在日落之处，人必敬畏耶和华的名； 在日出之地，人必敬畏他的荣耀。 他必如湍急的河流冲来， 耶和华的灵催逼他自己。
ISA|59|20|必有一位救赎主来到 锡安 ， 来到 雅各 族中离弃过犯的人那里； 这是耶和华说的。
ISA|59|21|耶和华说：“这就是我与他们所立的约：我加给你的灵，传给你的话，必不离你的口，也不离你后裔与你后裔之后裔的口，从今直到永远；这是耶和华说的。”
ISA|60|1|兴起，发光！因为你的光已来到！ 耶和华的荣光发出照耀着你。
ISA|60|2|看哪，黑暗笼罩大地， 幽暗遮盖万民， 耶和华却要升起照耀你， 他的荣光要显在你身上。
ISA|60|3|列国要来就你的光， 列王要来就你发出的光辉。
ISA|60|4|你举目向四围观看， 众人都聚集到你这里。 你的儿子从远方来， 你的女儿也被抱着带来。
ISA|60|5|那时，你看见就有光荣， 你的心兴奋欢畅 ； 因为大海那边的财富必归你， 列国的财宝也来归你。
ISA|60|6|成群的骆驼， 并 米甸 和 以法 的独峰驼遮满你； 示巴 的众人都必来到， 要奉上黄金和乳香， 又要传扬赞美耶和华的话。
ISA|60|7|基达 的羊群都聚集到你这里， 尼拜约 的公羊供你使用， 献在我坛上蒙悦纳； 我必荣耀我那荣耀的殿。
ISA|60|8|那些飞来如云、 又像鸽子飞向窗户的是谁呢？
ISA|60|9|众海岛必等候我 ， 他施 的船只领先， 将你的儿女，连同他们的金银从远方带来， 这都因 以色列 的圣者、耶和华－你上帝的名， 因为他已经荣耀了你。
ISA|60|10|外邦人要建造你的城墙， 他们的君王必服事你。 我曾发怒击打你， 如今却施恩怜悯你。
ISA|60|11|你的城门必时常开放， 昼夜不关， 使人将列国的财物带来归你， 他们的君王也被牵引而来。
ISA|60|12|不事奉你的那邦、那国要灭亡， 那些国家必全然荒废。
ISA|60|13|黎巴嫩 的荣耀， 就是松树、杉树、黄杨树， 都必一同归你， 用以装饰我圣所坐落之处； 我也要使我脚所踏之地得荣耀。
ISA|60|14|压制你的，他的子孙必来向你屈身； 藐视你的，都要在你脚前下拜。 人要称你为“耶和华的城”， 为“ 以色列 圣者的 锡安 ”。
ISA|60|15|你虽曾被抛弃，被恨恶， 甚至无人经过， 我却使你有永远的荣华， 成为世世代代的喜乐。
ISA|60|16|你要吃列国的奶， 吃列王的乳。 你就知道我－耶和华是你的救主， 是你的救赎主，是 雅各 的大能者。
ISA|60|17|我要赏赐金子代替铜， 赏赐银子代替铁， 铜代替木头， 铁代替石头。 我要以和平为你的官长， 以公义为你的监督。
ISA|60|18|你的地不再听闻残暴的事， 境内不再听见破坏与毁灭。 你必称你的墙为“拯救”， 称你的门为“赞美”。
ISA|60|19|白昼太阳不再作你的光， 月亮 也不再发光照耀你； 耶和华却要作你永远的光， 你的上帝要成为你的荣耀。
ISA|60|20|你的太阳不再落下， 月亮也不消失； 因为耶和华必作你永远的光。 你悲哀的日子定要结束。
ISA|60|21|你的居民全是义人， 永远得地为业； 他们是我栽的苗，是我手的工作， 为了彰显我的荣耀。
ISA|60|22|稀少的要成为大族， 弱小的要变为强国。 我－耶和华到了时候必速速成就这事。
ISA|61|1|主耶和华的灵在我身上， 因为耶和华用膏膏我， 叫我报好信息给贫穷的人， 差遣我医好伤心的人， 报告被掳的得释放， 被捆绑的得自由；
ISA|61|2|宣告耶和华的恩年 和我们的上帝报仇的日子； 安慰所有悲哀的人，
ISA|61|3|为 锡安 悲哀的人，赐华冠代替灰烬， 喜乐的油代替悲哀， 赞美为衣代替忧伤的灵； 称他们为“公义树”， 是耶和华所栽植的，为要彰显他的荣耀。
ISA|61|4|他们必修造久已荒凉的废墟， 建立先前凄凉之处， 重修历代荒凉之城。
ISA|61|5|那时，陌生人要伺候、牧放你们的羊群； 外邦人必为你们耕种田地， 修整你们的葡萄园。
ISA|61|6|但你们要称为“耶和华的祭司”， 称作“我们上帝的仆人”。 你们必享用列国的财物， 必承受他们的财富 。
ISA|61|7|因为他们所受双倍的羞辱， 凌辱被称为他们的命运， 因此，他们在境内必得双倍的产业， 永远之乐必归给他们。
ISA|61|8|因为我－耶和华喜爱公平， 恨恶抢夺与恶行 ； 我要凭诚实施行报偿， 与我的百姓立永约。
ISA|61|9|他们的后裔必在列国中为人所知， 他们的子孙在万民中为人所识； 凡看见他们的必承认他们是耶和华所赐福的后裔。
ISA|61|10|我因耶和华大大欢喜， 我的心因上帝喜乐； 因他以拯救为衣给我穿上， 以公义为外袍给我披上， 好像新郎戴上华冠， 又如新娘佩戴首饰。
ISA|61|11|地怎样使芽长出， 园子怎样使所栽种的生长， 主耶和华也必照样 使公义和赞美在万国中发出。
ISA|62|1|我因 锡安 必不静默， 为 耶路撒冷 必不安宁， 直到它的公义如光辉发出， 它的救恩如火把燃烧。
ISA|62|2|列国要看见你的公义， 列王要看见你的荣耀。 你必得新的名字， 是耶和华亲口起的。
ISA|62|3|你在耶和华的手中成为华冠， 在你上帝的掌上成为冠冕。
ISA|62|4|你不再称为“被撇弃的”， 你的地也不再称为“荒芜的”； 你要称为“我所喜悦的”， 你的地要称为“有归属的”。 因为耶和华喜悦你， 你的地必归属于他。
ISA|62|5|年轻人怎样娶童女， 你的百姓也要照样娶你； 新郎怎样因新娘而喜乐， 你的上帝也要如此以你为乐。
ISA|62|6|耶路撒冷 啊， 我在你城墙上设立守望者， 他们昼夜不停地呼喊。 呼求耶和华的啊，你们不要歇息，
ISA|62|7|也不要使他歇息， 直等他建立 耶路撒冷 ， 使 耶路撒冷 在地上为人所赞美。
ISA|62|8|耶和华指着自己的右手和大能的膀臂起誓说： “我必不再将你的五谷给仇敌作食物， 外邦人也必不再喝你劳碌得来的新酒。
ISA|62|9|惟有那收割的要吃，并赞美耶和华； 那储藏葡萄的要在我圣所院内喝。”
ISA|62|10|你们当从门经过，经过， 预备百姓的路。 你们要修筑，修筑大道， 清除石头， 为万民竖立大旗。
ISA|62|11|看哪，耶和华曾宣告到地极， 你们要对 锡安 说： “看哪，你的拯救者已来到。 看哪，他的赏赐在他那里， 他的报偿在他面前。”
ISA|62|12|人称他们为“圣民”，为“耶和华救赎的民”， 你也必称为“受眷顾的”，为“不被撇弃的城”。
ISA|63|1|这从 以东 的 波斯拉 来， 穿红衣服， 装扮华美， 能力广大， 大步向前迈进的是谁呢？ 就是我， 凭公义说话， 以大能施行拯救的。
ISA|63|2|你为何以红色装扮？ 你的衣服为何像踹醡酒池的人呢？
ISA|63|3|我独自踹醡酒池， 万民中并无一人与我同在。 我发怒，将他们踹下， 发烈怒将他们践踏。 他们的血溅在我的衣服上， 玷污了我一切的衣裳。
ISA|63|4|因为报仇之日在我心中， 救赎我民之年已经来到。
ISA|63|5|我仰望，见无人帮助； 我诧异，竟无人扶持。 因此，我的膀臂为我施行拯救； 我的烈怒将我扶持。
ISA|63|6|我发怒，踹下众民； 发烈怒，使他们喝醉， 又将他们的血倒在地上。
ISA|63|7|我要照耶和华一切所赐给我们的， 并他凭怜悯与丰盛的慈爱 所赐给 以色列 家的大恩， 述说他的慈爱和美德。
ISA|63|8|他说：“他们诚然是我的百姓， 未行虚假的子民。” 这样，他就作了他们的救主。
ISA|63|9|他们在一切苦难当中， 他也同受苦难， 并且他面前的使者拯救他们 。 他以慈爱和怜悯救赎他们， 在古时的日子时常抱他们，背他们。
ISA|63|10|他们竟然悖逆，使他的圣灵忧伤。 他就转变，成为他们的仇敌， 亲自攻击他们。
ISA|63|11|那时，他的百姓想起古时 摩西 的日子： “那将百姓和牧养群羊的人 从海里领上来的在哪里呢？ 那将圣灵降在他们中间，
ISA|63|12|以荣耀的膀臂在 摩西 右边行动， 在百姓面前将水分开， 为要建立自己永远的名，
ISA|63|13|又带领他们经过深处的在哪里呢？” 他们如马行走旷野，不致绊跌；
ISA|63|14|又如牲畜下到山谷， 耶和华的灵使他们得安息； 照样，你也引导你的百姓， 为要建立自己荣耀的名。
ISA|63|15|求你从天上， 从你神圣荣耀的居所垂顾观看。 你的热心和你大能的作为在哪里呢？ 你内心的关怀和你的怜悯向我们停止了。
ISA|63|16|亚伯拉罕 虽然不承认我们， 以色列 也不承认我们， 你却是我们的父。 耶和华啊，你是我们的父； 自古以来，你的名是“我们的救赎主”。
ISA|63|17|耶和华啊，你为何使我们偏离你的道， 使我们心里刚硬、不敬畏你呢？ 求你为你的仆人， 为你产业的支派而回转。
ISA|63|18|你的圣民暂时得你的圣所， 但我们的敌人践踏了它。
ISA|63|19|我们就成了你未曾治理的人， 成了未曾称为你名下的人。
ISA|64|1|愿你破天而降， 愿山在你面前震动，
ISA|64|2|好像火烧干柴， 又如火将水烧开， 使你敌人知道你的名， 列国必在你面前发颤！
ISA|64|3|你曾做我们不能逆料可畏的事； 那时你降临，山岭在你面前震动。
ISA|64|4|自古以来，人未曾听见，未曾耳闻，未曾眼见， 除你以外，还有上帝能为等候他的人行事。
ISA|64|5|你迎见那欢喜行义、记念你道的人； 看哪，你曾发怒，因我们犯了罪； 这景况已久，我们还能得救吗？
ISA|64|6|我们都如不洁净的人， 所行的义都像污秽的衣服。 我们如叶子渐渐枯干， 罪孽像风把我们吹走。
ISA|64|7|无人求告你的名， 无人奋力抓住你。 你转脸不顾我们， 你使我们因罪孽而融化 。
ISA|64|8|但耶和华啊，现在你仍是我们的父！ 我们是泥，你是陶匠； 我们都是你亲手所造的。
ISA|64|9|耶和华啊，求你不要大发震怒， 也不要永远记得罪孽； 看哪，求你垂顾我们， 因我们都是你的百姓。
ISA|64|10|你的圣城已变为旷野； 锡安 变为旷野， 耶路撒冷 成为废墟。
ISA|64|11|我们那神圣华美的殿， 就是我们祖先赞美你的地方，已被火焚烧； 我们所羡慕的美地尽都荒芜。
ISA|64|12|耶和华啊，有这些事，你还能忍受吗？ 你还静默，使我们大受苦难吗？
ISA|65|1|没有求问我的，我要让他们找到； 没有寻找我的，我要让他们寻见； 我对没有呼求我名的国 说： “我在这里！我在这里！”
ISA|65|2|我整天向那悖逆的百姓招手， 他们随自己的意念行不善之道。
ISA|65|3|这百姓时常当面惹我发怒， 在园中献祭， 在砖上烧香，
ISA|65|4|在坟墓间停留， 在隐密处过夜， 吃猪肉， 器皿中有不洁净之肉熬的汤；
ISA|65|5|且对人说：“你站开吧！ 不要挨近我，因为我对你来说太神圣了 。” 这些人惹我鼻中冒烟， 如终日燃烧的火。
ISA|65|6|看哪，这些都写在我面前。 我必不静默，却要施行报应， 将你们和你们祖先的罪孽 全都报应在后人身上； 因为他们在山上烧香， 在冈上亵渎我， 我要按他们先前所行的，报应在他们身上 ； 这是耶和华说的。
ISA|65|7|
ISA|65|8|耶和华如此说： “人在葡萄中寻得新酒时会说： ‘不要毁坏它，因为它还有用处’； 同样，我必因我仆人的缘故， 不将他们全然毁灭。
ISA|65|9|我必从 雅各 中领出后裔， 从 犹大 中领出那要继承我众山的； 我的选民要继承它， 我的仆人要在那里居住。
ISA|65|10|沙仑 必成为羊群的圈， 亚割谷 成为牛群躺卧之处， 都为寻求我的民所得。
ISA|65|11|但你们这些离弃耶和华， 就是忘记我的圣山、 为‘幸运之神’摆设筵席、 为‘命运之神’装满调和酒的，
ISA|65|12|我命定你们归于刀下， 你们都要屈身被杀； 因为我呼唤，你们不回应； 我说话，你们不听从； 反倒做我眼中看为恶的事， 选择我所不喜悦的事。”
ISA|65|13|所以，主耶和华如此说： “看哪，我的仆人必得吃，你们却饥饿； 看哪，我的仆人必得喝，你们却干渴； 看哪，我的仆人必欢喜，你们却蒙羞。
ISA|65|14|看哪，我的仆人因心中喜乐而欢呼， 你们却因心里悲痛而哀哭， 因灵里忧伤而哀号。
ISA|65|15|你们必留下自己的名 给我选民指着赌咒： 主耶和华必杀你们， 另起别名称呼他的仆人。
ISA|65|16|在地上为自己求福的， 必凭真实的上帝求福； 在地上起誓的， 必指着真实的上帝起誓。 因为从前的患难已被遗忘， 从我眼前消逝。”
ISA|65|17|“看哪，我造新天新地！ 从前的事不再被记念，也不被人放在心上；
ISA|65|18|当因我所造的欢喜快乐，直到永远； 看哪，因为我造 耶路撒冷 为人所喜， 造其中的居民为人所乐。
ISA|65|19|我必因 耶路撒冷 欢喜， 因我的百姓快乐， 那里不再听见哭泣和哀号的声音。
ISA|65|20|那里没有数日夭折的婴孩， 也没有寿数不满的老人； 因为百岁死的仍算孩童， 未达百岁而亡的 算是被诅咒的。
ISA|65|21|他们建造房屋，居住其中， 栽葡萄园，吃园中的果子；
ISA|65|22|并非造了给别人居住， 也非栽种给别人享用； 因为我百姓的日子必长久如树木， 我的选民必享受亲手劳碌得来的。
ISA|65|23|他们必不徒然劳碌， 所生产的，也不遭灾害， 因为他们和他们的子孙 都是蒙耶和华赐福的后裔。
ISA|65|24|他们尚未求告，我就应允； 正说话的时候，我就垂听。
ISA|65|25|野狼必与羔羊同食， 狮子必吃草，与牛一样， 蛇必以尘土为食物； 在我圣山的遍处， 它们都不伤人，也不害物； 这是耶和华说的。”
ISA|66|1|耶和华如此说： “天是我的座位； 地是我的脚凳。 你们能为我造怎样的殿宇呢？ 哪里是我安歇的地方呢？
ISA|66|2|这一切是我手所造的， 这一切就都存在了。 我所看顾的是困苦、灵里痛悔、 因我言语而战兢的人。 这是耶和华说的。
ISA|66|3|“至于那些宰牛，杀人， 献羔羊，打断狗颈项， 献猪血为供物， 烧乳香，称颂偶像的， 他们选择自己的道路， 心里喜爱可憎恶的事；
ISA|66|4|我也必选择苦待他们， 使他们所惧怕的临到他们； 因为我呼唤，无人回应； 我说话，他们不听从； 反倒做我眼中看为恶的事， 选择我所不喜悦的事。”
ISA|66|5|你们因耶和华言语而战兢的人哪，当听他的话： “你们的弟兄，就是恨恶你们， 因我名赶出你们的，曾说： ‘愿耶和华彰显荣耀 ， 好让我们看见你们的喜乐。’ 但蒙羞的终究是他们！
ISA|66|6|“有喧哗的声音出自城中！ 有声音来自殿里！ 是耶和华向仇敌施行报应的声音！
ISA|66|7|“ 锡安 未曾阵痛就生产， 疼痛尚未来到，就生出男孩。
ISA|66|8|国岂能一日而生？ 民岂能一时而产？ 但 锡安 一阵痛就生下儿女， 这样的事有谁听见， 有谁看见呢？
ISA|66|9|耶和华说：我使人临产， 岂不让她 生产呢？ 你的上帝说：我使人生产， 难道还让她关闭 不生吗？
ISA|66|10|“你们所有爱慕 耶路撒冷 的啊， 要与她一同欢喜，为她高兴； 你们所有为她悲哀的啊， 都要与她一同乐上加乐；
ISA|66|11|使你们在她安慰的怀中吃奶得饱， 尽情吸取她丰盛的荣耀，满心喜乐。”
ISA|66|12|耶和华如此说： “看哪，我要使平安临到她，好像江河； 使列国的荣耀及于她，如同涨溢的溪流。 你们要尽情吸吮； 你们必被抱在身旁 ，摇弄在膝上。
ISA|66|13|我要安慰你们，如同母亲安慰儿女； 你们也必在 耶路撒冷 得安慰。
ISA|66|14|你们看见，心里就喜乐， 你们的骨头必如草生长； 耶和华的手在他仆人身上彰显， 他却要向他的仇敌发怒。”
ISA|66|15|看哪，耶和华必在火中降临， 他的战车宛如暴风， 以烈怒施行报应， 以火焰施行责罚；
ISA|66|16|耶和华必以火与刀审判凡有血肉之躯的， 被耶和华所杀的很多。
ISA|66|17|那些洁净自己献给偶像，进入园内，跟随其中一个人去吃猪肉和鼠肉，并可憎之物的，他们必一同灭绝。这是耶和华说的。
ISA|66|18|我知道他们的行为和他们的意念。聚集万国万族 的时候到了 ，他们要来瞻仰我的荣耀；
ISA|66|19|我要在他们中间显神迹，差遣他们当中的幸存者到列国去，就是到 他施 、 普勒 、以善射闻名的 路德 、 土巴 、 雅完 ，和未曾听见我名声，未曾看见我荣耀的遥远海岛那里去；他们必在列国中传扬我的荣耀。
ISA|66|20|他们要将你们的弟兄从列国中带回，或骑马，或坐车，或乘蓬车，或骑骡子，或骑独峰驼，到我的圣山 耶路撒冷 ，作为供物献给耶和华。这是耶和华说的。正如 以色列 人用洁净的器皿盛供物奉到耶和华的殿中，
ISA|66|21|我也必从他们中间立人作祭司，作 利未 人。这是耶和华说的。
ISA|66|22|“我所造的新天新地在我面前长存， 你们的后裔和你们的名号也必照样长存。 这是耶和华说的。
ISA|66|23|每逢初一、安息日， 凡有血肉之躯的必前来，在我面前下拜； 这是耶和华说的。
ISA|66|24|“他们要出去观看那些违背我的人的尸首， 他们的虫是不死的， 他们的火是不灭的， 凡有血肉之躯的都必憎恶他们。”
JER|1|1|这些是 便雅悯 地 亚拿突城 的祭司， 希勒家 的儿子 耶利米 的话。
JER|1|2|亚们 的儿子 犹大 王 约西亚 在位第十三年，耶和华的话临到 耶利米 。
JER|1|3|从 约西亚 的儿子 犹大 王 约雅敬 在位的时候，直到 约西亚 的儿子 犹大 王 西底家 在位的末年，就是第十一年五月间 耶路撒冷 被掳时，耶和华的话也常临到 耶利米 。
JER|1|4|耶利米 说，耶和华的话临到我，说：
JER|1|5|“我尚未将你造在母腹中，就已认识你； 你未出母胎，我已将你分别为圣， 派你作列国的先知。”
JER|1|6|我就说：“唉，主耶和华！看哪，我不知道怎么说，因为我年轻。”
JER|1|7|耶和华对我说： “不要说：‘我年轻’， 因为我差遣你到谁那里去，你都要去； 我吩咐你说什么话，你都要说。
JER|1|8|你不要怕他们， 因为我与你同在，要拯救你。 这是耶和华说的。”
JER|1|9|于是耶和华伸手按住我的口， 对我说： “看哪，我已将我的话放在你口中。
JER|1|10|我今日立你在列邦列国之上， 为要拔出，拆毁，毁坏，倾覆， 又要建立，栽植。”
JER|1|11|耶和华的话临到我，说：“ 耶利米 ，你看见什么？”我说：“我看见一根杏树枝。”
JER|1|12|耶和华对我说：“你看得不错；因为我要看守 我的话，使它实现。”
JER|1|13|耶和华的话第二次临到我，说：“你看见什么？”我说：“我看见一个水烧开的锅，从北而倾。”
JER|1|14|耶和华对我说：“必有灾祸从北方发出，临到这地所有的居民。
JER|1|15|看哪，我要召北方列国的万族。这是耶和华说的。他们要来，各安宝座在 耶路撒冷 的城门口，周围攻击城墙，又要攻击 犹大 的一切城镇。
JER|1|16|这百姓离弃我，向别神烧香，跪拜自己手所造的，我要针对这一切恶行，向他们宣读我的判决。
JER|1|17|所以你当束腰，起来，将我所吩咐你的一切话都告诉他们；不要因他们惊惶，免得我使你在他们面前惊惶。
JER|1|18|看哪，我今日使你成为坚城、铁柱、铜墙，对抗全地和 犹大 的君王、官长、祭司，并这地的百姓。
JER|1|19|他们要攻击你，却不能胜过你，因为我与你同在，要拯救你。这是耶和华说的。”
JER|2|1|耶和华的话临到我，说：
JER|2|2|“你去向 耶路撒冷 居民的耳朵呼喊说，耶和华如此说： ‘你年轻时的恩爱， 新婚时的爱情， 你怎样在旷野， 在未耕种之地跟随我， 我都记得。
JER|2|3|那时 以色列 归耶和华为圣， 作为他初熟的土产； 凡吞吃它的必算为有罪， 灾祸必临到他们。 这是耶和华说的。’”
JER|2|4|雅各 家， 以色列 家的各族啊，当听耶和华的话，
JER|2|5|耶和华如此说： “你们的祖先看我有什么错处， 竟远离我，随从那虚无的神明 ， 自己成为虚无呢？
JER|2|6|他们并不问： ‘那领我们从 埃及 地上来， 引导我们走过旷野、沙漠有坑洞之地， 走过干旱死荫、无人经过、 无人居住之地的耶和华在哪里呢？’
JER|2|7|我领你们进入肥沃之地， 使你们得吃其中的果子和美物； 你们进入时，却使我的地玷污， 使我的产业成为可憎恶的。
JER|2|8|祭司从来不问：‘耶和华在哪里呢？’ 传讲律法的不认识我， 官长违背我， 先知藉 巴力 说预言， 随从无益的东西。”
JER|2|9|“我因此必与你们争辩， 也与你们的子孙争辩。 这是耶和华说的。
JER|2|10|你们且渡到 基提 海岛察看， 派人往 基达 去留心查考， 看可曾有过这样的事。
JER|2|11|岂有一国换了它的神明吗？ 其实那不是神明！ 但我的百姓将他们的荣耀换了那无益的东西。
JER|2|12|诸天哪，要因此震惊， 颤栗，极其凄凉！ 这是耶和华说的。
JER|2|13|因为我的百姓做了两件恶事： 离弃我这活水的泉源； 又为自己凿出水池， 却是破裂不能储水的池子。”
JER|2|14|“ 以色列 是仆人吗？ 是家中生的奴仆吗？ 为何成为掠物呢？
JER|2|15|少壮狮子向它咆哮，大声吼叫， 使它的地荒芜； 城镇烧毁，无人居住。
JER|2|16|挪弗 人和 答比匿 人打破你的头颅。
JER|2|17|这不是你自己招惹的吗？ 不是因耶和华－你上帝引导你行路时， 你离弃了他吗？
JER|2|18|现今你为何在 埃及 路上喝 西曷河 的水呢？ 为何在 亚述 路上喝 大河 的水呢？
JER|2|19|你自己的恶必惩治你， 你背道的事必责罚你。 由此可知可见，你离弃耶和华－你的上帝， 不存敬畏我的心， 实为恶事，为苦事； 这是万军之主耶和华说的。”
JER|2|20|“你 在古时折断你的轭，解开你的绳索， 说：‘我必不事奉耶和华 。’ 你在各高冈上、各青翠的树下屈身行淫。
JER|2|21|然而，我栽种你为上等的葡萄树， 全用纯正的种子； 你怎么向我变为外邦葡萄树的坏枝子呢？
JER|2|22|你虽用碱、多用皂荚清洗， 你罪孽的痕迹仍显在我面前。 这是主耶和华说的。
JER|2|23|你怎能说： ‘我没有玷污，没有随从 巴力 ’？ 看看你在谷中所做的，思想你自己的所作所为； 你是快行的独峰驼，狂奔乱闯。
JER|2|24|你是野驴，习惯旷野， 欲心发动时就呼吸急促， 发情时谁能使它转回呢？ 凡寻找它的必不费力， 在它的季节必能寻见它。
JER|2|25|你不要弄到赤足而行， 喉咙干渴。 你却说：‘没有用的， 我喜爱陌生人， 我必随从他们。’”
JER|2|26|“贼被捉拿，怎样羞愧， 以色列 家和他们的君王、官长、 祭司、先知也都照样羞愧。
JER|2|27|他们向木头说：‘你是我的父’； 向石头说：‘你是生我的。’ 他们以背向我， 不肯以面向我； 及至遭遇患难时却说： ‘起来拯救我们吧！’
JER|2|28|你为自己做的神明在哪里呢？ 你遭遇患难的时候， 让它们起来拯救你吧！ 犹大 啊，你神明的数目与你城的数目相等。
JER|2|29|“你们为何与我争辩呢？ 你们都违背了我。 这是耶和华说的。
JER|2|30|我责打你们的儿女是徒然的， 他们不受管教。 你们自己的刀吞灭你们的先知， 好像残害人的狮子。
JER|2|31|这世代的人哪， 你们要留意耶和华的话。 我向 以色列 岂是旷野， 或幽暗之地呢？ 我的百姓为何说： ‘我们脱离约束，不再归向你了’？
JER|2|32|少女岂能忘记她的妆饰呢？ 新娘岂能忘记她的美衣呢？ 我的百姓却在无数的日子里忘记了我！
JER|2|33|“你竟然如此精于求爱之道， 可把你的门径教邪恶的女人！
JER|2|34|你衣服的边上有无辜贫穷人的血， 其实你并未发现他们挖洞进屋偷窃 。 虽有这一切的事 ，
JER|2|35|你还说：‘我无辜； 耶和华的怒气必定转离我了。’ 看哪，我必审问你； 因你自己说：‘我没有犯罪。’
JER|2|36|你为何东奔西跑改变你的道路呢？ 你必因 埃及 蒙羞， 像从前因 亚述 蒙羞一样。
JER|2|37|你也必两手抱头离开这里； 因为耶和华已经弃绝你所倚靠的， 你不能因他们而得顺利。”
JER|3|1|耶和华说 ：“人若休妻， 妻离他而去，做了别人的妻子， 前夫岂能再回到她那里呢？ 那地岂不是大大污秽了吗？ 但你和许多情郎行淫， 还是可以回到我这里。 这是耶和华说的。
JER|3|2|你举目向光秃的高地观看， 何处没有你的淫行呢？ 你坐在道路旁等候， 好像 阿拉伯 人在旷野埋伏， 你的淫行和邪恶使全地污秽了。
JER|3|3|因此甘霖停止， 春雨不降。 你还是一副娼妓之脸， 不顾羞耻。
JER|3|4|你不是才向我呼叫说： ‘我父啊，你是我年轻时的密友，
JER|3|5|人岂永远怀恨，长久存怒吗？’ 看哪，你虽这样说，还是竭尽所能去行恶。”
JER|3|6|约西亚 王在位的时候，耶和华对我说：“你看见背道的 以色列 所做的吗？她上到各高山，在各青翠的树下行淫。
JER|3|7|我说：‘她行这些事以后会回转归向我’，她却不回转。她奸诈的妹妹 犹大 也看见了。
JER|3|8|我看见背道的 以色列 行淫，我为这缘故给她休书休了她，她奸诈的妹妹 犹大 还不惧怕，也去行淫。
JER|3|9|因 以色列 轻忽了她的淫乱，与石头和木头行奸淫 ，她和这地就都污秽了 。
JER|3|10|虽有这一切的事，她奸诈的妹妹 犹大 还不一心归向我，不过是假意归我。这是耶和华说的。”
JER|3|11|耶和华对我说：“背道的 以色列 比奸诈的 犹大 还显为义。
JER|3|12|你去向北方宣告这些话，说： ‘背道的 以色列 啊，回来吧！ 这是耶和华说的。 我必不怒目看你们， 因为我是慈爱的， 这是耶和华说的。 我必不永远怀怒；
JER|3|13|只要你承认你的罪孽， 就是违背耶和华－你的上帝， 在各青翠的树下追逐外族的神明 ， 没有听从我的话。 这是耶和华说的。
JER|3|14|背道的儿女啊，回来吧！ 这是耶和华说的。 因为我作你们的丈夫， 要将你们从一城取一人， 从一族取两人，带到 锡安 。
JER|3|15|“‘我必将合我心意的牧者赏赐给你们，他们要以知识和智慧牧养你们。
JER|3|16|你们在国中生养众多的时候，那些日子，人必不再提说耶和华的约柜，不追想，不记念，不觉缺少，也不再制造。这是耶和华说的。
JER|3|17|那时，人必称 耶路撒冷 为耶和华的宝座；万国聚集在那里，为耶和华的名来到 耶路撒冷 ，他们必不再随从自己顽梗的恶心行事。
JER|3|18|当那些日子， 犹大 家要和 以色列 家同行，从北方之地一同来到我所赐给你们祖先为业之地。’”
JER|3|19|我说，我多么乐意把你列在儿女之中， 赐给你美地， 就是万国中最美的产业。 我说，你会以“我父啊”称呼我， 不再转离而跟从我。
JER|3|20|以色列 家啊，你们向我行诡诈， 真像妻子行诡诈离开丈夫。 这是耶和华说的。
JER|3|21|有声音从光秃的高地传来， 就是 以色列 人哭泣恳求的声音， 因为他们走弯曲之道， 忘记耶和华－他们的上帝。
JER|3|22|“你们这背道的儿女啊，回来吧！ 我要医治你们背道的病。” “看哪，我们来到你这里， 因你是耶和华－我们的上帝。
JER|3|23|从小山来的真是枉然， 大山的喧嚷也是枉然 。 以色列 得救，诚然在乎耶和华－我们的上帝。
JER|3|24|“从我们幼年以来，那可耻之物 吞吃了我们祖先劳碌得来的，就是他们的羊群、牛群和他们的儿女。
JER|3|25|我们在羞耻中躺卧吧！愿惭愧将我们遮盖！因为从我们幼年以来，我们和我们的祖先都得罪了耶和华－我们的上帝，没有听从耶和华－我们上帝的话。”
JER|4|1|耶和华说：“ 以色列 啊， 你若回转，回转归向我， 若从我眼前除掉你可憎的偶像， 不再犹疑不定，
JER|4|2|凭诚实、公平、公义 指着永生的耶和华起誓； 列国就必因他蒙福， 也必因他夸耀。”
JER|4|3|耶和华对 犹大 人和 耶路撒冷 人如此说： “你们要为自己开垦荒地， 不要撒种在荆棘里。
JER|4|4|犹大 人和 耶路撒冷 的居民哪， 你们当自行割礼，归耶和华， 将你们心里的污秽 除掉； 免得我的愤怒因你们的恶行发作， 如火燃起， 甚至无人能熄灭！”
JER|4|5|你们要在 犹大 传扬， 在 耶路撒冷 宣告，说： “当在国中吹角，高声呼叫说： ‘你们当聚集！ 我们好进入坚固城！’
JER|4|6|应当向 锡安 竖立大旗。 逃吧，不要迟延， 因我必使灾祸与大毁灭从北方来到。
JER|4|7|有狮子从密林中上来， 是毁坏列国的。 它已动身出离本处， 要使你的地荒凉， 使你的城镇变为废墟，无人居住。
JER|4|8|因此，你们当腰束麻布，哭泣哀号， 因为耶和华的烈怒并未转离我们。”
JER|4|9|耶和华说：“到那时，君王和领袖的心要失丧，祭司都要惊奇，先知都要诧异。”
JER|4|10|我说：“哀哉！主耶和华啊，你真是大大欺哄这百姓和 耶路撒冷 ，说：‘你们必得平安。’其实刀剑已经抵住喉咙了！”
JER|4|11|那时，必有话对这百姓和 耶路撒冷 说：“来自旷野光秃高地的热风吹向我的百姓 ，不是为簸扬，也不是为扬净。
JER|4|12|又有一阵比这更大的风向我刮来；现在，我要向他们宣读我的判决。”
JER|4|13|看哪，他必如云涌上； 他的战车如旋风， 他的马比鹰更快。 我们有祸了！ 我们败落了！
JER|4|14|耶路撒冷 啊，你当洗去心中的恶， 使你可以得救。 恶念在你里面要存到几时呢？
JER|4|15|有声音从 但 传出， 有灾祸从 以法莲山 传来。
JER|4|16|你们当传给列国， 看哪，要向 耶路撒冷 报告： “有围攻的人从远方来到， 向 犹大 的城镇大声喊叫。
JER|4|17|他们包围 耶路撒冷 ， 好像看守田园的， 因为它背叛了我。 这是耶和华说的。
JER|4|18|你的作风和行为招惹这事； 这是你罪恶的结果， 实在是苦， 刺透了你的心！”
JER|4|19|我的肺腑啊，我的肺腑啊，我心疼痛！ 我的心在我里面烦躁不安。 我不能静默不言， 因我已听见角声和打仗的喊声。
JER|4|20|毁坏的信息不断传来， 因为全地荒废。 我的帐棚忽然毁坏， 我的幔子顷刻破裂。
JER|4|21|我看见大旗，听见角声， 要到几时呢？
JER|4|22|“我的百姓愚顽，不认识我； 他们是愚昧无知的儿女， 有智慧行恶，没有知识行善。”
JER|4|23|我观看地， 看哪，地是空虚混沌； 我观看天，天也无光。
JER|4|24|我观看大山，看哪，尽都震动， 小山也都摇来摇去。
JER|4|25|我观看，看哪，无人； 空中的飞鸟也都躲避。
JER|4|26|我观看，看哪，肥田变为荒地； 所有城镇在耶和华面前， 因他的烈怒都被拆毁。
JER|4|27|耶和华如此说：“全地必然荒凉， 我却不毁灭净尽。
JER|4|28|因此，地要悲哀， 天上也必黑暗； 因为我言已出，我意已定， 必不改变，也不由此转回。”
JER|4|29|各城的人因骑兵和弓箭手的响声就都逃跑， 进入密林，爬上磐石； 城镇都被抛弃， 无人住在其中。
JER|4|30|你这被毁灭的啊， 你要做什么呢？ 你穿上朱红衣服， 佩戴黄金饰物， 用眼影修饰眼睛， 徒然美化你自己。 恋慕你的却藐视你， 寻索你的性命。
JER|4|31|我听见仿佛妇人临产的声音， 好像生头胎疼痛的声音， 原来是 锡安 的声音； 她喘着气，伸开手： “我有祸了！ 在杀人者跟前，我的心灵发昏。”
JER|5|1|你们要走遍 耶路撒冷 的街市， 在广场寻找， 看是否有人行公平、求诚实； 若有，我就赦免这城。
JER|5|2|虽然他们说“我对永生的耶和华发誓”， 所起的誓实在是假的。
JER|5|3|耶和华啊，你的眼目不是在寻找诚实吗？ 你击打他们，他们却不伤恸； 你摧毁他们，他们仍不领受管教。 他们使脸刚硬过于磐石， 不肯回头。
JER|5|4|我说：“这些人实在是贫寒的， 他们是愚昧的， 因为不知道耶和华的作为， 也不知道他们上帝的法则。
JER|5|5|我要去见尊贵的人，向他们说话， 他们应该知道耶和华的作为， 知道他们上帝的法则。” 然而，这些人却齐心将轭折断， 挣开绳索。
JER|5|6|因此，林中的狮子必害死他们， 野地的狼必灭绝他们， 豹子在城外窥伺。 凡出城的必被撕碎， 因为他们的罪过极多， 背道的事也增加。
JER|5|7|我怎能赦免你呢？ 你的儿女离弃我， 又指着那不是上帝的起誓。 我使他们饱足， 他们就行奸淫， 居住 在娼妓家里。
JER|5|8|他们如喂饱的马，精力旺盛， 各向邻舍的妻子吹哨。
JER|5|9|我岂不因这些事施行惩罚吗？ 像这样的国家，我岂能不报复呢？ 这是耶和华说的。
JER|5|10|你们要上去毁坏它的葡萄园， 但不可毁坏净尽， 只可除掉其枝子， 因为不属耶和华。
JER|5|11|以色列 家和 犹大 家向我大行诡诈。 这是耶和华说的。
JER|5|12|关乎耶和华他们说了虚谎的话： “他不会的， 灾祸必不临到我们， 我们也不会遇见刀剑和饥荒。
JER|5|13|先知不过是一阵风， 道也不在他们里面； 这灾祸必临到他们身上。”
JER|5|14|所以耶和华－万军之上帝如此说： “因为他们说这话， 看哪，我必使我的话在你口中为火， 使这百姓为柴， 火便将他们烧灭。
JER|5|15|以色列 家啊， 看哪，我必使一国从远方来攻击你， 是强盛的国， 是古老的国； 他们的言语你不知道， 所说的话你不明白。 这是耶和华说的。
JER|5|16|他们的箭袋有如敞开的坟墓， 他们全都是勇士。
JER|5|17|他们必吃尽你的庄稼和粮食， 是你儿女该吃的 ； 必吃尽你的牛羊， 吃尽你的葡萄和无花果； 又必用刀剑毁坏你所倚靠的坚固城。
JER|5|18|“就是在那些日子，我也不会将你们毁灭净尽。这是耶和华说的。
JER|5|19|百姓若说：‘耶和华－我们的上帝为什么向我们行这一切事呢？’你就对他们说：‘你们怎样离弃我，在你们的地上事奉外邦神明，也必照样在不属你们的地上事奉外族人。’”
JER|5|20|当在 雅各 家传扬， 在 犹大 宣告，说：
JER|5|21|“愚昧无知的百姓啊， 你们有眼不看， 有耳不听， 现在当听这话。
JER|5|22|你们难道不惧怕我吗？ 在我面前还不战兢吗？ 这是耶和华说的。 我以沙为海的界限， 作永远的条例，使它不得越过。 波浪汹涌，却不能胜过； 怒涛澎湃，仍无法越过。
JER|5|23|但这百姓有背叛忤逆的心， 他们转离而去。
JER|5|24|他们心里并不说： ‘我们应当敬畏耶和华－我们的上帝； 他按时赐雨，就是秋雨和春雨， 又为我们定收割的季节。’
JER|5|25|你们的罪孽使这些转离你们， 你们的罪恶使你们不能得福。
JER|5|26|在我百姓当中有恶人， 他们埋伏，好像捕鸟的人在窥探 ； 他们设罗网陷害人。
JER|5|27|笼子怎样装满雀鸟， 他们的屋里也照样充满诡诈； 他们因此得以强大富足。
JER|5|28|他们肥胖光润，作恶过甚， 不为人伸冤， 不为孤儿伸冤，使他们胜诉， 也不为贫穷人辩护。
JER|5|29|我岂不因这些事施行惩罚吗？ 像这样的国家，我岂能不报复呢？ 这是耶和华说的。
JER|5|30|“国中有令人惊骇、 恐怖的事发生，
JER|5|31|先知说假预言， 祭司把权柄抓在自己手上， 我的百姓也喜爱这样， 到了结局你们要怎么办呢？”
JER|6|1|便雅悯 人哪，当逃离 耶路撒冷 ， 在 提哥亚 吹号角， 在 伯．哈基琳 升信号， 因为有灾祸与大毁灭从北方逼近。
JER|6|2|那秀美娇嫩的 锡安 ， 我必剪除。
JER|6|3|牧人必引领羊群到它那里， 在它周围支搭帐棚， 各在自己的地方放牧。
JER|6|4|“你们要准备攻击它。 起来吧，我们要趁正午上去。” “哀哉！日已渐斜， 黄昏的影子拖长了。”
JER|6|5|“起来吧，我们要在夜间上去， 毁坏它的宫殿。”
JER|6|6|万军之耶和华如此说： “你们要砍伐树木， 建土堆攻打 耶路撒冷 ， 就是那该受罚的城 ， 其中尽是欺压。
JER|6|7|井怎样涌出水来， 这城也照样涌出恶来； 其中常听闻残暴毁灭的事， 病痛损伤也常在我面前。
JER|6|8|耶路撒冷 啊，当受管教， 免得我心与你生疏， 免得我使你荒凉， 成为无人居住之地。”
JER|6|9|万军之耶和华如此说： “他们洗劫 以色列 剩下的民， 如摘净葡萄一样； 现你的手如采收葡萄的人，在树枝上采了又采 。”
JER|6|10|现在我可以向谁说话，警告谁，使他们听呢？ 看哪，他们的耳朵未受割礼，不能听见。 看哪，他们以耶和华的话为羞辱， 不以为喜悦。
JER|6|11|因此我被耶和华的愤怒充满，难以忍受。 “你要把它倒在街上孩童 和成群的年轻人身上， 他们连夫带妻， 年长者与高龄的人都必被擒拿。
JER|6|12|他们的房屋、田地， 和妻子都要一起转归别人， 我要伸手攻击这地的居民。” 这是耶和华说的。
JER|6|13|“因为他们从最小的到最大的都贪图不义之财， 从先知到祭司全都行事虚假。
JER|6|14|他们轻忽地医治我百姓的损伤， 说：‘平安了！平安了！’ 其实没有平安。
JER|6|15|他们行可憎之事，应当羞愧； 然而他们却一点也不觉得羞愧， 也不知羞耻。 因此，他们必与仆倒的人一同仆倒， 我惩罚他们的时候， 他们必跌倒。” 这是耶和华说的。
JER|6|16|耶和华如此说： “你们当站在路边察看， 寻访古老的路， 哪里是完善的道路，就行走在其上； 这样，你们自己必找到安息。 他们却说：‘我们不走。’
JER|6|17|我为你们设立守望的人， 要留心听角声。 他们却说：‘我们不听。’
JER|6|18|因此，列国啊，当听！ 会众啊，要知道他们必遭遇的事。
JER|6|19|地啊，当听！ 看哪，我必使灾祸临到这百姓， 是他们计谋所结的果子； 因为他们不肯留心听我的话， 至于我的律法，他们也厌弃。
JER|6|20|从 示巴 来的乳香， 从远方出的香菖蒲， 奉来给我有何用呢？ 你们的燔祭不蒙悦纳； 你们的祭物，我也不喜悦。”
JER|6|21|所以耶和华如此说： “看哪，我要将绊脚石放在这百姓面前； 父亲和儿子要一同跌在其上， 邻舍与朋友也都灭亡。”
JER|6|22|耶和华如此说： “看哪，有一民族从北方而来； 有一大国被激起，从地极来到。
JER|6|23|他们拿弓和枪， 性情残忍，不施怜悯； 他们的声音如海浪澎湃。 锡安 哪， 他们都骑马， 如上战场的人摆阵攻击你。”
JER|6|24|我们听见这样的风声，手就发软； 痛苦将我们抓住， 疼痛仿佛临产的妇人。
JER|6|25|你们不要出到田野去， 也不要行走在路上， 因四围有仇敌的刀剑和惊吓。
JER|6|26|我的百姓 啊，应当腰束麻布，滚在灰中。 要悲伤，如丧独子般痛痛哭号， 因为灭命的忽然临到我们。
JER|6|27|我使你作我百姓的测试者 和考验者 ， 使你知道并考验他们的行为。
JER|6|28|他们极其悖逆， 到处毁谤人， 他们是铜是铁， 全都败坏了。
JER|6|29|风箱吹火，铅被烧毁， 炼而又炼，终是徒然， 因为恶劣的还未除掉。
JER|6|30|人必称他们为被抛弃的银子， 因为耶和华已经抛弃了他们。
JER|7|1|耶和华的话临到 耶利米 ，说：
JER|7|2|“你当站在耶和华殿的门口，在那里宣讲这话说：所有从这些门进来敬拜耶和华的 犹大 人哪，当听耶和华的话。
JER|7|3|万军之耶和华－ 以色列 的上帝如此说：你们要改正你们的所作所为，我就使你们仍然居住这地 。
JER|7|4|不要倚靠虚谎的话，说：‘这是耶和华的殿，是耶和华的殿，是耶和华的殿！’
JER|7|5|“你们若实在改正你们的所作所为，彼此诚然施行公平，
JER|7|6|不欺压寄居的和孤儿寡妇，不在这地方流无辜人的血，也不随从别神陷害自己，
JER|7|7|我就使你们仍然居住这地 ，就是我从古时所赐给你们祖先的地，从永远到永远。
JER|7|8|“看哪，你们倚靠虚谎无益的话语。
JER|7|9|你们岂可偷盗，杀害，奸淫，起假誓，向 巴力 烧香，随从素不认识的别神，
JER|7|10|又来到这称为我名下的殿，在我面前敬拜，说‘我们平安无事’，为了要行这一切可憎的事呢？
JER|7|11|这称为我名下的殿在你们眼中岂可看为贼窝呢？看哪，我真的都看见了。这是耶和华说的。
JER|7|12|你们到我的地方 示罗 去，就是我先前在那里立为我名的居所，察看我因这百姓 以色列 的罪恶向那地方所行的事。
JER|7|13|现在，因你们行了这一切的事，我一再警戒你们，你们却不听从；我呼唤你们，你们也不回应。这是耶和华说的。
JER|7|14|所以我要向这称为我名下、你们所倚靠的殿，与我所赐给你们和你们祖先的地这样行，正如我从前向 示罗 所行的。
JER|7|15|我必将你们从我眼前赶出，正如赶出你们的众弟兄，就是所有 以法莲 的后裔。”
JER|7|16|“所以，你不要为这百姓祈祷；不要为他们呼求祷告，也不要为他们向我祈求，因我不听你。
JER|7|17|他们在 犹大 城镇和 耶路撒冷 街上所做的，你难道没有看见吗？
JER|7|18|孩子捡柴，父亲烧火，妇女揉面做饼，献给天后，又向别神献浇酒祭，惹我发怒。
JER|7|19|他们岂是惹我发怒呢？不是自己惹祸，以致脸上惭愧吗？这是耶和华说的。
JER|7|20|所以主耶和华如此说：看哪，我必将我的怒气和愤怒倾倒在这地方的人和牲畜身上、田野的树木和地里的出产上，它必燃烧，不会熄灭。”
JER|7|21|万军之耶和华－ 以色列 的上帝如此说：“你们要将燔祭加在你们的祭物上，又要吃肉；
JER|7|22|因为我将你们祖先从 埃及 地领出来的那日，燔祭和祭物的事我并没有提说，也没有吩咐他们。
JER|7|23|我只吩咐他们这一件事说：‘你们当听从我的话，我就作你们的上帝，你们也作我的子民。你们行走我所吩咐的一切道路，就可以得福。’
JER|7|24|他们却不听从，也不侧耳而听，竟随从自己的计谋和顽梗的恶心去行，不进反退。
JER|7|25|自从你们祖先出 埃及 地的那日，直到今日，我每日一再差遣我的仆人众先知到你们那里去。
JER|7|26|你们却不听我，不侧耳而听，竟硬着颈项行恶，比你们的祖先更甚。
JER|7|27|“你要将这一切的话告诉他们，他们却不听你；呼唤他们，他们却不回应。
JER|7|28|你要对他们说：‘这就是不听从耶和华－他们上帝的话、不领受训诲的国民；诚信已从他们口中消失殆尽了。
JER|7|29|耶路撒冷 啊，要剪头发，扔掉它， 在光秃的高地唱哀歌， 因为耶和华弃绝、离弃了惹他发怒的世代。’”
JER|7|30|“ 犹大 人行我眼中看为恶的事，将可憎之偶像立在称为我名下的殿里，玷污这殿。这是耶和华说的。
JER|7|31|他们在 欣嫩子谷 建造 陀斐特 的丘坛，要在火中焚烧自己的儿女。这并不是我所吩咐的，我心里也从来没有想过。
JER|7|32|因此，看哪，日子将到，这地方不再称为 陀斐特 和 欣嫩子谷 ，反倒称为 杀戮谷 。他们要在 陀斐特 埋葬尸首，甚至无处可葬。这是耶和华说的。
JER|7|33|并且这百姓的尸首要给空中的飞鸟和地上的走兽作食物，无人吓走它们。
JER|7|34|那时，我必止息 犹大 城镇和 耶路撒冷 街上欢喜和快乐的声音、新郎和新娘的声音，因为这地必然荒芜。”
JER|8|1|耶和华说：“那时，人必将 犹大 诸王和领袖的骸骨、祭司和先知的骸骨，以及 耶路撒冷 居民的骸骨，都从坟墓中取出来，
JER|8|2|散布在太阳、月亮和天上众星之下，就是他们从前所喜爱、所事奉、所随从、所求问、所敬拜的。这些骸骨不被收殓，不被埋葬，必在地面上成为粪土。
JER|8|3|这邪恶家族所幸存的余民，就是在我赶他们到的各处所剩下的 ，全都宁可选死不选活。这是万军之耶和华说的。”
JER|8|4|“你要对他们说，耶和华如此说： 人跌倒，不再起来吗？ 人转去，不再转回来吗？
JER|8|5|这 耶路撒冷 的百姓为何永久背道呢？ 他们抓住诡诈，不肯回头。
JER|8|6|我留心听，听见他们说不诚实的话。 无人懊悔自己的恶行，说： ‘我做的是什么呢？’ 他们全都转奔己路， 如马直闯战场。
JER|8|7|空中的鹳鸟知道自己的季节， 斑鸠、燕子与白鹤也守候当来的时令； 我的百姓却不知道耶和华的法则。
JER|8|8|“你们怎么说：‘我们有智慧， 耶和华的律法在我们这里’？ 看哪，其实文士的假笔舞弄虚假。
JER|8|9|智慧人惭愧，惊惶，被擒拿； 看哪，他们背弃耶和华的话， 还会有什么智慧呢？
JER|8|10|因此，我必将他们的妻子给别人， 将他们的田地给别人为业； 因为他们从最小的到最大的都贪图不义之财， 从先知到祭司全都行事虚假。
JER|8|11|他们轻忽地医治我百姓的损伤，说： ‘平安了！平安了！’ 其实没有平安。
JER|8|12|他们行可憎之事，应当羞愧； 然而他们却一点也不觉得羞愧， 又不知羞耻。 因此，他们必与仆倒的人一样仆倒； 我惩罚他们的时候， 他们必跌倒。 这是耶和华说的。
JER|8|13|我必使他们全然灭绝； 葡萄树上必没有葡萄 ， 无花果树上没有果子， 叶子也必枯干。 我所赐给他们的， 必离他们而去。 这是耶和华说的。”
JER|8|14|我们为何静坐不动呢？ 我们当聚集，进入坚固城， 在那里静默不言； 因为耶和华－我们的上帝使我们静默不言， 又将苦水给我们喝， 都因我们得罪了耶和华。
JER|8|15|我们指望平安， 却得不着福气； 指望痊愈的时刻， 看哪，受了惊惶。
JER|8|16|“从 但 那里传来敌人的马喷气的声音， 壮马发出嘶声， 全地就都震动； 因为他们来吞灭这地和其上所有的， 吞灭这城与其中的居民。
JER|8|17|看哪，我必派蛇进到你们中间， 就是法术无法驱除的毒蛇， 它们必咬你们。 这是耶和华说的。”
JER|8|18|忧愁时我寻找安慰 ， 我心在我里面发昏。
JER|8|19|听啊，是我百姓呼救的声音从远地传来： “耶和华不是在 锡安 吗？ 锡安 的王不是在其中吗？” “他们为什么以自己雕刻的偶像 和外邦虚无的神明 惹我发怒呢？”
JER|8|20|“秋收已过，夏季已完， 我们还未得救！”
JER|8|21|因我百姓的损伤， 我也受了损伤。 我哀恸，惊惶将我抓住。
JER|8|22|在 基列 岂没有乳香呢？ 在那里岂没有医生呢？ 我百姓 为何得不着医治呢？
JER|9|1|但愿我的头为水， 我的眼为泪水的泉源， 我好为我百姓 中被杀的人昼夜哭泣。
JER|9|2|惟愿在旷野有旅客的客栈， 我好离开我的百姓而去； 因他们全都行奸淫， 是行诡诈的一党。
JER|9|3|他们弯起舌头像弓， 为要说谎话； 他们在国中增长势力， 不是为诚信。 他们恶上加恶， 并不认识我。 这是耶和华说的。
JER|9|4|你们各人当谨防邻舍， 不可信赖弟兄； 因为弟兄尽行欺骗， 邻舍也都往来毁谤人。
JER|9|5|他们互相欺骗， 不说真话， 训练自己的舌头说谎， 竭尽所能地作恶。
JER|9|6|你居住在诡诈的人中； 他们因行诡诈 ，不愿意认识我。 这是耶和华说的。
JER|9|7|所以万军之耶和华如此说： “看哪，我要熬炼他们，考验他们； 不然，为了我的百姓 ，我该如何行呢？
JER|9|8|他们的舌头是毒箭，说话诡诈， 跟邻舍口说平安， 心却谋害他。
JER|9|9|我岂不因这些事向他们施行惩罚吗？ 像这样的国家，我岂能不报复呢？ 这是耶和华说的。”
JER|9|10|我要为山岭哭泣悲哀， 为旷野的草场扬声哀号； 因为都已枯焦，甚至无人经过。 牲畜的鸣叫听不见， 空中的飞鸟和地上的走兽也都逃离。
JER|9|11|我必使 耶路撒冷 成为废墟，为野狗的住处， 也必使 犹大 的城镇荒废，无人居住。
JER|9|12|谁是智慧人，可以明白这事？耶和华的口可向谁述说，使他传讲呢？这地为何毁灭，枯焦如旷野，无人经过呢？
JER|9|13|耶和华说：“因为这百姓离弃我在他们面前所设立的律法，不听从我的话，不肯遵行，
JER|9|14|反随从自己顽梗的心行事，照他们祖先所教训的随从诸 巴力 。”
JER|9|15|所以万军之耶和华－ 以色列 的上帝如此说：“看哪，我必将茵蔯给这百姓吃，又用苦水给他们喝。
JER|9|16|我要把他们分散在他们和他们祖宗所不认识的列国；我也要使刀剑追杀他们，直到将他们灭尽。”
JER|9|17|万军之耶和华如此说： “你们要考虑， 将唱哀歌的妇女召来， 差人召善哭的妇女前来，
JER|9|18|叫她们速速为我们举哀， 使我们泪眼汪汪， 使我们的眼皮涌出泪水。
JER|9|19|因为有哀声从 锡安 传来： ‘我们竟然败落！ 我们何等惭愧！ 我们撇下土地， 人拆毁了我们的房屋。’”
JER|9|20|妇女们哪，当听耶和华的话， 领受他口中的言语； 当教导你们的女儿举哀， 各人教导女伴唱哀歌。
JER|9|21|因为死亡从窗户进来， 进入我们的宫殿， 从外边剪除孩童， 从街上剪除少年。
JER|9|22|你当说，耶和华如此说： 人的尸首必倒在田野像粪土， 又像收割的人身后遗落的禾稼， 无人拾取。
JER|9|23|耶和华如此说：“智慧人不要因他的智慧夸口，勇士不要因他的力气夸口，财主也不要因他的财富夸口；
JER|9|24|夸口的却要夸自己有聪明，认识我是耶和华，知道我喜悦在世上施行慈爱、公平和公义。这是耶和华说的。
JER|9|25|“看哪，日子将到，这是耶和华说的，我要惩罚只在肉身受割礼的人，
JER|9|26|就是 埃及 、 犹大 、 以东 、 亚扪 人、 摩押 人，和住旷野所有剃鬓发的人；因为列国都未受割礼， 以色列 全家心中也未受割礼。”
JER|10|1|以色列 家啊，要听耶和华对你们所说的话，
JER|10|2|耶和华如此说： “不要效法列国的行为， 任凭列国因天象惊惶， 你们不要惊惶。
JER|10|3|万民的习俗是虚空的； 偶像 不过是从树林中砍来的木头， 是匠人用斧头做成的手工。
JER|10|4|人用金银妆饰它， 用钉子和锤子钉稳， 使它不动摇。
JER|10|5|偶像好像瓜田里的稻草人， 不能说话，不能行走， 必须有人抬着。 不要怕它们， 因它们不能降祸， 也无力降福。”
JER|10|6|耶和华啊，没有谁能与你相比！ 你本为大，你的名也大有能力。
JER|10|7|万国的王啊，谁不敬畏你？ 敬畏你本是合宜的； 列国所有的智慧人中， 在他们一切的国度里， 都没有能与你相比的。
JER|10|8|他们如同畜牲，尽都愚昧。 偶像的训诲算什么呢？ 偶像不过是木头，
JER|10|9|锤炼的银片是从 他施 来的， 金子则从 乌法 而来， 都是匠人和银匠的手工； 又有蓝色和紫色的衣服， 全都是巧匠的作品。
JER|10|10|惟耶和华是真上帝， 是活的上帝，是永远的王。 他一发怒，大地震动； 他一恼恨，列国担当不起。
JER|10|11|你们要对他们这样说：“那些不是创造天地的神明，必从地上、从天下被除灭！”
JER|10|12|耶和华以能力创造大地， 以智慧建立世界， 以聪明铺张穹苍。
JER|10|13|他一出声，天上就有众水澎湃； 他使云雾从地极上腾， 造电随雨而闪， 从仓库中吹出风来。
JER|10|14|人人都如同畜牲，毫无知识； 银匠都因偶像羞愧， 他所铸的偶像本是虚假， 它们里面并无气息。
JER|10|15|偶像都是虚无的， 是迷惑人的作品， 到受罚的时刻必被除灭。
JER|10|16|雅各 所得的福分不是这样， 因主 是那创造万有的， 以色列 是他产业的支派， 万军之耶和华是他的名。
JER|10|17|受围困的居民哪，当收拾你的行囊， 离开这地。
JER|10|18|因为耶和华如此说： “看哪，这一次，我必将此地的居民抛出去， 又必加害他们， 使他们觉悟 。”
JER|10|19|祸哉！我受损伤， 我的伤痕极其重大。 我却说：“这真的是我必须忍受的痛苦。”
JER|10|20|我的帐棚毁坏， 我的绳索折断， 我的儿女都离我而去，不在了。 再无人来支搭我的帐棚，挂起我的幔子。
JER|10|21|因为牧人如同畜牲， 没有寻求耶和华， 所以不得顺利； 他们的羊群也都分散了。
JER|10|22|有风声！看哪，来了！ 有大扰乱从北方而来， 要使 犹大 的城镇变为废墟， 成为野狗的住处。
JER|10|23|耶和华啊，我知道人的道路不由自己， 行路的人也不能定自己的脚步。
JER|10|24|耶和华啊，求你按公平管教我， 不要在你的怒中惩治我， 免得你使我归于无有。
JER|10|25|求你将愤怒倾倒在不认识你的列国中， 倾倒在不求告你名的各族上； 因为他们吞了 雅各 ，不但吞吃，而且灭绝， 使他的住处变为荒凉。
JER|11|1|耶和华的话临到 耶利米 ，说：
JER|11|2|“当听这约的话，告诉 犹大 人和 耶路撒冷 的居民，
JER|11|3|对他们说，耶和华－ 以色列 的上帝如此说：‘不听从这约之话的人必受诅咒。
JER|11|4|这约是我将你们祖先从 埃及 地领出来，脱离铁炉的那日所吩咐他们的，说：你们要听从我的话，照我所吩咐的一切去做。这样，你们作我的子民，我也作你们的上帝，
JER|11|5|我好坚定我向你们列祖所起的誓，赏赐他们流奶与蜜之地，正如今日一样。’”我就回应说：“耶和华啊，阿们！”
JER|11|6|耶和华对我说：“你要在 犹大 城镇和 耶路撒冷 街市宣告这一切话，说：‘当听从遵行这约的话，
JER|11|7|因为我将你们祖先从 埃及 地领出来的那日，直到今日，都一再切切告诫他们说：当听从我的话。
JER|11|8|他们却不听从，也不侧耳而听，竟随从自己顽梗的恶心去行。我就使这约中一切诅咒的话临到他们身上；这约是我吩咐他们遵行的，他们却不遵行。’”
JER|11|9|耶和华对我说：“在 犹大 人和 耶路撒冷 居民中有同谋背叛的事。
JER|11|10|他们转去效法他们祖先的恶行，不肯听我的话，竟随从别神，事奉它们。 以色列 家和 犹大 家违背了我与他们列祖所立的约。
JER|11|11|所以耶和华如此说：看哪，我必使灾祸临到他们，是他们不能逃脱的。他们向我哀求，我却不听。
JER|11|12|那时， 犹大 城镇的人和 耶路撒冷 的居民要哀求他们烧香所供奉的神明；只是遭难的时候，这些神明一点也不能拯救他们。
JER|11|13|犹大 啊，你神明的数目与你城镇的数目相等；你所筑可耻的坛，就是向 巴力 烧香的坛 ，也与 耶路撒冷 街道的数目相等。
JER|11|14|“所以你不要为这百姓祈祷，也不要为他们呼求祷告，因为他们遭难向我哀求的时候，我必不应允。
JER|11|15|我所亲爱的既多设恶谋，还能在我殿中做什么呢？你因作恶就喜乐，圣肉要离开你。
JER|11|16|从前耶和华给你起名叫青橄榄树，又华美又结好果子；如今他用一声巨响点火在其上，枝子就折断了。
JER|11|17|“原来栽培你的万军之耶和华已经说要降祸给你，是因 以色列 家和 犹大 家行恶。他们向 巴力 烧香，惹我发怒，是自作自受。”
JER|11|18|耶和华指示我，我才知道； 你将他们所做的给我指明。
JER|11|19|我像柔顺的羔羊被牵去宰杀， 并不知道他们设计谋害我： “我们把树连果子都灭了吧！ 把他从活人之地剪除， 使他的名不再被记得。”
JER|11|20|按公义判断、察验人肺腑心肠的万军之耶和华啊， 求你使我得见你在他们身上报仇， 因我已将我的案件向你禀明了。
JER|11|21|所以，耶和华论到寻索你命的 亚拿突 人如此说：“他们说：你不要奉耶和华的名说预言，免得你死在我们手中。
JER|11|22|所以万军之耶和华如此说：看哪，我必惩罚他们；他们的壮丁必被刀剑杀死，他们的儿女必因饥荒而死，
JER|11|23|他们当中必无任何幸存者；因为在他们受罚之年，我必使灾祸临到 亚拿突 人。”
JER|12|1|耶和华啊，我与你争辩的时候， 你总是显为义； 但有一件，我还要与你理论： 恶人的道路为何亨通呢？ 大行诡诈的为何得安逸呢？
JER|12|2|你栽培了他们， 他们也扎了根， 长大，而且结果。 他们的口与你相近， 心却与你远离。
JER|12|3|耶和华啊，你认识我，看见我， 你察验我向你的心如何。 求你将他们拉出来， 如将宰的羊， 为杀戮的日子分别出来。
JER|12|4|这地悲哀， 一切田野的青草枯干要到几时呢？ 因其上居民的恶行， 牲畜和飞鸟都灭绝了。 因为他们说：“他看不见 我们的结局 。”
JER|12|5|“你与步行的人同跑， 尚且觉得累， 怎能与马赛跑呢？ 你在安全之地尚且会跌倒 ， 在 约旦河 边的丛林要怎么办呢？
JER|12|6|因为连你兄弟和你父家都以诡诈待你， 甚至在你后边大声喊叫。 虽然他们向你说好话， 你也不要相信他们。”
JER|12|7|我离弃了我的殿宇， 撇弃了我的产业， 将我心里所亲爱的交在她 仇敌手中。
JER|12|8|我的产业向我如林中的狮子， 出声攻击我， 因此我恨恶她。
JER|12|9|我的产业向我如斑点的鸷鸟， 有鸷鸟在四围攻击她。 你们去聚集田野的百兽， 叫它们来吞吃吧！
JER|12|10|许多牧人毁坏我的葡萄园， 践踏我的地产， 使我美好的地产变为荒凉的旷野。
JER|12|11|他们使地荒凉； 地既荒凉，就向我哀哭。 全地荒凉，却无人在意。
JER|12|12|灭命的来到旷野中一切光秃的高地； 耶和华的刀从地这边直到地那边，尽行杀灭， 凡血肉之躯都不得平安。
JER|12|13|他们种的是麦子， 收的却是荆棘； 辛辛苦苦却无收获。 因耶和华的烈怒， 你们必为自己的收成感到羞愧。
JER|12|14|耶和华如此说：“看哪，我要将所有的恶邻拔出本地，他们曾占据了我赐给 以色列 百姓所承受的产业；我也要将 犹大 家从他们中间拔出来。
JER|12|15|我拔出他们以后，必回转过来怜悯他们，使他们归回，各归本业，各归故土。
JER|12|16|他们若殷勤学习我百姓的道，指着我的名起誓：‘我指着永生的耶和华起誓’，正如他们从前教我百姓指着 巴力 起誓，他们必在我百姓中得以建立。
JER|12|17|他们若是不听，我必拔出那国，不但拔出，还要毁灭。这是耶和华说的。”
JER|13|1|耶和华对我如此说：“你去买一条麻布带子，束在你腰上，不可把它泡在水里。”
JER|13|2|我就照耶和华的话，买了一条带子，束在我的腰上。
JER|13|3|耶和华的话第二次临到我，说：
JER|13|4|“要拿你所买、在你腰上的带子，起来往 幼发拉底河 去，把腰带藏在那里的磐石穴中。”
JER|13|5|我就去，照着耶和华命令我的，把腰带藏在 幼发拉底河 边。
JER|13|6|过了多日，耶和华对我说：“你起来往 幼发拉底河 去，把我命令你藏在那里的腰带取出来。”
JER|13|7|我就往 幼发拉底河 去，把那腰带从我所藏的地方挖出来。看哪，腰带已经破烂，毫无用处了。
JER|13|8|耶和华的话临到我，说：
JER|13|9|“耶和华如此说：我要照样败坏 犹大 的骄傲和 耶路撒冷 的狂傲。
JER|13|10|这恶民不肯听我的话，按自己顽梗的心而行，随从别神，事奉敬拜它们；这恶民必像这腰带，毫无用处。
JER|13|11|腰带怎样紧贴人的腰，照样，我也曾使 以色列 全家和 犹大 全家紧贴着我，归我为子民，使我得名声，得颂赞，得荣耀；他们却不肯听从。这是耶和华说的。”
JER|13|12|“所以你要对他们说：‘耶和华－ 以色列 的上帝如此说：各坛都要装满酒。’他们必对你说：‘我们岂不知道各坛都要装满酒吗？’
JER|13|13|你就对他们说：‘耶和华如此说：看哪，我必使这地所有的居民，就是坐 大卫 宝座的君王、祭司和先知，并 耶路撒冷 所有的居民，都酩酊大醉。
JER|13|14|我要使他们彼此冲突，连父与子也互相冲突；我必不可怜，不顾惜，不怜悯，以致将他们灭绝。这是耶和华说的。’”
JER|13|15|你们当听，当侧耳而听； 不可骄傲，因为耶和华已经吩咐了。
JER|13|16|当耶和华－你们的上帝 尚未使黑暗来临， 在昏暗的山上 你们的脚未绊跌以前， 要将荣耀归给他。 你们盼望光明， 他却使光明变为死荫， 成为幽暗。
JER|13|17|你们若不听这话， 我的心必因你们的骄傲暗自哭泣； 我的眼必痛哭流泪， 因为耶和华的羊群被掳去了。
JER|13|18|你要对君王和太后说： “你们当自卑，坐下； 因你们的王冠， 就是你们华美的冠冕已经掉落了 。”
JER|13|19|尼革夫 的城镇都被关闭， 无人打开； 犹大 全被掳掠， 掳掠净尽。
JER|13|20|你们要举目观看从北方来的人。 先前赐给你的羊群， 就是你所引以为荣的羊， 现今在哪里呢？
JER|13|21|耶和华立你自己所教导的盟友， 立他们为头来辖制你， 你还有什么话可说呢？ 痛苦岂不将你抓住像临产的妇人吗？
JER|13|22|你若心里说：“这一切的事为何临到我呢？” 是因你罪孽甚多。 你的下摆揭起， 你的脚跟受伤。
JER|13|23|古实 人岂能改变皮肤呢？ 豹岂能改变斑点呢？ 若能，你们这善于行恶的便能行善了。
JER|13|24|我必吹散他们， 如碎秸随旷野的风飘动。
JER|13|25|这是你所当得的， 是我量给你的报应 ； 因为你忘记了我， 倚靠虚假 。 这是耶和华说的。
JER|13|26|我要揭起你的下摆， 蒙在你脸上， 显露你的羞耻。
JER|13|27|你在田野的山上行奸淫， 发嘶声，谋淫乱， 这些可憎之事我都看见了。 耶路撒冷 啊，你有祸了！ 你不肯洁净 还要等到几时呢？
JER|14|1|耶和华的话临到 耶利米 ，论到旱灾的事：
JER|14|2|“ 犹大 悲哀，城门衰败； 众人坐在地上哀恸， 耶路撒冷 的哀声上达。
JER|14|3|他们的贵族打发童仆去打水； 他们来到水池， 找不到水，就拿着空器皿， 蒙羞惭愧，抱头而回。
JER|14|4|因为无雨降在地上，土地就干裂， 农夫为此蒙羞抱头。
JER|14|5|田野的母鹿因为无草 也撇弃才生的小鹿。
JER|14|6|野驴站在光秃的高地喘气，好像野狗； 它们的眼目因无草而失明。”
JER|14|7|耶和华啊，虽然我们的罪孽控告我们， 求你为你名的缘故行动吧！ 我们本是多次背道，得罪了你。
JER|14|8|以色列 所盼望，在患难时作他救主的啊， 你在这地为何像寄居的， 又如旅行的只住一夜呢？
JER|14|9|你为何像受惊吓的人， 像不能救人的勇士呢？ 耶和华啊，你在我们中间， 我们是称为你名下的人， 求你不要离开我们。
JER|14|10|耶和华论到这百姓如此说： “这百姓喜爱游荡， 不约束自己的脚步， 所以耶和华不悦纳他们。 现今他要记起他们的罪孽， 惩罚他们的罪恶。”
JER|14|11|耶和华又对我说：“不要为这百姓求福。
JER|14|12|他们禁食的时候，我不听他们的呼求；他们献燔祭和素祭，我也不悦纳。我却要用刀剑、饥荒、瘟疫灭绝他们。”
JER|14|13|我就说：“唉！主耶和华，看哪，那些先知常对他们说：‘你们必不见刀剑，也不遭饥荒；耶和华要在这地方赏赐你们真正的平安。’”
JER|14|14|耶和华对我说：“那些先知托我的名说假预言，我并未差遣他们，没有吩咐他们，也没有对他们说话；他们向你们预言的是虚假的异象、占卜、虚无，以及心中的诡诈。
JER|14|15|所以耶和华如此说：‘论到托我名说预言的那些先知，我并未差遣他们；他们说这地不会有刀剑、饥荒，其实那些先知自己必被刀剑、饥荒灭绝。
JER|14|16|听他们说预言的百姓必因饥荒、刀剑被扔在 耶路撒冷 的街道上，无人埋葬。他们连妻子带儿女，都是如此。我必将他们的恶倒在他们身上。’”
JER|14|17|你要向他们说这些话： 愿我眼泪汪汪， 昼夜不息， 因为少女─我百姓 受了重大的打击， 伤口极其严重。
JER|14|18|我若出到田间， 看哪，有被刀杀的； 我若进入城内， 看哪，有因饥荒患病的； 先知和祭司也在各地往来经商， 不知如何是好。
JER|14|19|你全然弃绝 犹大 吗？ 你的心厌恶 锡安 吗？ 你为何击打我们，使我们无法得医治呢？ 我们指望平安，却得不着福气； 指望痊愈，看哪，受了惊惶。
JER|14|20|耶和华啊，我们承认自己的罪恶 和我们祖先的罪孽， 因我们得罪了你。
JER|14|21|求你为你名的缘故， 不厌恶，不轻视你荣耀的宝座。 求你记念， 不要违背你与我们所立的约。
JER|14|22|外邦虚无的神明 中有能降雨的吗？ 天能自降甘霖吗？ 耶和华－我们的上帝啊，不是你吗？ 我们要等候你， 因为这一切都是你所造的。
JER|15|1|耶和华对我说：“虽有 摩西 和 撒母耳 站在我面前，我的心也不顾惜这百姓。你把他们从我眼前赶出，叫他们出去吧！
JER|15|2|他们若问你说：‘我们往哪里去呢？’你就告诉他们，耶和华如此说： ‘定为死亡的，必致死亡； 定为刀杀的，必被刀杀； 定为饥荒的，必遭饥荒； 定为掳掠的，必被掳掠。’”
JER|15|3|“我命定四样灾害临到他们，就是刀剑杀戮、群狗拖拉、空中的飞鸟和地上的走兽吞吃毁灭。这是耶和华说的。
JER|15|4|我必使地上万国因他们而惊骇，都因 希西家 的儿子 犹大 王 玛拿西 在 耶路撒冷 所做的事。”
JER|15|5|耶路撒冷 啊，有谁同情你呢？ 有谁为你悲伤呢？ 有谁转身问你安呢？
JER|15|6|你弃绝了我， 转身退后； 因此我伸手攻击你，毁灭你， 我已怜悯到厌烦了。 这是耶和华说的。
JER|15|7|我在境内各关口 用簸箕筛我的百姓， 使他们丧掉儿女， 又毁灭他们， 他们仍不转离所行的道。
JER|15|8|他们的寡妇在我面前比海沙更多； 我使灭命者在正午来到， 攻击年轻人的母亲， 使痛苦惊吓忽然临到她身上。
JER|15|9|生过七个孩子的妇人衰弱； 尚在白昼，太阳忽然落下， 她就抱愧蒙羞。 我必当着敌人的面， 将他们当中的幸存者交给刀剑。 这是耶和华说的。
JER|15|10|我的母亲哪，我有祸了！因你生我作全地争相指控的人。我素来没有借贷给人，人也没有借贷给我，人人却都咒骂我。
JER|15|11|耶和华说：“我必定释放 你，使你得福气。灾祸苦难来临时，我必使仇敌央求你。
JER|15|12|人岂能将铜与铁，就是北方的铁折断呢？
JER|15|13|“我必因你在四境之内所犯的一切罪，将你的货物财宝当掠物，白白地交出来 。
JER|15|14|我要使你的仇敌过去，到你所不认识的地方 ，因为你们要被我怒中所起的火焚烧。”
JER|15|15|耶和华啊，你是知道的； 求你记念我，眷顾我， 向迫害我的人为我报仇； 不要把我取去，因你不轻易发怒， 要知道我为你的缘故受了凌辱。
JER|15|16|耶和华－万军之上帝啊， 我得着你的话就把它们吃了， 你的话是我心中的欢喜快乐； 因我是称为你名下的人。
JER|15|17|我并未坐在享乐人的会中欢乐； 因你的手，我就独自静坐， 你使我满心愤慨。
JER|15|18|我的痛苦为何长久不止呢？ 我的伤痕为何无法可医，不能痊愈呢？ 难道你以诡诈待我，像流干的河道吗？
JER|15|19|所以耶和华如此说：“你若回转， 我就使你归回， 站在我面前。 你若能将宝物和无用之物分别出来， 你就可以当作我的口。 他们必归向你， 你却不可归向他们。
JER|15|20|我必使你向这百姓成为坚固的铜墙。 他们必攻击你，却不能胜过你； 因我与你同在，要拯救你，搭救你。 这是耶和华说的。
JER|15|21|我必搭救你脱离恶人的手， 救赎你脱离残暴之人的手。”
JER|16|1|耶和华的话又临到我，说：
JER|16|2|“你不可在这地方娶妻，为自己生儿育女。
JER|16|3|因为论到在这地方所生的儿女，又论到在这国中生他们的父母，耶和华如此说：
JER|16|4|他们必死于致命的疾病，无人哀哭，不得埋葬，在地上如粪土，因刀剑和饥荒而灭绝；他们的尸首必给空中的飞鸟和地上的走兽作食物。
JER|16|5|“耶和华如此说：不要进入丧家，不要去哀哭，也不要为他们悲伤，因我已使我的平安、慈爱、怜悯离开这百姓。这是耶和华说的。
JER|16|6|他们连大带小，都必在这地死亡，不得埋葬。人必不为他们哀哭，不为他们割划自己，也不剃光头。
JER|16|7|有丧事，人不为他们擘饼 ，也不因死人安慰他们；他们丧父丧母，人也不给他们一杯酒安慰他们。
JER|16|8|你不可进入宴乐的家，与人同坐又吃又喝，
JER|16|9|因为万军之耶和华－ 以色列 的上帝如此说：看哪，你们还活着的日子，我必在你们眼前止息这地方欢喜和快乐的声音、新郎和新娘的声音。
JER|16|10|“你将这一切的话指示这百姓，他们若问你说：‘耶和华为什么说，要降这大灾祸攻击我们呢？我们有什么罪孽呢？我们向耶和华－我们的上帝犯了什么罪呢？’
JER|16|11|你就对他们说：‘因为你们祖先离弃了我，随从别神，事奉敬拜它们，却离弃我，不遵守我的律法。这是耶和华说的。
JER|16|12|你们行恶比你们祖先更甚，看哪，各人随从自己顽梗的恶心行事，不听从我。
JER|16|13|所以我必将你们从这地赶出，直赶到你们和你们祖先素不认识之地。你们在那里昼夜必事奉别神，因为我必不再向你们施恩。’”
JER|16|14|“看哪，日子将到，人必不再指着那领 以色列 人从 埃及 地上来的永生耶和华起誓。这是耶和华说的。
JER|16|15|人却要指着那领 以色列 人离开北方之地，离开他们被赶到的各国之永生的耶和华起誓；并且我要领他们归回我从前赐给他们祖先之地。”
JER|16|16|“看哪，我要差派许多打鱼的捕获他们；以后，我也要派许多打猎的，从各山上、各冈上、各石穴中猎取他们。这是耶和华说的。
JER|16|17|因我的眼目察看他们一切的行为；他们不能在我面前遮掩，他们的罪孽也不能在我眼前隐藏。
JER|16|18|我要先加倍报应他们的罪孽和罪恶，因为他们以可憎之偶像的尸首使我的地玷污，使我的产业充斥可厌之物。”
JER|16|19|耶和华啊，你是我的力量， 是我的保障， 在患难之日是我的避难所。 列国的人必从地极来到你这里，说： “我们祖先所承受的， 不过是虚假，是虚空无益之物。
JER|16|20|人岂可为自己制造神明呢？ 其实它们不是神明。”
JER|16|21|“所以，看哪，我要使他们知道，就是这一次使他们知道我的手和我的能力。他们就知道我的名是耶和华了。”
JER|17|1|犹大 的罪是用铁笔、用金刚石记录的，铭刻在他们的心版和祭坛角上。
JER|17|2|他们的儿女思念他们在高冈上、青翠树旁的祭坛和 亚舍拉 。
JER|17|3|我田野的山哪，因你在全境内的丘坛所犯的罪，我必使你的财富和一切的财宝成为掠物。
JER|17|4|因自己所做的 ，你必失去我所赐给你的产业。我也必使你在你所不认识的地服侍你的仇敌；因你们激起了我的怒火，直烧到永远。
JER|17|5|耶和华如此说： “倚靠人，以血肉为膀臂， 心中离弃耶和华的， 那人该受诅咒！
JER|17|6|他必像沙漠里的矮树， 不见福乐来到； 他要住在旷野干旱之处， 无人居住的盐地。
JER|17|7|倚靠耶和华、以耶和华为他所仰赖的， 那人有福了！
JER|17|8|他必像树栽于水旁， 在河边扎根， 炎热来到，毫不察觉 ， 叶子仍必青翠； 在干旱之年，一无挂虑， 并且结果不止。
JER|17|9|“人心比万物都诡诈， 坏到极处， 谁能识透呢？
JER|17|10|我－耶和华是鉴察人心，考验人肺腑的， 要按各人所行的和他做事的结果报应他。”
JER|17|11|那不按正道得财富的， 好像鹧鸪孵不是自己生的； 到了中年，财富必离开他， 终久他必成为愚顽人。
JER|17|12|我们的圣所是荣耀的宝座， 从太初就在高处。
JER|17|13|耶和华－ 以色列 的盼望啊， 凡离弃你的必蒙羞。 离我而去的， 他们必被写在地里， 因为他们离弃耶和华，这活水的泉源。
JER|17|14|耶和华啊，求你医治我，我就痊愈， 拯救我，我便得救； 因你是我所赞美的。
JER|17|15|看哪，他们对我说： “耶和华的话在哪里呢？ 让它应验吧！”
JER|17|16|至于我，我并没有逃避作牧人跟随你 ， 也没有想望那灾殃的日子； 这是你所知道的。 我嘴唇所出的都在你面前。
JER|17|17|不要使我因你惊恐； 灾祸来临时，你是我的避难所。
JER|17|18|愿那些迫害我的蒙羞， 却不要使我蒙羞； 使他们惊惶， 却不要使我惊惶； 愿灾祸的日子临到他们， 以加倍的毁坏毁坏他们。
JER|17|19|耶和华对我如此说：“你去站在 犹大 君王出入的 平民门 ，和 耶路撒冷 的各城门口，
JER|17|20|对他们说：‘你们这 犹大 君王、 犹大 众人和 耶路撒冷 所有的居民，凡从这些城门进入的，都当听耶和华的话。
JER|17|21|耶和华如此说：你们要谨慎，不可在安息日挑什么担子进入 耶路撒冷 的城门，
JER|17|22|也不可在安息日从家中挑担子出去。无论何工都不可做，只要以安息日为圣日，正如我所吩咐你们祖先的。’
JER|17|23|他们却不听从，也不侧耳而听，竟硬着颈项不听，不肯领受训诲。
JER|17|24|“你们若留意听从我，在安息日不挑什么担子进入这城的各门，只以安息日为圣日，在那日不做任何工作，这是耶和华说的，
JER|17|25|就必有坐 大卫 宝座的君王和领袖，与 犹大 人，并 耶路撒冷 的居民，或坐车，或骑马，进入这城的各门，而且这城必存到永远。
JER|17|26|也必有人从 犹大 城镇和 耶路撒冷 四围的各处，从 便雅悯 地、 谢非拉 、山区，并 尼革夫 而来，都带燔祭和祭物，素祭和乳香，并感谢祭，到耶和华的殿去。
JER|17|27|你们若不听从我，不以安息日为圣日，仍在安息日挑担子进入 耶路撒冷 的各城门，我必在城门中点火；这火必烧毁 耶路撒冷 的宫殿，不会熄灭。”
JER|18|1|耶和华的话临到 耶利米 ，说：
JER|18|2|“你起来，下到陶匠的家里去，在那里我要使你听见我的话。”
JER|18|3|我就下到陶匠的家里去，看哪，他在转盘上做器皿。
JER|18|4|陶匠用泥做的器皿在他手中做坏了，他就用它另做别的器皿，照他看为好的去做。
JER|18|5|耶和华的话临到我，说：
JER|18|6|“ 以色列 家啊，我待你们岂不能像这陶匠弄泥吗？ 以色列 家，看哪，泥在陶匠的手中怎样，你们在我的手中也怎样。这是耶和华说的。
JER|18|7|我何时论到一邦或一国说，要拔出、拆毁、毁坏；
JER|18|8|我所说的那一邦若回转离开他们的恶，我就改变心意，不将我想要施行的灾祸降与他们。
JER|18|9|我何时论到一邦或一国说，要建立、栽植；
JER|18|10|他们若行我眼中看为恶的事，不听从我的话，我就改变心意，不将我所说的福气赐给他们。
JER|18|11|现在你要对 犹大 人和 耶路撒冷 的居民说：‘耶和华如此说：看哪，我捏塑灾祸降给你们，定意惩罚你们。你们各人当回转离开所行的恶道，改正你们的所作所为。’
JER|18|12|“他们却说：‘没有用的，我们要照自己的计谋去行，各人要随自己顽梗的恶心行事。’”
JER|18|13|“所以，耶和华如此说： 你们且往各国访问， 有谁听见这样的事？ 少女 以色列 行了一件极恐怖的事。
JER|18|14|黎巴嫩 的雪岂能从田野 的磐石上融化呢？ 从远处 流下的凉水岂能干涸呢？
JER|18|15|我的百姓竟忘记我， 向那虚无的神明 烧香， 它们使百姓在所行的路上、在古道上绊跌， 去行未修筑的斜路，
JER|18|16|他们的地就变为荒凉， 长久被人嘲笑； 凡经过这地的必惊骇摇头。
JER|18|17|在仇敌面前，我必如东风刮散他们， 遭难的日子，我要以背向他们， 不以脸看他们。”
JER|18|18|他们说：“来吧！让我们设计谋害 耶利米 ；因为我们有祭司讲律法，有智慧人设谋略，有先知说预言，都未曾断绝。来吧！让我们用舌头攻击他，不要理他一切的话。”
JER|18|19|耶和华啊，求你留心听我， 且听那些指控我的人的话。
JER|18|20|人岂可以恶报善呢？ 他们竟挖坑要害我的性命！ 求你记念我站在你面前为他们说好话， 要使你的愤怒转离他们。
JER|18|21|因此，愿他们的儿女忍受饥荒， 愿他们死于刀剑之手； 愿他们的妻无子，且作寡妇， 愿他们的男人被死亡所灭， 他们的壮丁在阵上被刀击杀。
JER|18|22|你使敌军忽然临到他们的时候， 愿人听见哀声从他们的屋内发出； 因他们挖坑要捉拿我， 暗设罗网要绊我的脚。
JER|18|23|耶和华啊，他们要杀我的那一切计谋， 你都知道。 求你不要赦免他们的罪孽， 也不要从你面前涂去他们的罪恶。 愿他们在你面前跌倒， 愿你在发怒的时候对付他们。
JER|19|1|耶和华如此说：“你去买陶匠的瓷瓶 ，你和 百姓中的长老、位尊的祭司
JER|19|2|出去到 欣嫩子谷 、 哈珥西 的门口，在那里宣告我所吩咐你的话，
JER|19|3|说：‘ 犹大 君王和 耶路撒冷 的居民哪，当听耶和华的话。万军之耶和华－ 以色列 的上帝如此说：看哪，我必使灾祸临到这地方，凡听见的人都必耳鸣；
JER|19|4|因为他们和他们祖先，并 犹大 君王都离弃我，使这地方与我疏远 ，在这里向素不认识的别神烧香，又使这地方遍满无辜人的血。
JER|19|5|他们建造 巴力 的丘坛，要在火中焚烧自己的儿女，作为燔祭献给 巴力 。这不是我命令的，不是我吩咐的，我心里也从来没有想过。
JER|19|6|因此，看哪，日子将到，这地方不再称为 陀斐特 和 欣嫩子谷 ，反倒称为 杀戮谷 。这是耶和华说的。
JER|19|7|我要在这地方使 犹大 和 耶路撒冷 的计谋落空，也必使他们在仇敌面前倒在刀下，倒在寻索其命的人手下。我要把他们的尸首给空中的飞鸟和地上的走兽作食物。
JER|19|8|我必使这城令人惊骇嘲笑；凡路过的，必因这城所遭的灾难惊骇嘲笑。
JER|19|9|仇敌和寻索其命的人追逼他们，使他们落在围困窘迫之中，我必使他们各人吃自己儿女的肉和朋友的肉。’
JER|19|10|“你要在跟你同去的人眼前打碎那瓶，
JER|19|11|对他们说：‘万军之耶和华如此说：我要打碎这百姓和这城，正如人打碎陶匠的器皿，不能再使其完整。他们要在 陀斐特 埋葬，甚至无处可葬。
JER|19|12|我必向这地方和其中的居民如此行，使这城与 陀斐特 一样。这是耶和华说的。
JER|19|13|耶路撒冷 的房屋和 犹大 君王的宫殿，就是他们在其上向天上的万象烧香、向别神献浇酒祭的宫殿房屋，都必被玷污，和 陀斐特 一样。’”
JER|19|14|耶利米 从耶和华差他去说预言的 陀斐特 回来，站在耶和华殿的院中对众百姓说：
JER|19|15|“万军之耶和华－ 以色列 的上帝如此说：‘看哪，我必使我所说的一切灾祸临到这城和属它的城镇，因为他们硬着颈项不听我的话。’”
JER|20|1|音麦 的儿子 巴施户珥 祭司作耶和华殿的总管，听见 耶利米 预言这些事，
JER|20|2|就打 耶利米 先知，用耶和华殿里 上便雅悯门 内的枷锁，把他锁在那里。
JER|20|3|次日， 巴施户珥 开枷释放 耶利米 。于是 耶利米 对他说：“耶和华不叫你的名为 巴施户珥 ，而叫你 玛歌珥．米撒毕 ，
JER|20|4|因耶和华如此说：‘看哪，我要使你和你的众朋友惊吓；你们要亲眼看见他们倒在仇敌的刀下。我必将 犹大 人全都交在 巴比伦 王的手中，他要把他们掳到 巴比伦 去，用刀杀他们。
JER|20|5|我要将这城中一切的货财和劳碌得来的，并一切的珍宝，以及 犹大 君王所有的宝物，都交在仇敌手中。仇敌要抢夺他们，抓住他们，把他们带到 巴比伦 去。
JER|20|6|你， 巴施户珥 ，和所有住在你家中的人都必被掳；你和你的朋友，就是你向他们说假预言的，都要到 巴比伦 去，死在那里，葬在那里。’”
JER|20|7|耶和华啊，你欺哄了我， 我也被你欺哄了。 你比我强，并且得胜。 我终日成为笑柄， 人人都戏弄我。
JER|20|8|我每逢讲话的时候，就哀叹， 我喊叫：“有暴力和毁灭！” 因为耶和华的话终日成了我的凌辱和讥刺。
JER|20|9|我若说：“我不再提耶和华， 也不再奉他的名讲论”， 我心里便觉得 似乎有烧着的火闷在我骨中， 我忍受不住，不能自禁。
JER|20|10|我听见许多的毁谤， 四围都是惊吓； 连我知己朋友都看着我跌倒： “告他吧，我们要告他！ 或者他被引诱， 我们就能胜他， 在他身上报仇。”
JER|20|11|然而，耶和华与我同在， 好像可怕的勇士。 因此，迫害我的都绊跌， 不能得胜； 他们大大蒙羞， 由于行事没有智慧， 必永远受那不能忘怀的羞辱。
JER|20|12|考验义人、察看人肺腑心肠的万军之耶和华啊， 求你使我得见你在他们身上报仇， 因我已将我的案件向你禀明了。
JER|20|13|你们要向耶和华唱歌！ 要赞美耶和华！ 因他救了穷人的性命 脱离恶人的手。
JER|20|14|愿我出生的那日受诅咒！ 愿我母亲生我的那天不蒙福！
JER|20|15|报信给我父亲说 “你得了儿子”， 使我父亲甚欢喜的， 愿那人受诅咒。
JER|20|16|愿那人像耶和华所倾覆而不怜惜的城镇； 愿他早晨听见哀声， 中午听见呐喊；
JER|20|17|因他没有在我未出胎就把我杀了， 以致我母亲成为我的坟墓， 她却一直怀着胎 。
JER|20|18|我为何出胎见劳碌愁苦， 在羞愧中度尽我的年日呢？
JER|21|1|耶和华的话临到 耶利米 。那时， 西底家 王差派 玛基雅 的儿子 巴施户珥 和 玛西雅 的儿子 西番雅 祭司到他那里去，说：
JER|21|2|“请你为我们求问耶和华，因为 巴比伦 王 尼布甲尼撒 前来攻击我们；或者耶和华照他一切奇妙的作为待我们，使 巴比伦 王离开我们而去。”
JER|21|3|耶利米 对他们说：“你们当对 西底家 这样说：
JER|21|4|‘耶和华－ 以色列 的上帝如此说：看哪，我要使你们手中的兵器，就是你们与城外围困你们的 巴比伦 王和 迦勒底 人打仗所用的兵器转回来，把它们聚集在这城中。
JER|21|5|我要在怒气、愤怒和大恼怒中，用伸出来的手和大能的膀臂，亲自攻击你们；
JER|21|6|又要击打这城的居民，他们连人带牲畜都必遭遇大瘟疫而死亡。
JER|21|7|以后，我要将 犹大 王 西底家 和他的臣仆百姓，就是在城内，从瘟疫、刀剑、饥荒中幸存的人，都交在 巴比伦 王 尼布甲尼撒 手中，交在仇敌和寻索其命的人手中。 巴比伦 王必用刀击杀他们，不顾惜，不同情，不怜悯。这是耶和华说的。’
JER|21|8|“你要对这百姓说：‘耶和华如此说：看哪，我将生命的路和死亡的路摆在你们面前。
JER|21|9|住在这城里的必遭刀剑、饥荒、瘟疫而死；但出去投降围困你们之 迦勒底 人的必得存活，保全自己的性命。
JER|21|10|我向这城板脸，降祸不降福；这城必交在 巴比伦 王的手中，他必用火焚烧。这是耶和华说的。’”
JER|21|11|“至于 犹大 王的家，你们当听耶和华的话。
JER|21|12|大卫 家啊，耶和华如此说： ‘每早晨你们要施行公平， 拯救被抢夺的脱离欺压者的手， 免得我的愤怒因你们的恶行发作， 如火燃起，无人能熄灭。’
JER|21|13|住在山谷和平原磐石上的居民啊， 看哪，我与你们为敌， 因为你们说：‘谁能下来攻击我们？ 谁能进入我们的住处呢？’ 这是耶和华说的。
JER|21|14|我必按你们行事的结果惩罚你们， 也必使火在 耶路撒冷 的林中燃起， 将四围所有的尽行烧灭。 这是耶和华说的。”
JER|22|1|耶和华如此说：“你要下到 犹大 王的宫中，在那里说这话，
JER|22|2|你要说：‘坐 大卫 宝座的 犹大 王啊，你和你的臣仆，并进入这些城门的百姓，都当听耶和华的话。
JER|22|3|耶和华如此说：你们要施行公平和公义，拯救被抢夺的脱离欺压者的手，不可亏负寄居的和孤儿寡妇，不可用残暴对待他们，也不可在这地方流无辜人的血。
JER|22|4|你们若切实遵行这话，就必有坐 大卫 宝座的君王和他的臣仆百姓，或坐车或骑马，从这王宫的各门进入。
JER|22|5|你们若不听这些话，我指着自己起誓，这王宫必变为废墟。这是耶和华说的。’
JER|22|6|耶和华论到 犹大 王的家如此说： “我看你如 基列 ， 如 黎巴嫩 的山顶； 然而，我必使你变为旷野， 成为无人居住的城镇。
JER|22|7|我要预备施行毁灭的人， 各人佩带兵器攻击你； 他们要砍伐你佳美的香柏树， 扔在火中。
JER|22|8|“许多国的百姓经过这城，就彼此谈论说：‘耶和华为何向这大城这样做呢？’
JER|22|9|必有人回答说：‘是因他们离弃了耶和华－他们上帝的约，事奉敬拜别神。’”
JER|22|10|不要为已死的人哀哭， 也不要为他悲伤， 却要为离家外出的人大大哀哭； 因为他不再回来见自己的出生地。
JER|22|11|因为论到离开这地方的 约西亚 之子 犹大 王 沙龙 ，就是接续他父亲 约西亚 作王的，耶和华这样说：“他必不再回到这里来，
JER|22|12|却要死在被掳去的地方，必不得再见这地。”
JER|22|13|祸哉！那以不公义盖房，以不公平造楼， 白白使邻舍做工，却不给工钱的人，
JER|22|14|他说：“我要为自己盖宽敞的房，盖高大的楼。” 他为它开窗户， 以香柏木为墙板， 漆上丹红色。
JER|22|15|难道你作王就是要盖香柏木楼房争胜的吗？ 你的父亲岂不是也吃也喝， 也施行公平和公义吗？ 那时他得了福乐。
JER|22|16|他为困苦和贫穷的人伸冤， 那时就得了福乐。 认识我不就在此吗？ 这是耶和华说的。
JER|22|17|你的眼和你的心却专顾不义之财， 流无辜人的血， 行欺压和残暴。
JER|22|18|所以，耶和华论到 约西亚 的儿子 犹大 王 约雅敬 如此说： 人必不为他举哀： “哀哉，我的哥哥！ 哀哉，我的姊姊！” 也不为他举哀： “哀哉，我的主！ 哀哉，我主的荣华！”
JER|22|19|他被埋葬好像埋驴子一样， 被拖出去，扔在 耶路撒冷 城门外。
JER|22|20|你要上 黎巴嫩 哀号， 在 巴珊 扬声， 从 亚巴琳 哀号， 因为你所亲爱的都毁灭了。
JER|22|21|你兴盛的时候，我对你说话； 你却说：“我不听。” 你从年轻时就是这样， 不肯听我的话。
JER|22|22|你的牧人要被风吞吃， 你所亲爱的必被掳去； 那时你必因你一切的恶行抱愧蒙羞。
JER|22|23|你这住 黎巴嫩 、在香柏树上搭窝的， 有痛苦临到你， 如疼痛临到临产的妇人， 那时你何等可怜 ！
JER|22|24|耶和华说：“ 约雅敬 的儿子 犹大 王 哥尼雅 ，虽是我右手上带印的戒指，我凭我的永生起誓，我必将你从其上摘下来。
JER|22|25|我要将你交在寻索你命的人和你所惧怕的人手中，就是 巴比伦 王 尼布甲尼撒 和 迦勒底 人手中。
JER|22|26|我也要将你和生你的母亲赶到别国，不是你们出生的地方；你们必死在那里，
JER|22|27|心中虽然很想归回那地，却不得归回。”
JER|22|28|哥尼雅 这人是被轻看、遭毁坏的罐子， 是无人喜爱的器皿吗？ 他和他的后裔为何被赶到素不认识之地呢？
JER|22|29|地啊，地啊，地啊，当听耶和华的话！
JER|22|30|耶和华如此说： “要把这人登记为无子， 是平生不得亨通的人； 因为他后裔中再无一人得亨通， 能坐在 大卫 的宝座上治理 犹大 。”
JER|23|1|耶和华说：“祸哉！那些残害、赶散我草场之羊的牧人！”
JER|23|2|耶和华－ 以色列 的上帝论到那些牧养他百姓的牧人如此说：“你们赶散我的羊群，并未看顾他们；看哪，我必惩罚你们的恶行。这是耶和华说的。
JER|23|3|我要从我赶他们到的各国召集我羊群中剩余的，领他们归回本处；他们必生养众多。
JER|23|4|我必设立牧人照管他们，牧养他们。他们不再惧怕，不再惊惶，没有一个失丧的。这是耶和华说的。
JER|23|5|“看哪，日子将到，我要为 大卫 兴起公义的苗裔； 他必掌王权，行事有智慧，在地上施行公平和公义。这是耶和华说的。
JER|23|6|在他的日子， 犹大 必得救， 以色列 也安然居住。他的名必称为‘耶和华－我们的义’。
JER|23|7|“看哪，日子将到，人必不再指着那领 以色列 人从 埃及 地上来的永生耶和华起誓。这是耶和华说的。
JER|23|8|人却要指着那领 以色列 家的后裔离开北方之地，离开我赶他们到的各国的永生耶和华起誓。他们必住在本地。”
JER|23|9|论到那些先知， 我心在我里面忧伤， 我的骨头全都发颤； 因耶和华和他的圣言， 我像醉酒的人， 像被酒所胜的人。
JER|23|10|全地满了犯奸淫的人！ 因妄自赌咒，地就悲哀， 旷野的草场都枯干了。 他们所行的道是恶的； 他们的权力用得不对。
JER|23|11|连先知带祭司都是亵渎的， 就是在我殿中，我也看见他们的恶行。 这是耶和华说的。
JER|23|12|因此，他们的道路必像黑暗中的滑地， 他们必被追赶，仆倒在其上； 因为在他们受罚之年， 我必使灾祸临到他们。 这是耶和华说的。
JER|23|13|我在 撒玛利亚 的先知中曾见狂妄的事； 他们藉 巴力 说预言， 使我的百姓 以色列 走迷了路。
JER|23|14|我在 耶路撒冷 的先知中曾见恐怖的事； 他们犯奸淫，行虚谎， 又坚固恶人的手， 无人回转离开自己的恶行。 他们在我面前都像 所多玛 ， 耶路撒冷 的居民都像 蛾摩拉 。
JER|23|15|因此，万军之耶和华论到先知如此说： “看哪，我必使他们吃茵蔯， 喝苦水； 因为亵渎的事出于 耶路撒冷 的先知，遍及各地。”
JER|23|16|万军之耶和华如此说：“你们不要听这些先知向你们所说的预言。他们使你们成为虚无，所说的异象是出于自己的心，不是出于耶和华的口。
JER|23|17|他们常对藐视我的人说：‘耶和华说：你们必享平安。’ 又对一切按自己顽梗之心而行的人说：‘灾祸必不临到你们。’”
JER|23|18|有谁站在耶和华的会中 察看并听见他的话呢？ 有谁留心听他的话呢？
JER|23|19|看哪！耶和华的暴风 在震怒中发出， 是旋转的暴风， 必转到恶人头上。
JER|23|20|耶和华的怒气必不转消， 直到他心中所定的成就了，实现了。 末后的日子，你们要全然明白。
JER|23|21|我并未差遣那些先知， 他们竟自奔跑； 我没有对他们说话， 他们竟自预言。
JER|23|22|他们若站在我的会中， 必使我的百姓听我的话， 又使他们回转离开恶道， 离开他们所行的恶。
JER|23|23|我是靠近你们的上帝，不是遥远的上帝，不是吗？ 这是耶和华说的。
JER|23|24|人岂能在隐密处藏身，使我看不见他呢？这是耶和华说的。我岂不遍满天和地吗？这是耶和华说的。
JER|23|25|我已听见那些先知所说的，他们托我的名说假预言：“我做了梦！我做了梦！”
JER|23|26|所言虚假、心存诡诈的先知，他们这样存心要到几时呢？
JER|23|27|他们彼此述说所做的梦，想要使我的百姓忘记我的名，正如他们祖先因 巴力 忘记我的名一样。
JER|23|28|得梦的先知可以述说那梦；领受我话的人可以诚实讲我的话。糠秕怎能与麦子比较呢？这是耶和华说的。
JER|23|29|我的话岂不像火，又像能打碎磐石的大锤吗？这是耶和华说的。
JER|23|30|看哪，那些先知各从邻舍偷窃我的话，因此我必与他们为敌。这是耶和华说的。
JER|23|31|那些先知用自己的舌头说是耶和华说的；看哪，我必与他们为敌。这是耶和华说的。
JER|23|32|那些以假梦为预言，又述说这梦，以谎言和鲁莽使我百姓走迷了路的，看哪，我必与他们为敌。这是耶和华说的。我并未差遣他们，也没有吩咐他们。他们对这百姓毫无益处。这是耶和华说的。
JER|23|33|无论是这百姓、是先知、是祭司，问你说：“耶和华有什么默示呢？”你就对他们说：“什么默示啊？ 我已撇弃你们了。这是耶和华说的。”
JER|23|34|凡说“耶和华的默示”的，无论是先知、是祭司、是百姓，我必惩罚那人和他的家。
JER|23|35|你们各人要对邻舍、对弟兄如此说：“耶和华回答了什么？耶和华说了什么呢？”
JER|23|36|你们不可再提“耶和华的默示”，因为各人所说的话必成为自己的重担 ；你们错用了永生上帝、万军之耶和华－我们上帝的话。
JER|23|37|你们要对先知如此说：“耶和华回答了你什么？耶和华说了什么呢？”
JER|23|38|你们若说“耶和华的默示”，耶和华就必如此说：“我曾差人到你们那里去，告诉你们不可说‘耶和华的默示’这几个字，你们却说‘耶和华的默示’；
JER|23|39|所以，看哪，我必忘记你们 ，将你们和我所赐给你们并你们祖先的城都撇弃了；
JER|23|40|又必使永远的凌辱和长久的羞耻临到你们，是不能忘记的。”
JER|24|1|巴比伦 王 尼布甲尼撒 将 约雅敬 的儿子 犹大 王 耶哥尼雅 和 犹大 的领袖，并工匠、铁匠从 耶路撒冷 掳去，带到 巴比伦 。这事以后，耶和华指给我看，看哪，有两筐无花果放在耶和华殿前。
JER|24|2|一筐是极好的无花果，像是初熟的；一筐是极坏的无花果，坏得不能吃。
JER|24|3|耶和华对我说：“ 耶利米 ，你看见什么？”我说：“我看见无花果，好的极好，坏的极坏，坏得不能吃。”
JER|24|4|于是耶和华的话临到我，说：
JER|24|5|“耶和华－ 以色列 的上帝如此说：‘被掳去的 犹大 人，就是我所打发离开这地到 迦勒底 人之地去的，我必看顾他们如这好的无花果，使他们得福乐。
JER|24|6|我要眷顾他们，使他们得福乐，领他们归回这地。我也要建立他们，必不拆毁；栽植他们，必不拔出。
JER|24|7|我要赐给他们认识我的心，认识我是耶和华。他们要作我的子民，我要作他们的上帝，他们要一心归向我。’”
JER|24|8|耶和华如此说：“我必将 犹大 王 西底家 和他的众领袖，以及留在这地 耶路撒冷 剩余的人，并住在 埃及 地的 犹大 人都交出来，好像那极坏、坏得不能吃的无花果。
JER|24|9|我必使他们在地上万国中成为恐惧，成为灾祸，在我赶逐他们到的各处成为凌辱、笑柄、讥笑、诅咒的对象。
JER|24|10|我必使刀剑、饥荒、瘟疫临到他们，直到他们从我所赐给他们和他们祖先之地灭绝。”
JER|25|1|约西亚 的儿子 犹大 王 约雅敬 第四年，就是 巴比伦 王 尼布甲尼撒 的元年，耶和华论 犹大 众百姓的话临到 耶利米 。
JER|25|2|耶利米 先知就将这些话对 犹大 众百姓和 耶路撒冷 所有的居民说：
JER|25|3|“从 亚们 的儿子 犹大 王 约西亚 十三年直到今日，在这二十三年中，常有耶和华的话临到我；我也一再对你们传讲，只是你们不听从。
JER|25|4|耶和华也曾一再差遣他的仆人众先知到你们这里来，只是你们不听从，也不侧耳而听，
JER|25|5|说：‘你们各人当回转离开恶道和恶行，就可居住耶和华从古时所赐给你们和你们祖先之地，直到永远。
JER|25|6|不可随从别神，事奉敬拜它们，以你们手所做的惹我发怒；这样，我就不会降灾祸给你们。
JER|25|7|然而你们不听从我，竟以手所做的惹我发怒，害了自己。这是耶和华说的。’”
JER|25|8|所以万军之耶和华如此说：“因为你们不听我的话，
JER|25|9|看哪，我必召北方的众族和我仆人 巴比伦 王 尼布甲尼撒 前来攻击这地和这地的居民，并四围所有的国民。我要将他们尽行灭绝，以致他们令人惊骇、嗤笑，并且永久荒凉 。这是耶和华说的。
JER|25|10|我又要止息他们欢喜和快乐的声音、新郎和新娘的声音、推磨的声音和灯的亮光。
JER|25|11|这全地必然荒凉，令人惊骇。这些国家要服事 巴比伦 王七十年。
JER|25|12|七十年满了以后，我必惩罚 巴比伦 王和那国，并 迦勒底 人之地，因他们的罪孽使那地永远荒凉。这是耶和华说的。
JER|25|13|我也必使我向那地所说的话，就是所有记在这书上， 耶利米 向这些国家说的预言，都临到那地。
JER|25|14|因为必有许多国家和大君王使 迦勒底 人作奴仆；我也必照他们的行为，按他们手所做的报应他们。”
JER|25|15|耶和华－ 以色列 的上帝对我如此说：“你从我手中拿这杯愤怒的酒，给我所差遣你去的各国的百姓喝。
JER|25|16|他们喝了就要东倒西歪，并要发狂，因我使刀剑临到他们中间。”
JER|25|17|我就从耶和华的手中拿了这杯，给耶和华所差遣我去的各国的百姓喝，
JER|25|18|其中有 耶路撒冷 和 犹大 的城镇，并 耶路撒冷 的君王与领袖；因此这城镇荒凉，令人惊骇、嗤笑、诅咒，正如今日一样。
JER|25|19|又有 埃及 王法老和他的臣仆、官长，以及他的众百姓，
JER|25|20|并混居的各族和 乌斯 地的诸王，与 非利士 人之地的诸王，包括 亚实基伦 、 迦萨 、 以革伦 ，以及 亚实突 剩下的人，
JER|25|21|还有 以东 、 摩押 、 亚扪 人，
JER|25|22|推罗 的诸王、 西顿 的诸王、海的那边沿海地区的诸王，
JER|25|23|底但 、 提玛 、 布斯 ，和所有剃鬓发的人，
JER|25|24|阿拉伯 的诸王、住旷野混居各族的诸王、
JER|25|25|心利 的诸王、 以拦 的诸王、 玛代 的诸王、
JER|25|26|北方远近的诸王，以及天下、地面上的万国也一个一个都喝了，以后 示沙克 王也要喝。
JER|25|27|“你要对他们说：‘万军之耶和华－ 以色列 的上帝如此说：你们要喝，且要喝醉，要呕吐，且要跌倒，不再起来，都因我使刀剑临到你们中间。’
JER|25|28|“他们若不肯从你手中拿这杯来喝，你就要对他们说：‘万军之耶和华如此说：你们一定要喝！
JER|25|29|看哪，我既从称为我名下的城起首施行灾祸，你们能免去惩罚吗？你们必不能免，因为我要命刀剑临到地上所有的居民。这是万军之耶和华说的。’
JER|25|30|“所以你要向他们预言这一切的话，对他们说： ‘耶和华从高天吼叫， 从圣所发出声音， 向自己的羊群大声吼叫； 他要向地上所有的居民呐喊， 像踹葡萄的人一样。
JER|25|31|必有响声达到地极， 因为耶和华与列国争辩。 凡有血肉之躯的，他必审问； 至于恶人，他必交给刀剑。 这是耶和华说的。’
JER|25|32|“万军之耶和华如此说： 看哪，必有灾祸发出，从这国到那国， 并有大暴风从地极刮起。
JER|25|33|“到那日，从地这边到地那边，都有耶和华所杀戮的人。必无人哀哭，不得收殓，不得埋葬，必在地面上成为粪土。
JER|25|34|“牧人哪，你们当哀号，呼喊； 羊群的领导者啊，你们要在灰中翻滚； 因为你们被宰杀、被分散 的日子已经来到。 你们要仆倒，好像珍贵的器皿打碎一样。
JER|25|35|牧人无路可逃， 羊群的领导者也无法逃脱。
JER|25|36|听啊，有牧人呼喊， 有羊群领导者哀号的声音， 因为耶和华摧毁他们的草场。
JER|25|37|因耶和华猛烈的怒气， 平安的羊圈都被肃清。
JER|25|38|他像狮子离开洞穴， 他们的地因凶猛的怒气 和他强烈的怒气，都变为荒凉。”
JER|26|1|约西亚 的儿子 犹大 王 约雅敬 登基时，有这话从耶和华临到 耶利米 ，说：
JER|26|2|“耶和华如此说：你要站在耶和华殿的院内，对 犹大 所有城镇的人，就是到耶和华的殿来礼拜的，传讲我所吩咐你的一切话，一字也不可删减。
JER|26|3|或者他们肯听从，各人回转离开恶道，我就改变心意，不将我因他们所行的恶、想要施行的灾祸降与他们。
JER|26|4|你要对他们说，耶和华如此说：‘你们若不听从我，不遵行我在你们面前所设立的律法，
JER|26|5|不听从我一再差遣我仆人众先知到你们那里去所说的话，你们果然没有听从，
JER|26|6|我就必使这殿如 示罗 ，使这城成为地上万国所诅咒的。’”
JER|26|7|耶利米 在耶和华殿中所说的这些话，祭司、先知与众百姓都听见了。
JER|26|8|耶利米 说完了耶和华吩咐他对众百姓说的一切话，祭司、先知与众百姓都来抓住他，说：“你该死！
JER|26|9|你为何假借耶和华的名预言，说这殿必如 示罗 ，这城必荒废无人居住呢？”于是众百姓都聚集在耶和华的殿中围住 耶利米 。
JER|26|10|犹大 的官长们听见这些事，就从王宫上到耶和华的殿，坐在耶和华殿 新门 的入口。
JER|26|11|祭司、先知对官长和众百姓说：“这人该死，因为他说预言攻击这城，正如你们亲耳听见的。”
JER|26|12|耶利米 就对官长和众百姓说：“耶和华差遣我预言攻击这殿和这城，传讲你们所听见的这一切话。
JER|26|13|现在，要改正你们的所作所为，听从耶和华－你们上帝的话，他就必改变心意，不把所说的灾祸降与你们。
JER|26|14|至于我，看哪，我在你们手中，你们眼里看什么是好的，是正确的，就那样待我吧！
JER|26|15|但你们要确实知道，你们若把我处死，就使流无辜人血的罪归给你们和这城，以及城里的居民了；因为耶和华确实差遣我到你们这里来，将这一切话传到你们耳中。”
JER|26|16|官长和众百姓对祭司和先知说：“这人是不该死的，因为他奉耶和华－我们上帝的名向我们说话。”
JER|26|17|国中的长老就有几个人起来，对聚集的众百姓说：
JER|26|18|“当 犹大 王 希西家 的日子，有 摩利沙 人 弥迦 对 犹大 众百姓预言说： ‘万军之耶和华如此说： 锡安 要被耕种像一块田地， 耶路撒冷 要变为废墟， 这殿的山必像丛林的高处。’
JER|26|19|“ 犹大 王 希西家 和 犹大 人岂是把他处死呢？ 希西家 岂不是敬畏耶和华，恳求耶和华施恩吗？耶和华就改变心意，不把所说的灾祸降与他们。若处死这人，我们就做了大恶，害死自己了。”
JER|26|20|有一个人，就是 示玛雅 的儿子 基列．耶琳 人 乌利亚 ，也奉耶和华的名说预言；他说预言攻击这城和这地，和 耶利米 所说的完全一样。
JER|26|21|约雅敬 王和他所有的勇士、官长听见了 乌利亚 的话，王想要把他处死。 乌利亚 听见就惧怕，逃往 埃及 去了。
JER|26|22|约雅敬 王差 亚革波 的儿子 以利拿单 ，带领几个人前往 埃及 。
JER|26|23|他们将 乌利亚 从 埃及 带出来，解送到 约雅敬 王那里；王用刀杀了他，把他的尸首抛在平民的坟地中。
JER|26|24|然而， 沙番 的儿子 亚希甘 保护 耶利米 ，不将他交在百姓手中，以免他们把他处死。
JER|27|1|约西亚 的儿子 犹大 王 约雅敬 登基时，有这话从耶和华临到 耶利米 ，说：
JER|27|2|“耶和华对我如此说：你要为自己做皮带和木轭，套在你的颈项上，
JER|27|3|然后托那些来到 耶路撒冷 ，到 犹大 王 西底家 那里的使节，把皮带和木轭送到 以东 王、 摩押 王、 亚扪 王、 推罗 王、 西顿 王那里，
JER|27|4|且嘱咐他们转达他们的主人。万军之耶和华－ 以色列 的上帝如此说，你们要对你们的主人这样说：
JER|27|5|我用大能和伸出来的膀臂创造大地和地上的人民、牲畜。我看给谁合适，就把地给谁。
JER|27|6|现在我将全地都交在我仆人 巴比伦 王 尼布甲尼撒 手中，也把野地的走兽给他使用。
JER|27|7|列国都要服事他和他的子孙，直到他本国遭报的日期来到；那时，许多国家和大君王要使他作奴隶。
JER|27|8|“无论哪一邦、哪一国，不肯服事 巴比伦 王 尼布甲尼撒 ，不把颈项放在他的轭下，我必用刀剑、饥荒、瘟疫惩罚那邦，直到我藉 巴比伦 王的手毁灭他们。这是耶和华说的。
JER|27|9|至于你们，不可听从你们的先知和占卜的、做梦的 、观星象的，以及行邪术的；他们对你们说：‘你们必不致服事 巴比伦 王。’
JER|27|10|他们向你们传的是假预言，要叫你们远离本地，以致我将你们赶出去，使你们灭亡。
JER|27|11|但哪一邦肯把颈项放在 巴比伦 王的轭下服事他，我必使那邦仍在本地存留，在那里耕种居住。这是耶和华说的。”
JER|27|12|我就照这一切话对犹大王 西底家 说：“你们要把颈项放在 巴比伦 王的轭下，服事他和他的百姓，就得存活。
JER|27|13|你和你的百姓何必因刀剑、饥荒、瘟疫而死亡，像耶和华所论不肯服事 巴比伦 王的国家呢？
JER|27|14|不可听那些先知对你们所说的话，他们说：‘你们必不致服事 巴比伦 王’，其实他们向你们传的是假预言。
JER|27|15|耶和华说：‘我并未差遣他们，他们却托我的名传假预言，使我将你们和向你们说预言的那些先知赶出去，一同灭亡。’”
JER|27|16|我又对祭司和这众百姓说：“耶和华如此说：你们不可听那先知对你们所说的预言，他们说：‘看哪，耶和华殿中的器皿快要从 巴比伦 带回来’；其实他们向你们传的是假预言。
JER|27|17|不可听从他们，只管服事 巴比伦 王，就得存活。何必使这城变为废墟呢？
JER|27|18|他们若真是先知，有耶和华的话临到他们，让他们祈求万军之耶和华，使耶和华殿中和 犹大 王宫内，并 耶路撒冷 剩下的器皿，不致被带到 巴比伦 去。
JER|27|19|万军之耶和华这样论柱子、铜海、盆座，并留在这城里剩下的器皿，
JER|27|20|就是 巴比伦 王 尼布甲尼撒 掳掠 约雅敬 的儿子 犹大 王 耶哥尼雅 ，并 犹大 、 耶路撒冷 所有贵族时，没有从 耶路撒冷 掠去 巴比伦 的器皿。
JER|27|21|论到那在耶和华殿中和 犹大 王宫内，并 耶路撒冷 剩下的器皿，万军之耶和华－ 以色列 的上帝如此说：
JER|27|22|它们必被带到 巴比伦 ，存放在那里，直到我眷顾 以色列 人，将这些器皿带回归还此地的日子。这是耶和华说的。”
JER|28|1|当年，就是 犹大 王 西底家 登基第四年五月， 押朔 的儿子 基遍 人 哈拿尼雅 先知，在耶和华的殿中当着祭司和众百姓的面对我说：
JER|28|2|“万军之耶和华－ 以色列 的上帝如此说：我已经折断 巴比伦 王的轭。
JER|28|3|二年之内，我要将 巴比伦 王 尼布甲尼撒 从这地掳掠到 巴比伦 的器皿，就是耶和华殿中的一切器皿，都带回此地。
JER|28|4|我又要将 约雅敬 的儿子 犹大 王 耶哥尼雅 和被掳到 巴比伦 所有的 犹大 人带回此地，因为我要折断 巴比伦 王的轭。这是耶和华说的。”
JER|28|5|耶利米 先知当着祭司和站在耶和华殿里众百姓的面，对 哈拿尼雅 先知说：
JER|28|6|“阿们！愿耶和华如此行，愿耶和华实现你所预言的话，将耶和华殿中的器皿和所有被掳去的人从 巴比伦 带回此地。
JER|28|7|然而我在你和众百姓耳中所要说的话，你应当听。
JER|28|8|从古以来，在你我以前的众先知，向多国和大邦说预言，论到战争、灾祸 、瘟疫的事。
JER|28|9|至于那预言平安的先知，到先知的话应验的时候，人就知道他真是耶和华所差来的。”
JER|28|10|哈拿尼雅 先知就取下 耶利米 先知颈项上的轭，把它折断。
JER|28|11|哈拿尼雅 又当着众百姓的面说：“耶和华如此说：二年之内我必照样从列国的颈项上折断 巴比伦 王 尼布甲尼撒 的轭。” 耶利米 先知就离开了。
JER|28|12|哈拿尼雅 先知折断 耶利米 先知颈项上的轭以后，耶和华的话临到 耶利米 ，说：
JER|28|13|“你去告诉 哈拿尼雅 说，耶和华如此说：你折断木轭，却换来铁轭！
JER|28|14|万军之耶和华－ 以色列 的上帝如此说：我已将铁轭加在这些国的颈项上，使他们服事 巴比伦 王 尼布甲尼撒 。他们总要服事他，我也把野地的走兽给了他。”
JER|28|15|于是 耶利米 先知对 哈拿尼雅 先知说：“ 哈拿尼雅 啊，你应当听！耶和华并没有差遣你，你竟使这百姓倚靠谎言。
JER|28|16|所以耶和华如此说：看哪，我要把你从地面上除掉，你今年必死，因为你向耶和华说了叛逆的话。”
JER|28|17|这样， 哈拿尼雅 先知当年七月间就死了。
JER|29|1|耶利米 先知从 耶路撒冷 送信给被掳幸存的长老，以及祭司、先知，和 尼布甲尼撒 从 耶路撒冷 掳到 巴比伦 去的众百姓。
JER|29|2|这是在 耶哥尼雅 王和太后、官员，并 犹大 和 耶路撒冷 的领袖，以及工匠、铁匠都离开 耶路撒冷 之后。
JER|29|3|他藉 沙番 的儿子 以利亚萨 和 希勒家 的儿子 基玛利 的手送去；他们二人是 犹大 王 西底家 差往 巴比伦 去见 巴比伦 王 尼布甲尼撒 的。
JER|29|4|信上说：“万军之耶和华－ 以色列 的上帝对所有被掳的，就是我使他们从 耶路撒冷 被掳到 巴比伦 去的人如此说：
JER|29|5|你们要建造房屋，住在其中；要开垦田园，吃园中所出产的；
JER|29|6|要娶妻生儿养女，为你们的儿子娶妻，使你们的女儿嫁人，生儿养女。你们要在那里生养众多，不可减少。
JER|29|7|我使你们被掳到的那城，你们要为那城求平安，为那城向耶和华祈求，因为那城得平安，你们也随着得平安。
JER|29|8|万军之耶和华－ 以色列 的上帝如此说：不要被你们中间的先知和占卜的所诱惑，也不要听信你们 所做的梦，
JER|29|9|因为他们托我的名对你们说假预言，我并未差遣他们。这是耶和华说的。
JER|29|10|“耶和华如此说：为 巴比伦 所定的七十年满了以后，我要眷顾你们，向你们实现我的恩言，使你们归回此地。
JER|29|11|我知道我向你们所怀的意念是赐平安的意念，不是降灾祸的意念，要叫你们末后有指望。这是耶和华说的。
JER|29|12|你们呼求我，向我祷告，我就应允你们。
JER|29|13|你们寻求我，若专心寻求我，就必寻见。
JER|29|14|我必被你们寻见，也必使你们被掳的人归回。这是耶和华说的。我必将你们从各国和我赶你们到的各处召集过来，又将你们带回我使你们被掳离开的地方。这是耶和华说的。
JER|29|15|“你们说：‘耶和华已在 巴比伦 为我们兴起先知。’
JER|29|16|所以耶和华如此论坐 大卫 宝座的君王和住在这城里所有的百姓，就是未曾与你们一同被掳的弟兄，
JER|29|17|万军之耶和华如此说：‘看哪，我必使刀剑、饥荒、瘟疫临到他们，使他们像极坏的无花果，坏得不能吃。
JER|29|18|我必用刀剑、饥荒、瘟疫追赶他们，使地上万国因他们而惊骇；在我赶他们到的各国，令人诅咒、惊骇、嗤笑、羞辱。
JER|29|19|这是因为他们不听从我先前一再差遣我仆人众先知说的话。这是耶和华说的。你们 也一样不听。这是耶和华说的。’
JER|29|20|所以你们所有被掳去的，就是我从 耶路撒冷 放逐到 巴比伦 去的，当听耶和华的话。
JER|29|21|万军之耶和华－ 以色列 的上帝论 哥赖雅 的儿子 亚哈 和 玛西雅 的儿子 西底家 如此说：‘他们托我的名向你们说假预言，看哪，我必把他们交在 巴比伦 王 尼布甲尼撒 的手中，他要在你们眼前杀害他们。
JER|29|22|在 巴比伦 所有被掳的 犹大 人必藉这二人赌咒说：愿耶和华使你像 巴比伦 王在火中焚烧的 西底家 和 亚哈 一样。
JER|29|23|这二人在 以色列 中做了丑事，与邻舍的妻行淫，又假托我的名说我未曾吩咐他们的话。我知道这一切，也作见证。这是耶和华说的。’”
JER|29|24|“你要对 尼希兰 人 示玛雅 说：
JER|29|25|万军之耶和华－ 以色列 的上帝如此说：你曾用自己的名送信给 耶路撒冷 的众百姓和 玛西雅 的儿子 西番雅 祭司，并众祭司，说：
JER|29|26|‘耶和华已经立你 西番雅 为祭司，代替 耶何耶大 祭司，使耶和华的殿中有总管，好把所有狂妄自称先知的人用枷枷住，用锁锁住。
JER|29|27|现在 亚拿突 人 耶利米 向你们自称先知，你为什么不责备他呢？
JER|29|28|他送信给我们在 巴比伦 的人说：被掳的事必长久，你们要建造房屋，住在其中；要开垦田园，吃园中所出产的。’”
JER|29|29|西番雅 祭司就把这信念给 耶利米 先知听。
JER|29|30|于是耶和华的话临到 耶利米 ，说：
JER|29|31|“你当送信给所有被掳的人，说：‘耶和华论到 尼希兰 人 示玛雅 说：因为 示玛雅 向你们说预言，使你们倚靠谎言，而我并没有差遣他，
JER|29|32|所以耶和华如此说：看哪，我必惩罚 尼希兰 人 示玛雅 和他的后裔，他必无一人存留住在这民中，也看不见我所要赏赐给我百姓的福乐，因为他向耶和华说了叛逆的话。这是耶和华说的。’”
JER|30|1|耶和华的话临到 耶利米 ，说：
JER|30|2|“耶和华－ 以色列 的上帝如此说：你要将我对你说过的一切话都写在书上。
JER|30|3|看哪，日子将到，我要使我的百姓 以色列 和 犹大 被掳的人归回。这是耶和华说的。耶和华说：我要使他们回到我所赐给他们祖先之地，他们就得这地为业。”
JER|30|4|以下是耶和华论到 以色列 和 犹大 所说的话：
JER|30|5|耶和华如此说： “我们听见颤抖的声音， 令人惧怕，没有平安。
JER|30|6|你们且访查看看， 男人会生孩子吗？ 我怎么看见人人都用手撑腰， 像临产的妇人， 脸都发白了呢？
JER|30|7|哀哉！ 那日为大， 无日可比； 这是 雅各 遭难的时刻， 但他必从患难中得拯救。”
JER|30|8|万军之耶和华说：“到那日，我必折断你颈项上仇敌的轭，拉断你的皮带。陌生人必不再使他作奴隶。
JER|30|9|他们却要事奉耶和华－他们的上帝，事奉我为他们所兴起的 大卫 王。”
JER|30|10|我的仆人 雅各 啊，不要惧怕； 以色列 啊，不要惊惶； 因我从远方拯救你， 从被掳之地拯救你的后裔； 雅各 必回来得享平静安逸， 无人能使他害怕。 这是耶和华说的。
JER|30|11|因我与你同在，要拯救你， 也要将那些国灭绝净尽， 就是我赶你去的那些国； 却不将你灭绝净尽， 倒要从宽惩治你， 但绝不能不罚你。 这是耶和华说的。
JER|30|12|耶和华如此说： “你的损伤无法医治， 你的伤痕极其重大。
JER|30|13|无人为你的伤痛辩护， 也没有可医治你的良药。
JER|30|14|你所亲爱的都忘记你， 不来探望你。 我因你罪孽甚大，罪恶众多， 曾藉仇敌加的伤害伤害你， 藉残忍者惩治你。
JER|30|15|你为何因所受的损伤哀号呢？ 你的痛苦无法医治。 我因你罪孽甚大，罪恶众多， 曾将这些加在你身上。
JER|30|16|因此，凡吞吃你的必被吞吃， 你的敌人个个都被掳去； 掳掠你的必成为掳物， 我使抢夺你的成为掠物。
JER|30|17|我必使你痊愈， 医好你的伤痕， 都因人称你为被赶散的， 这是 锡安 ，是无人来探望的！ 这是耶和华说的。”
JER|30|18|耶和华如此说： “看哪，我必使 雅各 被掳去的帐棚归回， 也必顾惜他的住处。 城必建造在原有的废墟上， 宫殿也必照样有人居住。
JER|30|19|必有感谢和欢乐的声音从其中发出， 我使他们增多，不致减少； 使他们尊荣，不致卑微。
JER|30|20|他们的儿女必如往昔； 他们的会众坚立在我面前； 凡欺压他们的，我必惩罚。
JER|30|21|他们的君王是他们自己的人， 掌权的必出自他们。 我要使他接近我， 他也要亲近我； 不然，谁敢放胆亲近我呢？ 这是耶和华说的。
JER|30|22|你们要作我的子民， 我要作你们的上帝。”
JER|30|23|看哪，耶和华的愤怒 如暴风已经发出； 是扫灭的暴风， 必转到恶人的头上。
JER|30|24|耶和华的烈怒必不转消， 直到他心中所定的成就了，实现了； 末后的日子你们就会明白。
JER|31|1|耶和华说：“那时，我必作 以色列 各家的上帝，他们必作我的子民。”
JER|31|2|耶和华如此说： “从刀剑生还的百姓 在旷野蒙恩； 以色列 寻找安歇之处。”
JER|31|3|耶和华从远方向我显现： “我以永远的爱爱你， 因此，我以慈爱吸引你。”
JER|31|4|少女 以色列 啊， 我要再建立你，你就得以建立； 你必再拿起手鼓， 随着欢乐的舞者而出。
JER|31|5|你必在 撒玛利亚 的山上栽葡萄园， 栽种的人栽种，而且享用。
JER|31|6|日子将到，守望的人必在 以法莲 山上呼叫： “起来吧！我们要上 锡安 ， 到耶和华－我们的上帝那里去。”
JER|31|7|耶和华如此说： “你们当为 雅各 欢乐歌唱， 为万国中为首的欢呼。 当传扬，颂赞说： ‘耶和华啊， 求你拯救你的百姓 ， 拯救 以色列 的余民。’
JER|31|8|看哪，我必将他们从北方之地领来， 从地极召集而来； 同他们来的有盲人、瘸子、孕妇、产妇； 他们必成群结队回到这里。
JER|31|9|他们要哭泣而来。 我要照他们恳求的引导他们， 使他们在河水旁行走正直的路， 他们在其上必不致绊跌； 因为我是 以色列 的父， 以法莲 是我的长子。
JER|31|10|列国啊，要听耶和华的话， 要在远方的海岛传扬，说： “赶散 以色列 的必召集他， 看守他，如牧人看守羊群。”
JER|31|11|因为耶和华救赎了 雅各 ， 救赎他脱离比他更强之人的手。
JER|31|12|他们来到 锡安 的高处歌唱， 因耶和华的宏恩而喜乐洋溢， 就是五谷、新酒和新的油， 并羔羊和牛犊。 他们必像有水浇灌的园子， 一点也不再有愁烦。
JER|31|13|那时，少女必欢乐跳舞； 年轻的、年老的，都一同欢乐； 因为我要使他们的悲哀变为欢喜， 并要安慰他们，使他们的愁烦转为喜乐。
JER|31|14|我必以肥油使祭司的心满足， 我的百姓也要因我的恩惠知足。 这是耶和华说的。
JER|31|15|耶和华如此说： “在 拉玛 听见号啕痛哭的声音， 是 拉结 哭她儿女，不肯因她儿女受安慰， 因为他们都不在了。”
JER|31|16|耶和华如此说： “不要出声哀哭， 你的眼目也不要流泪； 因你的辛劳必有报偿， 他们必从仇敌之地归回。 这是耶和华说的。
JER|31|17|你末后必有指望， 你的儿女必回到自己的疆土。 这是耶和华说的。
JER|31|18|我听见 以法莲 为自己悲叹说： ‘你管教我，我便受管教， 我如未驯服的牛犊。 求你使我回转，我便回转， 因为你是耶和华－我的上帝。
JER|31|19|我背离以后就懊悔， 受教以后就捶胸 ； 我因担当年轻时的凌辱就抱愧蒙羞。’
JER|31|20|以法莲 是我的爱子吗？ 是我喜欢的孩子吗？ 我每逢责备他，仍深顾念他。 因此，我的心肠牵挂着他， 我必要怜悯他。 这是耶和华说的。
JER|31|21|少女 以色列 啊， 当为自己设立路标， 为自己竖起指路牌。 要留心向着大道， 就是你曾走过的路； 你当回转，回到你自己的城镇。
JER|31|22|背道的女子啊， 你翻来覆去要到几时呢？ 耶和华在地上造了一件新事， 就是女子护卫男子。”
JER|31|23|万军之耶和华－ 以色列 的上帝如此说：“我使被掳之人归回的时候，他们在 犹大 地和其中的城镇必再这样说： 公义的居所啊，圣山哪， 愿耶和华赐福给你。
JER|31|24|犹大 和 犹大 城镇的人，耕地的和带着群畜游牧的人，都要一同住在其中。
JER|31|25|疲乏的人，我使他振作；愁烦的人，我使他满足。”
JER|31|26|于是我醒了，我看到我睡得香甜。
JER|31|27|“看哪，日子将到，我要使人的后代和牲畜的种，在 以色列 家和 犹大 家繁衍。这是耶和华说的。
JER|31|28|我先前怎样看守他们，为要拔出、拆毁、毁坏、倾覆、苦害，也必照样看守他们，为要建立、栽植。这是耶和华说的。
JER|31|29|当那些日子，人不再说： ‘父亲吃了酸葡萄， 儿子牙齿就酸倒。’
JER|31|30|但各人要因自己的罪死亡；凡吃酸葡萄的，自己的牙必酸倒。
JER|31|31|“看哪，日子将到，我要与 以色列 家和 犹大 家另立新的约。这是耶和华说的。
JER|31|32|这约不像我拉着他们祖宗的手，领他们出 埃及 地的时候与他们所立的约。我虽作他们的丈夫，他们却背了我的约。这是耶和华说的。
JER|31|33|那些日子以后，我与 以色列 家所立的约是这样：我要将我的律法放在他们里面，写在他们心上。我要作他们的上帝，他们要作我的子民。这是耶和华说的。
JER|31|34|他们各人不再教导自己的邻舍和弟兄说：‘你该认识耶和华’，因为他们从最小的到最大的都必认识我。我要赦免他们的罪孽，不再记得他们的罪恶。这是耶和华说的。”
JER|31|35|耶和华使太阳白昼发光， 按定例使月亮和星辰照耀黑夜， 又搅动大海，使海中波浪澎湃， 万军之耶和华是他的名， 他如此说：
JER|31|36|“这些定例若能在我面前废掉， 以色列 的后裔才会在我面前断绝， 永远不再成国。 这是耶和华说的。”
JER|31|37|耶和华如此说： “若有人能测量上面的天， 探索下面地的根基， 我才会因 以色列 后裔所做的一切弃绝他们。 这是耶和华说的。”
JER|31|38|看哪，日子将到，这城必为耶和华而造，从 哈楠业楼 直到 角门 。这是耶和华说的。
JER|31|39|丈量的绳子要往外拉出，直到 迦立山 ，又转到 歌亚 ；
JER|31|40|抛尸的全谷和倒灰之处，并一切田地，直到 汲沦溪 ，又到东边 马门 的角落，都要归耶和华为圣；不再拔出，不再倾覆，直到永远。
JER|32|1|犹大 王 西底家 第十年，就是 尼布甲尼撒 十八年，耶和华的话临到 耶利米 。
JER|32|2|那时 巴比伦 王的军队围困 耶路撒冷 ， 耶利米 先知被囚在 犹大 王宫中护卫兵的院内；
JER|32|3|因为 犹大 王 西底家 囚禁他，说：“你为什么预言耶和华如此说：‘看哪，我要把这城交在 巴比伦 王的手中，他必攻下这城。
JER|32|4|犹大 王 西底家 必不能逃脱 迦勒底 人的手，定要交在 巴比伦 王手中，他要亲眼看到 巴比伦 王，亲口跟他说话。
JER|32|5|巴比伦 王要将 西底家 带到 巴比伦 ； 西底家 必住在那里，直到我惩罚 他的时候。你们虽与 迦勒底 人争战，却不顺利。这是耶和华说的。’”
JER|32|6|耶利米 说：“耶和华的话临到我，说：
JER|32|7|‘看哪，你叔父 沙龙 的儿子 哈拿篾 必到你这里来，说：请你买我在 亚拿突 的那块地，因为你有代赎的责任。’
JER|32|8|我叔父的儿子 哈拿篾 果然照耶和华的话来到护卫兵的院内，对我说：‘请你买我在 便雅悯 境内、 亚拿突 的那块地；因为它应该由你来承受，而且你也有代赎的责任。请你买下它吧！’我就知道这确是耶和华的话。
JER|32|9|“我便向我叔父的儿子 哈拿篾 买了 亚拿突 的那块地，秤了十七舍客勒银子给他。
JER|32|10|我在契上签字，将契封缄，又请证人来，用天平把银子秤给他。
JER|32|11|我又将按照法定条例所立的买契，就是封缄的那一张和敞开的那一张，
JER|32|12|在我叔父的儿子 哈拿篾 和签字作证的人，并坐在护卫兵院内所有 犹大 人眼前，交给 玛西雅 的孙子 尼利亚 的儿子 巴录 。
JER|32|13|我在众人眼前嘱咐 巴录 说：
JER|32|14|‘万军之耶和华－ 以色列 的上帝如此说：你拿着这文件，就是封缄的和敞开的买契，把它们放在瓦器里，以便长久保存。
JER|32|15|因为万军之耶和华－ 以色列 的上帝如此说：将来在这地必有人再购置房屋、田地和葡萄园。’”
JER|32|16|“我将买契交给 尼利亚 的儿子 巴录 以后，就向耶和华祷告说：
JER|32|17|‘唉！主耶和华，看哪，你曾用大能和伸出来的膀臂创造天和地，在你没有难成的事。
JER|32|18|你施慈爱给千万人，又将祖先的罪孽报应在他后世子孙身上。至大全能的上帝啊，万军之耶和华是你的名，
JER|32|19|你谋事有大略，行事有大能，注目观看世人一切的举动，为要照各人所做的和他做事的结果报应他。
JER|32|20|你在 埃及 地显神迹奇事，直到今日在 以色列 和世人中间也是如此，建立了自己的名声，正如今日一样。
JER|32|21|你用神迹奇事、大能的手、伸出来的膀臂和大可畏的事，领你的百姓 以色列 出了 埃及 ，
JER|32|22|把这地赏赐给他们，就是你向他们列祖起誓应许要赐给他们的流奶与蜜之地。
JER|32|23|他们进入并取得这地，却不听从你的话，也不遵行你的律法。你吩咐他们所当行的，他们都不去行，因此你使这一切的灾祸临到他们。
JER|32|24|看哪，敌人已经来到，用土堆攻取这城；这城也因刀剑、饥荒、瘟疫被交在攻城的 迦勒底 人手中。你所说的话都应验了，看哪，你也看见了。
JER|32|25|主耶和华啊，你却对我说，要用银子为自己买那块地，又请人作证；其实这城已交在 迦勒底 人的手中了。’”
JER|32|26|耶和华的话临到 耶利米 ，说：
JER|32|27|“看哪，我是耶和华，是凡有血肉之躯者的上帝，在我岂有难成的事吗？
JER|32|28|耶和华如此说：看哪，我必将这城交给 迦勒底 人的手和 巴比伦 王 尼布甲尼撒 的手，他必攻取这城。
JER|32|29|攻城的 迦勒底 人必来放火焚烧这城和城里的房屋；人曾在这房顶上向 巴力 烧香，向别神献浇酒祭，惹我发怒。
JER|32|30|以色列 人和 犹大 人从年轻时，就专做我眼中看为恶的事。 以色列 人尽以手所做的惹我发怒。这是耶和华说的。
JER|32|31|这城自从建造的那日直到今日，常惹我的怒气和愤怒，以致我将这城从我面前除掉；
JER|32|32|这是因 以色列 人和 犹大 人一切的邪恶，就是他们和他们的君王、官长、祭司、先知，并 犹大 人，以及 耶路撒冷 居民所做的，惹我发怒。
JER|32|33|他们以背向我，不以面向我；我虽然一再教导他们，他们却不听从，不领受训诲，
JER|32|34|竟把可憎之偶像设立在称为我名下的殿中，玷污了这殿。
JER|32|35|他们在 欣嫩子谷 建造 巴力 的丘坛，把自己的儿女经火献给 摩洛 ；他们行这可憎的事，使 犹大 陷在罪里，这并不是我吩咐的，我心里也从来没有想过。”
JER|32|36|现在论到这城，就是你们所说，已经因刀剑、饥荒、瘟疫被交在 巴比伦 王手中的，耶和华－ 以色列 的上帝如此说：
JER|32|37|“看哪，我曾在怒气、愤怒和大恼怒中，将 以色列 人赶到各国；我必从那里将他们召集出来，领他们回到此地，使他们安然居住。
JER|32|38|他们要作我的子民，我要作他们的上帝。
JER|32|39|我要使他们彼此同心同道，好叫他们永远敬畏我，使他们和他们后世的子孙得享福乐。
JER|32|40|我要跟他们立永远的约，要施恩给他们，绝不转离；又要把敬畏我的心放在他们心里，不离弃我。
JER|32|41|我必欢喜施恩给他们，尽心尽意、真诚地将他们栽于此地。
JER|32|42|“因为耶和华如此说：我怎样使这一切大灾祸临到这百姓，也要照样使我所应许他们的一切福乐都临到他们。
JER|32|43|你们所说荒凉、无人、无牲畜，已交给 迦勒底 人手的这地，必有人购置田地。
JER|32|44|在 便雅悯 地、 耶路撒冷 四围的各处、 犹大 的城镇、山区的城镇、 谢非拉 的城镇，并 尼革夫 的城镇，人必用银子买田地，在契上签字，将契封缄，找人作证，因为我必使被掳的人归回。这是耶和华说的。”
JER|33|1|耶利米 还囚在护卫兵的院内，耶和华的话第二次临到他，说：
JER|33|2|“成事的耶和华，塑造它为要建立它的耶和华，名为耶和华的那位如此说：
JER|33|3|‘你求告我，我就应允你，并将你所不知道、又大又隐密的事指示你。
JER|33|4|论到这城中的房屋和 犹大 君王的宫殿，就是拆毁来挡围城工事和刀剑的，耶和华－ 以色列 的上帝如此说：
JER|33|5|他们与 迦勒底 人争战，用我在怒气和愤怒中所杀之人的尸首塞满这房屋；我因他们一切的恶，转脸不顾这城。
JER|33|6|看哪，我要使这城得以痊愈安舒，我要医治他们，将丰盛的平安与信实显明给他们。
JER|33|7|我也要使 犹大 被掳的和 以色列 被掳的人归回，并要建立他们，如起初一样。
JER|33|8|我要洗净他们干犯我的一切罪，赦免他们干犯我、违背我的一切罪。
JER|33|9|这城在地上万国面前要因我的缘故，以喜乐得名，得颂赞，得荣耀，因为他们听见我所赏赐的一切福乐。他们因我向这城所施的一切福乐平安，就惧怕战兢。”
JER|33|10|耶和华如此说：“你们论这地方，说是荒废、无人、无牲畜之地，但在这荒凉、无人、无居民、无牲畜的 犹大 城镇和 耶路撒冷 街上，必再听见
JER|33|11|欢喜和快乐的声音、新郎和新娘的声音，并听见有人说： 你们要称谢万军之耶和华， 因耶和华本为善， 他的慈爱永远长存！ 他们奉感谢祭到耶和华的殿中；因为我必使这地被掳的人归回，如起初一样。这是耶和华说的。”
JER|33|12|万军之耶和华如此说：“在这荒废、无人、无牲畜之地，并其中所有的城镇，必再有牧人的草场，可让羊群躺卧在那里。
JER|33|13|在山区的城镇、 谢非拉 的城镇、 尼革夫 的城镇、 便雅悯 地、 耶路撒冷 四围的各处和 犹大 的城镇，必再有羊群从数点的人手下经过。这是耶和华说的。
JER|33|14|“看哪，日子将到，我应许 以色列 家和 犹大 家的恩言必然实现。这是耶和华说的。
JER|33|15|在那些日子、那时候，我必使 大卫 公义的苗裔长起来；他必在地上施行公平和公义。
JER|33|16|在那些日子， 犹大 必得救， 耶路撒冷 必安然居住，他的名必称为‘耶和华－我们的义’。
JER|33|17|“因为耶和华如此说： 大卫 家必永远不断有人坐在 以色列 家的宝座上；
JER|33|18|利未 家的祭司也不断有人在我面前献燔祭、烧素祭，时常办理献祭的事。”
JER|33|19|耶和华的话临到 耶利米 ，说：
JER|33|20|“耶和华如此说：你们若能废弃我所立白日黑夜的约，使白日黑夜不按时轮转，
JER|33|21|就能废弃我与我仆人 大卫 所立的约，使他没有后裔在他的宝座上作王，并能废弃我与事奉我的 利未 家的祭司所立的约。
JER|33|22|正如天上的万象不能数算，海边的尘沙不能斗量，我必照样使我仆人 大卫 的后裔和事奉我的 利未 人多起来。”
JER|33|23|耶和华的话临到 耶利米 ，说：
JER|33|24|“你没有留意这百姓所说的话吗？他们说：‘耶和华所拣选的二族，他已经弃绝了。’他们这样藐视我的百姓，不把他们当作国来看待。
JER|33|25|耶和华如此说：除非我没有立白日黑夜之约，也未曾安排天和地的定例，
JER|33|26|否则我不会弃绝 雅各 的后裔和我仆人 大卫 的后裔，使 大卫 的后裔不再治理 亚伯拉罕 、 以撒 、 雅各 的后裔。我必使他们被掳的人归回，也必怜悯他们。”
JER|34|1|巴比伦 王 尼布甲尼撒 率领他的全军和地上他管辖的各国各邦，攻打 耶路撒冷 和 耶路撒冷 所有的城镇。那时，耶和华的话临到 耶利米 ，说：
JER|34|2|“耶和华－ 以色列 的上帝说，你去告诉 犹大 王 西底家 ，耶和华如此说：看哪，我要把这城交在 巴比伦 王的手中，他必用火焚烧。
JER|34|3|你必不能逃脱他的手，定被拿住，交在他手中。你要亲眼看到 巴比伦 王，他要亲口跟你说话，你也必到 巴比伦 去。
JER|34|4|犹大 王 西底家 啊，你一定要听耶和华的话。耶和华论到你如此说：你必不死于刀下；
JER|34|5|必平安而终，人要为你焚烧，好像为你祖先，就是在你以前早先的王焚烧一样。人要为你举哀说：‘哀哉！我主啊。’这话是我说的。这是耶和华说的。”
JER|34|6|于是， 耶利米 先知在 耶路撒冷 把这一切话告诉 犹大 王 西底家 。
JER|34|7|那时， 巴比伦 王的军队正攻打 耶路撒冷 ，又攻打 犹大 仅存的城镇，就是 拉吉 和 亚西加 ；原来 犹大 的坚固城只剩下这两座。
JER|34|8|西底家 王与 耶路撒冷 的众百姓立约，要他们宣告自由，叫各人释放自己的仆人和婢女，使 希伯来 的男人和女人得自由，谁也不可使他的 犹大 弟兄作奴仆。这事以后，耶和华的话临到 耶利米 。
JER|34|9|
JER|34|10|所有前来立约的领袖和众百姓都顺从，各人释放自己的仆人和婢女，使他们得自由，不再叫他们作奴仆。大家都顺从，将仆婢释放了。
JER|34|11|但后来他们又反悔，叫被释放得自由的仆人婢女回来，强迫他们仍为仆婢。
JER|34|12|因此耶和华的话临到 耶利米 ，说：
JER|34|13|“耶和华－ 以色列 的上帝如此说：我将你们祖先从 埃及 地为奴之家领出时，与他们立约说：
JER|34|14|‘你的一个 希伯来 弟兄若卖给你，服事你六年，到第七年你们各人就要释放他自由出去。’只是你们祖先不听我，不侧耳而听。
JER|34|15|如今你们回转，行我眼中看为正的事，各人向邻舍宣告自由，并且在我面前、在称为我名下的殿中立约。
JER|34|16|你们却反悔，亵渎我的名，各人叫所释放得自由的仆人婢女回来，强迫他们仍为仆婢。
JER|34|17|所以耶和华如此说：你们不听从我，各人不向弟兄邻舍宣告自由。看哪！我要向你们宣告自由，把你们自由地交给刀剑、饥荒、瘟疫，并且使地上万国因你们而惊骇。这是耶和华说的。
JER|34|18|那些违背我约的人，就是不遵守在我面前立约之话的，我要使他们成了那劈成两半的牛犊，使人从切块中经过：
JER|34|19|犹大 的领袖、 耶路撒冷 的领袖、官员、祭司，和从牛犊切块中经过的这地的众百姓，
JER|34|20|我必将他们交在仇敌和寻索其命的人手中；他们的尸首必给空中的飞鸟和地上的走兽作食物。
JER|34|21|我必将 犹大 王 西底家 和他的众领袖交在仇敌和寻索其命的人手中，与那暂时离你们而去的 巴比伦 王军队的手中。
JER|34|22|看哪，我要吩咐他们回到这城，攻打这城，将城攻取，用火焚烧；我也要使 犹大 的城镇变为废墟，无人居住。这是耶和华说的。”
JER|35|1|当 约西亚 的儿子 约雅敬 作 犹大 王的时候，耶和华的话临到 耶利米 ，说：
JER|35|2|“你去见 利甲 族的人，吩咐他们，领他们进入耶和华殿的一个房间，给他们酒喝。”
JER|35|3|我就带 哈巴洗尼雅 的孙子 雅利米雅 的儿子 雅撒尼亚 ，和他的兄弟，并他所有的儿子，以及 利甲 全族的人，
JER|35|4|领他们到耶和华的殿，进入 伊基大利 的儿子神人 哈难 儿子们的房间；那房间靠近官长的房间，在 沙龙 之子门口的守卫 玛西雅 的房间上面。
JER|35|5|于是我在 利甲 族的人面前摆设盛满了酒的碗和杯，对他们说：“请喝酒。”
JER|35|6|他们却说：“我们不喝酒，因为我们祖先 利甲 的儿子 约拿达 曾吩咐我们说：‘你们与你们的子孙永不可喝酒，
JER|35|7|不可盖房子，不可撒种，也不可栽葡萄园，连拥有都不可；但一生的年日要住帐棚，使你们的日子在寄居的地面上得以长久。’
JER|35|8|凡我们祖先 利甲 的儿子 约拿达 所吩咐我们的话，我们都听从了。我们和我们的妻子儿女一生的年日都不喝酒，
JER|35|9|不盖房子居住，我们也没有葡萄园、田地和种子；
JER|35|10|但住在帐棚里，听从并遵行我们祖先 约拿达 所吩咐我们的一切话。
JER|35|11|巴比伦 王 尼布甲尼撒 上来攻打这地的时候，我们说：‘来吧，我们到 耶路撒冷 去，躲避 迦勒底 的军队和 亚兰 的军队。’这样，我们才住在 耶路撒冷 。”
JER|35|12|耶和华的话临到 耶利米 ，说：
JER|35|13|“万军之耶和华－ 以色列 的上帝如此说：你去对 犹大 人和 耶路撒冷 的居民说，你们不肯领受训诲，听从我的话吗？这是耶和华说的。
JER|35|14|利甲 的儿子 约拿达 所吩咐他子孙不可喝酒的话，他们已经遵守了；他们因为听从祖先的吩咐，直到今日都不喝酒。至于我，我一再警戒你们，你们却不肯听从我。
JER|35|15|我一再差遣我的仆人众先知到你们那里去，说：‘你们各人当回头离开恶道，改正行为，不再随从事奉别神，如此，就必住在我所赐给你们和你们祖先的地上。’只是你们不侧耳而听，也不听我。
JER|35|16|利甲 的儿子 约拿达 的子孙能遵守祖先所吩咐他们的命令，这百姓却不肯听从我！
JER|35|17|因此，耶和华－万军之上帝、 以色列 的上帝如此说：看哪，我要使我所说的一切灾祸临到 犹大 人和 耶路撒冷 所有的居民。因为我向他们说话，他们不听从；我呼唤他们，他们也没有回应。”
JER|35|18|耶利米 对 利甲 族的人说：“万军之耶和华－ 以色列 的上帝如此说：因你们听从你们祖先 约拿达 的吩咐，谨守他的一切命令，照他所吩咐的去做，
JER|35|19|所以万军之耶和华－ 以色列 的上帝如此说： 利甲 的儿子 约拿达 必永远不断有人侍立在我面前。”
JER|36|1|约西亚 的儿子 犹大 王 约雅敬 第四年，有这话从耶和华临到 耶利米 ，说：
JER|36|2|“你要取一书卷，把我对你所说攻击 以色列 和 犹大 ，并各国的一切话，从我对你说话的那日，就是从 约西亚 的日子起直到今日，都写在其上；
JER|36|3|或者 犹大 家听见我想要降给他们的一切灾祸，各人就回转离开恶道，我就赦免他们的罪孽和罪恶。”
JER|36|4|耶利米 召了 尼利亚 的儿子 巴录 来； 巴录 就从 耶利米 口中，把耶和华对 耶利米 所说的一切话写在书卷上。
JER|36|5|耶利米 吩咐 巴录 说：“我被禁止，不能进耶和华的殿。
JER|36|6|所以你要趁禁食的日子进入耶和华的殿中，把耶和华的话，就是你从我口中写在书卷上的话，念给百姓和所有从各城镇前来的 犹大 人亲耳听；
JER|36|7|或者他们的恳求达到耶和华面前，各人回转离开恶道，因为耶和华向这百姓所说要发的怒气和愤怒实在很大。”
JER|36|8|尼利亚 的儿子 巴录 就照 耶利米 先知所吩咐的一切去做，在耶和华殿中宣读书卷上耶和华的话。
JER|36|9|约西亚 的儿子 犹大 王 约雅敬 第五年九月， 耶路撒冷 的众百姓和那从 犹大 城镇前来 耶路撒冷 的众百姓，在耶和华面前宣告禁食，
JER|36|10|巴录 就在耶和华殿的上院，靠近耶和华殿的 新门 口， 沙番 的儿子 基玛利雅 文士的房间里，宣读书卷上 耶利米 的话给众百姓亲耳听。
JER|36|11|沙番 的孙子 基玛利雅 的儿子 米该亚 听见书卷上耶和华的一切话，
JER|36|12|就下到王宫，进入书记的房间。看哪，所有的官长都坐在那里，包括 以利沙玛 文士、 示玛雅 的儿子 第莱雅 、 亚革波 的儿子 以利拿单 、 沙番 的儿子 基玛利雅 、 哈拿尼雅 的儿子 西底家 和其余的官长。
JER|36|13|米该亚 向他们述说他所听见的一切话，就是当 巴录 向众百姓宣读那书卷时亲耳听见的。
JER|36|14|官长们就派 犹底 ，就是 古示 的曾孙， 示利米雅 的孙子， 尼探雅 的儿子到 巴录 那里，对他说：“你把你所念给百姓听的书卷拿在手里，到我们这里来。” 尼利亚 的儿子 巴录 就手拿书卷到他们那里来。
JER|36|15|他们对他说：“请坐下，念给我们亲耳听。” 巴录 就念给他们亲耳听。
JER|36|16|他们听见这一切话就害怕，面面相觑，对 巴录 说：“我们必须将这一切话禀告王。”
JER|36|17|他们问 巴录 说：“请你告诉我们，你怎样从他口中写下这一切话呢？”
JER|36|18|巴录 回答说：“他向我口述这一切话，我就用笔墨把它写在书卷上。”
JER|36|19|众官长对 巴录 说：“你和 耶利米 要去躲起来，不可叫人知道你们躲在哪里。”
JER|36|20|众官长把书卷留在 以利沙玛 文士的房间里，然后进院见王，把这一切话说给王听。
JER|36|21|王就派 犹底 去拿这书卷来；他就从 以利沙玛 文士的房间内取来，念给王和侍立在王左右的众官长亲耳听。
JER|36|22|那时正是九月，王坐在过冬的房屋里，王前面有燃烧的火盆 。
JER|36|23|犹底 念了三、四段 ，王就用文士的刀把书卷割破，丢在火盆里，直到全卷在火中烧尽了。
JER|36|24|王和听见这一切话的臣仆都不惧怕，也不撕裂衣服。
JER|36|25|以利拿单 和 第莱雅 ，并 基玛利雅 恳求王不要烧这书卷，王却不听。
JER|36|26|王吩咐王 的儿子 耶拉篾 、 亚斯列 的儿子 西莱雅 和 亚伯叠 的儿子 示利米雅 ，去捉拿 巴录 文士和 耶利米 先知；耶和华却将他们隐藏起来。
JER|36|27|王烧了有 巴录 从 耶利米 口中所写之话的书卷以后，耶和华的话临到 耶利米 ，说：
JER|36|28|“你再取一书卷，将 犹大 王 约雅敬 所烧前一卷书上原有的一切话写在上面。
JER|36|29|论到 犹大 王 约雅敬 你要说，耶和华如此说：你烧了这书卷，说：‘你为什么在上面写着， 巴比伦 王必要来毁灭这地，使这地绝了人民和牲畜呢？’
JER|36|30|所以耶和华论到 犹大 王 约雅敬 说：他后裔中必没有人坐在 大卫 的宝座上；他的尸首必被抛弃，白天受炎热，黑夜受寒霜。
JER|36|31|我必因他和他后裔，并他臣仆的罪孽惩罚他们。我要使我所说的一切灾祸临到他们和 耶路撒冷 的居民，并 犹大 人；只是他们不肯听从。”
JER|36|32|于是， 耶利米 又取一书卷交给 尼利亚 的儿子 巴录 文士，他就从 耶利米 的口中写了 犹大 王 约雅敬 在火中所烧书卷上的一切话，另外又添了许多相仿的话。
JER|37|1|约西亚 的儿子 西底家 接续 约雅敬 的儿子 哥尼雅 作王，因为 巴比伦 王 尼布甲尼撒 立他在 犹大 地作王。
JER|37|2|但 西底家 、他的臣仆和这地的百姓都不听从耶和华藉 耶利米 先知所说的话。
JER|37|3|西底家 王派 示利米雅 的儿子 犹甲 和 玛西雅 的儿子 西番雅 祭司，去见 耶利米 先知，说：“求你为我们祈求耶和华－我们的上帝。”
JER|37|4|那时 耶利米 仍在百姓中进出，因为他们还没有把他囚在监里。
JER|37|5|法老的军队已经从 埃及 出来，那围困 耶路撒冷 的 迦勒底 人听见这风声，就拔营离开 耶路撒冷 去了。
JER|37|6|耶和华的话临到 耶利米 先知，说：
JER|37|7|“耶和华－ 以色列 的上帝如此说：你们要对派你们来求问我的 犹大 王如此说：‘看哪，那出来帮助你们的法老军队必回 埃及 本国去。
JER|37|8|迦勒底 人必再来攻打这城，并要攻下，用火焚烧。
JER|37|9|耶和华如此说：你们不要自欺说“ 迦勒底 人必定离开我们”，因为他们必不离开。
JER|37|10|你们即使击败与你们争战的 迦勒底 全军，他们当中剩下受伤的人也必各自从帐棚里起来，用火焚烧这城。’”
JER|37|11|迦勒底 的军队因躲避法老的军队，拔营离开 耶路撒冷 的时候，
JER|37|12|耶利米 离开 耶路撒冷 ，往 便雅悯 地去，要在那里从百姓当中取得自己的地产。
JER|37|13|他到了 便雅悯门 ，那里的守门官名叫 伊利雅 ，是 哈拿尼亚 的孙子， 示利米雅 的儿子，他逮捕 耶利米 先知，说：“你是去投降 迦勒底 人的！”
JER|37|14|耶利米 说：“你这是谎话，我并不是去投降 迦勒底 人。” 伊利雅 不听 耶利米 的话，就逮捕他，把他带到官长那里。
JER|37|15|官长们恼怒 耶利米 ，打了他，把他囚在 约拿单 文士的房屋中，因为他们把这屋子当作监牢。
JER|37|16|耶利米 来到地牢，进入牢房，在那里拘留多日。
JER|37|17|西底家 王差人提他出来，在自己的宫内私下问他说：“有什么话从耶和华临到没有？” 耶利米 说：“有！”又说：“你必被交在 巴比伦 王手中。”
JER|37|18|耶利米 又对 西底家 王说：“我在什么事上得罪你，或你的臣仆，或这百姓，你们竟将我囚在监里呢？
JER|37|19|对你们预言‘ 巴比伦 王必不来攻击你们和这地’的先知在哪里呢？
JER|37|20|主－我的王啊，现在求你垂听，允准我在你面前的恳求：不要把我送回 约拿单 文士的房屋中，免得我死在那里。”
JER|37|21|于是 西底家 王下令，他们就把 耶利米 交在护卫兵的院中，每天从饼店街取一个饼给他，直到城中所有的饼都用尽了。这样， 耶利米 仍拘留在护卫兵的院中。
JER|38|1|玛坦 的儿子 示法提雅 、 巴施户珥 的儿子 基大利 、 示利米雅 的儿子 犹甲 、 玛基雅 的儿子 巴示户珥 听见 耶利米 对众百姓所说的话，说：
JER|38|2|“耶和华如此说：留在这城里的必遭刀剑、饥荒、瘟疫而死，但归向 迦勒底 人的必得存活；至少能保全自己的性命，得以存活。
JER|38|3|耶和华如此说：这城必要交在 巴比伦 王军队的手中，他必攻下这城。”
JER|38|4|于是官长们对王说：“求你把这人处死，因他向城里剩下的士兵和众人说这样的话，使他们的手发软。这人不是为这百姓求平安，而是叫他们受灾祸。”
JER|38|5|西底家 王说：“看哪，他在你们手中，王不能反对你们所做的事。”
JER|38|6|他们就拿住 耶利米 ，把他丢在王 的儿子 玛基雅 的井里；那口井在护卫兵的院中。他们用绳子把 耶利米 缒下去，井里没有水，只有淤泥， 耶利米 就陷在淤泥中。
JER|38|7|在王宫里的太监 古实 人 以伯．米勒 ，听见他们把 耶利米 丢进井里，那时王坐在 便雅悯门 前。
JER|38|8|以伯．米勒 从王宫里出来，对王说：
JER|38|9|“主－我的王啊，这些人向 耶利米 先知一味地行恶，把他丢在井里；他在那里必因饥饿而死，因为城里不再有粮食了。”
JER|38|10|王就吩咐 古实 人 以伯．米勒 说：“你从这里带领三十人，趁 耶利米 先知还没死，把他从井里拉上来。”
JER|38|11|于是 以伯．米勒 带领这些人同去，进入王宫，到库房以下 ，从那里取了些碎布和破衣服，用绳子缒下去，到井里 耶利米 那里。
JER|38|12|古实 人 以伯．米勒 对 耶利米 说：“你用这些碎布和破衣服放在绳子上，垫你的腋下。” 耶利米 就照样做。
JER|38|13|这样，他们用绳子将 耶利米 从井里拉上来。 耶利米 仍在护卫兵的院中。
JER|38|14|西底家 王差人将 耶利米 先知带进耶和华殿的第三个门，到王那里去。王对 耶利米 说：“我要问你一件事，你一点都不可向我隐瞒。”
JER|38|15|耶利米 对 西底家 说：“我若告诉你，你岂不是一定要把我处死吗？我若劝你，你必不听我。”
JER|38|16|西底家 王就私下对 耶利米 说：“我指着那造我们生命之永生的耶和华起誓：我必不把你处死，也不将你交在寻索你命的人手中。”
JER|38|17|耶利米 对 西底家 说：“耶和华－万军之上帝、 以色列 的上帝如此说：你若归顺 巴比伦 王的官长，你的命就必存活，这城也不致被火焚烧，你和你的全家都必存活。
JER|38|18|你若不归顺 巴比伦 王的官长，这城必交在 迦勒底 人手中。他们必用火焚烧，你也不得脱离他们的手。”
JER|38|19|西底家 王对 耶利米 说：“我怕那些投降 迦勒底 人的 犹大 人，恐怕 迦勒底 人把我交在他们手中，他们就戏弄我。”
JER|38|20|耶利米 说：“ 迦勒底 人必不把你交出。求你听从我对你所说耶和华的话，这样对你有好处，你的命也必存活。
JER|38|21|你若不肯归顺，耶和华指示我的话是这样：
JER|38|22|看哪， 犹大 王宫里所留下来的妇女必被带到 巴比伦 王的官长那里。这些妇女要说： 你知己的朋友引诱你， 他们胜过你； 你的脚陷入淤泥， 他们却离弃你。
JER|38|23|“人必将你的后妃和你的儿女带到 迦勒底 人那里；你也不得脱离他们的手，必被 巴比伦 王的手捉住，这城也必被火焚烧 。”
JER|38|24|西底家 对 耶利米 说：“不要让人知道这些对话，你就不至于死。
JER|38|25|官长们若听见我跟你说话，到你那里对你说：‘告诉我们，你对王说了什么话，王又向你说了什么；不可向我们隐瞒，否则我们就要杀你。’
JER|38|26|你就对他们说：‘我在王面前恳求不要把我送回 约拿单 的房屋，免得我死在那里。’”
JER|38|27|随后官长们到 耶利米 那里，问他，他就照王所吩咐的一切话回答他们。他们就不再问他，因为事情没有泄漏。
JER|38|28|于是 耶利米 仍在护卫兵的院中，直到 耶路撒冷 被攻下的日子。当 耶路撒冷 被攻下时，他仍在那里。
JER|39|1|犹大 王 西底家 第九年十月， 巴比伦 王 尼布甲尼撒 率领全军前来围困 耶路撒冷 。
JER|39|2|西底家 十一年四月初九日，城被攻破。
JER|39|3|耶路撒冷 被攻下的时候， 巴比伦 王的众官长， 尼甲．沙利薛 、 三甲．尼波 、 撒西金 将军 、 尼甲．沙利薛 将军 ，并 巴比伦 王其余的官长都来坐在 中门 。
JER|39|4|犹大 王 西底家 和所有士兵看见他们，就在夜间从靠近王的花园、两城墙中间的门逃跑出城，往 亚拉巴 逃去。
JER|39|5|迦勒底 的军队追赶他们，在 耶利哥 的平原追上 西底家 ，将他逮住，带到 哈马 地的 利比拉 、 巴比伦 王 尼布甲尼撒 那里； 尼布甲尼撒 就判他的罪。
JER|39|6|在 利比拉 ， 巴比伦 王在 西底家 眼前杀了他的儿女； 巴比伦 王又杀了 犹大 所有的贵族，
JER|39|7|并且挖了 西底家 的眼睛，用铜链锁住他，要带到 巴比伦 去。
JER|39|8|迦勒底 人用火焚烧王宫和百姓的房屋，又拆毁 耶路撒冷 的城墙。
JER|39|9|那时， 尼布撒拉旦 护卫长把城里所剩下的百姓和投降他的降民，以及其余的百姓都掳到 巴比伦 去了。
JER|39|10|尼布撒拉旦 护卫长却把百姓中一无所有的穷人留在 犹大 地，当时就赏给他们葡萄园和田地 。
JER|39|11|巴比伦 王 尼布甲尼撒 为了 耶利米 ，嘱咐 尼布撒拉旦 护卫长：
JER|39|12|“你领他去，好好地看待他，切不可害他；他对你怎么说，你就向他怎样做。”
JER|39|13|尼布撒拉旦 护卫长和 尼布沙斯班 将军 、 尼甲．沙利薛 将军 ，并 巴比伦 王众官长，
JER|39|14|派人把 耶利米 从护卫兵的院中提出来，交给 沙番 的孙子， 亚希甘 的儿子 基大利 ，让他自由进出屋子；于是 耶利米 住在百姓中间。
JER|39|15|耶利米 还囚在护卫兵院中的时候，耶和华的话临到他，说：
JER|39|16|“你去告诉 古实 人 以伯．米勒 说，万军之耶和华－ 以色列 的上帝如此说：看哪，我说降祸不降福的话必临到这城，到那时必在你面前实现。
JER|39|17|到那日我必拯救你，你必不致交在你所怕的人手中。这是耶和华说的。
JER|39|18|我定要搭救你，你必不致倒在刀下，却要保全自己的性命，因你倚靠我。这是耶和华说的。”
JER|40|1|耶利米 被链子锁在 耶路撒冷 和 犹大 被掳到 巴比伦 的人中， 尼布撒拉旦 护卫长把他从 拉玛 提出来，释放他以后，耶和华的话临到 耶利米 。
JER|40|2|护卫长提 耶利米 来，对他说：“耶和华－你的上帝曾说要降这灾祸给此地。
JER|40|3|耶和华照他所说的做了，已使这灾祸临到；因你们得罪耶和华，不听从他的话，所以这事临到你们。
JER|40|4|看哪，现在我解开你手上的链子，你若看与我同往 巴比伦 去好，就可以去，我必厚待你；你若看与我同往 巴比伦 去不好，就不必去。看哪，全地在你面前，你以为哪里美好，哪里合宜，只管去吧
JER|40|5|─ 耶利米 尚未回去 ─你可以回到 巴比伦 王所立管理 犹大 城镇的 沙番 的孙子， 亚希甘 的儿子 基大利 那里去，在他那里住在百姓当中。不然，你看哪里合宜就可以去。”于是护卫长送他粮食和礼物，释放了他。
JER|40|6|耶利米 就来到 米斯巴 ， 亚希甘 的儿子 基大利 那里去，与他同住，住在留于境内的百姓当中。
JER|40|7|在乡间所有的军官和属他们的人，听见 巴比伦 王立了 亚希甘 的儿子 基大利 作当地的省长，并将没有掳到 巴比伦 的男人、妇女、孩童和当地极穷的人全交给他，
JER|40|8|于是 尼探雅 的儿子 以实玛利 ， 加利亚 的两个儿子 约哈难 和 约拿单 ， 单户篾 的儿子 西莱雅 ，并 尼陀法 人 以斐 的众子， 玛迦 人的儿子 耶撒尼亚 ，和属他们的人，都来到 米斯巴 的 基大利 那里。
JER|40|9|沙番 的孙子， 亚希甘 的儿子 基大利 向他们和属他们的人起誓说：“不要怕服事 迦勒底 人，只管住在这地，服事 巴比伦 王，就可以得福。
JER|40|10|至于我，我要住在 米斯巴 ，侍候那些到我们这里来的 迦勒底 人；只是你们当积蓄酒、油和夏天的果子，收藏在器皿里，并住在你们所占的城镇中。”
JER|40|11|在 摩押 地和 亚扪 人当中，在 以东 地和各国，所有的 犹大 人听见 巴比伦 王留下一些 犹大 人，并立 沙番 的孙子、 亚希甘 的儿子 基大利 管理他们，
JER|40|12|所有的 犹大 人就从被赶到的各处回来，到 犹大 地 米斯巴 的 基大利 那里。他们积蓄了许多的酒，并夏天的果子。
JER|40|13|加利亚 的儿子 约哈难 和在乡间的军官来到 米斯巴 的 基大利 那里，
JER|40|14|对他说：“ 亚扪 人的王 巴利斯 派 尼探雅 的儿子 以实玛利 来谋害你的命，你知道吗？” 亚希甘 的儿子 基大利 却不相信他们的话。
JER|40|15|加利亚 的儿子 约哈难 在 米斯巴 私下对 基大利 说：“求你容我去杀 尼探雅 的儿子 以实玛利 ，必无人知道。何必让他害你的命，使聚集到你这里来的 犹大 人都分散，以致 犹大 剩余的人都灭亡呢？”
JER|40|16|亚希甘 的儿子 基大利 对 加利亚 的儿子 约哈难 说：“你不可做这事，你所论 以实玛利 的话是假的。”
JER|41|1|七月中，王的大臣，就是王室后裔 以利沙玛 的孙子、 尼探雅 的儿子 以实玛利 带着十个人，来到 米斯巴 ， 亚希甘 的儿子 基大利 那里；他们在 米斯巴 一同吃饭。
JER|41|2|尼探雅 的儿子 以实玛利 和同他来的那十个人起来，用刀击杀 沙番 的孙子， 亚希甘 的儿子 基大利 ，就是 巴比伦 王所立为当地省长的，把他杀死。
JER|41|3|以实玛利 把所有在 米斯巴 与 基大利 一起的 犹大 人，以及他们在那里所遇见的 迦勒底 人和士兵都杀了。
JER|41|4|他杀了 基大利 的第二天，还没有人知道的时候，
JER|41|5|有八十人从 示剑 、 示罗 和 撒玛利亚 前来，胡须剃去，衣服撕裂，身体划破，手拿素祭和乳香，要奉到耶和华的殿。
JER|41|6|尼探雅 的儿子 以实玛利 从 米斯巴 出来迎接他们，随走随哭，遇见了他们，就对他们说：“你们可以到 亚希甘 的儿子 基大利 那里。”
JER|41|7|他们到了城中， 尼探雅 的儿子 以实玛利 和与他一起的人就把他们杀了，丢在坑里。
JER|41|8|只是他们中间有十个人对 以实玛利 说：“不要杀我们，因为我们有许多大麦、小麦、油和蜜藏在田间。”于是他住手，没有在弟兄中间杀他们。
JER|41|9|以实玛利 把那些因 基大利 事件所杀之人的尸首都丢在坑里；这坑是从前 亚撒 王因怕 以色列 王 巴沙 所挖的。 尼探雅 的儿子 以实玛利 把那些被杀的人填满了坑。
JER|41|10|以实玛利 把 米斯巴 剩下的人，就是众公主和仍住在 米斯巴 所有的百姓都掳去，他们原是 尼布撒拉旦 护卫长交给 亚希甘 的儿子 基大利 的。 尼探雅 的儿子 以实玛利 掳了他们，要到 亚扪 人那里去。
JER|41|11|加利亚 的儿子 约哈难 和与他一起的军官，听见 尼探雅 的儿子 以实玛利 所做的一切恶事，
JER|41|12|就带领众人前往，要和 尼探雅 的儿子 以实玛利 争战，他们在 基遍 的大水池 旁遇见他。
JER|41|13|在 以实玛利 那里的众人看见 加利亚 的儿子 约哈难 和与他一起的军官，就都欢喜。
JER|41|14|这样， 以实玛利 从 米斯巴 所掳去的众人都转而归向 加利亚 的儿子 约哈难 。
JER|41|15|尼探雅 的儿子 以实玛利 和八个人脱离 约哈难 的手，逃到 亚扪 人那里去。
JER|41|16|尼探雅 的儿子 以实玛利 杀了 亚希甘 的儿子 基大利 ，从 米斯巴 把所有幸存的百姓、士兵、妇女、孩童、太监掳到 基遍 之后， 加利亚 的儿子 约哈难 和与他一起的军官把他们都抢回来，
JER|41|17|带到靠近 伯利恒 的 基罗特金罕 住下，要到 埃及 去，
JER|41|18|躲避 迦勒底 人。他们惧怕 迦勒底 人，因为 尼探雅 的儿子 以实玛利 杀了 巴比伦 王所立管理那地的 亚希甘 的儿子 基大利 。
JER|42|1|众军官和 加利亚 的儿子 约哈难 ，并 何沙雅 的儿子 耶撒尼亚 以及众百姓，从最小的到最大的都进前来，
JER|42|2|对 耶利米 先知说：“请你准我们在你面前祈求，为我们这幸存的人向耶和华－你的上帝祷告。我们本来众多，现在剩下的极少，这是你亲眼看见的。
JER|42|3|愿耶和华－你的上帝指示我们当走的路，当做的事。”
JER|42|4|耶利米 先知对他们说：“我已经听见了，看哪，我必照你们的话向耶和华－你们的上帝祷告。耶和华无论回答什么，我都必告诉你们，绝不隐瞒。”
JER|42|5|于是他们对 耶利米 说：“我们若不照耶和华－你上帝差遣你说的一切话去做，愿耶和华在我们中间作真实可靠的见证。
JER|42|6|我们请你到耶和华－我们的上帝面前，他说的无论是好是歹，我们都必听从；因为我们听从耶和华－我们上帝的话，就可以得福。”
JER|42|7|过了十天，耶和华的话临到 耶利米 。
JER|42|8|他就将 加利亚 的儿子 约哈难 和与他一起所有的军官和百姓，从最小的到最大的都召来，
JER|42|9|对他们说：“你们请我到耶和华－ 以色列 的上帝面前为你们祈求，他如此说：
JER|42|10|‘你们若仍留在这地，我就建立你们，必不拆毁；栽植你们，必不拔出；因我为所降与你们的灾祸感到遗憾。
JER|42|11|不要怕你们所惧怕的 巴比伦 王。不要怕他！因为我与你们同在，要拯救你们脱离他的手。这是耶和华说的。
JER|42|12|我要向你们施怜悯，他 就怜悯你们，使你们归回本地。’
JER|42|13|倘若你们说：‘我们不留在这地’，不听从耶和华－你们上帝的话，
JER|42|14|说：‘我们不留在这地，却要进入 埃及 地，在那里我们看不见战争，听不见角声，也不致缺食挨饿；我们要住在那里。’
JER|42|15|幸存的 犹大 人哪，你们现在要听耶和华的话；万军之耶和华－ 以色列 的上帝如此说：‘你们若定意进入 埃及 ，在那里寄居，
JER|42|16|你们所惧怕的刀剑在 埃及 地必追上你们，你们所惧怕的饥荒在 埃及 要紧紧跟随你们，你们必死在那里。
JER|42|17|凡定意进入 埃及 在那里寄居的，必遭刀剑、饥荒、瘟疫而死，无一人存留，得以逃脱我所降与他们的灾祸。’
JER|42|18|“万军之耶和华－ 以色列 的上帝如此说：‘我怎样将我的怒气和愤怒倾倒在 耶路撒冷 的居民身上，你们进入 埃及 的时候，我也必照样将我的愤怒倾倒在你们身上，以致你们受辱骂、惊骇、诅咒、羞辱，并且不得再看见这地方。’
JER|42|19|幸存的 犹大 人哪，耶和华论到你们说：‘不要进入 埃及 。’你们要确实知道，我今日已警戒你们了。
JER|42|20|你们行诡诈害自己；因为你们请我到耶和华－你们上帝那里，说：‘请你为我们向耶和华－我们的上帝祷告，你把耶和华－我们上帝所说的一切告诉我们，我们就必遵行。’
JER|42|21|我今日把这话告诉你们，你们却不听耶和华－你们上帝为这一切事差我到你们那里所说的话。
JER|42|22|现在你们要确实知道，你们在所要去的寄居之地必遭刀剑、饥荒、瘟疫而死。”
JER|43|1|耶利米 向众百姓说完了耶和华－他们上帝一切的话，就是耶和华－他们上帝差他去说的这一切话，
JER|43|2|何沙雅 的儿子 亚撒利雅 和 加利亚 的儿子 约哈难 ，以及所有狂傲的人，就对 耶利米 说：“你说谎！耶和华－我们的上帝并没有差遣你说：‘你们不可进入 埃及 ，在那里寄居。’
JER|43|3|这是 尼利亚 的儿子 巴录 挑唆你害我们，要把我们交在 迦勒底 人手中，使我们被杀或被掳到 巴比伦 去。”
JER|43|4|加利亚 的儿子 约哈难 和所有的军官、百姓，都不肯听从耶和华的话留在 犹大 地。
JER|43|5|加利亚 的儿子 约哈难 和所有的军官却将幸存的 犹大 人，就是从被赶到的各国回来，在 犹大 地寄居的男人、妇女、孩童和众公主，并 尼布撒拉旦 护卫长留在 沙番 的孙子， 亚希甘 的儿子 基大利 那里的众人，与 耶利米 先知，以及 尼利亚 的儿子 巴录 ，
JER|43|6|
JER|43|7|都带入 埃及 地，到了 答比匿 ；这是因他们不肯听从耶和华的话。
JER|43|8|在 答比匿 ，耶和华的话临到 耶利米 ，说：
JER|43|9|“你要在 犹大 人眼前用手拿几块大石头，藏在 答比匿 法老的宫门砌砖的石墩上，
JER|43|10|对他们说：‘万军之耶和华－ 以色列 的上帝如此说：看哪，我必召我的仆人 巴比伦 王 尼布甲尼撒 前来，安置他的宝座在所藏的这些石头上；他要在其上支搭华丽的帐幕。
JER|43|11|他要来攻击 埃及 地： 定为死亡的，必致死亡； 定为掳掠的，必遭掳掠； 定为刀杀的，必被刀杀。
JER|43|12|我要用火点燃 埃及 众神明的庙宇， 巴比伦 王要焚烧庙宇，掳去神像；他要围住 埃及 地，好像牧人披上外衣，从那里安然而去。
JER|43|13|他必打碎 埃及 地 伯．示麦 的柱像，用火焚烧 埃及 众神明的庙宇。’”
JER|44|1|有话临到 耶利米 ，论到住 埃及 地所有的 犹大 人，就是住在 密夺 、 答比匿 、 挪弗 、 巴特罗 境内的 犹大 人，说：
JER|44|2|“万军之耶和华－ 以色列 的上帝如此说：我所降与 耶路撒冷 和 犹大 各城的一切灾祸，你们都看见了。看哪，那些城镇今日荒凉，无人居住；
JER|44|3|这是因居民所行的恶，去烧香事奉别神，就是他们和你们，以及你们列祖所不认识的神明，惹我发怒。
JER|44|4|我一再差遣我的仆人众先知去，说：你们切不可行我所厌恶这可憎之事。
JER|44|5|他们却不听从，不侧耳而听，也不转离恶事，仍向别神烧香。
JER|44|6|因此，我的怒气和愤怒都倾倒出来，在 犹大 城镇和 耶路撒冷 街市上燃起，以致它们都荒废凄凉，正如今日一样。
JER|44|7|现在耶和华－万军之上帝、 以色列 的上帝如此说：你们为何做这大恶自害己命，使你们的男人、妇女、孩童和吃奶的都从 犹大 剪除，不留一人呢？
JER|44|8|你们以手所做的，在寄居的 埃及 地向别神烧香，惹我发怒，使你们被剪除，在天下万国中受诅咒羞辱。
JER|44|9|你们祖先的恶行， 犹大 诸王和后妃的恶行，你们自己和你们妻子的恶行，就是在 犹大 地和 耶路撒冷 街市上所做的，你们都忘了吗？
JER|44|10|到如今你们还不懊悔，不惧怕，不肯遵行我在你们和你们祖先面前所设立的法度律例。
JER|44|11|“所以万军之耶和华－ 以色列 的上帝如此说：看哪，我必向你们变脸降灾，剪除 犹大 众人。
JER|44|12|我必使那定意进入 埃及 地、在那里寄居的，就是幸存的 犹大 人，尽都灭绝。他们必在 埃及 地仆倒，因刀剑饥荒灭绝，从最小的到最大的都必遭刀剑饥荒而死，甚至受辱骂、惊骇、诅咒、羞辱。
JER|44|13|我怎样用刀剑、饥荒、瘟疫惩罚 耶路撒冷 ，也必照样惩罚那些住在 埃及 地的 犹大 人。
JER|44|14|那进入 埃及 地、在那里寄居的，就是幸存的 犹大 人，都不得逃脱，也不得归回 犹大 地。他们心中很想归回，居住在那里；但除了少数逃脱的以外，都不得归回。”
JER|44|15|那些知道自己妻子向别神烧香的男人，与站在那里的一大群妇女，就是住 埃及 地 巴特罗 所有的百姓，回答 耶利米 说：
JER|44|16|“论到你奉耶和华的名向我们所说的话，我们必不听从。
JER|44|17|我们定要照我们口中所说的一切话去做，向天后烧香，献浇酒祭，按着我们与我们祖先、君王、官长在 犹大 城镇和 耶路撒冷 街市上素常所做的一样；因为那时我们得以吃饱、享福乐，并未遇见灾祸。
JER|44|18|自从我们停止向天后烧香，献浇酒祭，我们倒缺乏这一切，又因刀剑饥荒灭绝。”
JER|44|19|妇女们说 ：“我们向天后烧香，献浇酒祭，做天后像的饼供奉它，向它献浇酒祭，难道我们的丈夫没有参与吗？”
JER|44|20|耶利米 对这样回答他的男人和妇女说：
JER|44|21|“你们与你们祖先、君王、官长，以及这地的百姓，在 犹大 城镇和 耶路撒冷 街市上所烧的香，耶和华岂不记得，放在他心上吗？
JER|44|22|耶和华因你们所行的恶、所做可憎的事，不能再容忍，所以使你们的地荒凉，受惊骇诅咒，无人居住，正如今日一样。
JER|44|23|你们烧香，得罪耶和华，不听耶和华的话，不遵行他的律法、条例、法度，所以你们遭遇这灾祸，正如今日一样。”
JER|44|24|耶利米 又对众百姓和妇女说：“所有在 埃及 地的 犹大 人哪，当听耶和华的话。
JER|44|25|万军之耶和华－ 以色列 的上帝如此说：你们和你们的妻子口中说过、手里做到，说：‘我们定要向天后还愿，向它烧香，献浇酒祭。’现在你们尽管坚定所许的愿，去还愿吧！
JER|44|26|所有住 埃及 地的 犹大 人哪，当听耶和华的话。耶和华说：看哪，我指着我至大的名起誓，在 埃及 全地，我的名必不再被 犹大 任何人的口呼喊：‘我指着主－永生的耶和华起誓。’
JER|44|27|看哪，我看守他们，为要降祸不降福；在 埃及 地的 犹大 人必因刀剑、饥荒而灭亡，直到灭绝。
JER|44|28|从 埃及 地能脱离刀剑、归回 犹大 地的人数很少。那进入 埃及 地、在那里寄居的，就是幸存的 犹大 人，必知道是谁的话站得住，是我的话呢，还是他们的话。
JER|44|29|我在这地方惩罚你们，必有预兆，使你们知道我降祸给你们的话必站得住。这是耶和华说的。
JER|44|30|耶和华如此说：看哪，我必将 埃及 王 合弗拉 法老交在他仇敌和寻索其命的人手中，像我将 犹大 王 西底家 交在他仇敌和寻索其命的 巴比伦 王 尼布甲尼撒 手中一样。”
JER|45|1|约西亚 的儿子 犹大 王 约雅敬 第四年， 尼利亚 的儿子 巴录 把 耶利米 先知口中所说的话写在书上； 耶利米 对 巴录 说：
JER|45|2|“ 巴录 啊，耶和华－ 以色列 的上帝说：
JER|45|3|你曾说：‘哀哉！耶和华使我愁上加愁，我因呻吟而困乏，不得安歇。’
JER|45|4|你要这样告诉他，耶和华如此说：看哪，我所建立的，我必拆毁；我所栽植的，我必拔出；在全地我都如此行。
JER|45|5|你为自己图谋大事吗？不要图谋！看哪，我必使灾祸临到凡有血肉之躯的。但你无论往哪里去，我要保全你的性命。这是耶和华说的。”
JER|46|1|耶和华论列国的话临到 耶利米 先知。
JER|46|2|论到 埃及 ，关于 埃及 王 尼哥 法老的军队，这军队安营在 幼发拉底河 边的 迦基米施 ，是 巴比伦 王 尼布甲尼撒 在 约西亚 的儿子 犹大 王 约雅敬 第四年所打败的。
JER|46|3|你们要预备大小盾牌， 往前上阵，
JER|46|4|套上车， 骑上马！ 顶盔站立， 磨枪披甲！
JER|46|5|我为何看见他们惊惶， 转身退后呢？ 他们的勇士打败仗， 急忙逃跑，并不回头； 四围都有惊吓！ 这是耶和华说的。
JER|46|6|不要容快跑的逃避， 也不要容勇士逃脱 ； 在北方 幼发拉底河 边， 他们绊跌仆倒。
JER|46|7|这是谁，像 尼罗河 涨溢， 如江河的水翻腾呢？
JER|46|8|埃及 像 尼罗河 涨溢， 如江河的水翻腾。 它说：“我要涨溢遮盖全地； 我要毁灭城镇和其中的居民。
JER|46|9|马匹啊，上去吧！ 战车啊，要疾行！ 手拿盾牌的 古实 和 弗 的勇士， 擅长拉弓的 路德 人，前进吧！”
JER|46|10|那日是万军之主耶和华报仇的日子， 要向敌人报仇。 刀剑必吞吃饱足， 饮血满足； 因为在北方 幼发拉底河 边， 有祭物献给万军之主耶和华。
JER|46|11|少女 埃及 啊， 要上 基列 去取乳香； 你虽服用许多药， 还是徒然，不得治好。
JER|46|12|列国听见你的羞辱， 遍地满了你的哀声； 勇士与勇士彼此相撞， 二人一起跌倒。
JER|46|13|以下是耶和华对 耶利米 先知说的话，论到 巴比伦 王 尼布甲尼撒 要来攻击 埃及 地。
JER|46|14|你们要在 埃及 传扬，在 密夺 报告， 在 挪弗 、 答比匿 宣告说： “要摆好阵势，预备作战， 因为刀剑在你四围施行吞灭。”
JER|46|15|你的壮士为何被扫除呢？ 他们站立不住， 因为耶和华驱逐他们；
JER|46|16|他使多人绊跌，彼此撞倒。 他们说：“起来，让我们回到自己的同胞、 回到自己的出生地去， 好躲避欺压的刀剑。”
JER|46|17|他们在那里称 埃及 王法老 为 “错失良机的夸大者”。
JER|46|18|名为万军之耶和华的君王说： 我指着我的永生起誓： “ 尼布甲尼撒 来的时候， 必像众山之中的 他泊 ， 像海边的 迦密 。”
JER|46|19|住在 埃及 的啊， 要预备被掳时需用的物品； 因为 挪弗 必成为废墟， 被烧毁，无人居住。
JER|46|20|埃及 是肥美的母牛犊； 但来自北方的牛虻来到了！来到了！
JER|46|21|它的佣兵好像圈里的肥牛犊， 他们转身退后， 一齐逃跑，站立不住； 因为他们遭难的日子、 受罚的时刻已经来临。
JER|46|22|它的声音好像蛇在滑行。 敌人要成队而来，如砍伐树木的人， 手拿斧头攻击它。
JER|46|23|虽然它的树林不易穿过， 敌人却要砍伐， 因敌人比蝗虫还多，不可胜数。 这是耶和华说的。
JER|46|24|埃及 必然蒙羞， 被交在北方人的手中。
JER|46|25|万军之耶和华－ 以色列 的上帝说：“看哪，我要惩罚 挪 的 亚扪 和法老、 埃及 和它的神明，以及君王，也要惩罚法老和倚靠他的人。
JER|46|26|我要将他们交给寻索其命之人的手和 巴比伦 王 尼布甲尼撒 与他臣仆的手。但 埃及 日后必再有人居住，与从前一样。这是耶和华说的。”
JER|46|27|我的仆人 雅各 啊，不要惧怕！ 以色列 啊，不要惊惶！ 因我要从远方拯救你， 从被掳之地拯救你的后裔。 雅各 必回来，得享平静安逸， 无人令他害怕。
JER|46|28|我的仆人 雅各 啊，不要惧怕！ 因我与你同在。 我要将那些国灭绝净尽， 就是我赶你去的那些国； 却不将你灭绝净尽， 倒要从宽惩治你， 但绝不能不罚你。 这是耶和华说的。
JER|47|1|在法老攻击 迦萨 之前，耶和华论 非利士 人的话临到 耶利米 先知。
JER|47|2|耶和华如此说： 看哪，有水从北方涨起，成为涨溢的河， 要淹没全地和其中所充满的， 淹没城和城里的居民。 人必呼喊， 境内的居民都必哀号。
JER|47|3|一听见敌人壮马蹄踏的响声、 战车隆隆、车轮轰轰， 为父的手就发软， 不能回头看顾儿女。
JER|47|4|因为日子将到， 耶和华必毁灭所有 非利士 人， 剪除 推罗 、 西顿 仅存的帮助者； 他要毁灭 非利士 人、 迦斐托 海岛剩余的人。
JER|47|5|迦萨 成了光秃， 亚实基伦 归于无有。 平原 中所剩的啊， 你割划自己，要到几时呢？
JER|47|6|耶和华的刀剑哪，你要到几时才止息呢？ 要入鞘，安静不动。
JER|47|7|耶和华吩咐它攻击 亚实基伦 和海边之地， 既已派定它，你 怎能静止不动呢？
JER|48|1|论 摩押 。 万军之耶和华－ 以色列 的上帝如此说： 祸哉， 尼波 ！它要变为废墟。 基列亭 蒙羞被攻取， 米斯迦 蒙羞被毁坏，
JER|48|2|摩押 不再被称赞。 有人在 希实本 设计谋害它： “来吧！我们将它剪除，使它不再成国。” 玛得缅 哪，你也必静默无声； 刀剑必追赶你。
JER|48|3|从 何罗念 有哀号声： “荒凉！大毁灭！”
JER|48|4|“ 摩押 毁灭了！” 它的孩童哀号，使人听见。
JER|48|5|人上 鲁希坡 随走随哭， 因为在 何罗念 的下坡听见毁灭的哀声。
JER|48|6|你们要奔逃，自救己命， 使你们的性命如旷野里的矮树 。
JER|48|7|你因倚靠自己所做的 和自己的财宝，必被攻取。 基抹 和属它的祭司、官长也要一同被掳去。
JER|48|8|那行毁灭的要来到各城， 并无一城幸免。 山谷必败落， 平原必毁坏， 正如耶和华所说的。
JER|48|9|你们要将翅膀给 摩押 ， 使它可以飞去 。 它的城镇必荒凉， 无人居住。
JER|48|10|懒惰不肯为耶和华做事的，必受诅咒；禁止刀剑不见血的，必受诅咒。
JER|48|11|摩押 自幼年以来常享安逸， 如沉淀未被搅动的酒 ， 没有从这器皿倒在那器皿， 也未曾被掳掠过。 因此，它的原味尚存， 香气未变。
JER|48|12|看哪，日子将到，我必差倒酒的到它那里去，将它倒出来；他们要倒空器皿，打碎坛子。这是耶和华说的。
JER|48|13|摩押 必因 基抹 羞愧，像 以色列 家因倚靠 伯特利 羞愧一样。
JER|48|14|你们怎么说： “我们是勇士，是会打仗的壮士”呢？
JER|48|15|摩押 变为废墟， 敌人上去占它的城镇。 它精良的壮丁都下去遭杀戮； 这是名为万军之耶和华的君王说的。
JER|48|16|摩押 的灾殃临近， 灾难速速来到。
JER|48|17|凡在它四围的和认识它名的， 都要为它悲伤，说： 那结实的杖和美好的棍， 竟然折断了！
JER|48|18|底本 的居民哪， 要从你荣耀的座位上下来， 坐着忍受干渴； 因毁灭 摩押 的人上来攻击你， 毁坏了你的堡垒。
JER|48|19|住 亚罗珥 的啊， 要站在道路的边上观望， 问逃跑的男人和逃脱的女人说： “发生了什么事呢”？
JER|48|20|摩押 因毁坏蒙羞； 你们要哀号呼喊， 要在 亚嫩 报告： “ 摩押 已成废墟！”
JER|48|21|审判临到平原之地的 何伦 、 雅杂 、 米法押 、
JER|48|22|底本 、 尼波 、 伯．低比拉太音 、
JER|48|23|基列亭 、 伯．迦末 、 伯．米恩 、
JER|48|24|加略 、 波斯拉 和 摩押 地远近所有的城镇。
JER|48|25|摩押 的角砍断了，膀臂折断了。这是耶和华说的。
JER|48|26|你们要使 摩押 沉醉，因它向耶和华夸大。它要在自己所吐之物中打滚，又要被人嗤笑。
JER|48|27|以色列 不是你的笑柄吗？它难道是在贼中被逮到，使你每逢提到它就摇头的吗？
JER|48|28|摩押 的居民哪， 要离开城镇，住在山崖里， 像鸽子在峡谷口上搭窝。
JER|48|29|我们听闻 摩押 人的骄傲， 极其骄傲； 他们自高、自傲、 自我狂妄、居心自大。
JER|48|30|我知道他们的愤怒是虚空的， 他们夸大的话一无所成。 这是耶和华说的。
JER|48|31|因此，我要为 摩押 哀号， 为 摩押 全地呼喊； 人必为 吉珥．哈列设 人叹息。
JER|48|32|西比玛 的葡萄树啊，我为你哀哭， 甚于 雅谢 人的哀哭。 你的枝子蔓延过海， 直伸到 雅谢海 。 那行毁灭的已经临到你夏天的果子和葡萄。
JER|48|33|肥田和 摩押 地的欢喜快乐都被夺去， 我使酒池不再流出酒来， 无人踹酒欢呼； 呼喊的声音不再是欢呼。
JER|48|34|有哀声从 希实本 达到 以利亚利 ，他们发的哀声达到 雅杂 ；从 琐珥 达到 何罗念 ，达到 伊基拉．施利施亚 ，因为 宁林 的水必然干涸。
JER|48|35|我必在 摩押 地使那在丘坛献祭的，和那向他的神明烧香的都灭绝了。这是耶和华说的。
JER|48|36|因此，我的心为 摩押 哀鸣如箫，我的心为 吉珥．哈列设 人哀哭； 摩押 人所得的财物都毁灭了。
JER|48|37|各人头上光秃，胡须剪短，手有划伤，腰束麻布。
JER|48|38|在 摩押 的各房顶上和街市上到处有人哀哭，因我打碎 摩押 ，好像打碎无人喜爱的器皿。这是耶和华说的。
JER|48|39|打得粉碎了！他们要哀号了！ 摩押 要羞愧转背了！这样， 摩押 必受四围的人嗤笑惊骇。
JER|48|40|耶和华如此说： 看哪，仇敌必如鹰展翅快飞， 攻击 摩押 。
JER|48|41|加略 被攻取，堡垒也被占据。 到那日， 摩押 的勇士心中疼痛如临产的妇人。
JER|48|42|摩押 必被毁灭，不再成国， 因它向耶和华夸大。
JER|48|43|摩押 的居民哪， 惊吓、陷阱、罗网都临近你。 这是耶和华说的。
JER|48|44|躲过惊吓的必坠入陷阱， 逃离陷阱的又被罗网缠住， 因我必使惩罚之年临到 摩押 。 这是耶和华说的。
JER|48|45|逃难的人站在 希实本 的荫下，筋疲力尽， 因为有火从 希实本 发出， 有火焰出自 西宏 ， 烧尽 摩押 的鬓角和闹哄人的头顶。
JER|48|46|摩押 啊，你有祸了！ 属 基抹 的百姓灭亡了！ 因你的儿子都被掳去， 你的女儿也被掳去。
JER|48|47|到末后，我却要使 摩押 被掳的人归回。 摩押 受审判的话到此为止。 这是耶和华说的。
JER|49|1|论 亚扪 人。 耶和华如此说： 以色列 没有儿子吗？ 没有后嗣吗？ 米勒公 为何承受 迦得 为业呢？ 属它的百姓为何住其中的城镇呢？
JER|49|2|看哪，日子将到，我必使人听见打仗的喊声， 攻击 亚扪 人所住的 拉巴 的喊声。 拉巴 要成为废墟， 属它的乡镇 要被火焚烧。 这是耶和华说的。 先前承受 以色列 为业的， 此时 以色列 倒要承受他们为业。 这是耶和华说的。
JER|49|3|希实本 哪，要哀号， 因为 爱 地已成荒地。 拉巴 的乡镇哪，要呼喊， 以麻布束腰； 要哭号，在篱笆中往来奔跑； 因 米勒公 和它的祭司、 官长要一同被掳去。
JER|49|4|背道的民 哪， 你为何因有山谷， 因有水流的山谷夸耀呢？ 为何倚靠自己的财宝，说： “谁能来到我们这里呢？”
JER|49|5|万军之主耶和华说： 看哪，我要使惊吓从四围的邻邦临到你们； 你们必被赶出， 各人一直往前， 无人收容难民。
JER|49|6|但后来，我却要使被掳的 亚扪 人归回。这是耶和华说的。
JER|49|7|论 以东 。 万军之耶和华如此说： 提幔 不再有智慧了吗？ 聪明人的谋略都用尽了吗？ 他们的智慧尽归无有了吗？
JER|49|8|底但 的居民哪，要转身逃跑， 住在深密处； 因为我惩罚 以扫 的时候， 必使灾殃临到他。
JER|49|9|摘葡萄的若来到你那里， 岂不留下几串吗？ 贼若夜间来到， 岂不是只毁坏他们要毁坏的吗？
JER|49|10|我却使 以扫 赤裸， 暴露他的藏身处； 他不能隐藏自己。 他的后裔、弟兄、邻舍全都灭绝， 他也归于无有。
JER|49|11|你撇下孤儿，我必保全他们的性命； 你的寡妇可以倚靠我。
JER|49|12|耶和华如此说：“看哪，既然原不该喝那杯的一定要喝，你能免去惩罚吗？必不能免，一定要喝！
JER|49|13|我指着自己起誓， 波斯拉 必令人惊骇、受羞辱、被诅咒，并且全然荒废。它所有的城镇都要永远成为废墟。这是耶和华说的。”
JER|49|14|我从耶和华那里听见消息， 有使者被差往列国去，说： “你们要聚集前来攻击 以东 ， 要起来争战。”
JER|49|15|看哪，我使你在列国中为最小， 在世人中被藐视。
JER|49|16|住在山穴中盘据山顶的啊， 你被自己的声势与心中的狂傲所蒙蔽； 你虽如大鹰高高搭窝， 我却要从那里拉你下来。 这是耶和华说的。
JER|49|17|以东 必令人惊骇；凡经过的人都惊骇，又因它一切的灾祸嗤笑。
JER|49|18|耶和华说：它要像 所多玛 、 蛾摩拉 和邻近的城镇一样倾覆，必无人住在那里，也无人在其中寄居。
JER|49|19|看哪，就像狮子从 约旦河 边的丛林上来，攻击坚固的居所，我要在转眼之间使 以东 人逃跑，离开这地。我拣选谁，就派谁治理这地。谁能像我呢？谁能召我出庭呢？ 有哪一个牧人能在我面前站得住呢？
JER|49|20|你们要听耶和华攻击 以东 所定的计划和他攻击 提幔 居民所定的旨意。他们羊群当中微弱的定要被拖走，他们的草场定要变为荒凉。
JER|49|21|因他们仆倒的声音，地就震动，哀号的声音传到 红海 那里。
JER|49|22|看哪，仇敌必如大鹰飞起，展开翅膀攻击 波斯拉 。到那日， 以东 的勇士心中疼痛如临产的妇人。
JER|49|23|论 大马士革 。 哈马 和 亚珥拔 蒙羞， 因为他们听见凶恶的消息就融化； 焦虑像海浪汹涌，不得平静。
JER|49|24|大马士革 发软，转身逃跑； 战兢将它捉住， 痛苦忧愁将它抓住， 如临产的妇人一样。
JER|49|25|我所喜乐受称赞的城， 怎能被撇弃 呢？
JER|49|26|它的壮丁必仆倒在街上， 当那日，战士全都静默无声。 这是万军之耶和华说的。
JER|49|27|我必用火点燃 大马士革 的城墙， 烧灭 便．哈达 的宫殿。
JER|49|28|论 巴比伦 王 尼布甲尼撒 所攻打的 基达 和 夏琐 诸国。 耶和华如此说： 迦勒底 人哪，起来上 基达 去， 毁灭东方人。
JER|49|29|人要夺去他们的帐棚和羊群， 人要带走他们的幔子、一切器皿，和骆驼，占为己有。 人向他们喊着说： 四围都有惊吓。
JER|49|30|夏琐 的居民哪，要逃奔远方， 住在深远之处； 因为 巴比伦 王 尼布甲尼撒 设计谋害你们， 起意攻击你们。 这是耶和华说的。
JER|49|31|迦勒底 人哪，起来！ 上到安逸无虑的国民那里去， 他们是无门无闩、单独居住的。 这是耶和华说的。
JER|49|32|他们的骆驼必成为掠物， 他们众多的牲畜必成为掳物。 我要将剃鬓发的人分散四方 ， 使灾殃从四围临到他们。 这是耶和华说的。
JER|49|33|夏琐 必成为野狗的住处， 永远荒废； 无人住在那里， 也无人在其中寄居。
JER|49|34|犹大 王 西底家 登基的时候，耶和华论 以拦 的话临到 耶利米 先知，说：
JER|49|35|“万军之耶和华如此说：看哪，我必折断 以拦 人的弓，那是他们战斗的主力。
JER|49|36|我要使风从天的四方刮来，临到 以拦 ，将他们分散四方。 以拦 被赶散的人没有一国不到的。
JER|49|37|我必使 以拦 人在仇敌和寻索其命的人面前惊惶；我也必使灾祸，就是我的烈怒临到他们，又必使刀剑追杀他们，直到将他们灭尽。这是耶和华说的。
JER|49|38|我要在 以拦 设立我的宝座，在那里除灭君王和官长。这是耶和华说的。
JER|49|39|“到末后，我却要使被掳的 以拦 人归回。这是耶和华说的。”
JER|50|1|以下是耶和华藉 耶利米 先知论 巴比伦 和 迦勒底 人之地所说的话。
JER|50|2|你们要在万国中传扬，宣告， 竖立大旗； 要宣告，不可隐瞒，说： “ 巴比伦 被攻取， 彼勒 蒙羞， 米罗达 惊惶。 巴比伦 的神像都蒙羞， 它的偶像都惊惶。”
JER|50|3|因有一国从北方上来攻击它，使它的地荒凉，无人居住，连人带牲畜都逃走了。
JER|50|4|在那日、在那时， 以色列 人要和 犹大 人同来，随走随哭，寻求耶和华－他们的上帝。这是耶和华说的。
JER|50|5|他们要问到 锡安 之路，又面向那里，说：“来吧，他们要 在永不被遗忘的约中与耶和华联合。”
JER|50|6|我的百姓成了失丧的羊，牧人使他们走迷了路，转入丛山之间。他们从大山走到小山，竟忘了自己安歇之处。
JER|50|7|凡遇见他们的，就把他们吞灭。敌人说：“我们不算有罪；因他们得罪了那可作真正 居所的耶和华，就是他们祖先所仰望的耶和华。”
JER|50|8|“你们要逃离 巴比伦 ，要离开 迦勒底 人之地，像走在羊群前面的公山羊。
JER|50|9|看哪，因我必激起大国联盟，带领他们从北方来攻击 巴比伦 ，他们要摆阵攻击它，它必在那里被攻取。他们的箭好像善射 勇士的箭，绝不徒然返回。
JER|50|10|迦勒底 要成为掠物，凡掳掠它的都必心满意足。这是耶和华说的。”
JER|50|11|抢夺我产业的啊， 你们因欢喜快乐， 像踹谷 嬉戏的母牛犊， 又像发嘶声的壮马。
JER|50|12|你们的母亲极其抱愧， 生你们的必然蒙羞。 看哪，她要列在诸国之末， 成为旷野、旱地、沙漠；
JER|50|13|因耶和华的愤怒， 巴比伦 必无人居住， 全然荒凉， 凡经过的都要受惊骇， 又因它所遭的灾殃嗤笑。
JER|50|14|所有拉弓的啊，要在 巴比伦 的四围摆阵， 射箭攻击它， 不用爱惜箭枝， 因为它得罪了耶和华。
JER|50|15|要在它四围呐喊： “它已经投降， 堡垒坍塌了， 城墙拆毁了！” 这是耶和华所报的仇。 你们要向它报仇； 它怎样待人，你们也要怎样待它。
JER|50|16|你们要将 巴比伦 撒种的 和收割时拿镰刀的全都剪除。 他们各人因躲避欺压的刀剑， 必归回本族，逃到本土。
JER|50|17|以色列 是打散的羊，被狮子赶散。首先是 亚述 王将他吞灭，末后是 巴比伦 王 尼布甲尼撒 折断他的骨头。
JER|50|18|所以万军之耶和华－ 以色列 的上帝如此说：“看哪，我必惩罚 巴比伦 王和他的地，像我从前惩罚 亚述 王一样。
JER|50|19|我必领 以色列 回他自己的草场，他要在 迦密 和 巴珊 吃草，又在 以法莲 山上和 基列 境内得以饱足。
JER|50|20|在那日、在那时，你寻找 以色列 的罪孽，一无所有；寻找 犹大 的罪恶，也无所得；因为我所留下的人，我必赦免。这是耶和华说的。”
JER|50|21|你要上去攻击 米拉大翁 之地， 又攻击 比割 的居民。 将他们追杀灭尽， 照我所吩咐你的一切去做。 这是耶和华说的。
JER|50|22|境内有打仗和大毁灭的响声。
JER|50|23|全地的大锤竟然砍断破坏！ 巴比伦 在列国中竟然荒凉！
JER|50|24|巴比伦 哪，我为你设下罗网， 你被缠住，竟不自觉。 你被寻着，也被捉住， 因为你对抗耶和华。
JER|50|25|耶和华已经打开军械库， 拿出他恼恨的兵器； 这是万军之主耶和华 在 迦勒底 人之地要做的事。
JER|50|26|你们要从极远的边界前来攻击它 ， 要开它的仓廪， 将它堆起如高堆， 毁灭净尽，丝毫不留。
JER|50|27|要杀它一切的牛犊， 使它们下去遭杀戮。 他们有祸了， 因为他们的日子，就是他们受罚的时刻已经来到。
JER|50|28|从 巴比伦 之地逃出来的难民，在 锡安 扬声宣告耶和华－我们的上帝要报仇，为他的圣殿报仇。
JER|50|29|你们要招集一切弓箭手来攻击 巴比伦 ，在 巴比伦 四围安营，不容一人逃脱。要照着它所做的报应它；它怎样待人，你们也要怎样待它，因为它向耶和华－ 以色列 的圣者狂傲。
JER|50|30|所以它的壮丁必仆倒在街上。当那日，它的士兵全都静默无声。这是耶和华说的。
JER|50|31|“看哪，你这狂傲的啊，我与你为敌， 因为你的日子， 我惩罚你的时刻已经来到。 这是万军之主耶和华说的。
JER|50|32|狂傲的必绊跌仆倒，无人扶起。 我必用火点燃他的城镇， 将他四围所有的尽行烧灭。”
JER|50|33|万军之耶和华如此说：“ 以色列 人和 犹大 人一同受欺压；凡掳掠他们的都紧紧抓住他们，不肯释放。
JER|50|34|他们的救赎主大有能力，万军之耶和华是他的名。他必定为他们伸冤，使全地得享平静；他却要搅扰 巴比伦 的居民。”
JER|50|35|有刀剑临到 迦勒底 人和 巴比伦 的居民， 临到它的领袖与智慧人。 这是耶和华说的。
JER|50|36|有刀剑临到矜夸的人， 他们就变为愚昧； 有刀剑临到它的勇士， 他们就惊惶。
JER|50|37|有刀剑临到它的马匹、战车， 和其中混居的各族， 他们变成与妇女一样； 有刀剑临到它的宝物， 宝物就被抢夺。
JER|50|38|有干旱 临到它的众水， 它们就必干涸； 因为这是雕刻偶像之地， 人因偶像颠狂 。
JER|50|39|所以野兽和土狼必住在那里，鸵鸟也住在其中，永远无人居住，世世代代无人定居。
JER|50|40|巴比伦 要像上帝所倾覆的 所多玛 、 蛾摩拉 和邻近的城镇一样，必无人住在那里，也无人在其中寄居。这是耶和华说的。
JER|50|41|看哪，有一民族从北方而来， 有一大国和许多君王被激起，从地极来到。
JER|50|42|他们拿弓和枪， 性情残忍，毫不留情； 他们的声音像海浪澎湃。 巴比伦 啊， 他们骑着马， 如上战场的人摆列队伍， 要攻击你。
JER|50|43|巴比伦 王听见他们的风声， 手就发软， 痛苦将他抓住， 仿佛临产的妇人疼痛一般。
JER|50|44|“看哪，就像狮子从 约旦河 边的丛林上来，攻击坚固的居所，我要在转眼之间使 迦勒底 人逃跑，离开这地。我拣选谁，就派谁治理这地。谁能像我呢？谁能召我出庭呢？有哪一个牧人能在我面前站得住呢？
JER|50|45|你们要听耶和华攻击 巴比伦 所定的计划和他攻击 迦勒底 人之地所定的旨意。他们羊群当中微弱的定要被拖走，他们的草场定要变为荒凉。
JER|50|46|因 巴比伦 被攻下的声音，地就震动，人在列国都听见呼喊的声音。”
JER|51|1|耶和华如此说： 看哪，我必刮起毁灭的风， 攻击 巴比伦 和住在 立加米 的人。
JER|51|2|我要差陌生人 来到 巴比伦 ， 他们要簸扬它，使它的地空无一物。 在它遭祸的日子， 他们要四围攻击它。
JER|51|3|不要叫拉弓的拉弓， 不要叫他佩戴盔甲 ； 不要怜惜 巴比伦 的壮丁， 要灭尽它的全军。
JER|51|4|他们必在 迦勒底 人之地被杀仆倒， 在 巴比伦 的街市上被刺透。
JER|51|5|以色列 和 犹大 境内虽然充满违背 以色列 圣者的罪， 却没有被他的上帝－万军之耶和华所遗弃。
JER|51|6|你们要奔逃，离开 巴比伦 ， 各救自己的性命！ 不要陷在它的罪孽中一同灭亡， 因为这是耶和华报仇的时刻， 他必向 巴比伦 施行报应。
JER|51|7|巴比伦 素来是耶和华手中的金杯， 使全地沉醉， 列国喝了它的酒就颠狂。
JER|51|8|巴比伦 忽然倾覆毁坏； 要为它哀号， 拿乳香来止它的疼痛， 或者可以治好。
JER|51|9|我们想医治 巴比伦 ， 它却未获痊愈。 离开它吧！让我们各人归回本国， 因为它受的审判通于上天，达到穹苍。
JER|51|10|耶和华已经彰显出我们的义。 来吧！我们要在 锡安 传扬耶和华－我们上帝的作为。
JER|51|11|你们要磨尖箭头， 抓住盾牌。 论到 巴比伦 ，耶和华定意要毁灭它，所以激起 玛代 君王的心；这是耶和华报仇，为他的圣殿报仇。
JER|51|12|你们要竖立大旗， 攻击 巴比伦 的城墙； 要坚固了望台， 派定守望的设下埋伏； 因为耶和华指着 巴比伦 居民所说的， 他不但这样定意，也已成就。
JER|51|13|住在众水之上多有财宝的啊， 你的结局已到！ 你贪婪之量已满盈 ！
JER|51|14|万军之耶和华指着自己起誓说： 我必使人遍满各处像蝗虫一样， 他们必呐喊攻击你。
JER|51|15|耶和华以能力创造大地， 以智慧建立世界， 以聪明铺张穹苍。
JER|51|16|他一出声，天上就有众水澎湃； 他使云雾从地极上腾， 造电随雨而闪， 从仓库中吹出风来。
JER|51|17|人人都如同畜牲，毫无知识； 银匠都因偶像羞愧， 他所铸的偶像本为虚假， 它们里面并无气息。
JER|51|18|它们都是虚无的， 是迷惑人的东西， 到它们受罚的时刻必被除灭。
JER|51|19|雅各 所得的福分不是这样， 因主 是那创造万有的， 以色列 是他产业的支派， 万军之耶和华是他的名。
JER|51|20|你是我争战的斧子和打仗的兵器。 我要用你打碎列邦， 毁灭列国；
JER|51|21|用你打碎马和骑马的， 打碎战车和坐在其上的；
JER|51|22|用你打碎男人和女人， 打碎老人和少年， 打碎壮丁和少女；
JER|51|23|用你打碎牧人和他的羊群， 打碎农夫和他的一对耕牛， 打碎省长和官员。
JER|51|24|我必在你们眼前报复 巴比伦 人和 迦勒底 居民在 锡安 所做的一切恶事。这是耶和华说的。
JER|51|25|行毁灭的山，看哪，我与你为敌， 你毁灭全地， 我必伸手攻击你， 将你从山岩滚下去， 使你成为烧毁了的山。 这是耶和华说的。
JER|51|26|人必不从你那里取石头为房角石， 也不取石头来作根基， 因为你必永远荒废。 这是耶和华说的。
JER|51|27|你们要在境内竖立大旗， 在列邦中吹角， 使列邦预备攻击 巴比伦 。 要招集 亚拉腊 、 米尼 、 亚实基拿 各国前来攻击它， 派将军攻击它， 使马匹上来如粗暴的蝗虫；
JER|51|28|使列邦和 玛代 君王，省长和官员， 他们所管的全地，都预备攻击它。
JER|51|29|地必震动而移转； 因耶和华向 巴比伦 旨意已确定， 要使 巴比伦 土地荒凉，无人居住。
JER|51|30|巴比伦 的勇士停止争战， 躲在堡垒之中。 他们的力气耗尽， 他们变成与妇女一样。 巴比伦 的住处焚烧， 门闩都折断了。
JER|51|31|通报的彼此相遇， 送信的彼此相遇， 报告 巴比伦 王， 城的四方都被攻下了，
JER|51|32|渡口被占据了， 芦苇被火焚烧， 战士都惊慌。
JER|51|33|万军之耶和华－ 以色列 的上帝如此说： 巴比伦 好像踹谷的禾场； 再过片时，它收割的时候就到了。
JER|51|34|巴比伦 王 尼布甲尼撒 吞灭我，压碎我， 使我成为空器皿。 他如大鱼将我吞下， 以我的美物充满他的肚腹， 又把我赶出去。
JER|51|35|锡安 的居民要说： 愿我和我骨肉之亲所受的残暴 归给 巴比伦 。 耶路撒冷 人要说： 愿我们所流的血 归给 迦勒底 的居民。
JER|51|36|所以，耶和华如此说： 看哪，我必为你伸冤，为你报仇； 我必使 巴比伦 的海枯竭， 使它的泉源干涸。
JER|51|37|巴比伦 必成为废墟， 为野狗的住处， 令人惊骇、嗤笑， 并且无人居住。
JER|51|38|他们要像少壮狮子一同咆哮， 像小狮子吼叫。
JER|51|39|他们食欲一来的时候， 我必为他们摆设酒席， 使他们沉醉，好叫他们快乐； 他们睡了长觉，永不醒起。 这是耶和华说的。
JER|51|40|我必使他们像羔羊、 像公绵羊和公山羊被牵去宰杀。
JER|51|41|示沙克 竟然被攻取！ 全地所称赞的被占据！ 巴比伦 在列国中竟然变为荒凉！
JER|51|42|海水涨起，漫过 巴比伦 ； 澎湃的海浪遮盖了它。
JER|51|43|它的城镇变废墟， 地变干旱，成为沙漠， 成为无人居住、 无人经过之地。
JER|51|44|我要惩罚 巴比伦 的 彼勒 ， 使它吐出所吞之物。 列国必不再流归到它那里， 巴比伦 的城墙也必坍塌。
JER|51|45|我的子民哪，你们要离开 巴比伦 ！ 各人逃命，躲避耶和华的烈怒。
JER|51|46|不要因境内所听见的风声 心惊胆怯或惧怕； 因为这年有风声传来， 那年也有风声传来； 境内有残暴的事， 官长攻击官长。
JER|51|47|所以，看哪，日子将到， 我必惩罚 巴比伦 雕刻的偶像。 它的全地必然抱愧， 它被杀的人必仆倒在其上。
JER|51|48|那时，天地和其中所有的， 必因 巴比伦 欢呼， 因为行毁灭的要从北方来到它那里。 这是耶和华说的。
JER|51|49|巴比伦 要因 以色列 被杀的人而仆倒， 正如全地被刺杀的人是因 巴比伦 仆倒一般。
JER|51|50|你们躲避刀剑的要快走， 不要站住！ 要在远方怀念耶和华， 心中追想 耶路撒冷 。
JER|51|51|我们听见辱骂就蒙羞，满面惭愧， 因为外邦人进入耶和华殿的圣所。
JER|51|52|所以，看哪，日子将到， 我必惩罚 巴比伦 雕刻的偶像， 在全境内到处都有刺伤的人在呻吟。 这是耶和华说的。
JER|51|53|巴比伦 虽升到天上， 虽使它坚固的高处更坚固， 我也要差毁灭者到它那里。 这是耶和华说的。
JER|51|54|有哀号的声音从 巴比伦 出来， 有大毁灭从 迦勒底 人之地而来。
JER|51|55|耶和华使 巴比伦 变为废墟， 使其中喧哗的大声灭绝。 仇敌仿佛众水， 波浪澎湃，发出响声；
JER|51|56|这是行毁灭的临到 巴比伦 。 巴比伦 的勇士被捉住， 他们的弓折断了； 因为耶和华是施行报应的上帝， 他必施行报应。
JER|51|57|我必使 巴比伦 的领袖、 智慧人、省长、官员和勇士都喝醉， 使他们永远沉睡，不再醒起。 这是名为万军之耶和华的君王说的。
JER|51|58|万军之耶和华如此说： 巴比伦 宽阔的城墙要夷为平地， 它高大的城门必被火焚烧。 万民所劳碌的必致虚空， 万族所劳碌的被火焚烧， 他们都必困乏。
JER|51|59|犹大 王 西底家 在位第四年， 玛西雅 的孙子， 尼利亚 的儿子 西莱雅 与王同去 巴比伦 ， 西莱雅 是王宫的大臣， 耶利米 先知有话吩咐他。
JER|51|60|耶利米 把一切要临到 巴比伦 的灾祸，就是论到 巴比伦 的这一切话，写在一书卷上。
JER|51|61|耶利米 对 西莱雅 说：“你到了 巴比伦 ，务要宣读这一切话，
JER|51|62|说：‘耶和华啊，你曾论到这地方说：要剪除它，不再有人与牲畜居住此地，必永远荒凉。’
JER|51|63|你读完这书卷，就要把一块石头拴在其上，投入 幼发拉底河 中，
JER|51|64|说：‘ 巴比伦 因耶和华所要降与它的灾祸，必如此沉下去，不再浮起来，百姓也必困乏。’” 耶利米 的话到此为止。
JER|52|1|西底家 登基的时候年二十一岁，在 耶路撒冷 作王十一年。他母亲名叫 哈慕她 ，是 立拿 人 耶利米 的女儿。
JER|52|2|西底家 行耶和华眼中看为恶的事，像 约雅敬 所做的一切。
JER|52|3|因此，耶和华向 耶路撒冷 和 犹大 发怒，以致把他们从自己面前赶出去。 西底家 背叛 巴比伦 王，
JER|52|4|他作王第九年十月初十， 巴比伦 王 尼布甲尼撒 率领全军前来攻击 耶路撒冷 ，对着城安营，四围筑堡垒攻城，
JER|52|5|城被围困，直到 西底家 王十一年。
JER|52|6|四月初九，城里的饥荒非常严重，当地的百姓都没有粮食。
JER|52|7|城被攻破，士兵全都在夜间从靠近王园两城墙中间的门逃跑出城； 迦勒底 人正在四围攻城，他们就往 亚拉巴 逃去。
JER|52|8|迦勒底 的军队追赶 西底家 王，在 耶利哥 的平原追上他。他的全军都离开他溃散了。
JER|52|9|迦勒底 人就拿住王，带他到 哈马 地 利比拉 的 巴比伦 王那里； 巴比伦 王就判他的罪。
JER|52|10|巴比伦 王在 西底家 眼前杀了他的儿女，又在 利比拉 杀了 犹大 全体的官长，
JER|52|11|并且挖了 西底家 的眼睛，用铜链锁着他，带到 巴比伦 去，将他囚在监里，直到他死的日子。
JER|52|12|巴比伦 王 尼布甲尼撒 十九年五月初十，在 巴比伦 王面前侍立的 尼布撒拉旦 护卫长进入 耶路撒冷 ，
JER|52|13|他焚烧了耶和华的殿、王宫和 耶路撒冷 的房屋；用火焚烧所有大户人家的房屋。
JER|52|14|跟随护卫长的 迦勒底 全军拆毁了 耶路撒冷 四围的城墙。
JER|52|15|那时 尼布撒拉旦 护卫长将百姓中最穷的和城里所剩下的百姓，并那些投降 巴比伦 王的人，以及剩下的工匠，都掳去了。
JER|52|16|但 尼布撒拉旦 护卫长留下一些当地最穷的人，叫他们修整葡萄园，耕种田地。
JER|52|17|耶和华殿的铜柱并殿内的盆座和铜海， 迦勒底 人都打碎了，把那些铜运到 巴比伦 去；
JER|52|18|他们又带走锅、铲子、钳子、盘子、勺子，和供奉用的一切铜器；
JER|52|19|杯、火盆、碗、锅、灯台、勺子、酒杯，无论金的银的，护卫长都带走了；
JER|52|20|还有 所罗门 为耶和华殿所造的两根柱子、一面铜海，并座下的十二只铜牛，这些器皿的铜多得无法可秤。
JER|52|21|至于柱子，这一根柱子高十八肘，厚四指，周围十二肘，中间是空的；
JER|52|22|柱上有铜顶，每个铜顶高五肘；铜顶的周围有网子和石榴，也都是铜的。另一根柱子与此相同，也有石榴。
JER|52|23|柱子四面有九十六个石榴，在网子周围，总共有一百个石榴。
JER|52|24|护卫长拿住 西莱雅 大祭司、 西番亚 副祭司和门口的三个守卫，
JER|52|25|又从城中拿住一个管理士兵的官 ，并在城里找到王面前的七个亲信，和召募当地百姓之将军的书记官，以及在城中找到的六十个当地百姓。
JER|52|26|尼布撒拉旦 护卫长把这些人带到 利比拉 的 巴比伦 王那里。
JER|52|27|巴比伦 王击杀他们，在 哈马 地的 利比拉 把他们处死。这样， 犹大 人就被掳去离开本地。
JER|52|28|这是 尼布甲尼撒 所掳百姓的数目：他在位第七年掳去 犹大 人三千零二十三人；
JER|52|29|尼布甲尼撒 十八年从 耶路撒冷 掳去八百三十二人；
JER|52|30|尼布甲尼撒 二十三年， 尼布撒拉旦 护卫长掳去 犹大 人七百四十五人；共有四千六百人。
JER|52|31|巴比伦 王 以未．米罗达 作王的元年，就是 犹大 王 约雅斤 被掳后三十七年十二月二十五日，他使 犹大 王 约雅斤 抬起头来，提他出监，
JER|52|32|对他说好话，使他的位高过与他一同被掳、在 巴比伦 众王的位；
JER|52|33|又给他脱了囚服，使他终身常在 巴比伦 王面前吃饭。
JER|52|34|巴比伦 王赐给他日常需用的食物，日日一份，终身都是这样，直到他死的日子。
LAM|1|1|唉！先前人口稠密的城市， 现在为何独坐！ 先前在列国中为大的， 现在竟如寡妇！ 先前在各省中为王后的， 现在竟成为服苦役的人！
LAM|1|2|她 夜间痛哭，泪流满颊， 在所有亲爱的人中，找不到一个安慰她的。 她的朋友都以诡诈待她， 成为她的仇敌。
LAM|1|3|犹大 被掳， 遭遇苦难，多服劳役。 她住在列国中，得不着安息； 追逼她的在狭窄之地追上她。
LAM|1|4|锡安 的道路因无人前来过节就哀伤， 她的城门荒凉， 祭司叹息， 少女悲伤； 她自己充满痛苦。
LAM|1|5|她的敌人作主， 她的仇敌亨通； 耶和华因她过犯多而使她受苦， 她的孩童在敌人面前去作俘虏。
LAM|1|6|锡安 的威荣全都失去。 她的领袖如找不着草场的鹿， 在追赶的人面前无力行走。
LAM|1|7|耶路撒冷 在困苦窘迫之时， 就追想古时一切的荣华。 她的百姓落在敌人手中，无人帮助； 敌人看见，就因她的毁灭嗤笑。
LAM|1|8|耶路撒冷 犯了大罪， 因此成为不洁净； 素来尊敬她的，见她裸露就都藐视她， 她自己也叹息退后。
LAM|1|9|她的污秽是在下摆上； 她未曾思想自己的结局， 她的败落令人惊诧， 无人安慰她。 “耶和华啊，求你看顾我的苦难， 因为仇敌强大。”
LAM|1|10|敌人伸手夺取她的一切贵重物品； 她眼见列国侵入她的圣所， 你曾吩咐他们不可进入你的集会。
LAM|1|11|她的百姓都叹息，寻求食物； 他们用贵重物品换取粮食，要救性命。 “耶和华啊，求你观看， 留意我多么卑微。”
LAM|1|12|所有过路的人哪，愿这事不要发生在你们身上 。 你们要留意观看， 有像这样临到我的痛苦没有？ 耶和华在他发烈怒的日子使我受苦。
LAM|1|13|他从高处降火进入我的骨头， 克制了我； 他张开网，绊我的脚， 使我退后， 又令我终日凄凉发昏。
LAM|1|14|他用手绑我罪过的轭， 卷绕着加在我颈项上； 他使我力量衰败。 主将我交在我不能抵挡的人手中。
LAM|1|15|主弃绝我们当中所有的勇士， 聚集会众攻击我， 要压碎我的年轻人。 主踹下少女 犹大 ， 在醡酒池中。
LAM|1|16|我因这些事哭泣， 眼泪汪汪； 因为那安慰我、使我重新得力的， 离我甚远。 我的儿女孤苦， 因为仇敌得胜了。
LAM|1|17|锡安 伸出双手，却无人安慰。 论到 雅各 ，耶和华已经出令， 使四围的人作他的仇敌； 耶路撒冷 在他们中间成为不洁净。
LAM|1|18|耶和华是公义的！ 我违背了他的命令。 万民哪，请听， 来看我的痛苦； 我的少女和壮丁都被掳去。
LAM|1|19|我招呼我所亲爱的， 他们却欺骗了我。 我的祭司和长老寻找食物，要救性命的时候， 就在城中断了气。
LAM|1|20|耶和华啊，求你观看， 因为我在急难中； 我的心肠烦乱， 我心在我里面翻转， 因我大大背逆。 在外，刀剑使人丧亡； 在家，犹如死亡。
LAM|1|21|有人听见我叹息 ， 却无人安慰我！ 我所有的仇敌听见我的患难就喜乐， 因这是你所做的。 你使你所宣告的日子来临， 愿他们像我一样。
LAM|1|22|愿他们的恶行都呈现在你面前； 你怎样因我一切的罪过待我， 求你也照样待他们； 因我叹息甚多，心中发昏。
LAM|2|1|唉！主竟发怒，使黑云遮蔽 锡安 ！ 他将 以色列 的华美从天扔在地上， 在他发怒的日子并不顾念自己的脚凳。
LAM|2|2|主吞灭 雅各 一切的住处，并不顾惜。 他发怒倾覆 犹大 的堡垒， 将它们夷为平地， 凌辱这国与她的领袖。
LAM|2|3|他发烈怒，砍断 以色列 一切的角， 在仇敌面前收回右手。 他将 雅各 烧毁，如火焰四围吞灭。
LAM|2|4|他张弓好像仇敌， 他站立举起右手， 如同敌人杀戮我们眼目所喜爱的。 他在 锡安 的帐棚 倾倒愤怒，如火一般。
LAM|2|5|主如仇敌吞灭 以色列 ， 吞灭它一切的宫殿， 毁坏境内的堡垒； 在 犹大 加添悲伤和哭号。
LAM|2|6|他摧毁自己的帐幕如摧毁园子， 毁坏自己的会幕。 耶和华使节庆和安息日在 锡安 尽被遗忘， 又在极其愤怒中厌弃君王与祭司。
LAM|2|7|耶和华撇弃自己的祭坛， 憎恶自己的圣所， 把宫殿的墙交给仇敌。 他们在耶和华的殿中喧嚷， 如在节庆之日一样。
LAM|2|8|耶和华定意拆毁 锡安 的城墙； 他拉了准绳， 不将手收回，定要毁灭。 他使城郭和城墙都悲哀， 一同衰败。
LAM|2|9|锡安 的门陷入地里， 主毁坏，折断她的门闩。 她的君王和官长都置身列国中，没有律法； 她的先知也不再从耶和华领受异象。
LAM|2|10|锡安 的长老坐在地上，默默无声； 他们扬起尘土落在头上，腰束麻布； 耶路撒冷 的少女垂头至地。
LAM|2|11|我的眼睛流泪，以致失明； 我的心肠烦乱，肝胆落地， 都因我的百姓 遭毁灭， 又因孩童和吃奶的在城内的广场上昏厥。
LAM|2|12|他们如受伤的人在城内广场上昏厥， 在母亲的怀里将要丧命时， 就对母亲说：“饼和酒在哪里呢？”
LAM|2|13|耶路撒冷 啊，我可用什么向你证明 呢？ 我可用什么与你相比呢？ 少女 锡安 哪，我拿什么和你比较，好安慰你呢？ 因你的裂伤大如海； 谁能医治你呢？
LAM|2|14|你的先知为你看见虚假和粉饰的异象， 并未揭露你的罪孽， 使你被掳的归回； 却传给你虚假与误导人的默示。
LAM|2|15|凡过路的都向你拍掌。 他们向 耶路撒冷 嗤笑，摇头： “这就是人称为全美的、 称为全地所喜悦的城吗？”
LAM|2|16|你所有的仇敌 张口来攻击你； 他们嗤笑，切齿，说： “我们把她吞灭了， 这是我们所盼望的日子！ 我们终于等到了，亲眼看见了！”
LAM|2|17|耶和华成就了他所定的， 应验了他古时所命定的。 他倾覆，并不顾惜， 他使仇敌向你夸耀， 使你敌人的角高举。
LAM|2|18|他们的心哀求主。 锡安 的城墙啊， 愿你日夜泪流如河，不让自己休息， 你眼中的瞳人也不歇息。
LAM|2|19|夜间每逢时辰开始，要起来呼喊， 在主面前倾心吐意如水。 你的孩童在街头上挨饿昏厥， 你要为他们的性命向主举手。
LAM|2|20|耶和华啊，求你观看， 留意你向谁这样行。 妇人岂可吃自己所生、所抚育的婴孩吗？ 祭司和先知岂可在主的圣所中被杀吗？
LAM|2|21|年轻人和老年人躺卧在街上， 我的少女和壮丁都倒在刀下。 你在发怒的日子杀了他们， 你杀戮，并不顾惜。
LAM|2|22|你从四围招聚使我惊吓的人， 像在节庆的日子一样。 耶和华发怒的日子， 无人逃脱，无人生还。 我所抚育养大的， 仇敌都杀尽了。
LAM|3|1|因耶和华愤怒的杖， 我是遭遇困苦的人。
LAM|3|2|他驱赶我走入黑暗， 没有光明。
LAM|3|3|他反手攻击我， 终日不停。
LAM|3|4|他使我皮肉枯干， 折断我的骨头。
LAM|3|5|他筑垒攻击我， 以苦楚和艰难围困我；
LAM|3|6|使我住在幽暗之处， 像死了许久的人一样。
LAM|3|7|他围住我，使我无法脱身； 他使我的铜链沉重。
LAM|3|8|尽管我哀号求救， 他仍拦阻我的祷告。
LAM|3|9|他用凿过的石头挡住我的道路， 使我的路径弯曲。
LAM|3|10|他向我如埋伏的熊， 如在隐密处的狮子。
LAM|3|11|他使我转离正路， 把我撕碎 ，使我凄凉。
LAM|3|12|他拉弓，命我站立， 作为箭靶；
LAM|3|13|把箭袋中的箭 射入我的肺腑。
LAM|3|14|我成了全体百姓的笑柄， 成了他们终日的歌曲。
LAM|3|15|他使我受尽苦楚， 饱食茵蔯；
LAM|3|16|用沙石磨断我的牙， 以灰尘覆盖我。
LAM|3|17|你使我远离平安， 我忘了何为福乐。
LAM|3|18|于是我说：“我的力量衰败， 在耶和华那里我毫无指望！”
LAM|3|19|求你记得我的困苦和流离， 它如茵蔯和苦胆一般；
LAM|3|20|我心想念这些， 就在我里面忧闷 。
LAM|3|21|但我的心回转过来， 因此就有指望；
LAM|3|22|因耶和华的慈爱，我们不致灭绝 ， 因他的怜悯永不断绝，
LAM|3|23|每早晨，这些都是新的； 你的信实极其广大！
LAM|3|24|我心里说：“耶和华是我的福分， 因此，我要仰望他。”
LAM|3|25|凡等候耶和华，心里寻求他的， 耶和华必施恩给他。
LAM|3|26|人仰望耶和华， 安静等候他的救恩， 这是好的。
LAM|3|27|人在年轻时负轭， 这是好的。
LAM|3|28|他当安静独坐， 因为这是耶和华加在他身上的。
LAM|3|29|让他脸伏于地 吧！ 或者还会有指望。
LAM|3|30|让人打他耳光， 使他饱受凌辱吧！
LAM|3|31|主必不永远撇弃，
LAM|3|32|他虽使人忧愁， 还要照他丰盛的慈爱施怜悯；
LAM|3|33|他并不存心要人受苦， 令世人忧愁。
LAM|3|34|把世上所有的囚犯 踹在脚下，
LAM|3|35|在至高者面前 扭曲人的公正，
LAM|3|36|在人的诉讼上 颠倒是非， 这都是主看不中的。
LAM|3|37|若非主发命令， 谁能说了就成呢？
LAM|3|38|是祸，是福， 不都出于至高者的口吗？
LAM|3|39|人都有自己的罪， 活人有什么好发怨言的呢？
LAM|3|40|让我们省察，检讨自己的行为， 归向耶和华吧！
LAM|3|41|让我们献上我们的心， 向天上的上帝举手！
LAM|3|42|我们犯罪悖逆， 你并未赦免。
LAM|3|43|你浑身是怒气，追赶我们； 你施行杀戮，并不顾惜。
LAM|3|44|你以密云围着自己， 祷告不能穿透。
LAM|3|45|你使我们在万民中 成为污物和垃圾。
LAM|3|46|我们所有的仇敌 张口来攻击我们；
LAM|3|47|惊吓和陷阱临到我们， 残害和毁灭也临到我们。
LAM|3|48|因我百姓 遭毁灭， 我的眼睛泪流成河。
LAM|3|49|我的眼睛流泪不停， 流泪不止，
LAM|3|50|直等到耶和华垂顾， 从天上观看。
LAM|3|51|为我城中的百姓 ， 我眼所见的使我心痛。
LAM|3|52|无故与我为敌的追逼我， 像追捕雀鸟一样。
LAM|3|53|他们要在坑中了结我的性命， 丢石头在我身上。
LAM|3|54|众水淹没我的头， 我说：“我没命了！”
LAM|3|55|耶和华啊， 在极深的地府里，我求告你的名。
LAM|3|56|我的声音你听见了， 求你不要掩耳不听 我的呼声，我的求救。
LAM|3|57|我求告你的时候， 你临近我，说：“不要惧怕！”
LAM|3|58|主啊，你为我伸冤， 你救赎了我的命。
LAM|3|59|耶和华啊，你已看见我的委屈， 求你为我主持正义。
LAM|3|60|他们要报复，谋害我， 你都看见了。
LAM|3|61|耶和华啊，你听见他们的辱骂， 他们害我的一切计谋，
LAM|3|62|那些起来攻击我的人嘴唇所说的话 和他们终日攻击我的计谋。
LAM|3|63|求你留意！ 他们无论坐下或起来， 我都是他们的笑柄。
LAM|3|64|耶和华啊，求你照他们手所做的 向他们施行报应。
LAM|3|65|求你使他们心里刚硬， 使你的诅咒临到他们。
LAM|3|66|求你发怒追赶他们， 从耶和华的地上 除灭他们。
LAM|4|1|唉！黄金竟然无光！ 纯金竟然变色！ 圣所的石头散落在街上。
LAM|4|2|锡安 宝贝的孩子虽然好比精金， 现在竟当作陶匠手所做的瓦瓶！
LAM|4|3|野狗尚且哺乳其子， 我百姓 的妇人反倒残忍， 如旷野的鸵鸟一般；
LAM|4|4|吃奶孩子的舌头因干渴贴住上膛， 孩童求饼，却无人擘给他们。
LAM|4|5|素来吃美好食物的， 如今遭遗弃在街上； 素来穿着朱红衣裳长大的， 如今却拥抱粪堆。
LAM|4|6|我百姓的罪孽比 所多玛 的罪还大； 所多玛 虽无人伸手攻击， 转眼之间就被倾覆。
LAM|4|7|锡安 的拿细耳人 比雪纯净， 比奶更白； 他们的身体比宝石更红， 身躯之美如蓝宝石一般。
LAM|4|8|但如今他们的面貌比煤炭更黑， 在街上无人认识； 他们的皮肤紧贴骨头， 枯干形同槁木。
LAM|4|9|被刀剑刺杀的 胜过因饥饿而死 的； 饥饿者由于缺乏田里的出产 就消瘦而亡 。
LAM|4|10|当我百姓遭毁灭的时候， 慈心的妇人亲手烹煮自己的儿女为食物。
LAM|4|11|耶和华发尽他的愤怒， 倾倒他的烈怒， 用火焚烧 锡安 ， 烧毁 锡安 的根基。
LAM|4|12|地上的君王和世上的居民都不信 敌人和仇敌竟能进入 耶路撒冷 的城门。
LAM|4|13|这都因她先知的罪恶和祭司的罪孽， 他们在城中流了义人的血。
LAM|4|14|他们如盲人在街上徘徊， 又被血玷污， 以致人不敢摸他们的衣服。
LAM|4|15|人向他们喊着： “你这不洁净的，走开！ 走开！走开！不要摸我！” 他们逃走流浪的时候， 列国中有人说： “他们不可再寄居此地。”
LAM|4|16|耶和华亲自赶散他们， 不再眷顾他们； 不看重祭司，也不厚待长老。
LAM|4|17|我们的眼目徒然仰望帮助，以致失明， 我们从了望台所守望的，竟是一个不能救人的国！
LAM|4|18|仇敌追逐我们的脚踪， 使我们不敢在自己的街上行走。 我们的结局临近， 日子已满， 我们的结局已经来到。
LAM|4|19|追赶我们的比空中的鹰更快； 他们在山上追逼我们， 在旷野埋伏，等候我们。
LAM|4|20|耶和华的受膏者是我们鼻中的气， 被抓到他们的坑里， 论到他，我们曾说： “我们必在他荫下， 在列国中存活。”
LAM|4|21|住 乌斯 地的 以东 啊，尽管欢喜快乐， 苦杯必传到你那里； 你要喝醉，裸露自己。
LAM|4|22|锡安 哪，你罪孽的惩罚已经结束， 耶和华必不再使你被掳去。 以东 啊，耶和华必惩罚你的罪孽， 揭露你的罪恶。
LAM|5|1|耶和华啊，求你顾念我们所遭遇的， 留意看我们所受的凌辱。
LAM|5|2|我们的产业归陌生人， 我们的房屋归外邦人。
LAM|5|3|我们是无父的孤儿， 我们的母亲如同寡妇。
LAM|5|4|我们出银钱才得水喝， 我们的柴也是用钱买来的。
LAM|5|5|我们被追赶，迫及颈项， 疲乏却不得歇息。
LAM|5|6|我们束手投降 埃及 和 亚述 ， 为要得粮吃饱。
LAM|5|7|我们的祖先犯罪，而今他们不在了， 我们却担当他们的罪孽。
LAM|5|8|奴仆辖制我们， 无人救我们脱离他们的手。
LAM|5|9|因旷野有刀剑， 我们冒生命的危险才能得粮食。
LAM|5|10|因饥荒的干热， 我们的皮肤热如火炉。
LAM|5|11|他们在 锡安 玷污妇人， 在 犹大 城镇污辱少女。
LAM|5|12|他们吊起领袖的手， 使长老脸上无光。
LAM|5|13|年轻人扛磨石， 孩童背木柴而跌倒。
LAM|5|14|城门口不再有老年人， 年轻人也不再奏乐。
LAM|5|15|我们心中的快乐止息， 跳舞转为悲哀。
LAM|5|16|冠冕从我们的头上掉落； 我们有祸了，因为犯了罪。
LAM|5|17|因这些事我们心里发昏， 眼睛昏花。
LAM|5|18|锡安山 荒凉， 狐狸行在其上。
LAM|5|19|耶和华啊，你治理直到永远， 你的宝座万代长存。
LAM|5|20|你为何全然忘记我们？ 为何长久离弃我们？
LAM|5|21|耶和华啊，求你使我们回转归向你， 我们就得以回转。 求你更新我们的年日，像古时一样，
LAM|5|22|难道你全然弃绝了我们， 向我们大发烈怒？
EZEK|1|1|在三十年四月初五，我在 迦巴鲁河 边被掳的人当中，那时天开了，我看见上帝的异象。
EZEK|1|2|正是 约雅斤 王被掳的第五年四月初五，
EZEK|1|3|在 迦勒底 人之地的 迦巴鲁河 边，耶和华的话特地临到 布西 的儿子 以西结 祭司，耶和华的手按在他身上。
EZEK|1|4|我观看，看哪，狂风从北方刮来，有一朵大云闪烁着火，周围有光辉，其中的火好像闪耀的金属；
EZEK|1|5|又从其中显出四个活物的形像。他们的形状是这样：有人的形像，
EZEK|1|6|各有四张脸，四个翅膀。
EZEK|1|7|他们的腿是直的，脚掌好像牛犊的蹄，灿烂如磨亮的铜。
EZEK|1|8|在四面的翅膀以下有人的手。这四个活物的脸和翅膀是这样：
EZEK|1|9|翅膀彼此相接，行走时并不转弯，各自往前直行。
EZEK|1|10|至于脸的形像：四个活物各有人的脸，右面有狮子的脸，左面有牛的脸，也有鹰的脸；
EZEK|1|11|这就是他们的脸 。他们的翅膀向上张开，各有两个翅膀彼此相接，用另外两个翅膀遮体。
EZEK|1|12|他们各自往前直行。灵往哪里去，他们就往哪里去，行走时并不转弯。
EZEK|1|13|至于四活物的形像，就如烧着火炭的形状，又如火把的形状。有火在四活物中间来回移动，这火有光辉，从火中发出闪电。
EZEK|1|14|这些活物往来奔走，好像电光一闪。
EZEK|1|15|我观看活物，看哪，有四张脸的活物旁边各有一个轮子在地上。
EZEK|1|16|轮子的形状结构 好像耀眼的水苍玉。四轮都是一个样式，形状 结构好像轮中套轮。
EZEK|1|17|轮子行走的时候，向四方直行，行走时并不转弯。
EZEK|1|18|至于轮圈，高而可畏；四个轮圈周围布满眼睛。
EZEK|1|19|活物行走，轮子也在旁边行走；活物离地上升，轮子也上升。
EZEK|1|20|灵往哪里去，活物就往哪里去；轮子在活物旁边上升，因为活物的灵在轮中。
EZEK|1|21|活物行走，轮子也行走；活物站住，轮子也站住；活物离地上升，轮子也在旁边上升，因为活物的灵在轮中。
EZEK|1|22|活物的头上面有穹苍的形像，像耀眼惊人的水晶，铺张在活物的头顶上。
EZEK|1|23|穹苍之下，活物的翅膀伸直，彼此相对，每个活物用两个翅膀遮住自己；每个活物用两个翅膀遮住自己 ，就是自己的身体。
EZEK|1|24|活物行走的时候，我听见翅膀的响声，像大水的声音，像全能者的声音，又像军队闹哄的声音。活物站住的时候，翅膀垂下。
EZEK|1|25|在他们头上的穹苍之上有声音。他们站住的时候，翅膀垂下。
EZEK|1|26|在他们头上的穹苍之上有宝座的形像，仿佛蓝宝石的样子；宝座的形像上方有仿佛人的样子的形像。
EZEK|1|27|我见他的腰以上有仿佛闪耀的金属，周围有仿佛火的形状，又见他的腰以下有仿佛火的形状，周围也有光辉。
EZEK|1|28|下雨的日子，云中彩虹的形状怎样，周围光辉的形状也是怎样。 这就是耶和华荣耀形像的样式，我一看见就脸伏于地。我又听见一位说话者的声音。
EZEK|2|1|他对我说：“人子啊，你站起来，我要和你说话。”
EZEK|2|2|他对我说话的时候，灵进入我里面，使我站起来，我就听见他对我说话。
EZEK|2|3|他对我说：“人子啊，我差你往悖逆我的国家， 以色列 人那里去，他们是悖逆我的。他们和他们的祖先违背我，直到今日。
EZEK|2|4|这些人厚着脸皮，心里刚硬。我差你到他们那里去，你要对他们说：‘主耶和华如此说。’
EZEK|2|5|他们是悖逆之家，他们或听，或不听，必知道在他们中间有了先知。
EZEK|2|6|你，人子啊，虽有荆棘和蒺藜在你那里，你又住在蝎子中间，总不要怕他们，也不要怕他们的话；他们虽是悖逆之家，但你不要怕他们的话，也不要因他们的脸色惊惶。
EZEK|2|7|他们或听，或不听，你只管将我的话告诉他们；他们是极其悖逆的。
EZEK|2|8|“但是你，人子啊，要听我对你说的话，不要像那悖逆之家一样悖逆，要开口吃我所赐给你的。”
EZEK|2|9|我观看，看哪，有一只手向我伸来；看哪，手中有一书卷。
EZEK|2|10|他在我面前展开书卷，它内外都写着字，上面所写的有哀号、叹息、悲痛的话。
EZEK|3|1|他对我说：“人子啊，要吃你所得到的，吃下这书卷；然后要去，对 以色列 家宣讲。”
EZEK|3|2|于是我张开了口，他就使我吃这书卷。
EZEK|3|3|他对我说：“人子啊，要吃我所赐给你的这书卷，塞满你的肚腹。”我就吃了，口中觉得其甜如蜜。
EZEK|3|4|他对我说：“人子啊，你要到 以色列 家那里去，对他们传讲我的话。
EZEK|3|5|你奉差遣不是往那说话艰涩、言语难懂的民那里，而是往 以色列 家去；
EZEK|3|6|你不是往那说话艰涩、言语难懂的许多民族那里去，他们的话你不懂。然而，我若差你往他们那里去，他们会听从你。
EZEK|3|7|以色列 家却不肯听从你，因为他们不肯听从我；原来 以色列 全家是额头坚硬、心里刚愎的人。
EZEK|3|8|看哪，我使你的脸坚硬，对抗他们的脸；使你的额头坚硬，对抗他们的额头。
EZEK|3|9|我使你的额头像金刚石，比火石更坚硬。他们虽是悖逆之家，但你不要怕他们，也不要因他们的脸色而惊惶。”
EZEK|3|10|他又对我说：“人子啊，我对你说的一切话，你心里要领会，耳朵要听。
EZEK|3|11|要到被掳的人，到你本国百姓那里去，他们或听，或不听，你要对他们宣讲，告诉他们这是主耶和华说的。”
EZEK|3|12|那时，灵将我举起，我就听见在我身后有极大震动的声音：“耶和华的荣耀，从他所在之处，是应当称颂的！”
EZEK|3|13|有活物的翅膀相碰的声音，也有活物旁边轮子的声音，是极大震动的声音。
EZEK|3|14|于是灵将我举起，带着我走。我就去了，十分苦恼，我的灵火热；耶和华的手重重地按在我身上。
EZEK|3|15|我就来到 提勒．亚毕 那些住在 迦巴鲁河 边被掳的人那里，到他们住的地方 ，在他们中间惊愕地坐了七日。
EZEK|3|16|过了七日，耶和华的话临到我，说：
EZEK|3|17|“人子啊，我立你作 以色列 家的守望者，所以你要听我口中的话，替我警戒他们。
EZEK|3|18|我何时指着恶人说：‘他必要死’；你若不警戒他，也不劝告他，使他离开恶行，拯救他的性命，这恶人必死在罪孽之中；我却要从你手里讨他的血债。
EZEK|3|19|倘若你警戒恶人，他仍不转离罪恶，也不离开恶行，他必死在罪孽之中，你却救了自己的命。
EZEK|3|20|但是义人若转离他的义而作恶，我要把绊脚石放在他面前，他必死亡；因你没有警戒他，他必死在罪中，他素来所行的义不被记念；我却要从你手里讨他的血债。
EZEK|3|21|倘若你警戒义人，使他不犯罪，他就不犯罪；他因领受警戒就必存活，你也救了自己的命。”
EZEK|3|22|在那里耶和华的手按在我身上。他对我说：“起来，到平原去，我要在那里和你说话。”
EZEK|3|23|于是我起来，到平原去，看哪，耶和华的荣耀停在那里，正如我在 迦巴鲁河 边所见到的一样，我就脸伏于地。
EZEK|3|24|灵进入我里面，使我站起来。耶和华对我说：“你进屋里去，把门关上。
EZEK|3|25|你，人子，看哪，人要用绳索捆绑你，使你不能出去到他们中间。
EZEK|3|26|我必使你的舌头贴住上膛，以致你哑口，不能作责备他们的人；他们原是悖逆之家。
EZEK|3|27|但我对你说话的时候，必使你开口，你就要对他们说：‘主耶和华如此说。’听的，让他听；不听的，任他不听，因为他们是悖逆之家。”
EZEK|4|1|“你，人子啊，拿一块砖，摆在你面前，将一座城 耶路撒冷 画在上面。
EZEK|4|2|你要围攻这城，筑堡垒，建土堆，安营攻击，周围设撞城槌攻城，
EZEK|4|3|又要拿一个铁盘放在你和城的中间，作为铁墙。你要把你的脸对着这城，使城被困。你要围攻这城，这要成为 以色列 家的预兆。
EZEK|4|4|“你要向左侧卧，承担 以色列 家的罪孽；按你向左侧卧的日数，担当他们的罪孽。
EZEK|4|5|我已将他们作恶的年数定了日期，就是三百九十天，你要如此担当 以色列 家的罪孽。
EZEK|4|6|这些日子结束之后，你还要向右侧卧，担当 犹大 家的罪孽。我为你定了四十天，一天顶一年。
EZEK|4|7|你要把你的脸对着被困的 耶路撒冷 ，露出膀臂，说预言攻击这城。
EZEK|4|8|看哪，我用绳索捆绑你，使你不能从这边翻到那边，直等到你围困的日子结束。
EZEK|4|9|“你要取小麦、大麦、豆子、红豆、小米、粗麦，装在一个器皿里，为自己做饼；在你侧卧的三百九十天吃这饼。
EZEK|4|10|你所吃食物的量是每天二十舍客勒，要按时吃。
EZEK|4|11|你喝水的量是每天六分之一欣，要按时喝。
EZEK|4|12|你要吃这饼像大麦饼一样，在众人眼前用人的粪烤它。”
EZEK|4|13|耶和华说：“ 以色列 人在我赶他们到的列国中，也必这样吃不洁净的食物。”
EZEK|4|14|我说：“唉！主耶和华，看哪，我从来未曾被玷污，从幼年到如今没有吃过自然死的，或被野兽撕裂的，那不洁净的肉也未曾入我的口。”
EZEK|4|15|于是他对我说：“看，我给你牛粪代替人粪，你要在上面烤你的饼。”
EZEK|4|16|他又对我说：“人子，看哪，我必断绝 耶路撒冷 粮食的供应 。他们要带着忧虑限量吃饼；带着惊惶限量喝水。
EZEK|4|17|他们因缺粮缺水，彼此惊惶，在自己的罪孽中消灭。”
EZEK|5|1|“你，人子啊，拿一把快刀当作剃刀，用这刀剃你的头发和胡须，然后用天平将须发分成几份。
EZEK|5|2|围困的日子满了，你要把三分之一放在城中用火焚烧；三分之一放在城的四围用刀砍碎；三分之一任风吹散，我要拔刀追赶它们。
EZEK|5|3|你要从其中取几根须发，用衣服的边包起来，
EZEK|5|4|再从其中取一些扔在火里，在火中焚烧；必有火从其中出来烧尽 以色列 全家。
EZEK|5|5|主耶和华如此说：这就是 耶路撒冷 。我曾将它安置在列国中，列邦都在它的四围。
EZEK|5|6|耶路撒冷 行恶，违背我的典章，过于列国；干犯我的律例，过于四围的列邦。它弃绝我的典章，也没有遵行我的律例。
EZEK|5|7|所以主耶和华如此说：因为你们混乱，过于四围的列国，不遵行我的律例，不顺从我的典章，甚至也不顺从四围列国的规条 ，
EZEK|5|8|所以主耶和华如此说：看哪，我，我必与你为敌，必在列国眼前，在你中间施行审判；
EZEK|5|9|并且因你一切可憎的事，我要在你中间行未曾行过，将来也不会行的事。
EZEK|5|10|在你中间，父亲要吃儿子，儿子要吃父亲。我必向你施行审判，将你剩下的人分散四方 。
EZEK|5|11|主耶和华说：我指着我的永生起誓，因你用一切可憎之物、可厌的事玷污我的圣所，所以，我要把你剃光 ，我的眼必不顾惜你，也不可怜你。
EZEK|5|12|你的百姓三分之一必遭瘟疫而死，因饥荒在你们中间而消灭；三分之一必在你四围倒在刀下；我必将三分之一分散四方，要拔刀追赶他们。
EZEK|5|13|“我要这样发尽我的怒气；我向他们发的愤怒停止以后，自己就得到平息。当我向他们发尽我的愤怒时，他们就知道我─耶和华所说的是出于妒忌。
EZEK|5|14|在四围的列国中，我要使你成为荒凉，在所有过路人的眼前看为羞辱。
EZEK|5|15|这样，我必以怒气、愤怒和烈怒的责备，向你施行审判。那时，它 就在四围的列国中成为羞辱、讥刺、警戒、惊骇；这是我─耶和华说的。
EZEK|5|16|我向灭亡的人射出饥荒的恶箭，将它们射出，毁灭你们；那时，我要加重你们的饥荒，断绝你们粮食的供应。
EZEK|5|17|我要令饥荒和恶兽临到你，使你丧失儿女。瘟疫和流血的事必在你那里盛行，我也要使刀剑临到你。这是我─耶和华说的。”
EZEK|6|1|耶和华的话临到我，说：
EZEK|6|2|“人子啊，你要面向 以色列 的众山说预言。
EZEK|6|3|你要说： 以色列 的众山哪，要听主耶和华的话。主耶和华对大山、小冈、水沟、山谷如此说：看哪，我要使刀剑临到你们，也必毁坏你们的丘坛。
EZEK|6|4|你们的祭坛要荒废，香坛必打碎。我要使你们当中被杀的人仆倒在你们的偶像面前，
EZEK|6|5|将 以色列 人的尸首放在他们的偶像面前，把你们的骸骨抛散在祭坛的四周围。
EZEK|6|6|无论你们住在何处，城镇要变为废墟，丘坛也必毁坏，以至于你们的祭坛荒废，被定罪 ，偶像打碎消除，香坛砍倒；你们所做的被涂去。
EZEK|6|7|被杀的人必仆倒在你们中间，你们就知道我是耶和华。
EZEK|6|8|“我必留下一些人，你们中有人得以在列国中脱离刀剑，分散在列邦。
EZEK|6|9|那些逃脱的人，必在被掳所到的各国中记得我，我心里何等伤痛，因他们起淫心，离弃我，淫荡的眼追随偶像。他们因所做一切可憎的恶事，必厌恶自己。
EZEK|6|10|他们必知道我是耶和华；我说过要使这灾祸临到他们身上，并非空话。
EZEK|6|11|“主耶和华如此说：你当击掌顿足，说：哀哉！ 以色列 家做了这一切可憎的恶事，必仆倒在刀剑、饥荒、瘟疫之下。
EZEK|6|12|在远方的，必遭瘟疫而死；在近处的，必倒在刀剑之下；那存留被围困的，必因饥荒而死；我要在他们身上发尽我的愤怒。
EZEK|6|13|被杀的要仆倒在祭坛四围的偶像中，在各高冈、各山顶、各青翠的树下，和各茂密的橡树下，就是他们献馨香的祭给一切偶像的地方。那时，他们就知道我是耶和华。
EZEK|6|14|我必伸手攻击他们，使他们的地荒废，从 第伯拉他 的旷野起 ，一切的住处都荒凉。他们就知道我是耶和华。”
EZEK|7|1|耶和华的话又临到我，说：
EZEK|7|2|“你，人子啊，主耶和华对 以色列 地如此说：结局，结局临到了地的四境！
EZEK|7|3|现在你的结局已经来临；我要使我的怒气临到你，也要按你的行为审判你，照你所做一切可憎的事惩罚你。
EZEK|7|4|我的眼必不顾惜你，也不可怜你，却要按你所做的报应你，照你们中间可憎的事惩罚你；你就知道我是耶和华。
EZEK|7|5|“主耶和华如此说：灾难，惟一的灾难 ，看哪，临近了！
EZEK|7|6|结局到了，结局到了，它要醒起来攻击你。看哪，它已来到！
EZEK|7|7|境内的居民哪，厄运临到你；时候到了，日子近了，有闹哄，但不是山上欢呼的声音。
EZEK|7|8|我快要将我的愤怒倾倒在你身上，向你发尽我的怒气，按你的行为审判你，照你所做一切可憎的事惩罚你。
EZEK|7|9|我的眼必不顾惜你，也不可怜你，必按你所做的报应你，照你中间可憎的事惩罚你；你就知道击打你的是我─耶和华。
EZEK|7|10|“看哪，那日子！看哪，已来到！厄运已经发生！杖已开花，骄傲已发芽。
EZEK|7|11|残暴兴起，成了罚恶的杖。他们将一无所有，他们的富足 、他们的财宝 都不复存在；他们中间也不再有尊荣。
EZEK|7|12|时候到了，日子近了，买主不可欢喜，卖主也不用愁烦，因为烈怒已经临到他们众人身上。
EZEK|7|13|卖主即使存活，也不能讨回所卖的，因为这异象关乎他们众人；谁都不能讨回，也没有人能在罪孽中使自己的生命刚强。”
EZEK|7|14|“他们吹了角，预备齐全，却无一人出战，因为我的烈怒临到他们众人身上。
EZEK|7|15|外有刀剑，内有瘟疫、饥荒。在田野的，必因刀剑而死；在城中的，必遭饥荒、瘟疫吞灭。
EZEK|7|16|其中幸存的要逃脱，各人因自己的罪孽在山上发出悲声，如谷中的鸽子哀鸣；
EZEK|7|17|双手发软，膝盖软弱如水，
EZEK|7|18|腰束麻布，战栗笼罩他们；各人脸上羞愧，头上光秃。
EZEK|7|19|他们要把银子抛弃在街上，看金子如污秽之物。正当耶和华发怒的日子，金银不能拯救他们，不能满足食欲，也不能使肚腹饱满，反倒成了自己罪孽的绊脚石。
EZEK|7|20|他们用所夸耀华美的妆饰制造可憎可厌的偶像，所以我使他们看它如污秽之物。
EZEK|7|21|我必将它交给外邦人为掠物，交给地上的恶人为掳物；他们要亵渎它。
EZEK|7|22|他们亵渎我宝贵之所 ，强盗也进去亵渎它。我必转脸不顾 以色列 人 。
EZEK|7|23|“要制造锁链；因为遍地都有流血的罪，满城都是残暴的事。
EZEK|7|24|所以，我要使列国中最凶恶的人前来占据他们的房屋；我要止息残暴人的骄傲，他们的圣所也要被亵渎。
EZEK|7|25|毁灭来到；他们求平安，却没有平安。
EZEK|7|26|灾害加上灾害，风声接连风声；他们要向先知寻求异象，但祭司的教诲、长老的谋略都必断绝。
EZEK|7|27|君王要悲哀，官长要披绝望为衣，这地百姓的手都发颤。我必照他们所做的待他们，按他们所应得的审判他们，他们就知道我是耶和华。”
EZEK|8|1|第六年六月初五，我坐在家中； 犹大 的众长老坐在我面前。在那里主耶和华的手降在我身上。
EZEK|8|2|我观看，看哪，有形像仿佛火 的形状，从他腰部以下形状是火，从他腰部以上有光辉的形状，好像闪耀的金属。
EZEK|8|3|他伸出一只手的样式，抓住我的一绺头发，灵就将我举到天地中间；在上帝的异象中，他带我到 耶路撒冷 朝北的内院门口，在那里有惹动妒忌的偶像的座位，它惹动了妒忌。
EZEK|8|4|看哪，在那里有 以色列 上帝的荣耀，形状与我在平原所见的一样。
EZEK|8|5|上帝对我说：“人子啊，你举目向北观看。”我就举目向北观看，看哪，祭坛门北边的门口有那惹动妒忌的偶像。
EZEK|8|6|他又对我说：“人子啊，你看见 以色列 家所做的吗？他们在这里做了极其可憎的事，使我远离我的圣所。你还要看见另有极其可憎的事。”
EZEK|8|7|他领我到院子门口。我观看，看哪，墙上有一个洞。
EZEK|8|8|他对我说：“人子啊，你要挖墙。”我就挖墙。看哪，有一扇门。
EZEK|8|9|他说：“你进去，看他们在这里所做可憎的恶事。”
EZEK|8|10|于是我进去看。看哪，四面墙上刻着各样爬行的动物、可憎的走兽和 以色列 家各样的偶像。
EZEK|8|11|以色列 家的七十个长老站在这些像前， 沙番 的儿子 雅撒尼亚 也站在其中，各人手拿他的香炉，烟云的香气上腾。
EZEK|8|12|他对我说：“人子啊，你看见 以色列 家的长老，暗中在自己偶像的房间里所做的吗？因为他们说：‘耶和华看不见我们；耶和华已经离弃这地。’”
EZEK|8|13|他又说：“你还要看见他们所做另外极其可憎的事。”
EZEK|8|14|他领我到耶和华殿朝北的门口。看哪，在那里有妇女们坐着，为 搭模斯 哭泣。
EZEK|8|15|他对我说：“人子啊，你看见了吗？你还要看见比这更可憎的事。”
EZEK|8|16|然后他领我到耶和华殿的内院。看哪，在耶和华殿门口、走廊和祭坛中间，约有二十五个人背向耶和华的殿，面向东方，向东拜太阳。
EZEK|8|17|他对我说：“人子啊，你看见了吗？ 犹大 家在这里行可憎的事还算为小吗？他们遍地行残暴，再三惹我发怒。看哪，他们手拿枝条举向鼻前 ！
EZEK|8|18|因此，我也要以愤怒行事。我的眼必不顾惜，也不可怜他们；他们虽在我耳边大声呼求，我还是不听。”
EZEK|9|1|他在我耳边大声喊叫，说：“上前来啊，惩罚这城的人，手中要各拿毁灭的兵器。”
EZEK|9|2|看哪，有六个人从朝北的 上门 而来，各人手里拿着致命的兵器；他们当中有一人身穿细麻衣，腰间系着文士用的墨盒。他们进来，站在铜的祭坛旁。
EZEK|9|3|在基路伯之上， 以色列 上帝的荣耀从那里上升，到殿的入口处。上帝召那身穿细麻衣、腰间系着墨盒的人前来。
EZEK|9|4|耶和华对他说：“你去走遍 耶路撒冷 全城，那些为城中所做可憎之事叹息哀哭的人，你要在他们额上做记号。”
EZEK|9|5|我耳中听见耶和华对其余的人说：“要跟随他走遍全城去击杀。你们的眼不要顾惜，也不要可怜他们。
EZEK|9|6|要将年老的、年轻的、少女、孩童和妇女，从我的圣所开始全都杀尽，只是不可挨近凡有记号的人。”于是他们从殿前的长老杀起。
EZEK|9|7|他对他们说：“要使这殿污秽，使院中遍满被杀的人。你们出去吧！”他们就出去，在城中击杀。
EZEK|9|8|他们击杀的时候，只剩我一人，我就脸伏在地上，呼喊说：“唉！主耶和华啊，你将愤怒倾倒在 耶路撒冷 ，岂要把 以色列 所剩余的人都灭绝吗？”
EZEK|9|9|他对我说：“ 以色列 家和 犹大 家的罪孽极其重大。遍地都有流血的事，满城有冤屈，因为他们说：‘耶和华已经离弃这地，他看不见我们。’
EZEK|9|10|因此，我的眼必不顾惜，也不可怜他们，要照他们所做的报应在他们头上。”
EZEK|9|11|看哪，那身穿细麻衣、腰间系着墨盒的人回覆这事说：“我已经照你所吩咐的做了。”
EZEK|10|1|我观看，看哪，在穹苍之中，也就是基路伯的头上，有蓝宝石的形状，仿佛宝座的形像显在他们上面。
EZEK|10|2|耶和华对那身穿细麻衣的人说：“你进到基路伯下面旋转的轮子中，从基路伯之间取出火炭装满两手掌，撒在城上。” 我亲眼看见他进去。
EZEK|10|3|那人进去的时候，基路伯站在殿的南边，云彩充满了内院。
EZEK|10|4|耶和华的荣耀从基路伯那里上升，到殿的入口处；殿内满布云彩，院子也充满了耶和华荣耀的光辉。
EZEK|10|5|基路伯翅膀的响声传到外院，好像全能上帝说话的声音。
EZEK|10|6|耶和华吩咐那身穿细麻衣的人说：“要从基路伯之间旋转的轮子中取火。”那人就进去站在一个轮子旁边。
EZEK|10|7|基路伯中的一个基路伯伸手到基路伯中间的火那里，取一些放在那身穿细麻衣人的手掌中，那人拿了就出去。
EZEK|10|8|在基路伯翅膀以下，显出有人手的样式。
EZEK|10|9|我又观看，看哪，这些基路伯的旁边有四个轮子。一个基路伯旁有一个轮子，另一个基路伯旁也有一个轮子；轮子的形状好像水苍玉石。
EZEK|10|10|至于四轮的形状，都是一个样式，好像轮中套轮。
EZEK|10|11|轮子行走的时候，向四方都能直行，行走时并不转弯。头转向何方，它们也随着向何方行走，行走时并不转弯。
EZEK|10|12|基路伯的全身，连背带手和翅膀，并轮子周围都布满眼睛。他们四个的轮子都是如此。
EZEK|10|13|我耳中听见这些轮子称为“旋转的轮”。
EZEK|10|14|基路伯各有四张脸：第一是基路伯的脸，第二是人的脸，第三是狮子的脸，第四是鹰的脸。
EZEK|10|15|基路伯升上去了；这就是我在 迦巴鲁河 边所看见的活物。
EZEK|10|16|基路伯行走，轮子也在旁边行走。基路伯展开翅膀，离地上升，轮子也不转离他们的旁边。
EZEK|10|17|基路伯站住，轮子也站住；基路伯上升，轮子也跟着上升，因为活物的灵在轮中。
EZEK|10|18|耶和华的荣耀离开殿的入口处，停在基路伯之上。
EZEK|10|19|基路伯展开翅膀，在我眼前离地上升；他们离去的时候，轮子在旁边，都停在耶和华殿的东门口。在他们上面有 以色列 上帝的荣耀。
EZEK|10|20|这是我在 迦巴鲁河 边所见的活物，他们在 以色列 上帝之下；因此我知道他们是基路伯。
EZEK|10|21|他们各有四张脸、四个翅膀，翅膀以下有人手的样式。
EZEK|10|22|至于他们脸的模样，以及身体的形像 ，正是我从前在 迦巴鲁河 边所看见的。他们各自往前直行。
EZEK|11|1|灵将我举起，带我到耶和华圣殿面向东方的东门。看哪，门口有二十五个人。我见其中有百姓的领袖 押朔 的儿子 雅撒尼亚 和 比拿雅 的儿子 毗拉提 。
EZEK|11|2|耶和华对我说：“人子啊，他们就是图谋罪孽，在这城中设计恶谋的人。
EZEK|11|3|他们说：‘盖房屋的时候尚未临近；这城是锅，我们是肉。’
EZEK|11|4|人子啊，因此你当说预言，说预言攻击他们。”
EZEK|11|5|耶和华的灵降在我身上，对我说：“你当说，耶和华如此说： 以色列 家啊，你们所说的，你们心里所想的，我都知道。
EZEK|11|6|你们在这城里大行屠杀，被杀的人遍满街道。
EZEK|11|7|所以主耶和华如此说：你们在城中杀的人是肉，这城是锅；你们却要从其中被带出去。
EZEK|11|8|你们怕刀剑，我却要使刀剑临到你们。这是主耶和华说的。
EZEK|11|9|我要把你们从这城中带出去，交在外邦人的手里，且要在你们中间施行审判。
EZEK|11|10|你们要仆倒在刀下；我必在 以色列 的边界审判你们，你们就知道我是耶和华。
EZEK|11|11|这城必不作你们的锅，你们也不作锅中的肉。我要在 以色列 的边界审判你们，
EZEK|11|12|你们就知道我是耶和华；因为你们不遵行我的律例，也不顺从我的典章，却随从你们四围列国的规条。”
EZEK|11|13|我正说预言的时候， 比拿雅 的儿子 毗拉提 死了。于是我脸伏在地，大声呼叫说：“唉！主耶和华啊，你要把 以色列 剩余的人都灭绝净尽吗？”
EZEK|11|14|耶和华的话临到我，说：
EZEK|11|15|“人子啊， 耶路撒冷 的居民对你的兄弟、你的本家、你的亲属、 以色列 全家所有的人说：‘你们远离耶和华吧！这地是赐给我们为业的。’
EZEK|11|16|所以你当说：‘主耶和华如此说：我虽将 以色列 全家远远流放到列国，使他们分散在列邦，我却要在他们所到的列邦，暂时作他们的圣所。’
EZEK|11|17|你当说：‘主耶和华如此说：我必从万民中召集你们，从分散的列邦中聚集你们，又将 以色列 地赐给你们。’
EZEK|11|18|他们到了那里，必从其中除掉一切可憎之物、可厌的事。
EZEK|11|19|我要使他们有合一的心，也要将新灵放在你们 里面，又从他们的肉体中除掉石心，赐给他们肉心，
EZEK|11|20|使他们顺从我的律例，谨守遵行我的典章。他们要作我的子民，我要作他们的上帝。
EZEK|11|21|至于那些心中随从可憎之物、可厌的事的人，我必照他们所做的报应在他们头上。这是主耶和华说的。”
EZEK|11|22|于是，基路伯展开翅膀，轮子都在他们旁边；在他们上面有 以色列 上帝的荣耀。
EZEK|11|23|耶和华的荣耀从城中上升，停在城东的那座山上。
EZEK|11|24|灵将我举起，在异象中上帝的灵将我带回 迦勒底 地，到被掳的人那里；之后我所见的异象就离我上升去了。
EZEK|11|25|我就把耶和华指示我的一切事都说给被掳的人听。
EZEK|12|1|耶和华的话临到我，说：
EZEK|12|2|“人子啊，你住在悖逆之家中；他们有眼可看却看不见，有耳可听却听不到，因为他们是悖逆之家。
EZEK|12|3|所以人子啊，你要收拾被掳时需用的物件，白天在他们眼前离去，在他们眼前离开你所住的地方，移到别处去；他们虽是悖逆之家，或者可以领悟。
EZEK|12|4|你要白天在他们眼前拿出你被掳时需用的物件。到了晚上，要在他们眼前离去，像被掳的人离去一样。
EZEK|12|5|你要在他们眼前挖通墙壁，从其中将物件带出去 。
EZEK|12|6|到天黑时，在他们眼前背在肩上带走 ，并要蒙住脸看不见地，因为我要使你成为 以色列 家的预兆。”
EZEK|12|7|我就照着所吩咐的去做，白天拿出被掳时需用的物件。到了晚上，用手挖通墙壁；天黑的时候，在他们眼前背在肩上带走。
EZEK|12|8|次日早晨，耶和华的话临到我，说：
EZEK|12|9|“人子啊， 以色列 家，就是那悖逆之家，岂不是问你说：‘你在做什么呢？’
EZEK|12|10|你要对他们说：‘主耶和华如此说：这是关乎 耶路撒冷 君王和其中 以色列 全家的默示。’
EZEK|12|11|你要说：‘我是你们的预兆：我怎样做，他们所遭遇的也必这样，他们必被掳去，作俘虏。’
EZEK|12|12|他们中间的君王也必在天黑时把物件背在肩上带走。他们要挖通墙壁，从其中带出去 。他必蒙住脸，眼看不见地。
EZEK|12|13|我要把我的网撒在他身上，他就被我的罗网缠住。我要带他到 迦勒底 人之地的 巴比伦 ；他没有看见那地，就死在那里。
EZEK|12|14|我要把四围帮助他的和他所有的军队分散到四方 ，也要拔刀追赶他们。
EZEK|12|15|我把他们驱逐到列国，分散在列邦的时候，他们就知道我是耶和华。
EZEK|12|16|我却要留下他们当中几个人得免刀剑、饥荒、瘟疫，使他们在所到的列国述说自己所做一切可憎的事；他们就知道我是耶和华。”
EZEK|12|17|耶和华的话临到我，说：
EZEK|12|18|“人子啊，你吃饭时必战抖，喝水时必惊惶忧虑。
EZEK|12|19|你要对这地的百姓说：主耶和华论 以色列 地的 耶路撒冷 居民如此说，他们吃饭时必忧虑，喝水时必惊惶，因其中居民所行残暴的事，这地必然荒废，一无所存。
EZEK|12|20|有人居住的城镇必变为废墟，地必荒凉；你们就知道我是耶和华。”
EZEK|12|21|耶和华的话临到我，说：
EZEK|12|22|“人子啊，在 以色列 地你们怎么有这俗语说：‘日子延长，一切异象却落了空’呢？
EZEK|12|23|你要告诉他们说：‘主耶和华如此说：我必令这俗语止息， 以色列 中不再有人引用这俗语。’你却要对他们说：‘日子临近，一切的异象都必应验。’
EZEK|12|24|从此以后， 以色列 家不再有虚假的异象和奉承的占卜。
EZEK|12|25|我─耶和华说话，所说的必定实现，不再耽延。你们这悖逆之家啊，你们在世的日子，我所说的话必定实现。这是主耶和华说的。”
EZEK|12|26|耶和华的话临到我，说：
EZEK|12|27|“人子，看哪， 以色列 家的人说：‘他所见的异象是许多日子以后的事，所说的预言是指着遥远的时候。’
EZEK|12|28|所以你要对他们说：‘主耶和华如此说：我的话不再有一句耽延，我所说的话必定实现。’这是主耶和华说的。”
EZEK|13|1|耶和华的话临到我，说：
EZEK|13|2|“人子啊，你要说预言，攻击 以色列 中说预言的先知，对那些随心说预言的人说：‘你们当听耶和华的话。’”
EZEK|13|3|主耶和华如此说：“祸哉！那些愚顽的先知，随从自己的心意，却一无所见
EZEK|13|4|以色列 啊，你的先知好像废墟中的狐狸，
EZEK|13|5|没有上去堵住缺口，也没有为 以色列 家重修城墙，使它在耶和华的日子来临时，可以在战争中站得住。
EZEK|13|6|他们看见的是虚假，是谎诈的占卜，说是耶和华说的；其实耶和华并没有差遣他们，他们却指望那话必站立得住。
EZEK|13|7|你们岂不是见了虚假的异象吗？岂不是说了谎诈的占卜吗？你们说，这是耶和华说的，其实我没有说过。”
EZEK|13|8|所以主耶和华如此说：“因你们说的是虚假，见的是谎诈，所以，看哪，我要敌对你们。这是主耶和华说的。
EZEK|13|9|我的手必攻击那见虚假异象、用谎诈占卜的先知，他们必不列在我百姓的会中，不录在 以色列 家的名册上，也不能进入 以色列 地；你们就知道我是主耶和华。
EZEK|13|10|他们诱惑我的百姓，说：‘平安！’其实没有平安，就像有人筑墙壁，看哪，他们倒去粉刷它。
EZEK|13|11|所以你要对那些粉刷的人说：‘墙要倒塌，暴雨漫过。你们大冰雹啊，要降下 ，狂风要吹裂这墙。’
EZEK|13|12|看哪，这墙倒塌，人岂不是要问你们说：‘你们所粉刷的在哪里呢？’”
EZEK|13|13|所以主耶和华如此说：“我要发怒，使狂风吹裂它，在怒中令暴雨漫过，又发怒降下大冰雹，毁坏它。
EZEK|13|14|我要这样拆毁你们那粉饰的墙，把它夷为平地，以致根基露出；墙一倒塌，你们也要在其中灭亡。你们就知道我是耶和华。
EZEK|13|15|我要对墙和粉刷它的人发尽我的愤怒，我 要对你们说：‘墙没有了！粉刷它的人也没有了！’
EZEK|13|16|这就是 以色列 的先知，他们指着 耶路撒冷 说预言，见到这城平安的异象，其实没有平安。这是主耶和华说的。”
EZEK|13|17|“你，人子啊，要面向你百姓中随心说预言的妇女们，说预言攻击她们，
EZEK|13|18|说，主耶和华如此说：‘这些妇女有祸了！她们为众人的手腕缝驱邪带，替身材高矮不同的人做头巾，为要猎取人的性命。难道你们要猎取我百姓的性命，使自己存活吗？
EZEK|13|19|你们为几把大麦、几块饼，在我的百姓中亵渎我，对那肯听谎言的百姓说谎言，让不该死的人死，让不该活的人活。’”
EZEK|13|20|所以主耶和华如此说：“看哪，我要对付你们那用以猎取人，如猎飞鸟般的驱邪带。我要把驱邪带从你们的手腕扯去，释放那些如飞鸟被你们猎取的人。
EZEK|13|21|我也必撕裂你们的头巾，救我百姓脱离你们的手，使他们不再被猎取，落在你们手中；你们就知道我是耶和华。
EZEK|13|22|我未曾使义人伤心，你们却以谎话使他伤心，且又坚固恶人的手，不使他回转离开恶道得以存活。
EZEK|13|23|所以，你们必不再看见虚假的异象，也不再行占卜的事；我要救我的百姓脱离你们的手；你们就知道我是耶和华。”
EZEK|14|1|有几个 以色列 的长老到我这里来，坐在我面前。
EZEK|14|2|耶和华的话临到我，说：
EZEK|14|3|“人子啊，这些人在心中设立偶像，把陷自己于罪的绊脚石放在面前，我真的能让他们求问吗？
EZEK|14|4|所以你要告诉他们，对他们说：‘主耶和华如此说： 以色列 家的人，凡在心中设立偶像，把陷自己于罪的绊脚石放在面前，却来到先知那里的，我─耶和华在他所求的事上，必因他拜许多偶像向他施行报应 ，
EZEK|14|5|为要夺回 以色列 家的心，他们全都拜偶像，与我疏远了。’
EZEK|14|6|“所以你要对 以色列 家说：‘主耶和华如此说：回转吧！回转离开你们的偶像，转脸离开一切可憎的事。’
EZEK|14|7|因为 以色列 家的人，或在 以色列 中寄居的外人，凡与我隔绝，在心中设立偶像，把陷自己于罪的绊脚石放在面前，却来到先知那里，要为自己的事求问我的，我─耶和华必亲自报应他。
EZEK|14|8|我要向那人变脸，使他成为警戒和笑柄，并且我要把他从我民中剪除；你们就知道我是耶和华。
EZEK|14|9|先知若被骗说了一句预言，是我─耶和华骗了那先知，我要伸手攻击他，把他从我百姓 以色列 中除灭。
EZEK|14|10|他们必担当自己的罪孽。先知的罪孽和求问之人的罪孽都一样，
EZEK|14|11|使 以色列 家不再走迷离开我，也不再因各样的罪过玷污自己，却要作我的子民，我也作他们的上帝。这是主耶和华说的。”
EZEK|14|12|耶和华的话临到我，说：
EZEK|14|13|“人子啊，若有一国犯罪干犯我，我也伸手攻击它，断绝他们粮食的供应，使饥荒临到那地，将人与牲畜从其中剪除；
EZEK|14|14|虽有 挪亚 、 但以理 、 约伯 这三人在那里，他们只能因自己的义救自己的命。这是主耶和华说的。
EZEK|14|15|我若使恶兽经过那地，大肆蹂躏，使地荒凉，以致因这些兽，人都不得经过；
EZEK|14|16|虽有这三人在其中，主耶和华说：我指着我的永生起誓，他们不能救儿子女儿，只有他们自己可以得救，那地仍然荒凉。
EZEK|14|17|或者我使刀剑临到那地，说：‘让刀剑穿越那地’，以致我把人与牲畜从其中剪除；
EZEK|14|18|虽有这三人在其中，主耶和华说：我指着我的永生起誓，他们不能救儿子女儿，只有他们自己可以得救。
EZEK|14|19|或者我叫瘟疫流行那地，把我的愤怒带着血倾在其中，好使人与牲畜从其中剪除；
EZEK|14|20|虽有 挪亚 、 但以理 、 约伯 在那里，主耶和华说：我指着我的永生起誓，他们不能救儿子女儿，只能因自己的义救自己的命。
EZEK|14|21|“主耶和华如此说：我若将这四样大灾，就是刀剑、饥荒、恶兽、瘟疫降在 耶路撒冷 ，将人与牲畜从其中剪除，岂不是更严重吗？
EZEK|14|22|看哪，在那里必有幸免于难的人带着儿子女儿；看哪，他们来到你们这里；你们看见他们的所作所为，就会因我降给 耶路撒冷 的灾祸，因我降给它的一切，得到安慰。
EZEK|14|23|你们因看见他们的所作所为，得到安慰，就会知道我在 耶路撒冷 所做的并非毫无缘故。这是主耶和华说的。”
EZEK|15|1|耶和华的话临到我，说：
EZEK|15|2|“人子啊，葡萄树比一切其他的树，就是树林里众树木的树枝，有什么长处呢？
EZEK|15|3|可以从其中取木料来做工吗？人可以拿来做钉子，挂东西在上面吗？
EZEK|15|4|看哪，它已经抛在火中当柴烧，火既烧了两头，中间也烧焦了，它还有什么用处呢？
EZEK|15|5|看哪，它完整的时候尚且不能拿来做工，何况被火烧焦了，还能拿来做工吗？
EZEK|15|6|所以，主耶和华如此说：我怎样使林中树里的葡萄树在火中当柴烧，我也必照样对待 耶路撒冷 的居民。
EZEK|15|7|我必向他们变脸；他们虽从火中逃出来，火仍要烧灭他们。我向他们变脸的时候，你们就知道我是耶和华。
EZEK|15|8|我必使这地荒凉，因为他们做了背叛的事。这是主耶和华说的。”
EZEK|16|1|耶和华的话临到我，说：
EZEK|16|2|“人子啊，你要使 耶路撒冷 知道它那些可憎的事。
EZEK|16|3|你要说，主耶和华对 耶路撒冷 如此说：你的根源，你的出身，是在 迦南 地；你的父亲是 亚摩利 人，母亲是 赫 人。
EZEK|16|4|论到你出世的景况，在你出生的日子没有人为你断脐带，也没有用水清洗，使你洁净；没有人撒盐在你身上，也没有人用布包你。
EZEK|16|5|没有人顾惜你，为你做一件这样的事来可怜你。你却被扔在田野上面，因你出生的日子就被厌恶。
EZEK|16|6|“我从你旁边经过，见你在血中打滚，就对你说：‘你虽在血中，却要活下去！’我又说：‘你虽在血中，却要活下去！’
EZEK|16|7|我使你成长如田间所生长的；你就渐长，美而又美 ，两乳成形，头发秀长，但你仍然赤身露体。
EZEK|16|8|“我从你旁边经过看见你，看哪，正是你渴慕爱情的时候，我就用我衣服的边搭在你身上，遮盖你的赤体；又向你起誓，与你立约，你就归我。这是主耶和华说的。
EZEK|16|9|那时我用水洗你，洗净你身上的血，又用油抹你。
EZEK|16|10|我使你身穿锦绣衣裳，脚穿海狗皮鞋，用细麻布裹着你，精致衣料披在你身上。
EZEK|16|11|我用首饰打扮你：我把手镯戴在你手上，项链在你颈上，
EZEK|16|12|我也把环子戴在你鼻上，耳环在你耳上，华冠在你头上。
EZEK|16|13|这样，你就有金银的首饰，穿的是细麻衣和精致衣料，以及锦绣衣裳；吃的是细面、蜂蜜和油。你也极其美貌，配登王后之位。
EZEK|16|14|你美貌的名声传到列国，因我加给你荣华，使你完美。这是主耶和华说的。
EZEK|16|15|“只是你仗着自己美貌，又凭着你的名声行淫。你向路人纵情淫乱，你的美貌就属于他的了 。
EZEK|16|16|你拿你的衣服为自己做成彩色丘坛，在其上行淫。这样的事本不该有，以后也不该发生。
EZEK|16|17|你拿我所赐给你的那些美丽的金银宝物，为自己制造男性的偶像，与它们行淫；
EZEK|16|18|你拿你的锦绣衣裳为它们披上，把我的膏油和香料摆在它们面前；
EZEK|16|19|你把我赐给你的食物，就是我赐给你享用的细面、油和蜂蜜，都摆在它们面前作为馨香的供物。事情就是这样。这是主耶和华说的。
EZEK|16|20|你拿你为我所生的儿女献给它们吞噬。你的淫乱岂是小事？
EZEK|16|21|你竟把我的儿女杀了，使他们经火献给它们！
EZEK|16|22|你做这一切可憎和淫乱的事，并未追念你幼年的日子，那时你赤身露体，在血中打滚。”
EZEK|16|23|“你有祸了！你有祸了！这是主耶和华说的。你做这一切恶事之后，
EZEK|16|24|又为自己建造土墩，在各广场上筑起高台。
EZEK|16|25|你在各个街头建造高台，使你的美貌变为可憎；又向所有过路的人招手 ，多行淫乱。
EZEK|16|26|你也和你那放纵情欲的邻邦 埃及 人行淫，增添你的淫乱，惹我发怒。
EZEK|16|27|看哪，我伸手攻击你，减少你的福分，却将你交给恨恶你的 非利士 人 ，让他们任意待你。他们为你的淫行也感到羞耻。
EZEK|16|28|你尚且不满意，又与 亚述 人行淫，但与他们行淫之后，仍不满足；
EZEK|16|29|于是你与那称为贸易之地的 迦勒底 多行淫乱，即使这样，你仍不满足。
EZEK|16|30|“你的心何等脆弱！这是主耶和华说的。你做这一切事，都是不知羞耻的妓女所做的，
EZEK|16|31|在各个街头建造土墩，在各广场上筑高台；但你藐视行淫的赏金，又不像妓女。
EZEK|16|32|你这行淫的妻子啊，竟然接外人，替代丈夫。
EZEK|16|33|凡妓女都是得人赠礼，你反倒馈赠你所爱的人，倒贴他们，使他们从四围来与你行淫。
EZEK|16|34|你的淫行与其他妇女相反，不是人要求与你行淫；是你给人赏金，不是人给你赏金；你是相反的。”
EZEK|16|35|“你这妓女啊，要听耶和华的话。
EZEK|16|36|主耶和华如此说：因你放纵情欲，露出下体，与你所爱的行淫，因你敬拜一切可憎的偶像，就像 自己儿女的血献给它们，
EZEK|16|37|所以，看哪，我要聚集所有与你交欢的情人，不论是你所爱的或你所恨的，聚集他们从四围到你那里来；我要在他们面前暴露你的下体，使他们看尽你的下体。
EZEK|16|38|我也要审判你，如审判淫妇和流人血的妇女一样。我要在愤怒和妒忌中使流血的罪归到你身上。
EZEK|16|39|我要把你交在他们手中；他们必拆毁你的土墩，毁坏你的高台，剥去你的衣服，夺取你美丽的宝物，留下你赤身露体。
EZEK|16|40|他们必聚集众人攻击你，用石头打死你，用刀剑刺透你，
EZEK|16|41|用火焚烧你的房屋，在许多妇女眼前审判你。我必使你不再行淫，你也不再给赏金。
EZEK|16|42|我止息了向你所发的愤怒，我的妒忌也离开了你；这样，我就平静，不再恼怒。
EZEK|16|43|因你不追念幼年的日子，反而在这一切的事上惹我发烈怒，所以，看哪，我必照你所做的报应在你头上。在你一切可憎的事上，你不是还行了淫乱吗？这是主耶和华说的。”
EZEK|16|44|“看哪，凡说俗语的必用这俗语攻击你，说：‘有其母必有其女。’
EZEK|16|45|你实在是你母亲的女儿，厌弃丈夫和儿女；你也是你姊妹的姊妹，厌弃丈夫和儿女。你的母亲是 赫 人，父亲是 亚摩利 人。
EZEK|16|46|你的姊姊是 撒玛利亚 ，她和她的女儿们住在你北边；你的妹妹是 所多玛 ，她和她的女儿们住在你南边。
EZEK|16|47|你不只效法她们的行为，照她们可憎的事去做，不消多时 ，你所做的一切就比她们更恶。
EZEK|16|48|主耶和华说：我指着我的永生起誓，你的妹妹 所多玛 与她的女儿们并未做你和你女儿们所做的事。
EZEK|16|49|看哪，你的妹妹 所多玛 的罪孽是这样：她和她的女儿们都骄傲，粮源充足，大享安逸，却不扶持困苦和贫穷人的手。
EZEK|16|50|她们狂傲，在我面前做可憎的事，我看见了就把她们除掉。
EZEK|16|51|撒玛利亚 所犯的罪不及你的一半，你所做可憎的事比她更多；比起你所做这一切可憎的事，你的姊妹倒显为义。
EZEK|16|52|你既为你的姊妹辩护，就要担当自己的羞辱。因你所犯的罪比她们更可憎，她们比你倒显为义；你既使你的姊妹显为义，就要抱愧，担当自己的羞辱。”
EZEK|16|53|“我必使她们被掳的归回，使 所多玛 和她的女儿们、 撒玛利亚 和她的女儿们，并与你一起被掳的都归回；
EZEK|16|54|好使你担当自己的羞辱，为所做的一切抱愧，让她们得到安慰。
EZEK|16|55|你的妹妹 所多玛 和她的女儿们必回复原状； 撒玛利亚 和她的女儿们必回复原状；你和你的女儿们也必回复原状。
EZEK|16|56|在你骄傲的日子，你的妹妹 所多玛 岂不是你口中的笑柄吗？
EZEK|16|57|在你的恶行显露以前，那受了凌辱的 亚兰 女儿们和 亚兰 四围 非利士 的女儿们，都在四围藐视你。
EZEK|16|58|耶和华说：你的淫荡和可憎之事，你自己要担当。”
EZEK|16|59|“主耶和华如此说：你这轻看誓言而背约的，我必照你所做的报应你。
EZEK|16|60|然而我要追念在你幼年时我与你所立的约，也要与你立定永约。
EZEK|16|61|当你接纳你的姊姊和妹妹时，你要追念你所行的，自觉惭愧；并且我要将她们赏给你做女儿，却不是按着我与你所立的约。
EZEK|16|62|我要坚定与你所立的约，你就知道我是耶和华，
EZEK|16|63|使你在我赦免你一切恶行时，心中追念，自觉惭愧，又因羞辱就不再开口。这是主耶和华说的。”
EZEK|17|1|耶和华的话临到我，说：
EZEK|17|2|“人子啊，你要向 以色列 家出谜语，设比喻，
EZEK|17|3|说，主耶和华如此说：有一只大鹰，翅膀大，翎毛长，羽毛丰满，色彩缤纷；它飞到 黎巴嫩 ，啄去香柏树梢，
EZEK|17|4|啄断它顶端的嫩枝，叼到贸易之地，放在商业城中。
EZEK|17|5|它又从这地取了一些种子，种在肥沃的田里，栽于丰沛的水源旁，如种植柳树。
EZEK|17|6|它渐渐生长，成为低矮蔓生的葡萄树；树枝伸向那鹰，根部在它下面。这样，它就长成了一棵葡萄树，生出枝子，长出枝干。
EZEK|17|7|“有一只 大鹰，翅膀大，羽毛多。看哪，葡萄树从栽种它的苗圃向这鹰伸出根来，长出枝子，期盼从它得到浇灌。
EZEK|17|8|这棵树栽于肥田丰沛的水源旁，原是为了生枝、结果，成为佳美的葡萄树。
EZEK|17|9|你要说，主耶和华如此说：这棵葡萄树岂能发旺呢？鹰岂不拔出它的根来，摘光它的果子，使它枯干，连长出的嫩叶都枯萎了吗？要把它连根拔除，并不需要费大力或动用许多人。
EZEK|17|10|看哪，葡萄树虽然栽种了，岂能发旺呢？一经东风击打，岂不全然枯干了吗？它必在生长的苗圃中枯干了。”
EZEK|17|11|耶和华的话临到我，说：
EZEK|17|12|“你要对那悖逆之家说：你们不知道这些事是什么意思吗？你要这样说，看哪， 巴比伦 王曾到 耶路撒冷 ，把其中的君王和官长带到 巴比伦 去，
EZEK|17|13|又从 以色列 王室后裔中选取一人，与他立约，令他发誓，又掳走国中有势力的人，
EZEK|17|14|使王国衰弱，不再强盛，只能靠守盟约方得生存。
EZEK|17|15|他却背叛 巴比伦 王，差派使者前往 埃及 ，要求 埃及 人给他马匹和许多人。他岂能亨通呢？这样做的人岂能逃脱呢？他背了约岂能逃脱呢？
EZEK|17|16|主耶和华说：我指着我的永生起誓，他定要死在 巴比伦 ，就是 巴比伦 王所在之处；因为 巴比伦 王立他为王，他竟轻看向王所起的誓，背弃王与他所立的约。
EZEK|17|17|当敌人建土堆，筑堡垒，要歼灭许多人时，法老虽有强大军队和大批人马，在战场上还是不能帮助他。
EZEK|17|18|他轻看誓言，背弃盟约，看哪，虽已投降 ，却又做这一切的事，他必不能逃脱。
EZEK|17|19|所以主耶和华如此说：我指着我的永生起誓，他既轻看我的誓言，背弃我的约，我必使这罪归到他头上。
EZEK|17|20|我要把我的网撒在他身上，他就被我的罗网缠住。我要带他到 巴比伦 ，在那里因他背叛我的罪惩罚他。
EZEK|17|21|所有逃跑的 军队必倒在刀下；剩余的也必分散四方 。你们就知道说这话的是我─耶和华。”
EZEK|17|22|主耶和华如此说：“我要从香柏树高高的树梢摘取并栽上，从顶端的嫩枝中折下一嫩枝，栽于极高的山上，
EZEK|17|23|栽在 以色列 高处的山上。它就生枝、结果，成为高大的香柏树，各类飞禽中的鸟都来宿在其下，宿在枝子的荫下 。
EZEK|17|24|田野的树木因此就知道是我─耶和华使高树矮小，使矮树高大，使绿树枯干，使枯树发旺。我─耶和华说了这话，就必成就。”
EZEK|18|1|耶和华的话又临到我，说：
EZEK|18|2|“你们在 以色列 地何以有这俗语，‘父亲吃了酸葡萄，儿子牙齿就酸倒’呢？
EZEK|18|3|主耶和华说：我指着我的永生起誓，你们在 以色列 必不再引用这俗语。
EZEK|18|4|看哪，所有的生命都是属我的；父亲的生命怎样属我，儿子的生命也照样属我；然而犯罪的，他必定死。
EZEK|18|5|“人若是公义，行公平公义的事：
EZEK|18|6|未曾在山上吃祭物，未曾向 以色列 家的偶像举目；未曾污辱邻舍的妻，也未曾在妇人的经期间亲近她；
EZEK|18|7|未曾亏负人，而是将欠债之人的抵押品还给他；未曾抢夺人的物件，却把食物给饥饿的人吃，把衣服给赤身的人穿；
EZEK|18|8|未曾向人取利息，也未曾索取高利，反倒缩手不作恶，在人与人之间施行诚实的判断；
EZEK|18|9|遵行我的律例，谨守我的典章，按诚实行事 ；这人是公义的，必要存活。这是主耶和华说的。
EZEK|18|10|“他若生了儿子，儿子作强盗，流人的血，作父亲的 虽然未犯此过，儿子却对弟兄 行了以上所说的恶，在山上吃祭物，污辱邻舍的妻；
EZEK|18|11|
EZEK|18|12|亏负困苦和贫穷的人，抢夺别人的物件，不归还抵押品，却向偶像举目，做可憎的事；
EZEK|18|13|向人取利息，索取高利，这人岂能存活呢？他不能存活。他因做这一切可憎的事，必要死亡，他的血要归到自己身上。
EZEK|18|14|“看哪，他若生了儿子，儿子见父亲所犯的一切罪，他见了，却不照样去做；
EZEK|18|15|他未曾在山上吃祭物，未曾向 以色列 家的偶像举目，未曾污辱邻舍的妻；
EZEK|18|16|也未曾亏负人，未曾取人的抵押品，未曾抢夺人的物件，却把食物给饥饿的人吃，把衣服给赤身的人穿，
EZEK|18|17|缩手不害困苦人，未曾向人索取利息或高利；反倒顺从我的典章，遵行我的律例；如此，他必不因父亲的罪孽死亡，定要存活。
EZEK|18|18|至于他父亲，因为施行欺压，抢夺弟兄，在百姓中行不善，看哪，他必因自己的罪孽死亡。
EZEK|18|19|“你们还说：‘儿子为什么不担当父亲的罪孽呢？’儿子若行公平公义的事，谨守遵行我一切的律例，他必要存活。
EZEK|18|20|惟有犯罪的，却必死亡。儿子不担当父亲的罪孽，父亲也不担当儿子的罪孽。义人的善果要归自己，恶人的恶报也要归自己。
EZEK|18|21|“恶人若回转离开所做的一切罪恶，谨守我的一切律例，行公平公义的事，他必要存活，不致死亡。
EZEK|18|22|他所犯的一切罪过都不被记念；他因所行的义，必要存活。
EZEK|18|23|恶人死亡，岂是我所喜悦的呢？我岂不是喜悦他回转离开所行的道而存活吗？这是主耶和华说的。
EZEK|18|24|至于义人，他若转离义行而作恶，照着恶人所做一切可憎的事去做，岂能存活呢？他所行的一切义都不被记念；反而因所行的恶、所犯的罪死亡。
EZEK|18|25|“你们却说：‘主的道不公平！’ 以色列 家啊，你们要听，我的道不公平吗？你们的道不是不公平吗？
EZEK|18|26|义人若转离义行而作恶，他就因这些恶而死亡。他要死在他所作的恶中。
EZEK|18|27|恶人若回转离开所行的恶，行公平公义的事，他必救自己的命；
EZEK|18|28|因为他省察，回转离开所犯的一切罪过，他必要存活，不致死亡。
EZEK|18|29|以色列 家还说：‘主的道不公平！’ 以色列 家啊，我的道不公平吗？你们的道不是不公平吗？
EZEK|18|30|所以， 以色列 家啊，我必按你们各人所做的审判你们。当回转，回转离开你们一切的罪过，免得罪孽成为你们的绊脚石。这是主耶和华说的。
EZEK|18|31|你们要把所犯的一切罪过尽行抛弃，为自己造一个新的心和新的灵。 以色列 家啊，你们为什么要死呢？
EZEK|18|32|我不喜欢有任何人死亡，所以你们当回转，要存活！这是主耶和华说的。”
EZEK|19|1|你当为 以色列 的领袖们唱哀歌，
EZEK|19|2|说： 你的母亲在狮子中 是怎样的母狮呢？ 它蹲伏在少壮狮子中， 养育小狮子。
EZEK|19|3|它养大了其中一只小狮子， 成了少壮狮子， 学会抓食， 它就吃人。
EZEK|19|4|列国听见了就把它逮住在他们的坑里， 用钩子拉它到 埃及 地去。
EZEK|19|5|母狮见自己等候， 期望落空， 就从小狮子中取一只 ， 养为少壮狮子；
EZEK|19|6|它在众狮子中徜徉， 长大成为少壮狮子， 学会抓食， 它就吃人。
EZEK|19|7|它拆毁他们的宫殿 ， 使他们的城镇变为废墟； 因它咆哮的声音， 遍地和其中所充满的都荒废了。
EZEK|19|8|于是四围列国 从各省前来攻击它， 把网撒在它身上， 把它逮住在他们的坑里。
EZEK|19|9|他们又用钩子钩住它，把它放入笼中， 带到 巴比伦 王那里， 把它押进城堡， 以色列 山上就不再听见它的声音。
EZEK|19|10|你的母亲如葡萄树， 在葡萄园中 ， 栽于水边，因为水多， 就多结果子，多生枝子；
EZEK|19|11|它长出坚固的枝干， 可作统治者的权杖。 这枝干高举在茂密的树枝中， 可见树身高大，枝子繁多。
EZEK|19|12|但在烈怒中它被拔出，摔在地上； 东风吹干其果子， 那坚固的枝干因折断而枯干， 被火烧毁；
EZEK|19|13|如今这葡萄树移植于旷野， 在干旱无水之地，
EZEK|19|14|火从枝干中发出， 烧灭它的枝条和它的果子 ， 以致不再有坚固的枝干， 可作统治者的权杖。 这是哀伤之歌，成为一首哀歌。
EZEK|20|1|第七年五月初十，有 以色列 的几个长老前来求问耶和华，坐在我面前。
EZEK|20|2|耶和华的话临到我，说：
EZEK|20|3|“人子啊，你要告诉 以色列 的长老，对他们说，主耶和华如此说：你们来是为求问我吗？主耶和华说：我指着我的永生起誓，我必不让你们求问。
EZEK|20|4|人子啊，你要审问他们吗？你要审问吗？你当使他们知道他们祖先那些可憎的事；
EZEK|20|5|你要对他们说，主耶和华如此说：当日我拣选 以色列 ，对 雅各 家的后裔起誓，在 埃及 地向他们显现，起誓说：我是耶和华─你们的上帝；
EZEK|20|6|那日我向他们起誓，要领他们出 埃及 地，到我为他们所找到的流奶与蜜之地，就是全地中最美好之地。
EZEK|20|7|我对他们说，你们各人要抛弃眼中所喜爱的可憎之物，不可用 埃及 的偶像玷污自己。我是耶和华─你们的上帝。
EZEK|20|8|他们却悖逆我，不肯听从我，不抛弃他们眼中所喜爱的可憎之物，离弃 埃及 的偶像。 “我就说，在 埃及 地，我要把我的愤怒倾倒在他们身上，向他们发尽我的怒气。
EZEK|20|9|我这么做是为了我名的缘故，免得我的名在他们所居住之列国眼中被亵渎；我曾在这些列国眼前向他们显现，领他们出了 埃及 地。
EZEK|20|10|我领他们出 埃及 地，带他们到旷野。
EZEK|20|11|我将我的律例赐给他们，将我的典章指示他们；人若遵行就必因此存活。
EZEK|20|12|我将我的安息日赐给他们，在我与他们中间作记号，让他们知道我─耶和华是使他们分别为圣的。
EZEK|20|13|以色列 家却在旷野中悖逆我，不顺从我的律例，厌弃我的典章；人若遵行就必因此存活。他们却大大干犯我的安息日。 “因此我说，我要在旷野把我的愤怒倾倒在他们身上，灭绝他们。
EZEK|20|14|我这么做是为了我名的缘故，免得我的名在列国眼中被亵渎，因为在这些列国眼前我领了他们出来。
EZEK|20|15|并且我在旷野向他们起誓，必不领他们进入我所赐的流奶与蜜之地，就是全地中最美好之地；
EZEK|20|16|因为他们厌弃我的典章，不顺从我的律例，干犯我的安息日，他们的心随从自己的偶像。
EZEK|20|17|虽然如此，我的眼仍顾惜他们，不毁灭他们，不在旷野把他们灭绝净尽。
EZEK|20|18|“我在旷野对他们的儿女说：‘不要遵行你们祖先的律例，不要谨守他们的规条，也不要用他们的偶像玷污自己。
EZEK|20|19|我是耶和华─你们的上帝，你们要顺从我的律例，谨守遵行我的典章，
EZEK|20|20|且以我的安息日为圣。这日必在我与你们中间作记号，使你们知道我是耶和华─你们的上帝。’
EZEK|20|21|只是他们的儿女悖逆我，不顺从我的律例，也不谨守遵行我的典章；人若遵行就必因此存活。他们却干犯我的安息日。 “因此我说，我要在旷野把我的愤怒倾倒在他们身上，向他们发尽我的怒气。
EZEK|20|22|但我却缩手而未如此行；我这么做是为了我名的缘故，免得我的名在列国眼中被亵渎，因为在这些列国眼前我领了他们出来。
EZEK|20|23|并且我在旷野向他们起誓，要把他们驱散到列国，分散在列邦；
EZEK|20|24|因为他们不遵行我的典章，厌弃我的律例，干犯我的安息日，眼目向着他们祖先的偶像。
EZEK|20|25|我也任他们遵行那无益的律例，随从那不能使人存活的规条。
EZEK|20|26|他们使所有头生的经火，我就任凭他们在这供物上玷污自己；我令他们惊恐，他们就知道我是耶和华。
EZEK|20|27|“人子啊，你要告诉 以色列 家，对他们说，主耶和华如此说：你们的祖先在背叛我的事上再次亵渎了我；
EZEK|20|28|我领他们到我起誓应许赐给他们的地，他们看见各高冈、各茂密的树，就在那里献祭，献上惹我发怒的供物，也在那里焚烧馨香的祭，献浇酒祭。
EZEK|20|29|我就对他们说：你们去的那丘坛叫什么呢？它名叫 巴麻 ，直到今日。
EZEK|20|30|所以你要对 以色列 家说，主耶和华如此说：你们仍要照你们祖先所做的玷污自己吗？还要照他们可憎的事行淫吗？
EZEK|20|31|当你们献上供物，使你们儿子经火的时候，你们仍用各样的偶像玷污自己，直到今日。 以色列 家啊，我岂能让你们求问呢？主耶和华说：我指着我的永生起誓，我必不让你们求问。
EZEK|20|32|“你们说：‘我们要像列国和列邦的宗族一样，去事奉木头与石头。’你们所起的心意万不能成就。”
EZEK|20|33|“主耶和华说：我指着我的永生起誓，我要作王，用大能的手和伸出的膀臂，并倾倒出来的愤怒治理你们。
EZEK|20|34|我必用大能的手和伸出的膀臂，并倾倒出来的愤怒，把你们从万民中领出来，从被赶散到的列邦聚集你们。
EZEK|20|35|我必带你们到万民的旷野，在那里当面审判你们。
EZEK|20|36|我怎样在 埃及 地的旷野审判你们的祖先，也必照样审判你们。这是主耶和华说的。
EZEK|20|37|我要使你们从杖下经过，按着约的拘束 带领你们。
EZEK|20|38|我必从你们中间除尽叛逆和得罪我的人；我将他们从所寄居的地方领出来，他们却不得进入 以色列 地，你们就知道我是耶和华。
EZEK|20|39|“你们， 以色列 家啊，主耶和华如此说：你们若不听从我，从今以后就让各人去事奉他的偶像吧，只是不可再以你们的供物和偶像亵渎我的圣名。
EZEK|20|40|“在我的圣山，就是 以色列 高处的山， 以色列 全家，那地所有的人，都要在那里事奉我。在那里我悦纳他们，并要你们献供物和初熟的土产，以及一切的圣物。这是主耶和华说的。
EZEK|20|41|我把你们从万民中领出来，从被赶散到的列邦聚集你们，那时我必悦纳你们如同悦纳馨香之祭，我要在列国眼前，在你们中间显为圣。
EZEK|20|42|我领你们进入 以色列 地，就是我起誓应许赐给你们列祖之地，那时你们就知道我是耶和华。
EZEK|20|43|你们在那里要追念那玷污自己的所作所为，又要因所行的一切恶事厌恶自己。
EZEK|20|44|以色列 家啊，我为我名的缘故，没有照着你们的恶行和你们的败坏对待你们；你们就知道我是耶和华。这是主耶和华说的。”
EZEK|20|45|耶和华的话临到我，说：
EZEK|20|46|“人子啊，你要面向南方，向南方传讲 ，向 尼革夫 田野的树林说预言。
EZEK|20|47|你要对 尼革夫 的树林说，要听耶和华的话。主耶和华如此说：看哪，我要在你那里点火，烧灭你们中间所有的绿树和枯树，猛烈的火焰必不熄灭；从南到北，人的脸都被烧焦。
EZEK|20|48|凡血肉之躯都知道是我─耶和华点了火，这火必不熄灭。”
EZEK|20|49|于是我说：“唉！主耶和华啊，人都指着我说：他不是说比喻的人吗？”
EZEK|21|1|耶和华的话临到我，说：
EZEK|21|2|“人子啊，把你的脸正对着 耶路撒冷 ，对着圣所 传讲 ，向 以色列 地说预言。
EZEK|21|3|你要向 以色列 地说，耶和华如此说：看哪，我与你为敌，拔刀出鞘，把义人和恶人从你中间剪除。
EZEK|21|4|因为我要剪除你当中的义人和恶人，所以我的刀要出鞘，从南到北攻击所有的血肉之躯；
EZEK|21|5|凡血肉之躯都知道我─耶和华已拔刀出鞘，刀必不再入鞘。
EZEK|21|6|你，人子啊，要叹息，在他们眼前断了腰，愁苦地叹息。
EZEK|21|7|若有人对你说：‘你为什么叹息呢？’你就说：‘因为有风声传来，人心惶惶，双手发软，精神衰败，膝弱如水。看哪，它临近了，一定会发生。’这是主耶和华说的。”
EZEK|21|8|耶和华的话临到我，说：
EZEK|21|9|“人子啊，你要预言说，耶和华如此吩咐，你要说： 有刀，刀已磨快， 又擦亮了；
EZEK|21|10|磨快为要大大杀戮， 擦亮为要像闪电。 我们岂能快乐呢？ 它藐视我儿的权杖和一切的木头 。
EZEK|21|11|它已经交给人擦亮，可以掌握使用；这刀已经磨快擦亮，好交在行杀戮的人手中。
EZEK|21|12|人子啊，你要呼喊哀号，因为这刀将临到我的百姓，临到 以色列 所有的领袖身上。他们和我的百姓都要交在刀下，所以你要捶胸 。
EZEK|21|13|因为这是一个考验，若它藐视权杖，也不算一回事，又怎么样呢？这是主耶和华说的。”
EZEK|21|14|“人子啊，你要拍掌预言，使这刀三番两次临到；这是致人死伤的刀，就是包围人，使人大受死伤的刀。
EZEK|21|15|我设立这恐吓 的刀，攻击他们一切的城门，为要使他们的心惊慌害怕，许多人因而跌倒。唉！它 造得像闪电，磨得尖利 ，要行杀戮。
EZEK|21|16|刀啊，要行动一致 ，向右边，或指向左边；面向哪方，就向哪方。
EZEK|21|17|我也要拍掌，使我的愤怒平息。这是我─耶和华说的。”
EZEK|21|18|耶和华的话临到我，说：
EZEK|21|19|“人子啊，你要画定两条路线，使 巴比伦 王的刀过来，这两条路必从同一地分出来；要在通往城里的路口画手作指标。
EZEK|21|20|你要划定一条路，使刀来到 亚扪 人的 拉巴 ，来到 犹大 ，在坚固城 耶路撒冷 。
EZEK|21|21|因为 巴比伦 王站在岔路上，在两条路口占卜。他摇签 求问神像，察看肝脏；
EZEK|21|22|右手是 耶路撒冷 的占卜，以便安设撞城槌，张口喊杀 ，扬声呼叫，建土堆，筑堡垒，以撞城槌攻打城门。
EZEK|21|23|在那些曾郑重起誓的 犹大 人眼中，这是虚假的占卜；但 巴比伦 王要使他们想起自己的罪孽，以便俘掳他们。”
EZEK|21|24|于是，主耶和华如此说：“因你们的过犯显露，你们的罪孽被记得，以致你们的罪恶在你们一切的行为上都彰显出来；你们既被记得，就被掳在掌中。
EZEK|21|25|你这亵渎行恶的 以色列 王啊，你的日子，最后惩罚的时刻已来临。
EZEK|21|26|主耶和华如此说：当除掉荣冕，摘下华冠，景况已不复从前；要使卑者升为高，使高者降为卑。
EZEK|21|27|我要将这国倾覆，倾覆，再倾覆；这国必不存在，直等到那应得的人来到，我就将国赐给他。”
EZEK|21|28|“人子啊，你要说预言；你要说，论到 亚扪 人和他们的凌辱，主耶和华吩咐我如此说：有刀，拔出来的刀，已经擦亮，为了行杀戮；它亮如闪电以行吞灭。
EZEK|21|29|他们为你见虚假的异象，行谎诈的占卜，使你倒在亵渎之恶人的颈项上；他们的日子，最后惩罚的时刻已来临。
EZEK|21|30|你收刀入鞘吧！我要在你受造之处、生长之地惩罚你。
EZEK|21|31|我要把我的愤怒倾倒在你身上，把我烈怒的火喷在你身上；又将你交在善于杀灭、畜牲一般的人手中。
EZEK|21|32|你要成为火中之柴，你的血必在地里；你必不再被记得，因为这是我─耶和华说的。”
EZEK|22|1|耶和华的话临到我，说：
EZEK|22|2|“你，人子啊，你要审问，审问这流人血的城吗？要使它知道它一切可憎的事。
EZEK|22|3|你要说，主耶和华如此说：那在其中流人血的城啊，它的时刻已到，它制造偶像玷污了自己。
EZEK|22|4|你因流了人的血，算为有罪；因所制造的偶像，玷污自己；你使你的日子临近，你的年数已来到 。所以我使你承受列国的凌辱和列邦的讥诮。
EZEK|22|5|你这恶名昭彰、混乱的城啊，离你或远或近的国家都必讥诮你。
EZEK|22|6|“看哪， 以色列 的领袖在你那里，为了流人的血各逞其能。
EZEK|22|7|你那里有轻慢父母的，在你当中有欺压寄居者的，你那里也有亏负孤儿寡妇的。
EZEK|22|8|你藐视我的圣物，干犯我的安息日。
EZEK|22|9|你那里有为流人血而毁谤人的，你那里有在山上吃祭物的，在你当中也有行淫乱的，
EZEK|22|10|有露父亲下体的 ，有玷辱经期中不洁净之妇人的。
EZEK|22|11|这人与邻舍的妻子行可憎的事，那人行淫污辱媳妇，在你那里还有人污辱他的姊妹，父亲的女儿。
EZEK|22|12|你那里有收取报酬而流人血的。你取利息，又索取高利；欺压邻舍，夺取财物；你竟然忘了我。这是主耶和华说的。
EZEK|22|13|“看哪，我因你所得不义之财和你们中间所流的血，就击打手掌。
EZEK|22|14|到了我对付你的日子，你的心岂能忍受呢？你的手还能有力吗？我─耶和华说了这话，就必成就。
EZEK|22|15|我要把你驱散到列国，分散在列邦。我也必除掉你们中间的污秽。
EZEK|22|16|你在列国眼前因自己所做的被侮辱 ，你就知道我是耶和华。”
EZEK|22|17|耶和华的话临到我，说：
EZEK|22|18|“人子啊，我看 以色列 家为渣滓。他们是炉中的铜、锡、铁、铅，是炼银的渣滓 。
EZEK|22|19|所以主耶和华如此说：因你们全都成为渣滓，所以，看哪，我必将你们聚集在 耶路撒冷 中。
EZEK|22|20|人怎样把银、铜、铁、铅、锡聚在炉中，吹火使它镕化；照样，我也要在我的怒气和愤怒中聚集你们，把你们安置在城中，使你们镕化。
EZEK|22|21|我必聚集你们，把我烈怒的火吹在你们身上，你们就在其中镕化。
EZEK|22|22|银子怎样在炉中镕化，你们也必照样在城中镕化，因此就知道是我─耶和华把愤怒倾倒在你们身上。”
EZEK|22|23|耶和华的话临到我，说：
EZEK|22|24|“人子啊，你要向这地说：你是未被洁净 之地，在我盛怒的日子，没有雨水在其上。
EZEK|22|25|其中的先知同谋背叛 ，如咆哮的狮子抓撕掠物。他们吞灭人命，抢夺财宝，使这地寡妇增多。
EZEK|22|26|其中的祭司曲解我的律法，亵渎我的圣物，不分别圣与俗，也不使人分辨洁净和不洁净，又遮眼不顾我的安息日；在他们中间连我也被亵慢了。
EZEK|22|27|其中的领袖仿佛野狼抓撕掠物，流人的血，伤害人命，为得不义之财。
EZEK|22|28|其中的先知为他们粉刷，见虚假的异象，行谎诈的占卜，说：‘主耶和华如此说’，其实耶和华并没有说。
EZEK|22|29|这地的百姓惯行欺压抢夺之事，亏负困苦和贫穷的人，欺压寄居者，没有公平。
EZEK|22|30|我在他们中间寻找一人重修城墙，在我面前为这地站在缺口上，使我不致灭绝它，却连一个也找不着。
EZEK|22|31|所以我把愤怒倾倒在他们身上，用烈怒之火消灭他们，照他们所做的报应在他们头上。这是主耶和华说的。”
EZEK|23|1|耶和华的话临到我，说：
EZEK|23|2|“人子啊，有两个女子，是一母所生，
EZEK|23|3|她们在 埃及 行淫，年少时就开始行淫；在那里任人拥抱胸怀，抚弄她们少女的乳房。
EZEK|23|4|她们的名字，大的叫 阿荷拉 ，妹妹叫 阿荷利巴 。她们都归于我，生了儿女。论到她们的名字， 阿荷拉 是 撒玛利亚 ， 阿荷利巴 是 耶路撒冷 。
EZEK|23|5|“ 阿荷拉 归我之后却仍行淫，恋慕所爱的人，就是 亚述 人，都是战士 ，
EZEK|23|6|穿着蓝衣，作省长、副省长，全都是俊美的年轻人，骑着马的骑士。
EZEK|23|7|阿荷拉 与 亚述 人中所有的美男子放纵淫行，她因拜所恋慕之人的一切偶像，玷污了自己。
EZEK|23|8|她从 埃及 的时候，就没有离开过淫乱；因为她年轻时，有人与她同寝，抚弄她少女的乳房，和她纵欲行淫。
EZEK|23|9|因此，我把她交在她所爱的人手中，就是她所恋慕的 亚述 人手中。
EZEK|23|10|他们暴露她的下体，掳掠她的儿女，用刀杀了她；他们向她施行审判，使她在妇女中留下臭名。
EZEK|23|11|“她妹妹 阿荷利巴 虽然看见了，却还是纵欲，比姊姊更加腐败，行淫乱比姊姊更甚。
EZEK|23|12|她恋慕 亚述 人，就是省长和副省长，披挂整齐的战士，骑着马的骑士，全都是俊美的年轻人。
EZEK|23|13|我看见她被污辱，姊妹二人同行一路。
EZEK|23|14|阿荷利巴 又加增淫行，她看见墙上刻有人像，就是鲜红色的 迦勒底 人雕刻的像。
EZEK|23|15|它们腰间系着带子，头上有飘扬的裹头巾，都是将军的样子， 巴比伦 人的形像； 迦勒底 是他们的出生地。
EZEK|23|16|阿荷利巴 一看见就恋慕他们，派遣使者往 迦勒底 他们那里去。
EZEK|23|17|巴比伦 人来到她那里，上了她爱情的床，与她行淫污辱她。她被污辱，随后她的心却与他们生疏。
EZEK|23|18|这样，她既暴露淫行，暴露下体；我的心就与她生疏，像先前与她的姊姊生疏一样。
EZEK|23|19|她仍继续增添淫行，追念她年轻时在 埃及 地行淫的日子，
EZEK|23|20|恋慕情人的身壮精足，如驴似马。
EZEK|23|21|这样，你就渴望年轻时的淫荡；那时， 埃及 人因你年轻时的胸怀，抚弄你的乳房 。”
EZEK|23|22|阿荷利巴 啊，主耶和华如此说：“看哪，我要激起先前你喜爱，而后生疏的人前来攻击你。我必使他们前来，在你四围攻击你；
EZEK|23|23|有 巴比伦 人、 迦勒底 众人、 比割 人、 书亚 人、 哥亚 人，还有 亚述 众人与他们一起，都是俊美的年轻人。他们是省长、副省长、将军、有名声的，全都骑着马。
EZEK|23|24|他们用兵器、 战车、辎重车，率领大军前来攻击你。他们要拿大小盾牌，戴着头盔，在你四围摆阵攻击你。我要把审判交给他们，他们必按着自己的规条审判你。
EZEK|23|25|我要向你倾泄我的妒忌，使他们以愤怒对待你。他们必割去你的鼻子和耳朵，你剩余的人必倒在刀下。他们必掳去你的儿女，你所剩余的必被火焚烧。
EZEK|23|26|他们必剥去你的衣服，夺取你美丽的宝物。
EZEK|23|27|这样，我必止息你的淫行和你从 埃及 地就开始犯的淫乱，使你不再仰望 亚述 ，也不再追念 埃及 。
EZEK|23|28|主耶和华如此说：看哪，我必把你交在你所恨恶的人手中，就是你心与他生疏的人手中。
EZEK|23|29|他们要以恨恶对待你，夺取你劳碌得来的一切，留下你赤身露体。你淫乱的下体，连你的淫行和淫荡，都必显露。
EZEK|23|30|人必向你行这些事；因为你随从外邦人行淫，用他们的偶像玷污自己。
EZEK|23|31|你走了你姊姊的路，所以我必把她的杯交在你的手中。”
EZEK|23|32|主耶和华如此说： “你必喝你姊姊的杯， 那杯又深又广， 盛得很多， 使你遭受嗤笑讥刺。
EZEK|23|33|你必酩酊大醉， 满有愁苦。 你姊姊 撒玛利亚 的杯， 惊骇和凄凉的杯，
EZEK|23|34|你必喝它，并且喝干。 甚至咀嚼杯片， 撕裂自己的胸脯； 因为我曾说过。 这是主耶和华说的。”
EZEK|23|35|主耶和华如此说：“因你忘记我，将我丢在背后，所以你要担当你的淫行和淫荡。”
EZEK|23|36|耶和华对我说：“人子啊，你要审问 阿荷拉 与 阿荷利巴 吗？要指出她们所做可憎的事。
EZEK|23|37|她们行奸淫，手中有血。她们与偶像行奸淫，使她们为我所生的儿女经火，给它们当食物。
EZEK|23|38|此外，她们还向我这样做：同一天又玷污我的圣所，干犯我的安息日。
EZEK|23|39|她们杀了儿女献给偶像，当天又进入我的圣所，亵渎了它。看哪，这就是她们在我殿中所做的。
EZEK|23|40|“况且你们两姊妹派人从远方召人来。使者到了他们那里，看哪，他们就来了。为了他们，你们沐浴，画眼影，佩戴首饰，
EZEK|23|41|坐在华美的床上，前面摆设桌子，把我的香料和膏油放在其上。
EZEK|23|42|在那里有一群人欢乐的声音；有许多的平民，从旷野来的醉汉 ，把镯子戴在她们手上，把华冠戴在她们头上。
EZEK|23|43|“我论到这久行奸淫而色衰的妇人说：现在人们还要与她行淫，她也要与人行淫。
EZEK|23|44|人去到 阿荷拉 和 阿荷利巴 二淫妇那里 ，好像与妓女行淫。
EZEK|23|45|义人必按照审判淫妇和流人血之妇人的规条，审判她们；因为她们是淫妇，她们的手中有血。”
EZEK|23|46|主耶和华如此说：“我要让军队上来攻击她们，使她们惊骇，成为掳物。
EZEK|23|47|这军队必用石头打死她们，用刀剑杀害她们，又杀戮她们的儿女，用火焚烧她们的房屋。
EZEK|23|48|我必使这地不再有淫行，所有的妇女都受警戒，不再效法你们的淫行 。
EZEK|23|49|人必因你们的淫行报应你们；你们要担当拜偶像的罪，因此你们就知道我是主耶和华。”
EZEK|24|1|第九年十月初十，耶和华的话临到我，说：
EZEK|24|2|“人子啊，你要记录这一天的名称，这特别的一天， 巴比伦 王围困 耶路撒冷 ，就在这特别的一天。
EZEK|24|3|你要向这悖逆之家设比喻，对他们说，主耶和华如此说： 把锅放在火上， 放好了，倒水在其中；
EZEK|24|4|要将肉块，一切肥美的肉块， 腿和肩都放在锅里， 要装满上等的骨头；
EZEK|24|5|要取羊群中最好的， 把柴 堆在下面， 把它煮开， 骨头煮在其中。
EZEK|24|6|“主耶和华如此说：祸哉！这流人血的城，就是长锈的锅。它的锈未曾除掉，要将肉块从其中一一取出，不必抽签。
EZEK|24|7|这城所流的血还在城中，血倒在光滑的磐石上，没有倒在地上，用土掩盖；
EZEK|24|8|是我使这城所流的血倒在光滑的磐石上，不得掩盖，为要惹动愤怒，施行报应。
EZEK|24|9|所以主耶和华如此说：祸哉！这流人血的城，我必亲自加大柴堆。
EZEK|24|10|你要添上木柴，使火着旺，将肉煮烂，加上香料 ，烤焦骨头；
EZEK|24|11|你要把空锅放在炭火上，将锅烧热，把铜烧红，镕化其中的污秽，除净其上的锈。
EZEK|24|12|然而这一切劳碌无效 ，它厚厚的锈，即使用火也除不掉。
EZEK|24|13|虽然我想洁净你污秽的淫行，你却不洁净，你的污秽再也不能洁净，直等我止息了向你发的愤怒。
EZEK|24|14|我─耶和华说了这话，时候到了，就必成就；必不退缩，不顾惜，也不怜悯。人必照你的所作所为审判你。这是主耶和华说的。”
EZEK|24|15|耶和华的话临到我，说：
EZEK|24|16|“人子，看哪，我要以灾病夺取你眼中所喜爱的，你却不可悲哀哭泣，也不可流泪，
EZEK|24|17|只可叹息，不可出声，不可办理丧事；裹上头巾，脚上穿鞋，不可捂着胡须，也不可吃一般人的食物 。”
EZEK|24|18|到了早晨我把这事告诉百姓，晚上我的妻子就死了。次日早晨我就遵命而行。
EZEK|24|19|百姓对我说：“你这样做跟我们有什么关系，你不告诉我们吗？”
EZEK|24|20|我对他们说：“耶和华的话临到我，说：
EZEK|24|21|‘你告诉 以色列 家，主耶和华如此说：我要使我的圣所被亵渎，就是你们凭势力所夸耀、眼里所喜爱、心中所爱惜的；并且你们所遗留的儿女必倒在刀下。
EZEK|24|22|那时，你们要照我所做的去做。你们不可捂着胡须，也不可吃一般人的食物。
EZEK|24|23|你们头要裹上头巾，脚要穿上鞋；不可悲哀哭泣。你们必因自己的罪孽衰残，相对叹息。
EZEK|24|24|以西结 必这样成为你们的预兆；凡他所做的，你们也必照样做。那事来到，你们就知道我是主耶和华。’”
EZEK|24|25|“你，人子啊，那日当我除掉他们所倚靠的保障、所欢喜的荣耀，并眼中所喜爱的，心里所重看的儿女时，
EZEK|24|26|逃脱的人岂不来到你这里，使你耳闻这事吗？
EZEK|24|27|那日你要向逃脱的人开口说话，不再哑口无言。你必这样成为他们的预兆，他们就知道我是耶和华。”
EZEK|25|1|耶和华的话临到我，说：
EZEK|25|2|“人子啊，你要面向 亚扪 人说预言，攻击他们。
EZEK|25|3|你要对 亚扪 人说，当听主耶和华的话。主耶和华如此说：我的圣所遭亵渎， 以色列 地变荒凉， 犹大 家被掳掠；那时，你因这些事说‘啊哈’，
EZEK|25|4|所以，看哪，我要把你交给东方人为业；他们必在你中间安营居住，设立居所，吃你的果子，喝你的奶。
EZEK|25|5|我必使 拉巴 成为牧放骆驼之地，使 亚扪 成为羊群躺卧之处，你们就知道我是耶和华。
EZEK|25|6|主耶和华如此说：因你们拍手顿足，幸灾乐祸，藐视 以色列 地，
EZEK|25|7|所以，看哪，我要伸手攻击你，把你交给列国作为掳物。我必从万民中剪除你，从列邦中消灭你。我必除灭你，你就知道我是耶和华。”
EZEK|25|8|“主耶和华如此说：因 摩押 和 西珥 人说‘看哪， 犹大 家与列国无异’，
EZEK|25|9|所以，看哪，我要破开 摩押 边界的城镇，就是 摩押 人所夸耀的城镇， 伯．耶施末 、 巴力．免 、 基列亭 ，
EZEK|25|10|令东方人前来攻击 亚扪 人。我必将 亚扪 交给他们为业，使 亚扪 人在列国中不再被记念。
EZEK|25|11|我也必向 摩押 施行审判，他们就知道我是耶和华。”
EZEK|25|12|“主耶和华如此说：因为 以东 向 犹大 家报仇，因向他们报仇而大大显为有罪，
EZEK|25|13|所以主耶和华如此说：我要伸手攻击 以东 ，将人与牲畜剪除，使 以东 从 提幔 起，直到 底但 ，地变荒凉，人也都倒在刀下。
EZEK|25|14|我要藉我子民 以色列 的手报复 以东 ；他们必照我的怒气，按我的愤怒对待 以东 ， 以东 人就知道施报的是我。这是主耶和华说的。”
EZEK|25|15|“主耶和华如此说：因 非利士 人报仇，就是心存轻蔑报仇；他们永怀仇恨，意图毁灭，
EZEK|25|16|所以主耶和华如此说：看哪，我要伸手攻击 非利士 人，剪除 基利提 人，灭绝沿海剩余的居民。
EZEK|25|17|我要大大报复他们，发怒斥责他们。我报复他们的时候，他们就知道我是耶和华。”
EZEK|26|1|第十一年某月初一，耶和华的话临到我，说：
EZEK|26|2|“人子啊，因 推罗 向 耶路撒冷 说：‘啊哈！那众民之门已经破坏，向我敞开；它既变为废墟，我必丰盛。’
EZEK|26|3|所以，主耶和华如此说： 推罗 ，看哪，我与你为敌，使许多国家涌上攻击你，如同海洋使波浪涌上一样。
EZEK|26|4|他们要破坏 推罗 的城墙，拆毁它的城楼。我也要刮净它的尘土，使它成为光滑的磐石。
EZEK|26|5|推罗 必成为海中的晒网场，因为我曾说过， 这是主耶和华说的。它必成为列国的掳物，
EZEK|26|6|推罗 乡间邻近的城镇 必遭刀剑灭绝，他们就知道我是耶和华。”
EZEK|26|7|主耶和华如此说：“看哪，我必使诸王之王，就是 巴比伦 王 尼布甲尼撒 ，率领马匹、战车、骑兵、军队和许多人从北方来攻击 推罗 。
EZEK|26|8|他必用刀剑杀灭你乡间邻近的城镇，也必筑堡垒，建土堆，举盾牌攻击你。
EZEK|26|9|他要安设撞城槌攻破你的城墙，以刀剑拆毁你的城楼。
EZEK|26|10|因他马匹众多，尘土必扬起遮蔽你。他进入你的城门，如同进入已有缺口之城。那时，你的城墙必因骑兵、车轮和战车的响声震动。
EZEK|26|11|他的马蹄必践踏你所有的街道；他必用刀剑杀戮你的居民。你坚固的柱子 必倒在地上。
EZEK|26|12|人必掳获你的财宝，掠夺你的货财；他们要破坏你的城墙，拆毁你华美的房屋，将你的石头、木头、尘土都抛在水中。
EZEK|26|13|我要使你唱歌的声音止息；人不再听见你弹琴的声音。
EZEK|26|14|我必使你成为光滑的磐石，作晒网的场所。你不得再被建造，因为我─耶和华已这样说了。这是主耶和华说的。”
EZEK|26|15|主耶和华对 推罗 如此说：“在你中间行杀戮，受伤的人唉哼时，海岛岂不都因你倾倒的响声震动吗？
EZEK|26|16|那时沿海的君王都要从宝座下来，除去朝服，脱下锦衣，披上战兢，坐在地上，不停发抖，为你而惊骇。
EZEK|26|17|他们必为你作哀歌，向你说： ‘你这闻名之城， 航海之人居住， 海上最为坚固的， 你和居民使所有住在沿海的人 无不惊恐， 现在竟然毁灭了！
EZEK|26|18|如今在你倾覆的日子， 海岛都要战兢； 海中的群岛见你归于无有 就都惊惶。’”
EZEK|26|19|主耶和华如此说：“ 推罗 啊 ，我要使你变为荒凉，如无人居住的城镇；又使深水漫过你，大水淹没你。
EZEK|26|20|那时，我要使你和下到地府的人同去，到古时候的人那里；我要使你和下到地府的人一同住在地的深处，在久已荒废的地方，使你那里不再有人居住；我要在活人之地显荣耀 。
EZEK|26|21|我必叫你令人惊恐，使你不再存留于世；人虽寻找你，却永不寻见。这是主耶和华说的。”
EZEK|27|1|耶和华的话临到我，说：
EZEK|27|2|“人子啊，要为 推罗 作哀歌。
EZEK|27|3|你要对位于海口，跟许多海岛的百姓做生意的 推罗 说，主耶和华如此说： 推罗 啊，你曾说： ‘我全然美丽。’
EZEK|27|4|你的疆界在海的中心， 造你的使你全然美丽。
EZEK|27|5|他们用 示尼珥 的松树作你的甲板， 用 黎巴嫩 的香柏树作桅杆，
EZEK|27|6|用 巴珊 的橡树作你的桨， 用镶嵌象牙的 基提 海岛黄杨木 为舱板。
EZEK|27|7|你的帆是用 埃及 绣花细麻布做的， 可作你的大旗； 你的篷是用 以利沙岛 的蓝色和紫色布做的。
EZEK|27|8|西顿 和 亚发 的居民为你划桨； 推罗 啊，你们中间的智慧人为你掌舵。
EZEK|27|9|迦巴勒 的长者和智者 在你中间修补裂缝； 海上一切的船只和水手 都在你那里进行货物交易。
EZEK|27|10|“ 波斯 人、 路德 人、 弗 人在你的军营中作战士；他们在你们中间悬挂盾牌和头盔，彰显你的尊荣。
EZEK|27|11|亚发 人和你的军队都驻守在四围的城墙上，你的城楼上也有勇士；他们悬挂盾牌，成全你的美丽。
EZEK|27|12|“ 他施 因你多有财物，就作你的客商，他们带着银、铁、锡、铅前来换你的商品。
EZEK|27|13|雅完 、 土巴 、 米设 都与你交易，以人口和铜器换你的货物。
EZEK|27|14|陀迦玛 族用马匹、战马和骡子换你的商品。
EZEK|27|15|底但 人与你交易，许多海岛成为你的码头；他们拿象牙、黑檀木与你交换。
EZEK|27|16|亚兰 因你货品充裕，就作你的客商；他们用绿宝石、紫色布、刺绣、细麻布、珊瑚、红宝石换你的商品。
EZEK|27|17|犹大 和 以色列 地都与你交易；他们用 米匿 的小麦、饼、蜜、油、乳香换你的货物。
EZEK|27|18|大马士革 也因你货品充裕，多有各类财物，就带来 黑本 酒和白羊毛与你交易。
EZEK|27|19|威但 和从 乌萨 来的 雅完 人 为了你的货物，以加工的铁、桂皮、香菖蒲换你的商品。
EZEK|27|20|底但 以骑马用的座垫毯子与你交换。
EZEK|27|21|阿拉伯 和 基达 所有的领袖都作你的客商，用羔羊、公绵羊、公山羊与你交换。
EZEK|27|22|示巴 和 拉玛 的商人也来与你交易，他们用各类上好的香料、各类的宝石和黄金换你的商品。
EZEK|27|23|哈兰 、 干尼 、 伊甸 、 示巴 商人、 亚述 和 基抹 都与你交易。
EZEK|27|24|这些商人将美好的货物包在蓝色的绣花包袱内，又将华丽的衣服装在香柏木的箱子里，用绳索捆着，以此与你交易 。
EZEK|27|25|他施 的船只为你运货， 你在海中满载货物，极其沉重。
EZEK|27|26|划桨的把你划到水深之处， 东风在海中将你击破。
EZEK|27|27|你的财宝、商品、货物、 水手、掌舵的、 修补船缝的、进行货物交易的， 并你那里所有的战士 和你中间所有的军队， 在你倾覆的日子都必沉在海底。
EZEK|27|28|因掌舵者的呼声， 郊野就必震动。
EZEK|27|29|所有划桨的 都从他们的船下来； 水手和所有在海上掌舵的， 都要登岸。
EZEK|27|30|他们必为你放声痛哭， 撒尘土于头上， 在灰中打滚；
EZEK|27|31|又为你使头光秃， 用麻布束腰， 号啕痛哭， 痛苦至极。
EZEK|27|32|他们哀号的时候， 为你作哀歌， 为你痛哭： 有何城如 推罗 ， 在海中沉寂呢？
EZEK|27|33|你由海上运出商品， 使许多民族充裕； 你以许多财宝货物 令地上的君王丰富。
EZEK|27|34|在深水中被海浪打破的时候， 你的货物和你中间所有的军队都下沉。
EZEK|27|35|海岛所有的居民为你惊奇， 他们的君王都甚恐慌，面带愁容。
EZEK|27|36|万民中的商人向你发嘘声； 你令人惊恐， 不再存留于世，直到永远。”
EZEK|28|1|耶和华的话临到我，说：
EZEK|28|2|“人子啊，你要对 推罗 的君王说，主耶和华如此说： 你心里高傲，说：‘我是神明； 我在海中坐诸神之位。’ 虽然你把你的心比作神明的心， 你却不过是人，并不是神明！
EZEK|28|3|看哪，你比 但以理 更有智慧， 任何秘密都不能向你隐藏。
EZEK|28|4|你靠自己的智慧聪明得了财宝， 把金银收入库房；
EZEK|28|5|你靠自己的大智慧以贸易增添财宝， 又因你的财宝心里高傲；
EZEK|28|6|所以主耶和华如此说： 因你把你的心比作神明的心，
EZEK|28|7|所以，看哪，我必使外国人， 就是列国中凶暴的人临到你这里； 他们要拔刀摧毁你用智慧得来的美物， 污损你的荣光。
EZEK|28|8|他们必使你坠入地府； 你要像被刺杀之人的死，死在海中。
EZEK|28|9|在杀你的人面前， 你还能说‘我是神明’吗？ 在杀害你的人手中， 你不过是人，并不是神明。
EZEK|28|10|你要死在陌生人手中， 像未受割礼之人的死， 因为我曾说过， 这是主耶和华说的。”
EZEK|28|11|耶和华的话临到我，说：
EZEK|28|12|“人子啊，要为 推罗 王作哀歌，对他说，主耶和华如此说： 你曾是完美的典范， 智慧充足，全然美丽。
EZEK|28|13|你在 伊甸 ─上帝的园中， 佩戴各样宝石， 就是红宝石、红璧玺、金刚石、 水苍玉、红玛瑙、碧玉、 蓝宝石、绿宝石、红玉； 你的宝石有黄金的底座，手工精巧 ， 都是在你受造之日预备的。
EZEK|28|14|我指定你为受膏的基路伯， 看守保护； 你在上帝的圣山上； 往来在如火的宝石中。
EZEK|28|15|你从受造之日起行为正直， 直到后来查出你的不义。
EZEK|28|16|你因贸易发达， 暴力充斥其中，以致犯罪， 所以我污辱你，使你离开上帝的山。 守护者基路伯啊， 我已将你从如火的宝石中歼灭。
EZEK|28|17|你因美丽心中高傲， 因荣光而败坏智慧， 我已将你抛弃在地， 把你摆在君王面前， 好叫他们目睹眼见。
EZEK|28|18|你因罪孽众多，贸易不公， 亵渎了你的圣所； 因此我使火从你中间发出， 烧灭了你， 使你在所有观看的人眼前 变为地上的灰烬。
EZEK|28|19|万民中凡认识你的 都必为你惊奇。 你令人惊恐， 不再存留于世，直到永远。”
EZEK|28|20|耶和华的话临到我，说：
EZEK|28|21|“人子啊，你要面向 西顿 ，向它说预言。
EZEK|28|22|你要说，主耶和华如此说： ‘ 西顿 ，看哪，我与你为敌， 我要在你中间得荣耀。’ 我在它中间施行审判、显为圣的时候， 人就知道我是耶和华。
EZEK|28|23|我必令瘟疫进入 西顿 ， 使血流在街上。 刀剑从四围临到它， 被杀的要仆倒在其中； 人就知道我是耶和华。”
EZEK|28|24|“四围恨恶 以色列 家的人，对他们必不再如刺人的荆棘、伤人的蒺藜；他们就知道我是主耶和华。”
EZEK|28|25|主耶和华如此说：“我将分散在万民中的 以色列 家召集回来，在列国眼前向他们显为圣的时候，他们仍可在我所赐给我仆人 雅各 之地居住。
EZEK|28|26|他们要在这地上安然居住。我向四围恨恶他们的众人施行审判之后，他们要建造房屋，栽葡萄园，安然居住，他们就知道我是耶和华─他们的上帝。”
EZEK|29|1|第十年十月十二日，耶和华的话临到我，说：
EZEK|29|2|“人子啊，你要面向 埃及 王法老，向他和 埃及 全地说预言。
EZEK|29|3|你要说，主耶和华如此说： 埃及 王法老， 你这卧在自己江河中的海怪， 看哪，我与你为敌。 你曾说：‘我的 尼罗河 是我的， 是我为自己造的。’
EZEK|29|4|我必用钩子钩住你的腮颊， 令江河中的鱼贴住你的鳞甲； 我要把你和所有贴着鳞甲的鱼 从你的江河中拉上来。
EZEK|29|5|我要把你和江河中的鱼全都抛弃在旷野； 你必仆倒在田间， 无人收殓，无人掩埋。 我已将你给了地上的走兽、空中的飞鸟作食物。
EZEK|29|6|“ 埃及 所有的居民必定知道我是耶和华。因为你已成为 以色列 家芦苇的杖；
EZEK|29|7|他们用手掌一握，你就断裂，伤了他们的肩；他们靠着你，你却折断，闪了他们的腰 。
EZEK|29|8|所以主耶和华如此说：我必使刀剑临到你，把人与牲畜从你中间剪除。
EZEK|29|9|埃及 地必荒芜废弃，他们就知道我是耶和华。 “因为法老说‘ 尼罗河 是我的，是我所造的’，
EZEK|29|10|所以，看哪，我必与你和你的江河为敌，使 埃及 地，从 密夺 到 色弗尼 ，直到 古实 边界，全然废弃荒芜。
EZEK|29|11|人的脚不经过，兽的蹄也不经过，四十年之久无人居住。
EZEK|29|12|我要使 埃及 地成为荒芜中最荒芜的地，使它的城镇变为荒废中最荒废的城镇，共四十年之久。我必将 埃及 人分散到列国，四散在列邦。
EZEK|29|13|“主耶和华如此说：满了四十年后，我必招聚分散在万民中的 埃及 人。
EZEK|29|14|我要令 埃及 被掳的人归回，使他们回到本地 巴特罗 。在那里，他们必成为弱小的国家，
EZEK|29|15|成为列国中最低微的，不再自高于列邦之上。我必使他们变为小国，不再辖制列邦。
EZEK|29|16|埃及 必不再作 以色列 家的倚靠，却使 以色列 家想起他们仰赖 埃及 的罪。他们就知道我是主耶和华。”
EZEK|29|17|第二十七年正月初一，耶和华的话临到我，说：
EZEK|29|18|“人子啊， 巴比伦 王 尼布甲尼撒 令他的军兵大力攻打 推罗 ，以致头都光秃，肩都磨破；然而他和军兵虽然为攻打 推罗 花这么多力气，却没有从那里得到什么犒赏。
EZEK|29|19|所以主耶和华如此说：我要将 埃及 地赐给 巴比伦 王 尼布甲尼撒 ；他必掳掠 埃及 的财富，抢夺它的掳物，掳掠它的掠物，用以犒赏他的军兵。
EZEK|29|20|我将 埃及 地赐给他，犒赏他，因他们为我效劳。这是主耶和华说的。
EZEK|29|21|“当那日，我必使 以色列 家壮大 ，又必使你─ 以西结 在他们中间开口；他们就知道我是耶和华。”
EZEK|30|1|耶和华的话临到我，说：
EZEK|30|2|“人子啊，你要说预言；你要说，主耶和华如此说： 哀哉这日！你们应当哭号，
EZEK|30|3|因为日子近了， 耶和华的日子临近了； 那是密云之日， 是列国受罚 之期。
EZEK|30|4|必有刀剑临到 埃及 ； 被杀的人仆倒在 埃及 时， 古实 人颤惊不已。 埃及 的财富遭掳掠， 根基被拆毁。
EZEK|30|5|古实 人、 弗 人、 路德 人、混居的各族和 古伯 人，以及盟国的人都要与 埃及 人一同倒在刀下。”
EZEK|30|6|耶和华如此说： 扶助 埃及 的必倾倒， 埃及 骄傲的权势必降为卑， 从 密夺 到 色弗尼 ，人必倒在刀下。 这是主耶和华说的。
EZEK|30|7|埃及 成为荒凉中最荒凉的国， 它的城镇变为荒废中最荒废的城镇。
EZEK|30|8|我在 埃及 放火， 帮助 埃及 的，都遭灭绝； 那时，他们就知道我是耶和华。
EZEK|30|9|“到那日，必有使者从我面前乘船出去，使安逸无虑的 古实 人惊惧；当 埃及 遭难的日子，痛苦也必临到他们。看哪，这事临近了！
EZEK|30|10|主耶和华如此说： 我要藉 巴比伦 王 尼布甲尼撒 的手 除灭 埃及 的军队。
EZEK|30|11|他和随从他的人， 就是列国中凶暴的人， 要前来毁灭这地， 拔刀攻击 埃及 ， 使遍地布满被杀的人。
EZEK|30|12|我要使江河干涸， 将这地卖在恶人手中； 我要藉外国人的手， 使这地和其中所充满的变为荒芜； 这是我─耶和华说的。
EZEK|30|13|“主耶和华如此说： 我要毁灭偶像， 从 挪弗 除掉神像； 不再有君王出自 埃及 地， 我要使 埃及 地的人惧怕。
EZEK|30|14|我必令 巴特罗 荒凉， 在 琐安 放火， 向 挪 施行审判。
EZEK|30|15|我要将我的愤怒倾倒在 训 ， 埃及 的堡垒上， 要剪除 挪 的众民。
EZEK|30|16|我必在 埃及 放火， 训 必大大痛苦， 挪 被攻破， 挪弗 终日遭敌侵袭。
EZEK|30|17|亚文 和 比．伯实 的年轻人必倒在刀下， 这些城镇将被掳掠。
EZEK|30|18|我在 答比匿 折断 埃及 的轭 ， 使它骄傲的权势止息。 那时，日光必退去； 至于这城，必有密云遮蔽， 邻近的城镇 也遭掳掠。
EZEK|30|19|我要如此向 埃及 施行审判， 他们就知道我是耶和华。”
EZEK|30|20|第十一年正月初七，耶和华的话临到我，说：
EZEK|30|21|“人子啊，我已折断 埃及 王法老的一只膀臂；看哪，无人为他敷药，也无人为他包扎绷带，使他有力持刀。
EZEK|30|22|因此，主耶和华如此说：看哪，我与 埃及 王法老为敌，要折断他的膀臂，折断强壮的和已受伤的，使刀从他手中掉落。
EZEK|30|23|我必将 埃及 人分散到列国，四散在列邦。
EZEK|30|24|我要使 巴比伦 王的膀臂有力，把我的刀交在他手中；却要折断法老的膀臂，使他在 巴比伦 王面前呻吟，如同被杀的人一样。
EZEK|30|25|我要使 巴比伦 王的膀臂强壮，法老的膀臂却要下垂；当我把我的刀交在 巴比伦 王手中时，他要举刀攻击 埃及 地，他们就知道我是耶和华。
EZEK|30|26|我必将 埃及 人分散到列国，四散在列邦；他们就知道我是耶和华。”
EZEK|31|1|第十一年三月初一，耶和华的话临到我，说：
EZEK|31|2|“人子啊，你要对 埃及 王法老和他的军队说： 论到你的强盛，谁能与你相比呢？
EZEK|31|3|看哪， 亚述 是 黎巴嫩 的香柏树， 枝条荣美，荫密如林， 极其高大，树顶高耸入云。
EZEK|31|4|众水使它生长， 深水使它长高； 所栽之地有江河环绕， 汊出的水道流至田野的树木。
EZEK|31|5|所以它高大超过田野的树木； 生长时因水源丰沛， 枝子繁多，枝条增长。
EZEK|31|6|空中所有的飞鸟在枝子上搭窝， 野地所有的走兽在枝条下生子， 所有的大国也在它的荫下居住。
EZEK|31|7|它树大枝长，极为荣美， 因它的根在众水之旁。
EZEK|31|8|上帝园中的香柏树不能遮蔽它； 松树不及它的枝子， 枫树不及它的枝条， 上帝园中的树都没有它荣美。
EZEK|31|9|我使它枝条繁多， 极为荣美； 在上帝的园中， 伊甸 所有的树都嫉妒它。”
EZEK|31|10|所以主耶和华如此说：“因它 高大，树顶高耸入云，心高气傲，
EZEK|31|11|我要把它交给 列国中强人的手里，他们必定按它的罪恶惩治它。我已经驱逐它。
EZEK|31|12|外国人，就是列国中凶暴的人，已把它砍断抛弃。它的枝条掉落山间和一切谷中，枝子折断，落在地上一切河道。地上的万民都离开它的遮荫，抛弃了它。
EZEK|31|13|空中的飞鸟都栖身在掉落的树干上，野地的走兽也都躺卧在它的枝条中。
EZEK|31|14|为了要使水边的树木枝干不再长高，树顶也不再高耸入云；那些得水滋润的，不再屹立于其中。因为它们和下到地府的人一起，都被交与死亡，到了地底下。”
EZEK|31|15|主耶和华如此说：“它坠落阴间的那日，我为它遮盖深渊，拦住江河，使众水停流，以表哀悼。我使 黎巴嫩 为它悲哀，田野的树木都因它枯萎。
EZEK|31|16|我把它扔到阴间，与下到地府的人一同坠落。那时，列国听见坠落的响声就震惊； 伊甸 一切的树木，就是 黎巴嫩 中得水滋润、最佳最美的树，在地底下都得了安慰。
EZEK|31|17|这些树也要与它同下阴间，到被刀所杀的人那里；它们曾作它的膀臂 ，在列国中曾居住在它的荫下。
EZEK|31|18|在这样的荣耀与威势中， 伊甸 树木有谁能与你相比呢？然而你要与 伊甸 的树木一同到地底下；在未受割礼的人中，与被刀所杀的人一同躺下。 “法老和他的军队正是如此。这是主耶和华说的。”
EZEK|32|1|第十二年十二月初一，耶和华的话临到我，说：
EZEK|32|2|“人子啊，你要为 埃及 王法老作哀歌，说： 你在列国中，如同少壮狮子， 却像海里的海怪， 冲出江河， 以爪搅动诸水， 使江河浑浊。
EZEK|32|3|主耶和华如此说： 许多民族聚集时， 我要将我的网撒在你身上， 他们要把你拉上来。
EZEK|32|4|我要把你丢在地上， 抛在田野， 使空中的飞鸟落在你身上， 遍地的野兽因你得以饱足。
EZEK|32|5|我要将你的肉丢在山间， 用你巨大的尸首 填满山谷。
EZEK|32|6|我要以你所流的血 浸透大地， 漫过山顶， 溢满河道。
EZEK|32|7|我毁灭你时， 要遮蔽诸天， 使众星昏暗； 我必以密云遮掩太阳， 月亮也不放光。
EZEK|32|8|我要使天上发亮的光体 在你上面变为昏暗， 使你的地也变为黑暗。 这是主耶和华说的。
EZEK|32|9|“我使你在列国，在你所不认识的列邦中灭亡 。那时，我必使许多民族的心因你愁烦。
EZEK|32|10|当我在他们面前举起我的刀，我要使许多民族因你惊恐，他们的君王也必因你极其恐慌。在你仆倒的日子，他们各人为自己的性命时时战兢。
EZEK|32|11|主耶和华如此说： 巴比伦 王的刀必临到你。
EZEK|32|12|我必藉勇士的刀使你的军队仆倒；这些勇士都是列国中凶暴的人。 他们必使 埃及 的骄傲归于无有， 埃及 的军队必被灭绝。
EZEK|32|13|我要除灭众水旁一切的走兽， 人的脚必不再搅浑这水， 兽的蹄也不搅浑这水。
EZEK|32|14|那时，我必使他们的水澄清， 使他们的江河像油缓流。 这是主耶和华说的。
EZEK|32|15|我使 埃及 地荒废， 使这地空无一物， 又击杀其中所有的居民； 那时，他们就知道我是耶和华。
EZEK|32|16|“这是一首为人所吟唱的哀歌；列国的女子要唱这哀歌，她们要为 埃及 和它的军队唱这哀歌。这是主耶和华说的。”
EZEK|32|17|第十二年某月 十五日，耶和华的话临到我，说：
EZEK|32|18|“人子啊，你要为 埃及 的军队哀号，把他们和强盛之国 一同扔到地底下，与那些下到地府的人在一起。
EZEK|32|19|‘你的美丽胜过谁呢？ 坠落吧，与未受割礼的人躺在一起！’
EZEK|32|20|他们要仆倒在被刀所杀的人当中。 埃及 被交给刀剑，人要把它和它的军队拉走。
EZEK|32|21|强壮的勇士要在阴间对 埃及 王和他的盟友说话；他们未受割礼，被刀剑所杀，已经坠落躺下。
EZEK|32|22|“ 亚述 和它的全军在那里，四围都是坟墓；他们全都是被杀倒在刀下的人。
EZEK|32|23|他们的坟墓在地府极深之处，它的众军环绕它的坟墓，他们全都是被杀倒在刀下的人，曾在活人之地使人惊恐。
EZEK|32|24|“ 以拦 在那里，它的全军环绕它的坟墓；他们全都是被杀倒在刀下、未受割礼而到地底下的，曾在活人之地使人惊恐；他们与下到地府的人一同担当羞辱。
EZEK|32|25|人为它和它的军队在被杀的人中设立床榻，四围都是坟墓；他们都是未受割礼被刀所杀的，曾在活人之地使人惊恐；他们与下到地府的人一同担当羞辱。 以拦 已列在被杀的人中。
EZEK|32|26|“ 米设 、 土巴 和他们的全军都在那里，四围都是坟墓；他们都是未受割礼被刀所杀的，曾在活人之地使人惊恐。
EZEK|32|27|他们不得与那未受割礼 仆倒的勇士躺在一起；这些勇士带着兵器下到阴间，头枕着刀剑，骨头带着本身的罪孽，曾在活人之地使人惊恐。
EZEK|32|28|法老啊，你必与未受割礼的人一起毁灭，与被刀所杀的人躺在一起。
EZEK|32|29|“ 以东 在那里，它的君王和所有官长虽然英勇，还是与被刀所杀的人同列；他们必与未受割礼的和下到地府的人躺在一起。
EZEK|32|30|“在那里有北方的众王子和所有的 西顿 人，全都与被杀的人一同下去。他们虽然英勇，使人惊恐，还是蒙羞。他们未受割礼，和被刀所杀的人躺在一起，与下到地府的人一同担当羞辱。
EZEK|32|31|“法老看见他们，就为他的军兵，就是被刀所杀属法老的人和他的全军感到安慰。这是主耶和华说的。
EZEK|32|32|我任凭法老在活人之地使人惊恐，法老和他的军兵必躺在未受割礼和被刀所杀的人中。这是主耶和华说的。”
EZEK|33|1|耶和华的话临到我，说：
EZEK|33|2|“人子啊，你要吩咐本国的百姓，对他们说：我使刀剑临到哪一国，哪一国的百姓从他们中间选立一人，作为守望者。
EZEK|33|3|守望者见刀剑临到那地，若吹角警戒百姓，
EZEK|33|4|有人听见角声却不受警戒，刀剑来除灭了他，这人的血必归到自己头上。
EZEK|33|5|他听见角声，不受警戒，他的血必归到自己身上；他若受警戒，就救了自己的命。
EZEK|33|6|倘若守望者见刀剑临到，却不吹角，以致百姓未受警戒，刀剑来杀了他们中间的一个人，这人虽然因自己的罪孽而死，我却要从守望者的手里讨他的血债。
EZEK|33|7|“人子啊，我照样立你作 以色列 家的守望者；你要听我口中的话，替我警戒他们。
EZEK|33|8|我对恶人说：‘恶人哪，你必要死！’你若不开口警戒恶人，使他离开所行的道，这恶人必因自己的罪孽而死，我却要从你手里讨他的血债。
EZEK|33|9|但是你，你若警戒恶人，叫他离弃所行的道，他仍不转离，他必因自己的罪孽而死，你却救了自己的命。”
EZEK|33|10|“人子啊，你要对 以色列 家说：你们曾这样说：‘我们的过犯罪恶在自己身上，我们必因此消灭，怎能存活呢？’
EZEK|33|11|你要对他们说，主耶和华说：我指着我的永生起誓，我断不喜悦恶人死亡，惟喜悦恶人转离他所行的道而存活。 以色列 家啊，你们回转，回转离开恶道吧！何必死亡呢？
EZEK|33|12|人子啊，你要对本国的百姓说：义人的义，在他犯罪之日不能救他；至于恶人的恶，在他转离恶行之日不会使他倾倒；义人在他犯罪之日不能因自己的义存活。
EZEK|33|13|我对义人说：‘你必存活！’他若倚靠自己的义作恶，所行的义就不被记念；他必因所作的恶死亡。
EZEK|33|14|我对恶人说：‘你必死亡！’他若转离他的罪恶，行公平公义的事；
EZEK|33|15|恶人若归还抵押品，归回所抢夺的东西，遵行生命的律例，不再作恶；他必存活，不致死亡。
EZEK|33|16|他所犯的一切罪必不被记念；他行了公平公义的事，必要存活。
EZEK|33|17|“你本国的百姓说：‘主的道不公平。’其实他们，他们的道才是不公平。
EZEK|33|18|义人转离自己的义作恶，他必因此而死亡。
EZEK|33|19|恶人转离他的恶，行公平公义的事，他必因此而存活。
EZEK|33|20|你们还说：‘主的道不公平。’ 以色列 家啊，我必按你们各人所行的审判你们。”
EZEK|33|21|我们被掳后第十二年的十月初五，有人从 耶路撒冷 逃到我这里，说：“城已被攻破。”
EZEK|33|22|逃来的人到的前一天晚上，耶和华的手按在我身上，开我的口。第二天早晨，等那人来到我这里，我的口就开了，不再说不出话来。
EZEK|33|23|耶和华的话临到我，说：
EZEK|33|24|“人子啊，住在 以色列 荒废之地的人说：‘ 亚伯拉罕 一人能得这地为业，我们人数众多，这地更是给我们为业的。’
EZEK|33|25|所以你要对他们说，主耶和华如此说：你们吃带血的食物，向偶像举目，并且流人的血，你们还能得这地为业吗？
EZEK|33|26|你们倚靠自己的刀剑行可憎的事，人人污辱邻舍的妻，你们还能得这地为业吗？
EZEK|33|27|你要对他们这样说，主耶和华如此说：我指着我的永生起誓，在废墟的，必倒在刀下；在田野的，必交给野兽吞吃；在堡垒和洞中的，必遭瘟疫而死。
EZEK|33|28|我必使这地荒废荒凉，它骄傲的权势也必止息； 以色列 的山都必荒废，无人经过。
EZEK|33|29|我因他们所做一切可憎的事，使地荒废荒凉；那时，他们就知道我是耶和华。”
EZEK|33|30|“你，人子啊，你本国的百姓在城墙旁边、在房屋门口谈论你。弟兄对弟兄彼此说：‘来吧！听听有什么话从耶和华而出。’
EZEK|33|31|他们如同百姓前来，来到你这里，坐在你面前仿佛是我的子民。他们听了你的话，却不实行；因为他们口里说爱，心却追随财利。
EZEK|33|32|看哪，他们看你如同一个唱情歌的人 ，声音优雅、善于奏乐；他们听了你的话，却不实行。
EZEK|33|33|看哪，这话就要应验；应验时，他们就知道在他们中间有了先知。”
EZEK|34|1|耶和华的话临到我，说：
EZEK|34|2|“人子啊，你要向 以色列 的牧人说预言，对他们说，主耶和华如此说：祸哉！ 以色列 的牧人只知牧养自己。牧人岂不当牧养群羊吗？
EZEK|34|3|你们吃肥油 、穿羊毛、宰杀肥羊，却不牧养群羊。
EZEK|34|4|瘦弱的，你们不调养；有病的，你们不医治；受伤的，你们未包扎；被逐的，你们不去领回；失丧的，你们不寻找；却用暴力严严地辖制它们 。
EZEK|34|5|它们因无牧人就分散；既分散，就成为一切野兽的食物。
EZEK|34|6|我的羊流落众山之间和各高冈上，分散在全地，无人去寻，无人去找。
EZEK|34|7|“所以，你们这些牧人要听耶和华的话。
EZEK|34|8|主耶和华说：我指着我的永生起誓，我的羊因无牧人就成为掠物，也作了一切野兽的食物。我的牧人不寻找我的羊；这些牧人只知喂养自己，并不喂养我的羊。
EZEK|34|9|所以你们这些牧人要听耶和华的话。
EZEK|34|10|主耶和华如此说：看哪，我必与牧人为敌，从他们手里讨回我的羊，使他们不再牧放群羊；牧人也不再喂养自己。我必救我的羊脱离他们的口，不再作他们的食物。”
EZEK|34|11|“主耶和华如此说：‘看哪，我必亲自寻找我的羊，将它们寻见。
EZEK|34|12|牧人在羊群四散的日子怎样寻找他的羊，我必照样寻找我的羊。这些羊在密云黑暗的日子散在各处，我要从那里救回它们。
EZEK|34|13|我要从万民中领出它们，从各国聚集它们，引领它们归回故土。我要在 以色列 山上，在一切溪水旁边，在境内所有可居住的地牧养它们。
EZEK|34|14|我要在肥美的草场牧养它们。它们的圈必在 以色列 高处的山上，它们必躺卧在佳美的圈内，在 以色列 山肥美的草场上吃草。
EZEK|34|15|我要亲自牧养我的群羊，使它们得以躺卧。这是主耶和华说的。
EZEK|34|16|失丧的，我必寻找；被逐的，我必领回；受伤的，我必包扎；有病的，我必医治；只是肥的壮的，我要除灭 ；我必秉公牧养它们。’
EZEK|34|17|“我的羊群哪，论到你们，主耶和华如此说：看哪，我要在羊与羊中间、公绵羊与公山羊中间施行审判。
EZEK|34|18|你们在肥美的草场上吃草还以为是小事吗？竟用你们的脚践踏剩下的草；你们喝了清水，竟用你们的脚搅浑剩下的水。
EZEK|34|19|至于我的羊，只能吃你们所践踏的，喝你们所搅浑的。
EZEK|34|20|“所以，主耶和华对它们如此说：看哪，我要亲自在肥羊和瘦羊中间施行审判。
EZEK|34|21|因为你们用侧边用肩推挤一切瘦弱的羊，又用角抵撞，使它们四散在外；
EZEK|34|22|所以，我要拯救我的群羊，它们必不再作掠物；我也要在羊和羊中间施行审判。
EZEK|34|23|我必在他们之上立一牧人 ，就是我的仆人 大卫 ，牧养它们；他必牧养他们，作他们的牧人。
EZEK|34|24|我─耶和华必作他们的上帝，我的仆人 大卫 要在他们中间作王。这是我─耶和华说的。
EZEK|34|25|“我要与他们立平安的约，使恶兽从境内断绝；他们在旷野也能安然居住，在树林也能躺卧。
EZEK|34|26|我要使他们和我山冈的四围蒙福；我也必叫时雨落下，使福如甘霖降下。
EZEK|34|27|田野的树木必结果子，地也必有出产；他们要在自己的土地安然居住。我折断他们所负的轭，救他们脱离奴役他们之人的手；那时，他们就知道我是耶和华。
EZEK|34|28|他们必不再作外邦人的掠物，地上的野兽也不再吞吃他们；他们却要安然居住，无人使他们惊吓。
EZEK|34|29|我必为他们建立闻名的 栽种之地；他们在境内就不再为饥荒所灭，也不再受列国的羞辱。
EZEK|34|30|他们必知道我─耶和华他们的上帝与他们同在，并知道他们， 以色列 家，是我的子民。这是主耶和华说的。
EZEK|34|31|你们这些人，你们是我的羊，我草场上的羊；我是你们的上帝。这是主耶和华说的。”
EZEK|35|1|耶和华的话临到我，说：
EZEK|35|2|“人子啊，你要面向 西珥山 ，向它说预言，
EZEK|35|3|对它说，主耶和华如此说： 西珥山 ，看哪，我与你为敌，必伸手攻击你，使你荒凉荒废。
EZEK|35|4|我必使你的城镇变为废墟，使你成为荒凉；你就知道我是耶和华。
EZEK|35|5|因为你永怀仇恨，在 以色列 人遭遇灾难、罪孽到了尽头时，把他们交给刀剑，
EZEK|35|6|所以主耶和华说：我指着我的永生起誓，我必使你遭遇血的报应，血必追赶你；你既不恨恶血，血必追赶你。
EZEK|35|7|我要使 西珥山 荒凉荒废，把来往经过的人从它那里剪除。
EZEK|35|8|我要使 西珥山 布满被杀的人。被刀杀的要倒在小山和山谷，并一切的溪水中。
EZEK|35|9|我必使你永远荒凉，使你的城镇无人居住，你们就知道我是耶和华。
EZEK|35|10|“因为你曾说‘这二国、这二邦必归我，我们必得为业’，其实耶和华仍在那里；
EZEK|35|11|所以主耶和华说：我指着我的永生起誓，我必照你因仇恨向他们发的怒气和嫉妒对待你；我审判你的时候，要在他们中间显明自己。
EZEK|35|12|你必知道我─耶和华已听见你一切凌辱的话，是针对 以色列 群山说的：‘这些山荒凉了，它们是给我们作食物的。’
EZEK|35|13|你们用口向我说夸大的话，增多与我敌对的话，我都听见了。
EZEK|35|14|主耶和华如此说：全地欢乐的时候，我必使你荒凉。
EZEK|35|15|你怎样因 以色列 家的地业荒凉而喜乐，我也要照你所做的对待你。 西珥山 哪，你和 以东 全地都必荒凉；人就知道 我是耶和华。”
EZEK|36|1|“人子啊，你要对 以色列 群山说预言： 以色列 群山哪，要听耶和华的话。
EZEK|36|2|主耶和华如此说，因仇敌说：‘啊哈！这古老的丘坛都归我们为业了！’
EZEK|36|3|所以你要预言，说：主耶和华如此说：因为敌人使你荒凉，四围践踏你，要叫你归其余的列国为业，使你们成为各族的话柄与百姓的笑谈；
EZEK|36|4|因此， 以色列 群山哪，要听主耶和华的话。对那遭四围其余列国占据、讥刺的大山小冈、水沟山谷、荒废之地、被弃之城，主耶和华如此说；
EZEK|36|5|所以，主耶和华如此说：我因妒火中烧，就责备其余的列国和 以东 的众人。他们快乐满怀，心存恨恶，将我的地占为己有，视为被抛弃的掠物。
EZEK|36|6|所以，你要指着 以色列 地说预言，对大山小冈、水沟山谷说，主耶和华如此说：看哪，我在妒忌和愤怒中宣布：因你们曾受列国的羞辱，
EZEK|36|7|所以我起誓说，你们四围的列国要担当自己的羞辱。这是主耶和华说的。
EZEK|36|8|“ 以色列 群山哪，要长出枝条，为我子民 以色列 结出果子，因为他们即将来到。
EZEK|36|9|看哪，我是帮助你们的，我要转向你们，使你们得以耕作栽种。
EZEK|36|10|我要使 以色列 全家在你们那里人数增多，城镇有人居住，废墟重新建造。
EZEK|36|11|我要使人丁和牲畜在你们那里加增，他们必生养众多。我要使你们那里像以前一样有人居住，并要赐福，比先前更多；你们就知道我是耶和华。
EZEK|36|12|我要使我的子民 以色列 在你们那里行走，他们必得你为业；你就成为他们的产业，不再使他们丧失儿女。
EZEK|36|13|主耶和华如此说，因为人对你们说‘你是吞吃人的，又使国民丧失儿女’，
EZEK|36|14|所以你必不再吞吃人，也不再使国民丧失儿女。这是主耶和华说的。
EZEK|36|15|我使你不再听见列国的羞辱；你必不再受万民的辱骂，也不再使国民绊跌。这是主耶和华说的。”
EZEK|36|16|耶和华的话临到我，说：
EZEK|36|17|“人子啊， 以色列 家住本地的时候，所作所为使那地玷污。他们的行为在我面前，好像妇人在经期中那样污秽。
EZEK|36|18|所以我因他们在那地流人的血，且以偶像使那地玷污，就把我的愤怒倾倒在他们身上。
EZEK|36|19|我将他们分散到列国，四散在列邦，按他们的所作所为惩罚他们。
EZEK|36|20|他们到了 所去的列国，使我的圣名被亵渎；因为人谈论他们说，这是耶和华的子民，却从耶和华的地出来。
EZEK|36|21|但我顾惜我的圣名，就是 以色列 家在所到的列国中亵渎的。
EZEK|36|22|“所以，你要对 以色列 家说，主耶和华如此说： 以色列 家啊，我做这事不是为你们，而是为了我的圣名，就是你们在所到的列国中亵渎的。
EZEK|36|23|我要使我至大的名显为圣；这名在列国中已遭亵渎，是你们在他们中间亵渎的。我在他们眼前，在你们身上显为圣的时候，他们就知道我是耶和华。这是主耶和华说的。
EZEK|36|24|我必从列国带领你们，从列邦聚集你们，领你们回到本地。
EZEK|36|25|我必洒清水在你们身上，你们就洁净了。我要洁净你们，使你们脱离一切的污秽，弃绝一切的偶像。
EZEK|36|26|我也要赐给你们一颗新心，将新灵放在你们里面，又从你们的肉体中除掉石心，赐给你们肉心。
EZEK|36|27|我必将我的灵放在你们里面，使你们顺从我的律例，谨守遵行我的典章。
EZEK|36|28|你们必住在我所赐给你们祖先之地；你们要作我的子民，我要作你们的上帝。
EZEK|36|29|我要救你们脱离一切的污秽，也要令五谷丰登，使你们不再遭遇饥荒。
EZEK|36|30|我要使树木多结果子，田地多出土产，好叫你们不再因饥荒被列国凌辱。
EZEK|36|31|那时，你们必追念自己的恶行和不好的作为，就因你们的罪孽和可憎的事厌恶自己。
EZEK|36|32|你们要知道，我这样做不是为你们。 以色列 家啊，你们当为自己的行为抱愧蒙羞。这是主耶和华说的。
EZEK|36|33|“主耶和华如此说：我洁净你们，使你们脱离一切罪孽的日子，必使城镇有人居住，废墟重新建造。
EZEK|36|34|这荒芜的土地，曾被过路的人看为荒芜，现今却得以耕种。
EZEK|36|35|他们必说：‘这荒芜之地，现在成了像 伊甸园 一样；这荒凉、荒废、毁坏的城镇，现今坚固，有人居住。’
EZEK|36|36|那时，在你们四围其余的列国必知道，我─耶和华修造那毁坏之处，开垦那荒芜之地。我─耶和华说了这话，就必成就。
EZEK|36|37|“主耶和华如此说：我要回应 以色列 家的求问，成全他们，增添他们的人数，使他们多如羊群。
EZEK|36|38|在 耶路撒冷 守节时，作为祭物所献的羊群有多少，照样，荒凉的城镇必为人群所充满；他们就知道我是耶和华。”
EZEK|37|1|耶和华的手按在我身上。耶和华藉着他的灵带我出去，把我放在平原中，平原遍满骸骨。
EZEK|37|2|他使我从骸骨的四围经过，看哪，平原上面的骸骨甚多，看哪，极其枯干。
EZEK|37|3|他对我说：“人子啊，这些骸骨能活过来吗？”我说：“主耶和华啊，你是知道的。”
EZEK|37|4|他又对我说：“你要向这些骸骨说预言，对它们说：枯干的骸骨啊，要听耶和华的话。
EZEK|37|5|主耶和华对这些骸骨如此说：‘看哪，我必使气息 进入你们里面，你们就要活过来。
EZEK|37|6|我要给你们加上筋，长出肉，又给你们包上皮，使气息进入你们里面，你们就要活过来；你们就知道我是耶和华。’”
EZEK|37|7|于是，我遵命说预言。正说预言的时候，有响声，看哪，有地震；骨与骨彼此接连。
EZEK|37|8|我观看，看哪，骸骨上面有筋，长了肉，又包上皮，只是里面还没有气息。
EZEK|37|9|耶和华对我说：“人子啊，你要说预言，向风 说预言。你要说，耶和华如此说：气息啊，要从四方 而来，吹在这些被杀的人身上，使他们活过来。”
EZEK|37|10|于是我遵命说预言，气息就进入骸骨，骸骨就活过来，并且用脚站起来，成为极大的军队。
EZEK|37|11|他对我说：“人子啊，这些骸骨就是 以色列 全家。他们说：‘看哪，我们的骨头枯干了，我们的指望失去了，我们灭绝净尽了！’
EZEK|37|12|所以你要说预言，对他们说，主耶和华如此说：我的子民，看哪，我要打开你们的坟墓，把你们带出坟墓，领你们进入 以色列 地。
EZEK|37|13|我的子民哪，我打开你们的坟墓，把你们带出坟墓时，你们就知道我是耶和华。
EZEK|37|14|我必将我的灵放在你们里面，你们就要活过来。我把你们安置在本地，你们就知道我─耶和华说了这话，就必成就。这是耶和华说的。”
EZEK|37|15|耶和华的话临到我，说：
EZEK|37|16|“人子啊，你要取一根木杖，在其上写‘为 犹大 和他的盟友 以色列 人’；又取一根 木杖，在其上写‘为 约瑟 ，就是 以法莲 的杖，和他的盟友 以色列 全家’。
EZEK|37|17|你要将这两根木杖彼此相接，连成一根，使它们在你手中合而为一。
EZEK|37|18|当你本国的子民对你说：‘你这是什么意思，你不指示我们吗？’
EZEK|37|19|你就对他们说，主耶和华如此说：看哪，我要将 约瑟 和他的盟友 以色列 支派的杖，就是在 以法莲 手中的那根，与 犹大 的杖接连成为一根，在我手中合而为一。
EZEK|37|20|你要在他们眼前，把写了字的那两根杖拿在手中，
EZEK|37|21|对他们说，主耶和华如此说：看哪，我要从 以色列 人所到的列国带领他们，从四围聚集他们，领他们回到本地。
EZEK|37|22|我要使他们在这地，在 以色列 群山上成为一国，必有一王作他们全体的王。他们不再成为二国，绝不再分为二国。
EZEK|37|23|他们不再因偶像和可憎的物，并一切的罪过玷污自己。我却要救他们离开一切犯罪所住的地方 ；我要洁净他们，如此，他们要作我的子民，我要作他们的上帝。’
EZEK|37|24|“我的仆人 大卫 要作他们的王；他们全体必归一个牧人。他们必顺从我的典章，谨守遵行我的律例。
EZEK|37|25|他们要住在我赐给我仆人 雅各 的地上，就是你们列祖所住之地。他们和他们的子孙，并子孙的子孙，都永远住在那里。我的仆人 大卫 要作他们的王，直到永远；
EZEK|37|26|并且我要与他们立平安的约，作为永约。我要安顿他们，使他们人数增多，又在他们中间设立我的圣所，直到永远。
EZEK|37|27|我的居所必在他们中间；我要作他们的上帝，他们要作我的子民。
EZEK|37|28|我的圣所在 以色列 人中间直到永远，列国就知道是我─耶和华使 以色列 分别为圣。”
EZEK|38|1|耶和华的话临到我，说：
EZEK|38|2|“人子啊，你要面向 玛各 地的 歌革 ，就是 米设 和 土巴 的大王，向他说预言。
EZEK|38|3|你要说，主耶和华如此说： 米设 和 土巴 的大王 歌革 ，看哪，我与你为敌。
EZEK|38|4|我要把你掉转过来，用钩子钩住你的腮颊，把你和你的军兵、马匹、骑兵都带走。他们全都披挂整齐，成为大军，佩带大小盾牌，各人拿着刀剑；
EZEK|38|5|他们当中有 波斯 人、 古实 人和 弗 人，都带着盾牌和头盔；
EZEK|38|6|还有 歌篾 人和他的军队，北方极远的 陀迦玛 族和他的军队，这许多民族都跟着你。
EZEK|38|7|“你和聚集到你那里的军队都要预备，预备妥当，你要作他们的守卫。
EZEK|38|8|过了多日，你必被差派；到末后之年，你要来到那脱离刀剑、从列国召集回来的人所住之地，来到 以色列 常久荒凉的山上；他们都从列国中被领出，在那里安然居住。
EZEK|38|9|你和你的全军，并跟随你的许多民族都要上来，如暴风刮来，如密云遮盖地面。
EZEK|38|10|“主耶和华如此说：那时，你的心必起意念，图谋恶计，
EZEK|38|11|说：‘我要上那无墙的乡村之地，到那安静的居民那里，他们无墙，无门、无闩，安然居住。
EZEK|38|12|我去那里要抢财为掳物，夺货为掠物，反手攻击那从前荒凉、现在有人居住之地，又攻击那从列国招聚出来、得了牲畜财货、住在地的高处的百姓。’
EZEK|38|13|示巴 人、 底但 人、 他施 的商人和他们的少壮狮子都对你说：‘你来是要抢财为掳物吗？你聚集军队是要夺货为掠物，夺取金银，掳去牲畜、财货，抢夺许多财宝为掳物吗？’
EZEK|38|14|“人子啊，你要因此说预言，对 歌革 说，主耶和华如此说：我的子民 以色列 安然居住时，你是知道的。
EZEK|38|15|你从你的地方，从北方极远处率领许多民族前来，他们都骑着马，是一队强而多的军兵。
EZEK|38|16|歌革 啊，你必上来攻击我的子民 以色列 ，如密云遮盖地面。末后的日子，我必领你来攻击我的地，我藉你在列国眼前显为圣的时候，他们就要认识我。
EZEK|38|17|主耶和华如此说：我在古时藉我仆人 以色列 众先知所说的，不就是你吗？ 他们在那些日子，多年说预言，我必领你来攻击 以色列 人。”
EZEK|38|18|“主耶和华说： 歌革 上来攻击 以色列 地的时候，我的怒气要从鼻孔里发出。
EZEK|38|19|我在妒忌和如火的烈怒中说：那日在 以色列 地必有大震动，
EZEK|38|20|甚至海中的鱼、天空的鸟、野地的兽，和地上爬的各种爬行动物，并地面上的众人，因见我的面就都震动；山岭崩裂，陡岩塌陷，一切的墙都必坍塌。
EZEK|38|21|我必令刀剑在我的众山攻击 歌革 ；人要用刀剑杀害弟兄。这是主耶和华说的。
EZEK|38|22|我要用瘟疫和血惩罚他。我也必降暴雨、大冰雹、火及硫磺在他和他的军队，并跟随他的许多民族身上。
EZEK|38|23|我必显为大，显为圣，在许多国家眼前显明自己；他们就知道我是耶和华。”
EZEK|39|1|“你，人子啊，要向 歌革 说预言。你要说，主耶和华如此说： 米设 和 土巴 的大王 歌革 ，看哪，我与你为敌。
EZEK|39|2|我要把你调转过来，带领你，从北方极远的地方上来，带你到 以色列 的群山上。
EZEK|39|3|我要打落你左手的弓，打掉你右手的箭。
EZEK|39|4|你和你的全军，并跟随你的列国的人，都必倒在 以色列 的群山上。我要将你给各类攫食的飞鸟和野地的走兽作食物。
EZEK|39|5|你必倒在田野，因为我曾说过，这是主耶和华说的。
EZEK|39|6|我要降火在 玛各 和海岛安然居住的人身上，他们就知道我是耶和华。
EZEK|39|7|“我要在我的子民 以色列 中彰显我的圣名，不容我的圣名再被亵渎，列国就知道我─耶和华是 以色列 中的圣者。
EZEK|39|8|看哪，时候到了，必然成就，这就是我曾说过的日子。这是主耶和华说的。
EZEK|39|9|“住 以色列 城镇的人要出去生火，用军器燃烧，就是大小盾牌、弓箭、棍棒、枪矛；用它们来烧火，直烧了七年。
EZEK|39|10|他们不必从田野捡柴，也不必从森林伐木，因为他们要用这些军器烧火。他们要抢夺那抢夺他们的人，掳掠那掳掠他们的人。这是主耶和华说的。”
EZEK|39|11|“当那日，我要把 以色列 境内、海东边的 旅人谷 给 歌革 在那里作坟地 ，阻挡了旅行的人 。在那里，人要埋葬 歌革 和他的军兵，称那地为 哈们．歌革谷 。
EZEK|39|12|以色列 家的人要用七个月埋葬他们，好使那地洁净。
EZEK|39|13|那地所有的百姓都来埋葬他们。当我得荣耀的日子，这事必叫百姓得名声。这是主耶和华说的。
EZEK|39|14|他们要分派人专职巡查遍地，埋葬那遗留在地面上入侵者的尸首，好洁净全地。过了七个月，他们还要再巡查。
EZEK|39|15|巡查的人要遍行全地，见有人的骸骨，就在旁边立一标记，等埋葬的人来将骸骨葬在 哈们．歌革谷 ，
EZEK|39|16|且有一城要取名为 哈摩那 。他们必这样洁净那地。
EZEK|39|17|“你，人子啊，主耶和华如此说：你要向各类的飞鸟和野地的走兽说：你们要聚集，来吧，从四方聚集来吃我为你们准备的祭物，就是在 以色列 的群山上丰盛的祭物，叫你们吃肉、喝血。
EZEK|39|18|你们要吃勇士的肉，喝地上领袖的血，如吃公绵羊、羔羊、公山羊、公牛；他们全都是 巴珊 的肥畜。
EZEK|39|19|你们吃我为你们准备的祭物，必吃油脂直到饱了，喝血直到醉了。
EZEK|39|20|你们要因我席上的马匹、骑兵、勇士和所有的战士而饱足。这是主耶和华说的。”
EZEK|39|21|“我要在列国中彰显我的荣耀，万国就必看见我怎样把手加在他们身上，施行审判。
EZEK|39|22|从那日以后， 以色列 家就知道我是耶和华─他们的上帝，
EZEK|39|23|列国也必知道， 以色列 家被掳掠是因他们的罪孽。他们得罪我，我就转脸不顾他们，将他们交在敌人手中，使他们全都倒在刀下。
EZEK|39|24|我照他们的污秽和罪过待他们，转脸不顾他们。
EZEK|39|25|“所以主耶和华如此说：现在，我要使 雅各 被掳的人归回，要怜悯 以色列 全家，又为我的圣名发热心。
EZEK|39|26|我将他们从万民中领回，从仇敌之地召来，在许多国家的眼前，在他们身上显为圣，他们在本地安然居住，无人使他们惊吓，那时，他们要担当 自己的羞辱和干犯我的一切罪。
EZEK|39|27|
EZEK|39|28|我使他们被掳到列国，后又聚集他们回到本地，不再留一人在那里，那时他们就知道我是耶和华─他们的上帝。
EZEK|39|29|我不再转脸不顾他们，因我已将我的灵浇灌 以色列 家。这是主耶和华说的。”
EZEK|40|1|我们被掳的第二十五年， 耶路撒冷城 攻破后十四年，正在年初，某月初十，就在那一天，耶和华的手按在我身上，把我带到那里。
EZEK|40|2|在上帝的异象中，他带我到 以色列 地，把我安置在一座极高的山上；在山的南边有仿佛一座城的建筑物。
EZEK|40|3|他带我到那里，看哪，有一人面貌 如铜，手拿麻绳和丈量的芦苇竿，站在门口。
EZEK|40|4|那人对我说：“人子啊，凡我所指示你的，你都要用眼看，用耳听，并要放在心上。我带你到这里来，为要指示你；凡你所见的，都要告诉 以色列 家。”
EZEK|40|5|看哪，殿外四围有墙。那人手拿丈量的芦苇竿，长六肘，每肘再加一掌。他量围墙，宽一竿，高一竿。
EZEK|40|6|他到了朝东的门，就上台阶，量这门的门槛，宽一竿；这门槛宽一竿。
EZEK|40|7|又有守卫房，每间长一竿，宽一竿，守卫房之间相隔五肘。挨着通往殿之门走廊的门槛，一竿。
EZEK|40|8|他量通往殿之门的走廊，一竿。
EZEK|40|9|他量门的走廊，八肘；墙柱，二肘；门的走廊通往殿那里。
EZEK|40|10|往东的门有守卫房：这旁三间，那旁三间，大小都一样；这边和那边的墙柱，大小也一样。
EZEK|40|11|他量门的入口，宽十肘，门长十三肘。
EZEK|40|12|守卫房前有矮墙，一肘，那边的矮墙也是一肘；守卫房这边六肘，那边也是六肘。
EZEK|40|13|他量门，从守卫房这边的房顶到那边的房顶，宽二十五肘；入口与入口相对。
EZEK|40|14|他量墙柱，六十肘，院子的四周围有挨着墙柱的门。
EZEK|40|15|从大门入口到里面门的走廊，五十肘。
EZEK|40|16|守卫房和四围挨着墙柱的门，都有嵌壁式的窗户，廊子也有；里面到处都有窗户，墙柱上雕刻着棕树。
EZEK|40|17|他带我到外院，看哪，院子的四围有房间，有石板地；石板地上有三十个房间。
EZEK|40|18|沿着门侧边的石板地，就是下面的石板地，与门的长度相同。
EZEK|40|19|他量宽度，从下门的前面到内院外的前面，东向北向一百肘。
EZEK|40|20|他量外院朝北的门的长和宽。
EZEK|40|21|门的守卫房，这旁三间，那旁三间；墙柱和廊子，与第一个门的大小一样。长五十肘，宽二十五肘。
EZEK|40|22|其窗户和廊子，并雕刻的棕树，与朝东的门大小一样。要登七个台阶才能上到这门，前面 有廊子。
EZEK|40|23|内院有门与这门相对，北面东面都是如此。他从这门量到那门，共一百肘。
EZEK|40|24|他带我往南去，看哪，朝南有门，他量门的墙柱 和廊子，大小与先前一样。
EZEK|40|25|门两旁与廊子的周围都有窗户，和先前量的窗户一样。门长五十肘，宽二十五肘。
EZEK|40|26|要登七个台阶才能上到这门，前面 有廊子；墙柱上雕刻着棕树，这边一棵，那边一棵。
EZEK|40|27|内院朝南也有门，从这门量到朝南的那门，共一百肘。
EZEK|40|28|他带我从南门到内院，他量南门，大小与先前一样。
EZEK|40|29|守卫房和墙柱、廊子，大小与先前一样。门两旁与廊子的周围都有窗户。门长五十肘，宽二十五肘。
EZEK|40|30|周围有廊子，长二十五肘，宽五肘。
EZEK|40|31|廊子朝着外院，墙柱上雕刻着棕树。要登八个台阶才能上到这门。
EZEK|40|32|他带我到内院的东边，他量那门，大小与先前一样。
EZEK|40|33|守卫房和墙柱、廊子，大小与先前一样。门两旁与廊子的周围都有窗户。长五十肘，宽二十五肘。
EZEK|40|34|廊子朝着外院。墙柱两边都雕刻着棕树。要登八个台阶才能上到这门。
EZEK|40|35|他带我到北门，他量了，大小与先前一样，
EZEK|40|36|就是量守卫房和墙柱、廊子。门的周围都有窗户；门长五十肘，宽二十五肘。
EZEK|40|37|墙柱 朝着外院。墙柱两边都雕刻着棕树。要登八个台阶才能上到这门。
EZEK|40|38|有房间和它的入口在门的墙柱 旁，那里是洗燔祭牲的地方。
EZEK|40|39|在门的走廊内，这边有两张桌子，那边也有两张桌子，其上可宰杀燔祭牲、赎罪祭牲和赎愆祭牲。
EZEK|40|40|上到北门的入口，朝向外面的这边有两张桌子，门的走廊那边也有两张桌子。
EZEK|40|41|门这边有四张桌子，那边也有四张桌子，共八张，在其上宰杀祭牲。
EZEK|40|42|为燔祭牲的四张桌子是用石头凿成的，长一肘半，宽一肘半，高一肘。宰杀燔祭牲和其他祭牲所用的器皿可放在其上。
EZEK|40|43|有钩子，宽一掌，挂在廊内的四周围。桌子上可放祭牲的肉。
EZEK|40|44|从外面进到内门，内院里有房间，为歌唱的人而设 ；一间在北门旁，朝南，又有一间在南 门旁，朝北。
EZEK|40|45|他对我说：“这朝南的房间是为了圣殿供职的祭司，
EZEK|40|46|那朝北的房间是为了祭坛前供职的祭司；这些祭司是 利未 人中 撒督 的子孙，近前来事奉耶和华的。”
EZEK|40|47|他又量内院，长一百肘，宽一百肘，是正方的。祭坛就在殿前。
EZEK|40|48|于是他带我到殿前的走廊，量走廊的墙柱。这面宽五肘，那面宽五肘。 门的两旁，这边三肘，那边三肘。
EZEK|40|49|走廊长二十肘，宽十一肘 。要登台阶 才能上到走廊。靠近墙柱又有柱子，这边一根，那边一根。
EZEK|41|1|他带我到殿那里，他量墙柱：这面宽六肘，那面宽六肘，宽窄与会幕相同 。
EZEK|41|2|门口宽十肘。门的两旁，这边五肘，那边五肘。他又量了殿，长四十肘，宽二十肘。
EZEK|41|3|他到内殿量门的墙柱，二肘，门口六肘，门的两旁各宽七肘。
EZEK|41|4|他量内殿，长二十肘，宽二十肘。他对我说：“这是至圣所。”
EZEK|41|5|他又量殿的墙，六肘；围着殿有厢房，各宽四肘。
EZEK|41|6|厢房有三层，层叠而上，每层排列三十间。殿的墙四周有凸出的墙支撑厢房，厢房就不必以殿的墙为支柱。
EZEK|41|7|这围绕着殿的厢房越高越宽；厢房围着殿悬叠而上，所以越上面越宽，从下一层，到中一层，到上一层。
EZEK|41|8|我又见有高台围绕着殿，作为厢房的根基，高足足有一竿，就是六大肘。
EZEK|41|9|厢房的外墙宽五肘。殿的厢房和那边的房间中间还有空地，宽二十肘，围绕着殿。
EZEK|41|10|
EZEK|41|11|厢房的门口向着空地：一门向北，一门向南。周围的空地宽五肘。
EZEK|41|12|在西边空地之后有房子，宽七十肘，长九十肘，墙四围厚五肘。
EZEK|41|13|这样，他量了殿，长一百肘，又量空地和那房子并墙，共长一百肘。
EZEK|41|14|殿的前面和东边的空地，宽一百肘。
EZEK|41|15|他量了空地后面的那房子，并两旁的楼廊，共长一百肘。 内殿、院的走廊、
EZEK|41|16|门槛 、嵌壁式的窗户，并对着门槛的三层楼廊，周围都镶上木板；地板到窗户，窗户都关着，
EZEK|41|17|直到门以上，就是到内殿和外殿内外四围墙壁，都这样测量。
EZEK|41|18|墙上雕刻基路伯和棕树，基路伯和基路伯之间有一棵棕树，每基路伯有两张脸；
EZEK|41|19|人的脸向着这边的棕树，狮子的脸向着那边的棕树，殿内四周围都是如此。
EZEK|41|20|从地板到门的上面，都有基路伯和棕树。殿的墙就是这样。
EZEK|41|21|殿的门柱是方的。至圣所的前面有个东西形状像
EZEK|41|22|木头做的坛，高三肘，长二肘 。坛角和底座 ，并四面，都是木头做的。他对我说：“这是耶和华面前的供桌。”
EZEK|41|23|殿和圣所各有一个双层门。
EZEK|41|24|每个门有两扇，每扇又有两个摺叠页；这一扇有两页，另一扇也有两页。
EZEK|41|25|殿的门扇上雕刻着基路伯和棕树，与刻在墙上的一样。在外面门的走廊前有木头做的飞檐。
EZEK|41|26|门的走廊这边和那边都有嵌壁式的窗户和棕树；殿的厢房和飞檐也是这样。
EZEK|42|1|他带我出来往北，到外院，又带我进入一个房间，一面对着空地，一面对着北边的房子。
EZEK|42|2|前面长一百肘，宽五十肘，有门向北；
EZEK|42|3|对着内院那二十肘 ，又对着外院的石板地，在第三层楼有楼廊对着楼廊。
EZEK|42|4|那些房间前有一条走道，宽十肘，往里面有宽一肘的通道 。房门都向北。
EZEK|42|5|房间因为楼廊占掉一些地方，所以房子的上层比中下两层窄。
EZEK|42|6|房间分三层，却不像外院的屋子用柱子支撑，而是从地面往上，所以一层比一层更窄。
EZEK|42|7|外面有一道墙，长五十肘，在房间前面，与朝外院的房间平行。
EZEK|42|8|靠着外院的房间长五十肘，看哪，朝圣殿的长一百肘。
EZEK|42|9|这些房间下面的东边有一个入口，从外院可由此进入；
EZEK|42|10|其宽如院墙。朝东 也有房间，一面对着空地，一面对着房子。
EZEK|42|11|这些房间前的通道与北边房间的通道一样；长、宽、出口、样式和入口都相同。
EZEK|42|12|在东边通道的开端，正对着那道墙有门可以进入，与向南边房间的门一样。
EZEK|42|13|他对我说：“面对空地南边的房间和北边的房间，都是圣的房间；亲近耶和华的祭司当在那里吃至圣的东西，也当在那里存放至圣的东西，就是素祭、赎罪祭和赎愆祭，因此处为圣。
EZEK|42|14|祭司进圣所，出来的时候，不可直接到外院，要在那里放下他们供职的衣服，因为这是圣衣；要穿上别的衣服才可以到百姓所在之处。”
EZEK|42|15|他量完了内殿的大小，就带我出朝东的门，去量院的四周围。
EZEK|42|16|他用丈量的芦苇竿量东面，五百竿 ；又转去
EZEK|42|17|用丈量的芦苇竿量北面，五百竿；又转去
EZEK|42|18|用丈量的芦苇竿量南面，五百竿。
EZEK|42|19|他又转到西面，用丈量的芦苇竿去量，五百竿。
EZEK|42|20|他量四面，长五百，宽五百，四周围有墙，为要分别圣与俗。
EZEK|43|1|以后，他带我到一座门，就是朝东的门。
EZEK|43|2|看哪， 以色列 上帝的荣光从东而来，他的声音如同众水的响声，地因他的荣耀发光。
EZEK|43|3|我所见的异象如同从前我 来灭城的时候所见的异象，又如我在 迦巴鲁河 边所见的异象，我就脸伏于地。
EZEK|43|4|耶和华的荣光从朝东的门照入殿中。
EZEK|43|5|灵将我举起，带入内院，看哪，耶和华的荣光充满了殿。
EZEK|43|6|我听见有一位从殿中向我说话，有一人站在我旁边。
EZEK|43|7|他对我说：“人子啊，这是我宝座之地，是我脚掌所踏之地。我要住在这里，住在 以色列 人中间直到永远。 以色列 家和他们的君王不可再以淫行，或在高处以君王的尸首 玷污我的圣名。
EZEK|43|8|因他们使自己的门槛挨近我的门槛，使自己的门框挨近我的门框，又使他们与我之间仅隔一墙，并且行可憎的事，玷污我的圣名，所以我发怒灭绝他们。
EZEK|43|9|现在，他们当从我面前远离淫行和君王的尸首，我就要住在他们中间，直到永远。
EZEK|43|10|“你，人子啊，要将这殿指示 以色列 家，让他们量殿的大小 ，使他们因自己的罪孽羞愧。
EZEK|43|11|他们若因自己所做的一切感到羞愧，你就要将殿的规模、样式、出口、入口，以及有关整体规模的条例、礼仪、律法指示他们 ，在他们眼前写下，使他们遵照殿整体的规模和条例去做。
EZEK|43|12|这是殿的律法：山顶上四周围的全地界都称为至圣；看哪，这就是殿的律法 。”
EZEK|43|13|这些是祭坛的大小，以肘来量，这肘是一肘一掌。底座高一肘，边宽一肘，四周围有边，高一虎口；这是祭坛的座 。
EZEK|43|14|从底座到下层的台座，二肘，边宽一肘。从小台座到大台座，四肘，边宽一肘。
EZEK|43|15|坛上的炉台，高四肘，从炉台向上突起四个角。
EZEK|43|16|这炉台长十二肘，宽十二肘，四面见方。
EZEK|43|17|台座长十四肘，宽十四肘，四面见方。四周围有边，高半肘，底座四围的边宽一肘。有台阶朝东。
EZEK|43|18|他对我说：“人子啊，主耶和华如此说：这些是建造祭坛，为要在其上献燔祭，把血洒在上面的条例：
EZEK|43|19|你要将一头公牛犊作为赎罪祭，交给那近前来事奉我的 利未 家的祭司 撒督 的后裔；这是主耶和华说的。
EZEK|43|20|你要取那公牛犊的一些血，抹在坛的四角和台座的四角，并周围的边上。你要这样洁净坛，为坛赎罪。
EZEK|43|21|你又要将那作赎罪祭的公牛烧在圣所外面，殿的预定之处。
EZEK|43|22|次日，要将无残疾的公山羊献为赎罪祭；要洁净坛，像用公牛洁净一样。
EZEK|43|23|你洁净了坛，就要将一头无残疾的公牛犊和羊群中一只无残疾的公绵羊
EZEK|43|24|奉到耶和华面前。祭司要撒盐在其上，献给耶和华为燔祭。
EZEK|43|25|七日内，你要每日献一只公山羊为赎罪祭，也要献一头公牛犊和羊群中的一只公绵羊，都要没有残疾的。
EZEK|43|26|七日内祭司要为坛赎罪，使它洁净，把它分别为圣。
EZEK|43|27|满了七日，自八日以后，祭司要在坛上献你们的燔祭和平安祭；我必悦纳你们。这是主耶和华说的。”
EZEK|44|1|他又带我回到圣所朝东的外门，那门关闭了。
EZEK|44|2|耶和华对我说：“这门必须关闭，不可敞开，谁也不可由其中进入；因为耶和华─ 以色列 的上帝已经由其中进入，所以必须关闭。
EZEK|44|3|至于君王，他必按君王的位分坐在其内，在耶和华面前吃饼。他必由这门的走廊而入，也必由此而出。”
EZEK|44|4|他又带我由北门来到殿前。我观看，看哪，耶和华的荣光充满耶和华的殿，我就脸伏于地。
EZEK|44|5|耶和华对我说：“人子啊，我对你所说耶和华殿中一切的条例和律法，你要留心，用眼看，用耳听，要留心殿的入口和圣所一切的出口。
EZEK|44|6|你要对那悖逆的 以色列 家说，主耶和华如此说： 以色列 家啊，你们行这一切可憎的事，够了吧！
EZEK|44|7|你们把我的食物，就是脂肪和血献上的时候，竟把心和肉体未受割礼的外邦人领进我的圣所，玷污我的殿；你们行这一切可憎的事，违背了我的约。
EZEK|44|8|你们未尽看守我圣物的职责，竟派别人在我的圣所替你们尽看守之责。
EZEK|44|9|“主耶和华如此说：所有心和肉体未受割礼的外邦人，就是住在 以色列 中间的任何外邦人，都不可进入我的圣所。”
EZEK|44|10|“ 以色列 人走迷的时候， 利未 人远离我，随从他们的偶像走迷离开我，他们必担当自己的罪孽。
EZEK|44|11|他们必在我的圣所当仆役，照管殿门，在殿里伺候；他们要为百姓宰杀燔祭牲和其他祭牲，站在百姓面前伺候他们。
EZEK|44|12|因为这些 利未 人曾在偶像前伺候他们，成了 以色列 家罪孽的绊脚石，所以我向他们起誓：他们必担当自己的罪孽。这是主耶和华说的。
EZEK|44|13|他们不可亲近我，作事奉我的祭司，也不可挨近我任何一件圣物，就是至圣的物；他们却要担当自己的羞辱和所行可憎之事的报应。
EZEK|44|14|我要指派他们在殿里看守，办理殿中一切事务，做一切当做的工。”
EZEK|44|15|“ 以色列 人走迷离开我的时候， 利未 家的祭司 撒督 的子孙仍然尽看守我圣所的职责；因此他们必亲近我，事奉我，并且侍立在我面前，把脂肪与血献给我。这是主耶和华说的。
EZEK|44|16|只有他们可以进我的圣所，来到我的桌前事奉我，守我吩咐的职责。
EZEK|44|17|他们进内院的门要穿细麻衣，在内院门和殿内供职时不可穿羊毛衣服。
EZEK|44|18|他们要头戴细麻布的头巾，腰穿细麻布的裤子；不可穿容易出汗的衣服。
EZEK|44|19|他们出到外院，到外院 百姓那里，要脱下供职所穿的衣服，放在圣的房间内，换上别的衣服，免得因他们的衣服使百姓成为圣。
EZEK|44|20|他们不可剃头，也不可留长发，头发一定要修剪。
EZEK|44|21|祭司进内院时不可喝酒。
EZEK|44|22|他们不可娶寡妇或被休的妇人为妻，只可娶 以色列 后裔中的处女，或祭司的寡妇。
EZEK|44|23|他们要教导我的子民分辨圣与俗，使他们知道洁净和不洁净的分别。
EZEK|44|24|有争讼的事，他们应当审判，按我的典章审判。他们要在我的节期守我的律法和条例，也当以我的安息日为圣日。
EZEK|44|25|祭司不可挨近死尸使自己不洁净，只可为父亲、母亲、儿子、女儿、兄弟和未出嫁的姊妹使自己不洁净。
EZEK|44|26|他洁净之后，他们必须再为他计算七天。
EZEK|44|27|当他进内院，入圣所，在圣所中事奉的日子，要为自己献上赎罪祭。这是主耶和华说的。
EZEK|44|28|“祭司必有产业，我就是他们的产业。不可在 以色列 中给他们基业，我就是他们的基业。
EZEK|44|29|素祭、赎罪祭和赎愆祭他们都可以吃， 以色列 中一切永献的祭物都归他们。
EZEK|44|30|各样上好的初熟之物和所献的供物，都要归祭司。你们也要将最先的面团给祭司；这样，福气就必临到你们的家。
EZEK|44|31|无论是鸟是兽，凡自然死去的，或是被撕裂的，祭司都不可吃。”
EZEK|45|1|你们抽签分地为业，要献上一份作为献给耶和华的圣地，长二万五千肘 ，宽二万 肘。整个地区都作为圣地。
EZEK|45|2|再从其中划出一块作为圣所，长五百肘，宽五百肘，四面见方；四围再加五十肘的空地。
EZEK|45|3|从这整个范围要划出长二万五千肘，宽一万肘的地，其中要有圣所，是至圣的。
EZEK|45|4|这是地上的一块圣地，要归给在圣所供职、亲近事奉耶和华的祭司，作为他们房屋用地与圣所的圣地。
EZEK|45|5|其余长二万五千肘，宽一万肘，要归给在殿中供职的 利未 人，作为他们二十间房屋 的地业。
EZEK|45|6|在那块献上的圣地旁边，你们要划分造城的地业，宽五千肘，长二万五千肘，归 以色列 全家。
EZEK|45|7|划归君王的地要在献上的圣地和城用地的两旁，面对着圣地，又面对城的用地，西至西边的疆界，东至东边的疆界，从西到东，长度与每支派所分得的一样。
EZEK|45|8|这地要在 以色列 中归君王为业。我所立的君王必不再欺压我的子民，却要按支派把地分给 以色列 家。
EZEK|45|9|主耶和华如此说：“ 以色列 的王啊，你们够了吧！要除掉残暴和抢夺的事，行公平和公义，不可再勒索我的百姓。这是主耶和华说的。
EZEK|45|10|“你们要用公道的天平、公道的伊法、公道的罢特。
EZEK|45|11|伊法要与罢特等量；一罢特为贺梅珥的十分之一，一伊法也是贺梅珥的十分之一，都以贺梅珥为计算单位。
EZEK|45|12|一舍客勒是二十季拉；二十舍客勒，二十五舍客勒，十五舍客勒，合起来为你们的一弥那。
EZEK|45|13|“你们当献的供物是这样：一贺梅珥麦子要献六分之一伊法，一贺梅珥大麦也要献六分之一伊法。
EZEK|45|14|献油的条例是这样，按油的罢特：每一歌珥油，即十罢特或一贺梅珥，要献十分之一罢特，原来十罢特等于一贺梅珥。
EZEK|45|15|从 以色列 水源丰沛的草场上，每二百只羊中要献一只羔羊。这都可作素祭、燔祭、平安祭，来为民赎罪。这是主耶和华说的。
EZEK|45|16|这地所有的百姓都要带这些供物到 以色列 王那里。
EZEK|45|17|王的本分是在节期、初一、安息日，就是 以色列 家一切的盛会，奉上燔祭、素祭、浇酒祭。他要献上赎罪祭、素祭、燔祭和平安祭，为 以色列 家赎罪。”
EZEK|45|18|主耶和华如此说：“正月初一，你要取无残疾的公牛犊，洁净圣所。
EZEK|45|19|祭司要取一些赎罪祭牲的血，抹在殿的门柱上和祭坛台座的四角上，并内院的门框上。
EZEK|45|20|本月初七，你也要为误犯罪的和因无知而犯罪的这样做；你们要为圣殿赎罪。
EZEK|45|21|“正月十四日，你们要守逾越节，七天的节期都要吃无酵饼。
EZEK|45|22|当日，王要为自己和全国百姓预备一头公牛作赎罪祭。
EZEK|45|23|节期的七天内，每天他要预备无残疾的七头公牛、七只公绵羊，给耶和华为燔祭；每天又要预备一只公山羊为赎罪祭。
EZEK|45|24|他也要预备素祭，为一头公牛同献一伊法细面，为一只公绵羊同献一伊法细面，每一伊法加一欣油。
EZEK|45|25|七月十五日守节的时候，七天他都要像这样预备赎罪祭、燔祭、素祭和油。”
EZEK|46|1|主耶和华如此说：“内院朝东的门，在六个工作的日子必须关闭；惟有安息日和初一要敞开。
EZEK|46|2|王从外面要由门的走廊进入，站在门框旁边；祭司要为他预备燔祭和平安祭，王要在门的门槛那里敬拜，然后退出。这门直到晚上不可关闭。
EZEK|46|3|安息日和初一，这地的百姓要在这门口，在耶和华面前敬拜。
EZEK|46|4|安息日，王要用六只无残疾的羔羊、一只无残疾的公绵羊，献给耶和华为燔祭；
EZEK|46|5|同献的素祭，要为公绵羊献一伊法细面，为羔羊则按照他的力量献，一伊法要加一欣油。
EZEK|46|6|初一，他要献一头无残疾的公牛犊、六只羔羊、一只公绵羊，全都要用无残疾的。
EZEK|46|7|他也要预备素祭，为公牛献一伊法细面，为公绵羊献一伊法细面，为羔羊则按照他的力量献，一伊法要加一欣油。
EZEK|46|8|王进入的时候要由这门的走廊而入，也要从原路出去。
EZEK|46|9|“在各节期，这地的百姓朝见耶和华的时候，从北门进入敬拜的，要由南门而出；从南门进入的，要由北门而出。不可从进入的门出去，要往前直行，从对面的门出去。
EZEK|46|10|他们进入时，王也跟他们一同进入；他们出去，他也要出去。
EZEK|46|11|“在节期和盛会的日子同献的素祭，要为一头公牛献一伊法细面，为一只公绵羊献一伊法细面，为羔羊则按照各人的力量献，一伊法要加一欣油。
EZEK|46|12|王奉献甘心祭，就是向耶和华甘心献的燔祭或平安祭时，当有人为他开朝东的门。他就献上燔祭和平安祭，与安息日所献的一样，然后退出。他出去之后，当有人将门关闭。”
EZEK|46|13|“每日，你要取一只无残疾一岁的羔羊献给耶和华为燔祭；要每天早晨献上。
EZEK|46|14|每天早晨你也要预备同献的素祭，六分之一伊法细面，并三分之一欣油，调和细面。这素祭要经常献给耶和华，作为永远的定例。
EZEK|46|15|每天早晨要这样献上羔羊、素祭和油，为经常献的燔祭。”
EZEK|46|16|主耶和华如此说：“王若将礼物赐给他的任何一个儿子，这就成为儿子的产业，可留给子孙，是他们所承受的地业。
EZEK|46|17|倘若王将他产业的一份赐给他的一个臣仆，这就成为他臣仆的产业，直到自由之年，然后地要归还王；王的产业终究要归自己的儿子。
EZEK|46|18|王不可夺取百姓的产业，以致赶逐他们离开自己的地业；他应该从自己的地业中将产业赐给子孙，免得我的子民离开自己的地业，四散各处。”
EZEK|46|19|他带领我从大门旁边的入口，进到朝北为祭司所预备圣的房间，看哪，西边尽头有一块土地。
EZEK|46|20|他对我说：“这是祭司煮赎愆祭牲、赎罪祭牲，烤素祭的地方，免得带出外院，使百姓成为圣。”
EZEK|46|21|他又带我出到外院，使我经过院子的四个角落，看哪，院子的每个角落都有一个小院子。
EZEK|46|22|院子四个角落有小院子，周围有墙，每个小院子长四十肘 ，宽三十肘；四个角落的小院子大小都一样，
EZEK|46|23|小院子周围各有一排石墙，每排石墙下面有炉灶。
EZEK|46|24|他对我说：“这些是煮肉用的屋子，殿内的仆役要在这里煮百姓的祭物。”
EZEK|47|1|他带我回到殿门，看哪，有水从殿的门槛下面往东流出，因为这殿是朝东的。水从殿的侧面，就是右边，从祭坛的南边往下流。
EZEK|47|2|他带我出北门，又领我从外边转到朝东的外门，看哪，水从右边流出。
EZEK|47|3|他手拿绳子往东出去，量了一千肘，使我涉水而过，水到脚踝。
EZEK|47|4|他又量了一千，使我涉水而过，水就到膝；再量了一千，使我过去，水就到腰；
EZEK|47|5|又量了一千，水已成河，无法过去；因为水势高涨成河，只能游泳，无法走过。
EZEK|47|6|他对我说：“人子啊，你看见了吗？” 他带我回到河边。
EZEK|47|7|我回到河边时，看哪，河这边与那边的岸上有极多的树木。
EZEK|47|8|他对我说：“这水往东方流，下到 亚拉巴 ，直到海。所流出来的水，一入海 就使水变淡 。
EZEK|47|9|这两条河 所到之处，凡滋生的动物都必存活；这水流到那里，使那里的水变淡，因此里面有极多的鱼。这河水所到之处，百物都必存活。
EZEK|47|10|必有渔夫站在河边，从 隐．基底 直到 隐．以革莲 ，全都成了晒 网的场所。那里的鱼各从其类，好像大海的鱼甚多。
EZEK|47|11|但是沼泽与池塘的水无法变淡，只能作产盐之用。
EZEK|47|12|河这边与那边的岸上必生长各类树木，可作食物；叶子不枯干，果子不断绝。每月必结新果子，因为这水是从圣所流出来的。树上的果子必作食物，叶子可以治病。”
EZEK|47|13|主耶和华如此说：“这是你们按 以色列 十二支派分地为业的地界， 约瑟 要得两份。
EZEK|47|14|你们承受这地为业，要彼此均分；我曾起誓应许将这地赐给你们的列祖，这地必归你们为业。
EZEK|47|15|“这地的疆界如下：北界从 大海 往 希特伦 ，直到 西达达 口；
EZEK|47|16|又往 哈马 、 比罗他 、 西伯莲 ( 西伯莲 在 大马士革 的边界与 哈马 的边界中间)，到 浩兰 边界的 哈撒．哈提干 。
EZEK|47|17|这样，疆界是从 大海 往 大马士革 地界上的 哈萨．以难 ，北边以 哈马 为界。这是北界。
EZEK|47|18|“东界在 浩兰 和 大马士革 中间， 基列 和 以色列 地的中间，以 约旦河 为界。你们要量疆界直到东海 。这是东界。
EZEK|47|19|“南界是从 他玛 到 加低斯 的 米利巴 水，经 埃及 溪谷 ，直到 大海 。这是南界。
EZEK|47|20|“西界就是 大海 ，从南界直到 哈马口 对面。这是西界。
EZEK|47|21|“你们要为自己按 以色列 的支派分这地。
EZEK|47|22|要抽签分这地为业，归自己和那在你们中间寄居，生儿育女的外人。你们要看他们如本地出生的 以色列 人，他们要在 以色列 支派中与你们同得地业。
EZEK|47|23|外人寄居在哪个支派，你们就在哪里将地业分给他们。这是主耶和华说的。”
EZEK|48|1|众支派的名字如下：从北边尽头，由 希特伦 往 哈马 口，到 大马士革 地界上的 哈萨．以难 。北边靠着 哈马 地，从东到西是 但 的一份。
EZEK|48|2|靠着 但 的地界，从东到西，是 亚设 的一份。
EZEK|48|3|靠着 亚设 的地界，从东到西，是 拿弗他利 的一份。
EZEK|48|4|靠着 拿弗他利 的地界，从东到西，是 玛拿西 的一份。
EZEK|48|5|靠着 玛拿西 的地界，从东到西，是 以法莲 的一份。
EZEK|48|6|靠着 以法莲 的地界，从东到西，是 吕便 的一份。
EZEK|48|7|靠着 吕便 的地界，从东到西，是 犹大 的一份。
EZEK|48|8|靠着 犹大 的地界，从东到西，必有你们所当献的圣地，宽二万五千肘 ；长短与各族从东到西所分的地相同，圣所当在其中。
EZEK|48|9|你们献给耶和华的圣地要长二万五千肘，宽一万肘。
EZEK|48|10|这圣地要归祭司，北长二万五千肘，西宽一万肘，东宽一万肘，南长二万五千肘。耶和华的圣所当在其中。
EZEK|48|11|这地要归 撒督 的子孙中成为圣的祭司，他们谨守我所吩咐的；当 以色列 人走迷的时候，他们不像那些 利未 人走迷了。
EZEK|48|12|在圣地中要特别保留一份归他们，为至圣，紧邻着 利未 人的地界。
EZEK|48|13|利未 人所得的地长二万五千肘，宽一万肘，与祭司的地界相等，都长二万五千肘，宽一万肘。
EZEK|48|14|这地不可卖，不可换；这上好的部分不可转让给别人，因为它归耶和华为圣。
EZEK|48|15|剩下的地长二万五千肘、宽五千肘，要作公用，为造城、盖房、空地之用；城要在中间。
EZEK|48|16|以下是城的大小：北面四千五百肘，南面四千五百肘，东面四千五百肘，西面四千五百肘。
EZEK|48|17|城要有空地，向北二百五十肘，向南二百五十肘，向东二百五十肘，向西二百五十肘。
EZEK|48|18|靠着圣地并排剩余的，东长一万肘，西长一万肘；它与圣地并排，其中所出产的要作城内工人的食物。
EZEK|48|19|以色列 支派中所有在城内做工的，都要耕种这地。
EZEK|48|20|你们要将整块四方的圣地，长二万五千肘，宽二万五千肘，连同城的用地都献作圣地。
EZEK|48|21|圣地和城的用地两边剩余的要归给王。地的东边，南北二万五千肘，东至东界；西边，南北二万五千肘，西至西界；靠着各支派所分的地，都要归给王。圣地和殿的圣所要在其中。
EZEK|48|22|利未 人的地与城的用地都在王的地中间， 犹大 边界和 便雅悯 边界之间，要归给王。
EZEK|48|23|论到其余的支派，从东到西，是 便雅悯 的一份。
EZEK|48|24|靠着 便雅悯 的地界，从东到西，是 西缅 的一份。
EZEK|48|25|靠着 西缅 的地界，从东到西，是 以萨迦 的一份。
EZEK|48|26|靠着 以萨迦 的地界，从东到西，是 西布伦 的一份。
EZEK|48|27|靠着 西布伦 的地界，从东到西，是 迦得 的一份。
EZEK|48|28|靠着 迦得 南边的地界，界限从 他玛 到 加低斯 的 米利巴 水，经 埃及 溪谷 ，直到 大海 。
EZEK|48|29|这就是你们要抽签分给 以色列 支派为业之地，是他们各支派所得的份。这是主耶和华说的。
EZEK|48|30|以下是城的出口：北面四千五百肘，
EZEK|48|31|城的各门要按 以色列 的支派命名。北面有三个门，一为 吕便 门，一为 犹大 门，一为 利未 门。
EZEK|48|32|东面四千五百肘，有三个门，一为 约瑟 门，一为 便雅悯 门，一为 但 门。
EZEK|48|33|南面四千五百肘，有三个门，一为 西缅 门，一为 以萨迦 门，一为 西布伦 门。
EZEK|48|34|西面四千五百肘，有三个门，一为 迦得 门，一为 亚设 门，一为 拿弗他利 门。
EZEK|48|35|城的周围共一万八千肘。从此以后，这城的名字必称为“耶和华的所在”。
DAN|1|1|犹大 王 约雅敬 在位第三年， 巴比伦 王 尼布甲尼撒 来到 耶路撒冷 ，将城围困。
DAN|1|2|主将 犹大 王 约雅敬 和上帝殿中的一些器皿交在他的手中。他就把他们带到 示拿 地他神明的庙里，将器皿收入他神明的库房中。
DAN|1|3|王吩咐太监长 亚施毗拿 ，从 以色列 人的王室后裔和贵族中带进几个人来，
DAN|1|4|就是没有残疾、相貌俊美、通达各样学问 、知识聪明俱备、足能在王宫侍立的少年，要教他们 迦勒底 的文字和语言。
DAN|1|5|王从自己所用的膳和所饮的酒中，派给他们每日的分量，养育他们三年，好叫他们期满以后侍立在王面前。
DAN|1|6|他们中间有 犹大 人 但以理 、 哈拿尼雅 、 米沙利 和 亚撒利雅 。
DAN|1|7|太监长给他们另外起名，称 但以理 为 伯提沙撒 ，称 哈拿尼雅 为 沙得拉 ，称 米沙利 为 米煞 ，称 亚撒利雅 为 亚伯尼歌 。
DAN|1|8|但以理 却立志，不以王的膳和王所饮的酒玷污自己，于是恳求太监长容他不使自己玷污。
DAN|1|9|上帝使 但以理 在太监长眼前蒙恩，得怜悯。
DAN|1|10|太监长对 但以理 说：“我惧怕我主我王，他已经派给你们饮食，何必让他见你们的面貌比你们同年龄的少年憔悴呢？这样，你们就使我的头在王那里不保了。”
DAN|1|11|但以理 对太监长所派监管 但以理 、 哈拿尼雅 、 米沙利 、 亚撒利雅 的管理者说：
DAN|1|12|“请你考验仆人们十天，给我们素菜吃，清水喝，
DAN|1|13|然后你亲自观察我们的面貌和那用王膳的少年的面貌；就照你所观察的待你的仆人吧！”
DAN|1|14|管理者准许他们这件事，考验他们十天。
DAN|1|15|过了十天，他们的身材看来比所有享用王膳的少年更加俊美健壮，
DAN|1|16|于是管理者撤去王派给他们用的膳和所饮的酒，只给他们素菜。
DAN|1|17|这四个少年，上帝在各样文字学问上赐给他们知识和聪明； 但以理 又明白各样异象和梦兆。
DAN|1|18|王吩咐带他们进宫的日子到了，太监长就把他们带到 尼布甲尼撒 面前。
DAN|1|19|王与他们谈论，在所有少年中找不到人能与 但以理 、 哈拿尼雅 、 米沙利 、 亚撒利雅 相比，于是他们就在王面前侍立。
DAN|1|20|王考问他们一切智慧和聪明的事，发现他们比全国所有的术士和巫师胜过十倍。
DAN|1|21|到 居鲁士 王元年， 但以理 还健在。
DAN|2|1|尼布甲尼撒 在位第二年，他做了很多梦，心里烦乱，不能睡觉。
DAN|2|2|王吩咐人将术士、巫师、行邪术的和 迦勒底 人召来，要他们把王的梦告诉王；他们就来，站在王面前。
DAN|2|3|王对他们说：“我做了一个梦，心里烦乱，想要知道这是什么梦。”
DAN|2|4|迦勒底 人用 亚兰 话对王说：“愿王万岁！请将梦告诉仆人，我们就可以讲解。”
DAN|2|5|王回答 迦勒底 人说：“这事我已决定，你们若不把梦和梦的解释告诉我，就必被凌迟，你们的房屋必成粪堆；
DAN|2|6|但你们若能说出这个梦和梦的解释，就必从我得到礼物、赏赐和殊荣。现在，你们要把梦和梦的解释告诉我。”
DAN|2|7|他们再一次回答说：“请王将梦告诉仆人，我们就可以讲解。”
DAN|2|8|王回答说：“我确实知道你们是故意拖延，因为你们知道这事我已决定。
DAN|2|9|你们若不将梦告诉我，只有一个办法对待你们；因为你们彼此串通，向我胡言乱语，要等候情势改变。现在，你们要将梦告诉我，让我知道你们真能为我解梦。”
DAN|2|10|迦勒底 人回答王说：“世上没有人能解释王的事情；从来没有君王、大臣、掌权者向术士、巫师，或 迦勒底 人问过这样的事。
DAN|2|11|王所问的事很难，除了不与血肉之躯同住的上帝，没有人能在王面前解释。”
DAN|2|12|王因这事生气，大大震怒，吩咐灭绝 巴比伦 所有的智慧人。
DAN|2|13|命令发出，智慧人将要被杀，人就寻找 但以理 和他的同伴，要杀他们。
DAN|2|14|王的护卫长 亚略 奉命去杀 巴比伦 的智慧人， 但以理 用婉言和智慧回应，
DAN|2|15|向王的大臣 亚略 说：“王的命令为何这样紧急呢？” 亚略 就把事情告诉 但以理 。
DAN|2|16|于是 但以理 进去求王宽限，好为王解梦。
DAN|2|17|但以理 回到他的居所，把这事告诉他的同伴 哈拿尼雅 、 米沙利 、 亚撒利雅 ，
DAN|2|18|要他们祈求天上的上帝施怜悯，将这奥秘指明，免得 但以理 和他的同伴与 巴比伦 其余的智慧人一同灭亡。
DAN|2|19|这奥秘就在夜间异象中显明给 但以理 ， 但以理 就称颂天上的上帝。
DAN|2|20|但以理 说： “上帝的名是应当称颂的，从亘古直到永远！ 因为智慧和能力都属乎他。
DAN|2|21|他改变时间、季节， 他废王，立王； 将智慧赐给智慧人， 将知识赐给聪明人。
DAN|2|22|他显明深奥隐秘的事， 洞悉幽暗中的一切， 光明也与他同住。
DAN|2|23|我列祖的上帝啊，我感谢你，赞美你， 因你将智慧才能赐给我， 我们所求问的现在你已指明给我， 把王的事给我们指明。”
DAN|2|24|于是， 但以理 进到王所派灭绝 巴比伦 智慧人的 亚略 那里去，对他这样说：“不要灭绝 巴比伦 的智慧人，求你领我到王面前，我可以为王解梦。”
DAN|2|25|亚略 就急忙领 但以理 到王面前，对王这样说：“我在被掳的 犹大 人中找到一人，能将梦的解释告诉王。”
DAN|2|26|王对那称为 伯提沙撒 的 但以理 说：“你能将我所做的梦和梦的解释告诉我吗？”
DAN|2|27|但以理 回答王说：“王所问的那奥秘，智慧人、巫师、术士、观兆的都不能告诉王，
DAN|2|28|只有那在天上的上帝能显明奥秘。他已把日后将要发生的事指示 尼布甲尼撒 王。你在床上做的梦和你脑中的异象是这样：
DAN|2|29|你，王啊，你在床上所思想的是关乎日后的事，那显明奥秘的主已把将来要发生的事指示你。
DAN|2|30|至于我，那奥秘显明给我，并非因我智慧胜过一切活着的人，而是为了让王知道梦的解释，知道你心里的意念。
DAN|2|31|“你，王啊，你正观看，看哪，有一个很大的像，这像甚高，极其光耀，立在你面前，形状非常可怕。
DAN|2|32|这像的头是纯金的，胸膛和膀臂是银的，腹部和腰是铜的，
DAN|2|33|腿是铁的，脚是半铁半泥的。
DAN|2|34|你正观看，见有一块非人手凿出来的石头打在它半铁半泥的脚上，把脚砸碎；
DAN|2|35|于是铁、泥、铜、银、金都一同砸得粉碎，如夏天禾场上的糠秕，被风吹散，无处可寻。打碎这像的石头成了一座大山，覆盖全地。
DAN|2|36|“这就是那梦；我们要在王面前讲解那梦。
DAN|2|37|你，王啊，你是诸王之王。天上的上帝已将国度、权势、能力、尊荣都赐给你。
DAN|2|38|世人和走兽，并天空的飞鸟，不论居住何处，他都交在你的手中，令你掌管这一切。你就是那金的头。
DAN|2|39|在你以后必兴起另一国，不及于你；又有第三国如铜，必掌管全地。
DAN|2|40|第四国必坚壮如铁，就像铁能打碎砸碎一切；铁怎样压碎一切，那国也必照样打碎压碎。
DAN|2|41|你既看见像的脚和脚趾头，一半是陶匠的泥，一半是铁，那国将来也必分裂。你既看见铁和泥搀杂，那国也必有铁的力量。
DAN|2|42|那脚趾头既是半铁半泥，那国也必半强半弱。
DAN|2|43|你既看见铁和泥搀杂，他们必有混杂的后裔，却不能彼此相合，正如铁和泥不能相合。
DAN|2|44|当诸王在位的时候，天上的上帝必另立一个永不败坏的国度，这国度必不归给其他百姓，却要打碎灭绝所有的国度，存立到永远。
DAN|2|45|你既看见非人手凿出来的一块石头从山而出，打碎铁、铜、泥、银、金，那就是至大的上帝把将来要发生的事给王指明。这梦是确实的，这解释也是准确的。”
DAN|2|46|当时， 尼布甲尼撒 王脸伏于地，向 但以理 下拜，并且吩咐人给他奉上供物和香。
DAN|2|47|王对 但以理 说：“你既能讲明这奥秘，你们的上帝诚然是万神之神、万王之主，是奥秘的启示者。”
DAN|2|48|于是王使 但以理 高升，赏赐他极多的礼物，派他管理 巴比伦 全省，又立他为总理，掌管 巴比伦 所有的智慧人。
DAN|2|49|但以理 求王，王就派 沙得拉 、 米煞 、 亚伯尼歌 管理 巴比伦 省的事务，只是 但以理 仍在朝中侍立。
DAN|3|1|尼布甲尼撒 王造了一个金像，高六十肘，宽六肘，立在 巴比伦 省的 杜拉 平原。
DAN|3|2|尼布甲尼撒 王差人将总督、钦差、省长、参谋、财务、法官、地方官和各省的官员都召了来，为 尼布甲尼撒 王所立的像行开光礼。
DAN|3|3|于是总督、钦差、省长、参谋、财务、法官、地方官和各省的官员都聚集，站在 尼布甲尼撒 所立的像前，要为 尼布甲尼撒 王所立的像行开光礼。
DAN|3|4|那时传令的大声呼叫说：“各方、各国、各族 的人哪，有命令传给你们：
DAN|3|5|你们一听见角、号、琴、瑟、三角琴、鼓和各样乐器的声音，就当俯伏，拜 尼布甲尼撒 王所立的金像。
DAN|3|6|凡不俯伏下拜的，必立刻扔在烈火的窑中。”
DAN|3|7|因此百姓一听见角、号、琴、瑟、三角琴 和各样乐器的声音，各方、各国、各族的人就都俯伏，拜 尼布甲尼撒 王所立的金像。
DAN|3|8|在那时，有几个 迦勒底 人进前来控告 犹大 人。
DAN|3|9|他们对 尼布甲尼撒 王说：“愿王万岁！
DAN|3|10|你，王啊，你曾降旨，凡听见角、号、琴、瑟、三角琴、鼓和各样乐器声音的，都当俯伏拜这金像。
DAN|3|11|凡不俯伏下拜的，必扔在烈火的窑中。
DAN|3|12|现在有几个 犹大 人，就是王所派管理 巴比伦 省事务的 沙得拉 、 米煞 、 亚伯尼歌 ；王啊，这些人不理你的谕旨，不事奉你的神明，也不拜你所立的金像。”
DAN|3|13|当时， 尼布甲尼撒 大发烈怒，命令把 沙得拉 、 米煞 、 亚伯尼歌 带过来；他们就把这几个人带到王面前。
DAN|3|14|尼布甲尼撒 对他们说：“ 沙得拉 、 米煞 、 亚伯尼歌 ，你们不事奉我的神明，不拜我所立的金像，是真的吗？
DAN|3|15|现在，你们若准备好，一听见角、号、琴、瑟、三角琴、鼓和各样乐器的声音，就俯伏拜我所造的像；若不下拜，必立刻扔在烈火的窑中，有哪一个神明能救你们脱离我的手呢？”
DAN|3|16|沙得拉 、 米煞 、 亚伯尼歌 对王说：“ 尼布甲尼撒 啊，这件事我们不必回答你，
DAN|3|17|即便如此，我们所事奉的上帝能将我们从烈火的窑中救出来。王啊，他必救我们脱离你的手；
DAN|3|18|即或不然，王啊，你当知道，我们绝不事奉你的神明，也不拜你所立的金像。”
DAN|3|19|当时， 尼布甲尼撒 怒气填胸，向 沙得拉 、 米煞 、 亚伯尼歌 变了脸色，命令把窑烧热，比平常热七倍；
DAN|3|20|又命令他军中的几个壮士，把 沙得拉 、 米煞 、 亚伯尼歌 捆起来，扔在烈火的窑中。
DAN|3|21|这三人穿着内袍、外衣、头巾和其他的衣服，被捆起来扔在烈火的窑中。
DAN|3|22|因为王的命令紧急，窑又非常热，那抬 沙得拉 、 米煞 、 亚伯尼歌 的人都被火焰烧死。
DAN|3|23|但是这三个人， 沙得拉 、 米煞 、 亚伯尼歌 被捆绑着，掉进烈火的窑中。
DAN|3|24|那时， 尼布甲尼撒 王惊奇，急忙站起来，对谋士说：“我们捆起来扔在火里的不是三个人吗？”他们回答王说：“王啊，是的。”
DAN|3|25|王说：“看哪，我看见有四个人，并没有捆绑，在火中行走，也没有受伤；那第四个的相貌好像神明的儿子。”
DAN|3|26|于是 尼布甲尼撒 靠近烈火窑门，说：“至高上帝的仆人 沙得拉 、 米煞 、 亚伯尼歌 ，出来，来吧！” 沙得拉 、 米煞 、 亚伯尼歌 就从火中出来。
DAN|3|27|那些总督、钦差、省长和王的谋士一同聚集来看这三个人，见火不能伤他们的身体，头发没有烧焦，衣裳也没有变色，都没有火烧过的气味。
DAN|3|28|尼布甲尼撒 说：“ 沙得拉 、 米煞 、 亚伯尼歌 的上帝是应当称颂的！他差遣使者救护倚靠他的仆人，他们不遵王的命令，甚至舍身，在他们上帝以外不肯事奉敬拜别神。
DAN|3|29|现在我降旨，无论何方、何国、何族，凡有人毁谤 沙得拉 、 米煞 、 亚伯尼歌 的上帝，他必被凌迟，他的房屋必成粪堆，因为没有别神能像这样施行拯救。”
DAN|3|30|那时王在 巴比伦 省使 沙得拉 、 米煞 、 亚伯尼歌 高升。
DAN|4|1|尼布甲尼撒 王对住在全地各方、各国、各族的人说：“愿你们大享平安！
DAN|4|2|我乐意宣扬至高上帝向我所行的神迹奇事。
DAN|4|3|他的神迹何其大！ 他的奇事何其盛！ 他的国度存到永远； 他的权柄存到万代！
DAN|4|4|“我－ 尼布甲尼撒 安居在家中，在宫里享受荣华。
DAN|4|5|我做了一个梦，使我惧怕。我在床上的意念和脑中的异象，使我惊惶。
DAN|4|6|因此我降旨召 巴比伦 的智慧人全都到我面前，要他们将梦的解释告诉我。
DAN|4|7|于是那些术士、巫师、 迦勒底 人、观兆的都进来，我将那梦告诉他们，他们却不能把梦的解释告诉我。
DAN|4|8|最后， 但以理 ，就是按照我神明的名字称为 伯提沙撒 的，来到我面前，他里头有神圣神明的灵，我将梦告诉他：
DAN|4|9|‘术士的领袖 伯提沙撒 啊，我知道你里头有神圣神明的灵，什么奥秘都不能为难你。现在你要把我梦中所见的异象和梦的解释告诉我 。’
DAN|4|10|“我在床上脑中的异象是这样：我观看，看哪，大地中间有一棵树，极其高大。
DAN|4|11|那树渐长，而且茁壮，高得顶天，从地极都能看见，
DAN|4|12|叶子华美，果子甚多，可作所有动物的食物；野地的走兽卧在荫下，天空的飞鸟宿在枝上，凡有血肉的都从这树得食物。
DAN|4|13|“我观看，我在床上脑中的异象是这样，看哪，有守望者，就是神圣的一位，从天而降，
DAN|4|14|大声呼叫说：‘砍倒这树！砍下枝子！拔掉叶子！抛散果子！使走兽逃离树下，飞鸟躲开树枝。
DAN|4|15|树的残干却要留在地里，在田野的青草中用铁圈和铜圈套住。任他让天上的露水滴湿，和地上的走兽一同吃草，
DAN|4|16|使他的心改变，不再是人的心，而给他一个兽心，使他经过七个时期 。
DAN|4|17|这是众守望者所发的命令，是众圣者所作的决定，好叫世人知道至高者在人的国中掌权，要将国赐给谁就赐给谁，并且立极卑微的人执掌国权。’
DAN|4|18|“这是我－ 尼布甲尼撒 王所做的梦。 伯提沙撒 啊，你要说明这梦的解释；我国中所有的智慧人都不能把梦的解释告诉我，惟独你能，因你里头有神圣神明的灵。”
DAN|4|19|于是称为 伯提沙撒 的 但以理 惊骇片时，心意惊惶。王说：“ 伯提沙撒 啊，不要因梦和梦的解释惊惶。” 伯提沙撒 回答说：“我主啊，愿这梦归给恨恶你的人，这梦的解释归给你的敌人。
DAN|4|20|你所见的树渐长，而且茁壮，高得顶天，全地都能看见，
DAN|4|21|叶子华美，果子甚多，可作所有动物的食物；野地的走兽住在其下，天空的飞鸟宿在枝上。
DAN|4|22|“王啊，这成长又茁壮的树就是你。你的威势成长及于天，你的权柄达到地极。
DAN|4|23|王既看见一位神圣的守望者从天而降，说：‘将这树砍倒毁坏，树的残干却要留在地里，在田野的青草中用铁圈和铜圈套住。任他让天上的露水滴湿，与野地的走兽一同吃草，直到经过七个时期。’
DAN|4|24|“王啊，梦的解释就是这样：临到我主我王的事是出于至高者的命令。
DAN|4|25|你必被赶出离开世人，与野地的走兽同住，吃草如牛，让天上的露水滴湿，且要经过七个时期，直等到你知道至高者在人的国中掌权，要将国赐给谁就赐给谁。
DAN|4|26|这使树的残干存留的命令，是要等你知道天在掌权，你的国必定归你。
DAN|4|27|王啊，求你悦纳我的谏言，以施行公义除去罪过，以怜悯穷人除掉罪恶，或者你的平安可以延长。”
DAN|4|28|这些事都临到 尼布甲尼撒 王。
DAN|4|29|过了十二个月，他在 巴比伦 王宫顶上散步。
DAN|4|30|王说：“这大 巴比伦 岂不是我用大能大力建为首都，要显示我威严的荣耀吗？”
DAN|4|31|这话还在王口中的时候，有声音从天降下，说：“ 尼布甲尼撒 王啊，有话对你说，你的国离开你了。
DAN|4|32|你必被赶出离开世人，与野地的走兽同住，吃草如牛，且要经过七个时期；等你知道至高者在人的国中掌权，要将国赐给谁就赐给谁。”
DAN|4|33|当时这话就应验在 尼布甲尼撒 身上，他被赶出离开世人，吃草如牛，身体被天上的露水滴湿，头发长得像鹰的羽毛，指甲长得像鸟爪。
DAN|4|34|“时候到了，我－ 尼布甲尼撒 举目望天，我的知识复归于我，我就称颂至高者，赞美尊敬活到永远的上帝。 他的权柄存到永远， 他的国度存到万代。
DAN|4|35|地上所有的居民都算为虚无； 在天上万军和地上居民中， 他都凭自己的旨意行事。 无人能拦住他的手， 或问他说，你在做什么呢？
DAN|4|36|“那时，我的知识复归于我，威严和光荣也复归于我，使我的国度得荣耀，我的谋士和大臣也来朝见我。我又重建我的国度，更大的权势加添在我身上。
DAN|4|37|现在我－ 尼布甲尼撒 赞美、尊崇、恭敬天上的王，因为他所行的全都信实，他所做的尽都公平。那行事骄傲的，他能降为卑。”
DAN|5|1|伯沙撒 王为他的一千大臣摆设盛筵，与这一千人饮酒。
DAN|5|2|伯沙撒 在欢饮之间，吩咐人将他父 尼布甲尼撒 从 耶路撒冷 圣殿所掳掠的金银器皿拿来，好使王与大臣、王后、妃嫔用这器皿饮酒。
DAN|5|3|于是他们把圣殿，就是 耶路撒冷 上帝殿中所掳掠的金器皿拿来，王和大臣、王后、妃嫔就用这器皿饮酒。
DAN|5|4|他们饮酒，赞美金、银、铜、铁、木、石造的神明。
DAN|5|5|当时，忽然有人的指头出现，在灯台对面王宫粉刷的墙上写字。王看见写字的指头，
DAN|5|6|就变了脸色，心意惊惶，腰骨好像脱节，双膝彼此相碰，
DAN|5|7|大声吩咐将巫师、 迦勒底 人和观兆的领进来。王对 巴比伦 的智慧人说：“谁能读这文字，并且向我讲解它的意思，他必身穿紫袍，项带金链，在我国中位列第三。”
DAN|5|8|于是王所有的智慧人都进前来，他们却不能读那文字，也不能为王讲解它的意思。
DAN|5|9|伯沙撒 王就甚惊惶，脸色改变，他的大臣也都困惑。
DAN|5|10|太后 因王和他大臣所说的话，就进入宴会厅，说：“愿王万岁！你的心不要惊惶，脸不要变色。
DAN|5|11|在你国中有一人，他里头有神圣神明的灵，你父在世的日子，这人心中光明，又有聪明智慧，好像神明的智慧。你父 尼布甲尼撒 王，就是王的父，曾立他为术士、巫师、 迦勒底 人和观兆者的领袖，
DAN|5|12|都因他有美好的灵性，又有知识聪明，能解梦，释谜语，解疑惑。这人名叫 但以理 ， 尼布甲尼撒 王又称他为 伯提沙撒 ，现在可以召他来，他必解明这意思。”
DAN|5|13|于是 但以理 被领到王面前。王问 但以理 说：“你就是我父王从 犹大 带来、被掳的 犹大 人 但以理 吗？
DAN|5|14|我听说你里头有神明的灵，心中有光，又有聪明和高超的智慧。
DAN|5|15|现在智慧人和巫师都被带到我面前，要叫他们读这文字，为我讲解它的意思；无奈他们都不能讲解它的意思。
DAN|5|16|我听说你能讲解，能解疑惑；现在你若能读这文字，为我讲解它的意思，就必身穿紫袍，项戴金链，在我国中位列第三。”
DAN|5|17|但以理 回答王说：“你的礼物可以归你自己，你的赏赐可以归给别人；我却要为王读这文字，讲解它的意思。
DAN|5|18|你，王啊，至高的上帝曾将国度、大权、荣耀、威严赐给你父 尼布甲尼撒 ；
DAN|5|19|因上帝所赐给他的大权，各方、各国、各族的人都在他面前恐惧战兢，因他要杀就杀，要人活就活，要升就升，要降就降。
DAN|5|20|但他的心高傲，灵也刚愎，以致行事狂傲，就被革去国度的王位，夺走荣耀。
DAN|5|21|他被赶出离开世人，他的心变为兽心，与野驴同住，吃草如牛，身体被天上的露水滴湿，直到他知道，至高的上帝在人的国中掌权，凭自己的旨意立人治国。
DAN|5|22|伯沙撒 啊，你是他的儿子 ，你虽知道这一切，却不谦卑自己，
DAN|5|23|竟向天上的主自高，差人将他殿中的器皿拿到你面前，你和大臣、王后、妃嫔用这器皿饮酒。你又赞美那不能看、不能听、无知无识，用金、银、铜、铁、木、石造的神明，没有将荣耀归与那手中掌管你气息，管理你一切行动的上帝。
DAN|5|24|于是从他那里显出指头写这文字。
DAN|5|25|“所写的文字是：‘弥尼，弥尼，提客勒，乌法珥新 。’
DAN|5|26|解释是这样：弥尼就是上帝数算你国的年日到此完毕。
DAN|5|27|提客勒就是你被秤在天平上，秤出你的亏欠来。
DAN|5|28|毗勒斯 就是你的国要分裂，归给 玛代 人和 波斯 人。”
DAN|5|29|于是 伯沙撒 下令，人就把紫袍给 但以理 穿上，把金链给他戴在颈项上，又传令使他在国中位列第三。
DAN|5|30|当夜， 迦勒底 王 伯沙撒 被杀。
DAN|5|31|玛代 人 大流士 年六十二岁，取了 迦勒底 国。
DAN|6|1|大流士 随心所愿，立了一百二十个总督，治理全国，
DAN|6|2|又在他们以上立总长三人， 但以理 也在其中；使总督在他们三人面前呈报，免得王受亏损。
DAN|6|3|这 但以理 因有卓越的灵性，超乎其余的总长和总督，王想立他治理全国。
DAN|6|4|那时，总长和总督在治国的事务上寻找 但以理 的把柄，为要控告他；只是找不到任何的把柄和过失，因他忠心办事，毫无错误过失。
DAN|6|5|那些人就说：“我们要找 但以理 的把柄，若不从他上帝的律法中下手，就寻不着。”
DAN|6|6|于是，总长和总督纷纷聚集来见王，说：“ 大流士 王万岁！
DAN|6|7|国中的总长、钦差、总督、谋士和省长彼此商议，求王下旨，立一条禁令，三十天之内，不拘何人，若在王以外，或向神明或向人求什么，就必扔在狮子坑中。
DAN|6|8|王啊，现在求你立这禁令，在这文件上签署，使它不能更改；照 玛代 人和 波斯 人的例，绝不更动。”
DAN|6|9|于是 大流士 王在这禁令的文件上签署。
DAN|6|10|但以理 知道这文件已经签署，就进自己的家，他家楼上的窗户开向 耶路撒冷 。他一天三次，双膝跪着，在他的上帝面前祷告感谢，像平常一样。
DAN|6|11|于是，那些人纷纷聚集，发现 但以理 在他上帝面前祈祷恳求。
DAN|6|12|他们就进到王面前，向王提及禁令，说：“三十天之内不拘何人，若在王以外，或向神明或向人求什么，必被扔在狮子坑中，王不是在这禁令上签署了吗？”王回答说：“确有这事，照 玛代 人和 波斯 人的例是不可更改的。”
DAN|6|13|他们对王说：“王啊，那被掳的 犹大 人 但以理 不理会你，也不遵守你签署的禁令，竟一天三次祈祷。”
DAN|6|14|王听见这话，就甚愁烦，一心要救 但以理 ，直到日落的时候，他还在筹划解救他。
DAN|6|15|那些人就纷纷聚集到王那里，对王说：“王啊，当知道 玛代 人和 波斯 人有例，凡王所立的禁令和律例都不可更改。”
DAN|6|16|于是王下令，人就把 但以理 带来，扔在狮子坑中。王对 但以理 说：“你经常事奉的上帝，他必拯救你。”
DAN|6|17|有人搬来一块石头放在坑口，王用自己的玺和大臣的印，封闭那坑，使惩办 但以理 的事绝不更改。
DAN|6|18|王回到宫里，终夜禁食，不让人带乐器 到他面前，他也失眠了。
DAN|6|19|次日黎明，王起来，急忙往狮子坑那里去，
DAN|6|20|临近坑边，哀声呼叫 但以理 。王对 但以理 说：“永生上帝的仆人 但以理 啊，你经常事奉的上帝能救你脱离狮子吗？”
DAN|6|21|但以理 对王说：“愿王万岁！
DAN|6|22|我的上帝差遣使者封住狮子的口，叫狮子不伤我，因我在上帝面前无辜。王啊，在你面前我也没有做过任何亏损的事。”
DAN|6|23|王因此就甚喜乐，吩咐把 但以理 从坑里拉上来。于是 但以理 从坑里被拉上来，身上毫无损伤，因为他信靠他的上帝。
DAN|6|24|王下令，把那些控告 但以理 的人和他们的妻子儿女都带来，扔在狮子坑中。他们还没有到坑底，狮子就制伏他们，咬碎他们的骨头。
DAN|6|25|于是， 大流士 王传旨给住在全地各方、各国、各族的人说：“愿你们大享平安！
DAN|6|26|现在我降旨，我所统辖全国的人民，都要在 但以理 的上帝面前战兢畏惧。 因为他是活的上帝， 永远长存， 他的国度永不败坏， 他的权柄永存无极！
DAN|6|27|他庇护，搭救， 在天上地下施行神迹奇事， 救了 但以理 脱离狮子的口。”
DAN|6|28|如此，这 但以理 ，当 大流士 在位的时候和 波斯 的 居鲁士 在位的时候，大享亨通。
DAN|7|1|巴比伦 王 伯沙撒 元年， 但以理 在床上做梦，脑中看见异象，就记录这梦，述说其中的大意。
DAN|7|2|但以理 说： 我在夜间的异象中观看，看哪，天上四风，突然刮在大海之上。
DAN|7|3|有四只巨兽从海里上来，它们各不相同：
DAN|7|4|头一个像狮子，有鹰的翅膀；我正观看的时候，它的翅膀被拔去，它从地上被扶起来，用两脚站立，像人一样，还给了它人的心。
DAN|7|5|看哪，另有一兽如熊，就是第二兽，半身侧立，口里的牙齿中有三根獠牙 。有人吩咐这兽说：“起来，吞吃许多的肉。”
DAN|7|6|其后，我观看，看哪，另有一兽如豹，背上有四个鸟的翅膀；这兽有四个头，还给了它权柄。
DAN|7|7|其后，我在夜间的异象中观看，看哪，第四兽可怕可惧，极其强壮，有大铁牙，吞吃嚼碎，剩下的用脚践踏。这兽与前面所有的兽不同，它有十只角。
DAN|7|8|我正思考这些角的时候，看哪，其中又长出另一只小角；先前的角中有三只角在它面前连根被拔出。看哪，这角有眼，像人的眼，有口说夸大的话。
DAN|7|9|我正观看的时候， 有宝座设立， 上面坐着亘古常在者。 他的衣服洁白如雪， 头发如纯净的羊毛。 宝座是火焰， 其轮为烈火。
DAN|7|10|有火如河涌出， 从他面前流出来； 事奉他的有千千， 在他面前侍立的有万万； 他坐着要行审判 ， 案卷都展开了。
DAN|7|11|于是我观看，因这角说夸大的话，我正观看的时候，那兽被杀，身体被毁，扔在火中焚烧。
DAN|7|12|其余的兽，权柄都被夺去，生命却得以延续，直到所定的时候和日期。
DAN|7|13|我在夜间的异象中观看， 看哪，有一位像人子的， 驾着天上的云而来， 被领到亘古常在者面前。
DAN|7|14|他得了权柄、荣耀、国度， 使各方、各国、各族的人都事奉他。 他的权柄是永远的，不能废去， 他的国度必不败坏。
DAN|7|15|至于我－ 但以理 ，我的灵在我里面忧伤，我脑中的异象使我惊惶。
DAN|7|16|我走近其中一位侍立者，问他这一切的实情。他就告诉我，使我知道这事的解释：
DAN|7|17|这四只巨兽就是将要在世上兴起的四个王 。
DAN|7|18|然而，至高者的众圣者必要得到这国度，并且拥有它，直到永远，永永远远。
DAN|7|19|于是我想要更清楚知道第四兽的实情，它与一切的兽不同，甚是可怕，有铁牙铜爪，吞吃嚼碎，剩下的用脚践踏；
DAN|7|20|头上有十只角和那另长出的一角，三只角在这角面前掉落；这角有眼，有口说夸大的话，形状比它的同类更强。
DAN|7|21|我观看，这角与众圣者争战，胜了他们，
DAN|7|22|直到亘古常在者来到，为至高者的众圣者伸冤，众圣者得到国度的时候就到了。
DAN|7|23|那侍立者这样说： 第四兽就是世上要兴起的第四国， 与其他各国不同， 它要并吞全地， 并且践踏嚼碎。
DAN|7|24|至于那十只角，就是从这国中兴起的十个王； 后来又兴起另一王， 与先前的不相同， 他要制伏三个王。
DAN|7|25|他说话抵挡至高者， 折磨至高者的众圣者， 又改变节期和律法。 众圣者要交在他手中一年 、两年、又半年。
DAN|7|26|然而，他坐着要行审判； 他的权柄要被夺去， 毁坏，灭绝，一直到底。
DAN|7|27|国度、权柄和天下诸国的大权 必赐给至高者的众圣民。 他的国是永远的国， 所有掌权的都必事奉他，顺从他。
DAN|7|28|这事到此结束。我－ 但以理 因这些念头甚是惊惶，脸色也变了，却将这事记在心里。
DAN|8|1|伯沙撒 王在位第三年，有异象向我－ 但以理 显现，是在先前所见的异象之后。
DAN|8|2|我在异象中观看，见自己在 以拦 省 书珊 的城堡中；我在异象中又见自己在 乌莱河 边。
DAN|8|3|我举目观看，看哪，有一只公绵羊站在河边，它有两只角，这两角都高，一角高过另一角，后长出来的比较高。
DAN|8|4|我见那公绵羊向西、向北、向南抵撞，没有任何兽在它面前站立得住，没有能逃脱它手的；它任意而行，自高自大。
DAN|8|5|我正思想的时候，看哪，有一只公山羊从西而来，遍行全地，脚不着地。这山羊两眼当中有一只显眼的角。
DAN|8|6|它往我先前所见、站在河边、有双角的公绵羊那里，以猛烈的怒气向它直闯。
DAN|8|7|我见公山羊靠近公绵羊，向它发怒，攻击它，折断它的两角。公绵羊在公山羊面前站立不住；它把公绵羊撞倒在地，用脚践踏，没有能救公绵羊脱离它手的。
DAN|8|8|这公山羊长得极其高大，正强壮的时候，那大角折断了，从角的下面向天的四方 长出四只显眼的角来。
DAN|8|9|从四角中的一角又长出另一只小角，向南、向东、向佳美之地，日渐壮大。
DAN|8|10|它渐壮大，高及诸天万象，把一些天象和星辰摔落在地，用脚践踏。
DAN|8|11|它自高自大 ，自以为高及万象之君，它除掉经常献给君的祭，毁坏君的圣所。
DAN|8|12|因罪过的缘故，有军队和经常献的祭交给它。它把真理抛在地上，任意而行 ，无往不利。
DAN|8|13|我听见有一位圣者说话，又有一位圣者向那说话的圣者说：“这经常献的祭、带来荒凉的罪过、圣所与军队被践踏的异象，要持续到几时呢？”
DAN|8|14|他对我 说：“要到二千三百日，圣所就必洁净 。”
DAN|8|15|我－ 但以理 见了这异象，想要明白其中的意思。看哪，有一位形状像人的站在我面前。
DAN|8|16|我听见 乌莱河 中有人声呼叫说：“ 加百列 啊，要使这人明白这异象。”
DAN|8|17|他就来到我所站的地方。他一来，我就惊慌，脸伏于地。他对我说：“人子啊，你要明白，因为这是关乎末后时期的异象。”
DAN|8|18|他对我说话的时候，我正沉睡，脸伏于地。他就摸我，扶我站起来。
DAN|8|19|他说：“看哪，我要指示你恼怒结束的时候必成的事，因为这是关乎末后指定的时期。
DAN|8|20|你所看见那有双角的公绵羊就是 玛代 王和 波斯 王。
DAN|8|21|那公山羊就是 希腊 王；两眼当中的大角就是第一个王。
DAN|8|22|至于角折断了，又从角的下面长出四只角，意思就是有四个国要从这国兴起，只是权势都不及它。
DAN|8|23|这四国末期，恶贯满盈的时候，必有一王兴起，面貌凶恶，诡计多端。
DAN|8|24|他的权柄极大，却不是因自己的能力；他要施行惊人的毁灭，无往不利，任意而行，又要毁灭强有力的人和众圣民。
DAN|8|25|他用权术使手中的诡计成功；他的心自高自大，趁人无备的时候毁灭多人。他又起来攻击万君之君，至终却非因人的手而遭毁灭。
DAN|8|26|所说二千三百日 的异象是真的，但你要将这异象封住，因为它关乎未来许多的日子。”
DAN|8|27|于是我－ 但以理 昏倒，病了数日，然后起来办理王的事务。我因这异象惊骇不已，但还是不能了解。
DAN|9|1|玛代 族 亚哈随鲁 的儿子 大流士 被立为王，统治 迦勒底 国元年，
DAN|9|2|就是他在位第一年，我－ 但以理 从书上得知，耶和华的话临到 耶利米 先知，论 耶路撒冷 荒凉期满的年数为七十年。
DAN|9|3|我面向主上帝，禁食，披麻蒙灰，恳切祷告祈求。
DAN|9|4|我向耶和华－我的上帝祈祷、认罪，说：“主啊，你是大而可畏的上帝，向爱主、守主诫命的人守约施慈爱。
DAN|9|5|我们犯罪作恶，行恶叛逆，偏离你的诫命典章，
DAN|9|6|没有听从你仆人众先知奉你的名向我们君王、官长、祖先和这地所有百姓所说的话。
DAN|9|7|主啊，你是公义的，但我们 犹大 人和 耶路撒冷 的居民，并你所赶到各国的 以色列 众人，不论远近，因为背叛了你，脸上蒙羞，正如今日一样。
DAN|9|8|耶和华啊，我们和我们的君王、官长、祖先因得罪了你，脸上就都蒙羞。
DAN|9|9|主－我们的上帝是怜悯饶恕人的，我们却违背了他，
DAN|9|10|没有听从耶和华－我们上帝的话，没有遵行他藉仆人众先知向我们颁布的律法。
DAN|9|11|以色列 众人都犯了你的律法，偏离、不听从你的话；因此，你仆人 摩西 律法上所写的诅咒和誓言倾倒在我们身上，因我们得罪了上帝。
DAN|9|12|上帝使大灾祸临到我们，实现了警戒我们和审判我们官长的话；原来 耶路撒冷 所遭遇的灾祸是普天之下未曾有过的。
DAN|9|13|这一切灾祸临到我们，是照 摩西 律法上所写的，我们却没有求耶和华－我们上帝的恩惠，使我们回转离开罪孽，明白你的真理。
DAN|9|14|所以耶和华特意使这灾祸临到我们，耶和华－我们的上帝在他所行的事上都是公义的；我们并没有听从他的话。
DAN|9|15|主－我们的上帝啊，你曾用大能的手领你的子民出 埃及 地，使自己得了名声，正如今日一样，现在，我们犯了罪，作了恶。
DAN|9|16|主啊，求你按你丰盛的公义，使你的怒气和愤怒转离你的城 耶路撒冷 ，就是你的圣山。因我们的罪恶和我们祖先的罪孽， 耶路撒冷 和你的子民被四围的人羞辱。
DAN|9|17|我们的上帝啊，现在求你垂听你仆人的祈祷恳求，为你自己的缘故使你的脸向荒凉的圣所发光。
DAN|9|18|我的上帝啊，求你侧耳而听，睁眼而看，眷顾我们那荒凉之地和称为你名下的城。我们在你面前恳求，不是因自己的义，而是因你丰富的怜悯。
DAN|9|19|主啊，求你垂听！主啊，求你赦免！主啊，求你侧耳，求你实行！为你自己的缘故不要迟延。我的上帝啊，因这城和这民都是称为你名下的。”
DAN|9|20|我正说话、祷告，承认我的罪和我百姓 以色列 的罪，为我上帝的圣山，在耶和华－我的上帝面前恳求；
DAN|9|21|我正在祷告中说话，先前在异象中所见的那位 加百列 ，约在献晚祭的时候迅速飞到我这里来。
DAN|9|22|他指教我说 ：“ 但以理 啊，现在我来要使你有智慧，有聪明。
DAN|9|23|你刚开始恳求的时候，就有命令发出。现在我来告诉你，因你是蒙爱的；所以你要思想这事，明白这异象。
DAN|9|24|“为你百姓和你圣城，已经定了七十个七，要止住罪过，除净罪恶，赎尽罪孽，引进永恒的公义，封住异象和预言，并膏至圣所 。
DAN|9|25|你当知道，当明白，从发出命令恢复并重建 耶路撒冷 ，直到受膏的君出现，必有七个七和六十二个七。 耶路撒冷城 连街带濠都必在艰难中恢复并重建。
DAN|9|26|过了六十二个七，那受膏者 被剪除，一无所有；必有一王的百姓来毁灭这城和圣所，它的结局 必如洪水冲没。必有战争，一直到末了，荒凉的事已经定了。
DAN|9|27|在一七之期，他必与许多人坚立盟约；一七之半，他必使献祭与供献止息。那施行毁灭的可憎之物必立在圣殿里 ，直到所定的结局倾倒在那行毁灭者的身上。”
DAN|10|1|波斯 王 居鲁士 第三年，有话指示那称为 伯提沙撒 的 但以理 。这话是确实的，指着大战争； 但以理 明白这话，明白这异象。
DAN|10|2|那时，我－ 但以理 悲伤了三个七日；
DAN|10|3|美味我没有吃，酒和肉没有入我的口，也没有用油抹我的身，直到满了三个七日。
DAN|10|4|正月二十四日，我在 大河 ，就是 底格里斯河 边，
DAN|10|5|举目观看，看哪，有一人身穿细麻衣，腰束 乌法 的纯金腰带。
DAN|10|6|他的身体如水苍玉，面貌如闪电，眼目如火把，手臂和脚如明亮的铜，说话的声音像众人的声音。
DAN|10|7|我－ 但以理 一人看见这异象，跟我一起的人没有看见，却有极大的战兢落在他们身上，他们就逃跑躲避，
DAN|10|8|只剩下我一人。我看见这大异象就浑身无力，面容变色，毫无气力。
DAN|10|9|我听见他说话的声音；一听见他说话的声音，我就沉睡，脸伏于地。
DAN|10|10|看哪，有一只手摸我，使我膝盖和手掌战抖。
DAN|10|11|他对我说：“蒙爱的 但以理 啊，要思想我对你所说的话，只管站起来，因为我现在奉差遣来到你这里。”他对我说这话，我就战战兢兢地站起来。
DAN|10|12|他说：“ 但以理 啊，不要惧怕！因为自从第一日你立志要明白，又在你上帝面前刻苦自己，你的话已蒙应允；我就是因你的话而来。
DAN|10|13|但 波斯 国的领袖拦阻了我二十一天。看哪，天使长 中的一位 米迦勒 来帮助我，因为我被留在 波斯 诸王那里。
DAN|10|14|现在我来，要使你明白你百姓日后必遭遇的事，因为这异象关乎未来的日子。”
DAN|10|15|他向我这样说，我就脸面朝地，哑口无声。
DAN|10|16|看哪，有一位形状像人的，摸我的嘴唇，我就开口说话，向那站在我面前的说：“我主啊，因这异象使我感到剧痛，毫无气力。
DAN|10|17|我主的仆人怎能跟我主说话呢？我现在浑身无力，毫无气息。”
DAN|10|18|有一位形状像人的再一次摸我，使我有力量。
DAN|10|19|他说：“蒙爱的人哪，不要惧怕，愿你平安！你要刚强！要刚强！ ”他一对我说话，我就觉得有力量，说：“我主请说，因你使我有力量。”
DAN|10|20|他说：“你知道我为什么到你这里来吗？现在我要回去与 波斯 的领袖争战，我去了之后，看哪， 希腊 的领袖必来。
DAN|10|21|但我要将那记录在真理之书上的话告诉你。除了你们的天使 米迦勒 之外，没有人帮助我抵挡他们。”
DAN|11|1|“至于我，当 玛代 的 大流士 元年，我曾起来扶助 米迦勒 ，使他坚强。
DAN|11|2|现在我要指示你确实的事。” “看哪， 波斯 还有三个王要兴起，第四王必富足远胜诸王。他因富足成为强盛，就煽动各国攻击 希腊 国。
DAN|11|3|必有一个勇敢的王兴起，执掌大权，随意而行。
DAN|11|4|他正兴起的时候，他的国必瓦解，向天的四方 裂开，却不归他的后裔，也不如他当年统治的权威；他的国必被拔出，归给他后裔之外的人。
DAN|11|5|“南方的王必强盛，他的将帅中必有一个比他更强，执掌权柄，权柄甚大。
DAN|11|6|过了几年，他们必结盟，南方王的女儿必来到北方王那里，使约生效；但这女子不能保留实力，王的力量 也未能存留。这女子、带她来的、生她的 和当时扶助她的必被杀害 。
DAN|11|7|但从这女子的本家必另有一子 接续王位，他要率领军队进入北方王的堡垒，攻击他们，而且得胜，
DAN|11|8|把他们的神像和铸成的偶像，与金银宝器都掳掠到 埃及 去。数年之内，他不去攻击北方的王。
DAN|11|9|北方的王必侵入南方王的国土，但却要撤回本地。
DAN|11|10|“北方王的儿子们必动干戈，招聚许多军兵。他要前进，如洪水泛滥；要再度争战，直捣南方王的堡垒。
DAN|11|11|南方王必发烈怒，出来与北方王争战，摆列大军；北方王的军兵必败在南方王的手下。
DAN|11|12|这大军既被扫荡，南方王的心就自高；他虽使万人仆倒，却不能保持胜利。
DAN|11|13|“北方王要再度摆列大军，比先前更多。过了几年，他必率领大军，带极多的装备而来。
DAN|11|14|那时，必有许多人起来攻击南方王，并且你百姓中的残暴人要兴起，应验异象，他们却要败亡。
DAN|11|15|北方王必来建土堆攻取坚固城，南方的军兵抵挡不住，就是精选的部队也无力抵挡；
DAN|11|16|前来攻击南方王的必任意而行，无人在北方王面前站立得住。他要站在那佳美之地，用手施行毁灭。
DAN|11|17|“他必定意倾全国之力而来，与南方王订约，把自己的女儿 给南方王为妻，企图败坏他的国度。这计谋却未得逞，自己也得不到好处。
DAN|11|18|其后北方王必转头，夺取许多海岛。但有一将帅除掉北方王对人的羞辱，并且使羞辱归到他自己身上。
DAN|11|19|他必转头回到本地的堡垒，却要绊跌仆倒，归于无有。
DAN|11|20|“那时，有一人兴起接续他的王位，他为了王国的荣华，差官员横征暴敛。这王过不多时就死了，不是因怒气 ，也不是因战役。”
DAN|11|21|“后来，有一个卑鄙的人兴起接续他的王位，人未曾将国的尊荣给他，他却趁人无备的时候前来，用诡诈夺取政权。
DAN|11|22|势如洪水般的军兵在他面前被冲没，遭击溃；立约的领袖也是如此。
DAN|11|23|他与人结盟之后，却行诡诈。跟随他的人虽不多，他却日渐强盛。
DAN|11|24|他趁人无备的时候，来到国中极肥沃之地，做他祖宗和祖宗的祖宗未曾做过的事，瓜分掳物、掠物和财宝，又策划进攻堡垒；然而这都是暂时的。
DAN|11|25|“他必奋勇向前，率领大军攻击南方王；南方王以极强的大军迎战，却抵挡不住，因为有人设计谋害南方王。
DAN|11|26|吃王饷的使王败坏，王的军队必被冲没，仆倒被杀的甚多。
DAN|11|27|至于这二王，他们心怀恶计，同席吃饭却彼此说谎，但计谋不成，因为结局要在指定的时期来到。
DAN|11|28|北方王必带许多财宝回本地，但他的心反对圣约；他恣意横行，回到本地。
DAN|11|29|“到了指定的时期，他必返回，侵入南方。这一次却不像前一次，
DAN|11|30|因为 基提 的战船要来攻击他，他就丧胆而退。他恼恨圣约，恣意横行，要回来善待那些背弃圣约的人。
DAN|11|31|他要兴兵，这兵必亵渎圣所，就是堡垒，除掉经常献的祭，设立那施行毁灭的可憎之物。
DAN|11|32|他必用巧言奉承违背圣约的恶人；惟独认识上帝的子民必刚强行事。
DAN|11|33|民间的智慧人必训诲许多人，然而在一段日子里，他们必因刀剑、火烧、掳掠、抢夺而仆倒。
DAN|11|34|他们仆倒的时候，会得到少许援助，却有许多人用诡诈加入他们。
DAN|11|35|智慧人中有些人仆倒，为要使他们受熬炼，成为洁净、洁白，直到末了；因为还有一段日子才到所定的时期。
DAN|11|36|“王必任意而行，自高自大，超过所有的神明，又用荒谬的话攻击万神之神。他必行事亨通，直到主的愤怒结束，因为所定的事必然实现。
DAN|11|37|他不顾他祖宗的神明，也不顾妇女所仰慕的神明，任何神明他都不顾；因为他自大，高过一切，
DAN|11|38|以敬奉堡垒的神明取而代之，用金、银、宝石和珍宝敬奉他祖宗所不认识的神明。
DAN|11|39|他靠外邦神明的帮助，攻破最坚固的堡垒。凡承认他的，他要给他们许多尊荣，使他们管辖许多人，又分封土地作为报偿。
DAN|11|40|“到末了，南方王要与北方王交战。北方王要用战车、骑兵和许多战船，势如暴风来攻击他，又要侵入列国，如洪水泛滥。
DAN|11|41|他要侵入那佳美之地，许多国就被倾覆 ，但 以东 人、 摩押 人和大半的 亚扪 人必逃离他的手。
DAN|11|42|他要伸手攻击列国，连 埃及 地也不得逃脱。
DAN|11|43|他要掌管 埃及 的金银财宝和各样珍宝， 路比 人和 古实 人都跟从他的脚步。
DAN|11|44|但从东方和北方必有消息传来扰乱他，他就大发烈怒出去，要将许多人杀灭净尽。
DAN|11|45|他要在海和荣美的圣山之间搭起王宫的帐幕；然而他的结局到了，无人能帮助他。”
DAN|12|1|“那时，保佑你百姓的天使长 米迦勒 必站起来，并且有大艰难，自从有国以来直到此时，未曾有过这样的事。那时，你的百姓凡记录在册上的，必得拯救。
DAN|12|2|睡在地里尘埃中的必有多人醒过来；其中有得永生的，有受羞辱永远被憎恶的。
DAN|12|3|智慧人要发光，如同天上的光；那领许多人归于义的必发光如星，直到永永远远。
DAN|12|4|但以理 啊，你要隐藏这话，封闭这书，直到末时。必有许多人往来奔跑 ，知识 就必增长。”
DAN|12|5|我－ 但以理 观看，看哪，另有两个人站立：一个在河这边，一个在河那边。
DAN|12|6|其中一个对那在河水之上、穿细麻衣的说：“这奇异的事要到几时才应验呢？”
DAN|12|7|我听见那在河水之上、穿细麻衣的，向天举起左右手，指着那活到永远的起誓说：“要到一年 、两年，又半年，粉碎圣民力量结束的时候，这一切的事就要应验。”
DAN|12|8|我听了却不明白，就说：“我主啊，这些事的结局是怎样呢？”
DAN|12|9|他说：“ 但以理 ，去吧！因为这话已经隐藏封闭，直到末时。
DAN|12|10|必有许多人使自己洁净、洁白，且受熬炼；但恶人仍必行恶，没有一个恶人明白，惟独智慧人能明白。
DAN|12|11|从除掉经常献的祭，设立那施行毁灭的可憎之物的时候起，必有一千二百九十日。
DAN|12|12|那等候，直到一千三百三十五日的有福了。
DAN|12|13|“至于你，你要去等候结局。你必安息，到了末期，你必起来，享受你的福分。”
HOS|1|1|当 乌西雅 、 约坦 、 亚哈斯 、 希西家 作 犹大 王， 约阿施 的儿子 耶罗波安 作 以色列 王的时候，耶和华的话临到 备利 的儿子 何西阿 。
HOS|1|2|耶和华初次向 何西阿 说话。耶和华对他说：“你去娶一个淫荡的女子为妻，收那从淫乱所生的儿女；因为这地行大淫乱，离弃耶和华。”
HOS|1|3|于是， 何西阿 去娶了 滴拉音 的女儿 歌篾 。她就怀孕，为 何西阿 生了一个儿子。
HOS|1|4|耶和华对 何西阿 说：“给他起名叫 耶斯列 ；因为再过片时，我要惩罚 耶户 家在 耶斯列 流人血的罪，也必终结 以色列 家的王朝。
HOS|1|5|到那日，我必在 耶斯列 平原折断 以色列 的弓。”
HOS|1|6|歌篾 又怀孕，生了一个女儿，耶和华对 何西阿 说：“给她起名叫 罗．路哈玛 ；因为我必不再怜悯 以色列 家，绝不赦免他们。
HOS|1|7|我却要怜悯 犹大 家，使他们靠耶和华－他们的上帝得救；我必不让他们靠弓、刀、战争、马匹与骑兵得救。”
HOS|1|8|歌篾 在 罗．路哈玛 断奶以后，又怀孕生了一个儿子。
HOS|1|9|耶和华说：“给他起名叫 罗．阿米 ；因为你们不是我的子民，我也不是你们的上帝 。”
HOS|1|10|然而， 以色列 的人数必多如海沙，不可量，不可数。从前在什么地方对他们说“你们不是我的子民”，将来就在那里称他们为“永生上帝的儿子”。
HOS|1|11|犹大 人和 以色列 人要一同聚集，为自己设立一个“头”，从这地上来，因为 耶斯列 的日子必为大日。
HOS|2|1|你们要称你们的众弟兄 为 阿米 ，称你们的众姊妹 为 路哈玛 。
HOS|2|2|要跟你们的母亲理论，理论， ─因为她不是我的妻子， 我也不是她的丈夫─ 叫她除掉脸上的淫相 和胸间的淫态，
HOS|2|3|免得我剥光她，使她赤身， 如刚出生的时候一样， 使她如旷野，如干旱之地， 干渴而死。
HOS|2|4|我必不怜悯她的儿女， 因为他们是从淫乱生的儿女。
HOS|2|5|他们的母亲行了淫乱， 怀他们的做了可羞耻的事； 因为她说：“我要跟随我所爱的， 我的饼、水、羊毛、麻、油、酒， 都是他们给的。”
HOS|2|6|因此，看哪，我要用荆棘堵塞她 的道， 筑墙挡住她， 使她找不着路；
HOS|2|7|以致她追随所爱的人，却追不上， 寻找他们，却寻不着， 就说：“我要回到前夫那里去， 因我那时比现在还好。”
HOS|2|8|她不知道是我给她五谷、新酒和新的油， 又加添她的金银； 他们却用来供奉 巴力 。
HOS|2|9|因此，我要在收割的日子收回我的五谷， 在当令的季节收回我的新酒， 我要夺回她用以遮体的羊毛和麻。
HOS|2|10|如今我必在她所爱的人眼前显露她的羞耻 ， 无人能救她脱离我的手。
HOS|2|11|我必使她的宴乐、节期、初一、安息日， 她一切的盛会都止息。
HOS|2|12|我要毁坏她的葡萄树和无花果树， 就是她所说“我所爱的给我为赏赐”的； 我要使它们变为荒林， 为野地的走兽所吞吃。
HOS|2|13|我要惩罚她素日给诸 巴力 烧香的罪； 那时她佩戴耳环和珠宝， 跟随她所爱的，却忘记我。 这是耶和华说的。
HOS|2|14|因此，看哪，我要诱导她，领她到旷野， 我要说动她的心。
HOS|2|15|在那里，我必赐她葡萄园， 又赐她 亚割谷 作为指望的门。 她必在那里回应， 像在年轻时从 埃及 地上来的时候一样。
HOS|2|16|那日你必称呼我 伊施 ，不再称呼我 巴力 。这是耶和华说的。
HOS|2|17|因为我必从她口中除掉诸 巴力 的名号，不再有人提这名号。
HOS|2|18|当那日，我必为我的百姓，与野地的走兽、天空的飞鸟和地上爬行的动物立约；又要在国中折断弓和刀，止息战争，使他们安然躺卧。
HOS|2|19|我必聘你永远归我为妻，以公义、公平、慈爱、怜悯聘你归我；
HOS|2|20|又以信实聘你归我，你就必认识耶和华。
HOS|2|21|耶和华说：那日我必应允， 我必应允天，天必应允地，
HOS|2|22|地必应允五谷、新酒和新的油； 这些都必应允在 耶斯列 身上。
HOS|2|23|我为自己必将她种在这地。 我必怜悯 罗．路哈玛 ； 对 罗．阿米 说： “你是我的子民”； 他必说：“我的上帝。”
HOS|3|1|耶和华又对我说：“你去爱那情人所爱却犯奸淫的妇人，正如耶和华爱那偏向别神、喜爱葡萄饼 的 以色列 人。”
HOS|3|2|于是我用十五舍客勒银子和一贺梅珥半大麦买她归我。
HOS|3|3|我对她说：“你当多日与我同住，不可行淫，不可归与别人，我对你也一样。”
HOS|3|4|因为 以色列 人必多日过着无君王，无领袖，无祭祀，无柱像，无以弗得，无家中神像的生活。
HOS|3|5|后来 以色列 人必归回 ，寻求耶和华─他们的上帝和他们的王 大卫 。在末后的日子，他们必敬畏耶和华，领受他的恩惠。
HOS|4|1|以色列 人哪，当听耶和华的话。 耶和华指控这地的居民， 因为在这地上无诚信， 无慈爱，无人认识上帝；
HOS|4|2|惟起誓、欺骗、杀害、 偷盗、奸淫、残暴、 流血又流血。
HOS|4|3|因此，这地悲哀， 其上的居民、野地的走兽、 天空的飞鸟都日趋衰微， 海中的鱼也必消灭。
HOS|4|4|然而，人都不必争辩，也不必指责。 你的百姓与抗拒祭司的人一样。
HOS|4|5|日间你必跌倒， 夜间先知也要与你一同跌倒； 我要灭绝你的母亲。
HOS|4|6|我的百姓因无知识而灭亡。 你抛弃知识， 我也必抛弃你， 使你不再作我的祭司。 你既忘了你上帝的律法， 我也必忘记你的儿女。
HOS|4|7|祭司越发增多，就越发得罪我； 我必使他们的荣耀变为羞辱。
HOS|4|8|他们吞吃我百姓的赎罪祭 ， 满心愿意我的子民犯罪。
HOS|4|9|将来百姓所受的， 祭司也必承受； 我必因他们所行的惩罚他们， 照他们所做的报应他们。
HOS|4|10|他们吃，却不得饱足； 行淫，却不繁衍； 因为他们离弃耶和华， 常行
HOS|4|11|淫乱。 酒和新酒夺去人的心。
HOS|4|12|我的百姓求问木头， 以为木杖能指示他们； 淫乱的心使他们失迷， 以致行淫离弃他们的上帝，
HOS|4|13|在各山顶献祭，在各高冈上烧香， 在橡树、杨树、大树之下， 因为那里树影美好。 所以，你们的女儿行淫， 你们的媳妇 犯奸淫。
HOS|4|14|我不因你们的女儿行淫 或你们的媳妇犯奸淫惩罚她们； 因为人自己转去与娼妓同居， 与神庙娼妓一同献祭。 这无知的百姓必致倾倒。
HOS|4|15|以色列 啊，你虽然行淫， 犹大 却不可犯罪； 不要往 吉甲 去， 不要上到 伯．亚文 ， 也不要指着永生的耶和华起誓。
HOS|4|16|以色列 倔强， 犹如倔强的母牛； 现在耶和华能牧放他们， 如在宽阔之地牧放羔羊吗？
HOS|4|17|以法莲 亲近偶像， 任凭他吧！
HOS|4|18|他们喝完了酒， 荒淫无度， 他们的官长甚爱羞耻的事。
HOS|4|19|风把他们卷在翅膀里， 他们必因所献的祭 蒙羞。
HOS|5|1|众祭司啊，要听这话！ 以色列 家啊，要留心听！ 王室啊，要侧耳而听！ 审判将临到你们， 因你们在 米斯巴 如罗网， 在 他泊山 如张开的网。
HOS|5|2|这些悖逆的人大行杀戮， 我要斥责他们众人。
HOS|5|3|至于我，我认识 以法莲 ， 以色列 不能向我隐藏。 以法莲 哪，现在你竟然行淫 ， 以色列 竟然被污辱。
HOS|5|4|他们所做的使他们不能归向上帝， 因有淫乱的心在他们里面； 他们不认识耶和华。
HOS|5|5|以色列 的骄傲使自己脸面无光 ； 以色列 和 以法莲 必因自己的罪孽跌倒， 犹大 也必与他们一同跌倒。
HOS|5|6|他们牵着牛羊去寻求耶和华， 却寻不着； 因他已转去离开他们。
HOS|5|7|他们不忠于耶和华， 生了私生子。 现在新月必吞灭他们和他们的地业。
HOS|5|8|你们当在 基比亚 吹角， 在 拉玛 吹号， 在 伯．亚文 发出警报； 便雅悯 哪，留意你的背后！
HOS|5|9|到了惩罚的日子， 以法莲 必变为废墟； 我在 以色列 众支派中，已指示将来必成的事。
HOS|5|10|犹大 的领袖如同挪移地界的人， 我必把我的愤怒如水倾倒在他们身上。
HOS|5|11|以法莲 因喜爱遵从荒谬的命令 就受欺压，在审判中被压碎。
HOS|5|12|我对 以法莲 竟如蛀虫， 向 犹大 家竟如朽烂。
HOS|5|13|以法莲 见自己有病， 犹大 见自己有伤， 以法莲 就前往 亚述 ， 差遣人去见大王 ； 他却不能医治你们， 不能治好你们的伤。
HOS|5|14|我必向 以法莲 如狮子， 向 犹大 家如少壮狮子。 我要撕裂，并且离去， 我必夺去，无人搭救。
HOS|5|15|我要去，我要回到原处， 等他们自觉有罪，寻求我的面； 急难时他们必切切寻求我。
HOS|6|1|来，我们归向耶和华吧！ 他撕裂我们，也必医治； 打伤我们，也必包扎。
HOS|6|2|过两天他必使我们苏醒， 第三天他必使我们兴起， 我们就在他面前得以存活。
HOS|6|3|我们要认识，要追求认识耶和华。 他如黎明必然出现， 他必临到我们像甘霖， 像滋润土地的春雨。
HOS|6|4|以法莲 哪，我可以向你怎样行呢？ 犹大 啊，我可以向你怎样做呢？ 因为你们的慈爱如同早晨的云雾， 又如速散的露水。
HOS|6|5|因此，我藉先知砍伐他们， 以我口中的话杀戮他们； 对你的审判 如光发出。
HOS|6|6|我喜爱慈爱 ，不喜爱祭物； 喜爱人认识上帝，胜于燔祭。
HOS|6|7|他们却如 亚当 背约， 在那里向我行诡诈。
HOS|6|8|基列 是作恶之人的城， 被血沾染。
HOS|6|9|成群的祭司如强盗埋伏等候， 在 示剑 的路上杀戮， 行了邪恶。
HOS|6|10|在 以色列 家我看见可憎的事， 在 以法莲 那里有淫行， 以色列 被污辱了。
HOS|6|11|犹大 啊，我使被掳之民归回的时候， 必有为你所预备的丰收。
HOS|7|1|我正要医治 以色列 的时候， 以法莲 的罪孽 和 撒玛利亚 的邪恶就显露出来。 他们行事虚谎， 内有贼人入侵， 外有群盗劫掠。
HOS|7|2|他们以为我不在意他们一切的恶行； 现在，他们所做的在我面前缠绕他们。
HOS|7|3|他们行恶使君王欢喜， 说谎使官长快乐。
HOS|7|4|他们全都犯奸淫， 如同烤热的火炉， 师傅在揉面到发面时 暂时停止煽火。
HOS|7|5|在我们君王宴乐的日子， 官长因酒的烈性而生病 ， 王与亵慢的人握手。
HOS|7|6|他们临近，心里如火炉一般， 他们等待，如烤饼的整夜睡觉， 到了早晨却如火焰熊熊。
HOS|7|7|他们全都热如火炉， 吞灭他们的审判官。 他们的君王都仆倒， 他们中间无一人求告我。
HOS|7|8|以法莲 混居在万民中 ， 以法莲 是没有翻过的饼。
HOS|7|9|外邦人消耗他的力量，他却不知道； 头发斑白，他也不觉得。
HOS|7|10|以色列 的骄傲使自己脸面无光。 他们虽遭遇这一切， 仍不归向耶和华－他们的上帝， 也不寻求他。
HOS|7|11|以法莲 好像鸽子愚蠢无知， 他们求告 埃及 ，投奔 亚述 。
HOS|7|12|他们去的时候，我要把我的网撒在他们身上； 我要捕获他们如同空中的鸟。 我必按他们会众所听到的 惩罚他们。
HOS|7|13|他们因离弃我，必定有祸； 因违背我，必遭毁灭。 我虽想要救赎他们，他们却向我说谎。
HOS|7|14|他们在床上呼号， 却不诚心哀求我； 他们为求五谷新酒而聚集 ， 却背叛我。
HOS|7|15|我虽管教他们，坚固他们的膀臂， 他们却图谋邪恶抗拒我。
HOS|7|16|他们归向，但不是归向至上者 ； 终究必如松弛的弓。 他们的领袖必因舌头的狂傲倒在刀下， 这在 埃及 地必成为人的笑柄。
HOS|8|1|你用口吹角吧！ 敌人如鹰攻打耶和华的家； 因为他们违背了我的约， 干犯了我的律法。
HOS|8|2|他们必呼求我： “我的上帝啊，我们 以色列 认识你了 。”
HOS|8|3|以色列 丢弃良善 ； 仇敌必追逼他。
HOS|8|4|他们立君王，并非出于我； 立官长，我却不知道。 他们用金银为自己制造偶像， 以致被剪除。
HOS|8|5|撒玛利亚 啊，耶和华已抛弃你的牛犊； 我的怒气向拜牛犊的人发作。 他们要到几时方能无罪呢？
HOS|8|6|因这牛犊是出于 以色列 ， 是匠人所造的， 并不是上帝。 撒玛利亚 的牛犊必被打碎。
HOS|8|7|他们所栽种的是风， 所收割的是暴风； 禾稼不长穗， 无以制成面粉； 即便制成， 外邦人也必吞吃它。
HOS|8|8|以色列 被吞吃， 如今在列国中像人所不喜爱的器皿。
HOS|8|9|他们投奔 亚述 如独行的野驴。 以法莲 雇用情人，
HOS|8|10|他们雇用列国； 如今我要聚集他们， 他们必因君王和官长所加的重担开始衰微 。
HOS|8|11|以法莲 为赎罪增添许多祭坛， 这些祭坛却使他犯罪。
HOS|8|12|我为他写了许多条 律法， 他却以为与他毫无关系。
HOS|8|13|他们献祭物作为给我的供物， 却自食其肉， 耶和华并不悦纳他们。 现在他必记起他们的罪孽， 惩罚他们的罪恶； 他们必返回 埃及 。
HOS|8|14|以色列 忘记造他的主，建造宫殿， 犹大 增添许多坚固的城； 我却要降火在他的城镇， 吞灭其堡垒。
HOS|9|1|以色列 啊，不要欢喜， 像 万民一样快乐； 因为你行淫离弃你的上帝， 喜爱各禾场上卖淫所得的赏金。
HOS|9|2|禾场和压酒池都不足以喂养他们， 它的新酒也必缺乏。
HOS|9|3|他们必不得住耶和华的地； 以法莲 却要返回 埃及 ， 在 亚述 吃不洁净的食物。
HOS|9|4|他们必不得向耶和华献浇酒祭， 所献的祭也不蒙悦纳。 他们的祭物如居丧者的食物， 凡吃的必使自己玷污； 因为他们的食物只为自己的口腹， 必不得入耶和华的殿。
HOS|9|5|到盛会的日子，在耶和华的节期， 你们要怎样行呢？
HOS|9|6|看哪，他们要逃避灾难； 埃及 人要收殓他们， 摩弗 人要埋葬他们。 蒺藜盘踞他们贵重的银器， 荆棘必占据他们的帐棚。
HOS|9|7|降罚的日子近了， 报应的时候已经来到。 以色列 必知道， 先知愚昧， 受灵感动的人狂妄， 皆因你多多作恶，大怀怨恨。
HOS|9|8|以法莲 替我的上帝守望； 至于先知，他所到之处都有捕鸟人的罗网， 在他上帝的家中也遭人怀恨。
HOS|9|9|他们深深败坏， 如在 基比亚 的日子一样。 耶和华必记起他们的罪孽， 惩罚他们的罪恶。
HOS|9|10|我发现 以色列 ， 如在旷野的葡萄； 我看见你们的祖先， 如春季无花果树上初熟的果子。 他们却来到 巴力．毗珥 ， 献上自己做羞耻的事， 成为可憎恶的， 与他们所爱的一样。
HOS|9|11|以法莲 ，他们的荣耀如鸟飞去， 必不生产，不怀胎，不成孕；
HOS|9|12|他们纵然将儿女养大， 我却要使他们丧子，一个也不留。 我离弃他们， 他们就有祸了。
HOS|9|13|我看 以法莲 如 推罗 栽于美地。 以法莲 却要将自己的儿女带出来， 交给行杀戮的人。
HOS|9|14|耶和华啊，求你加给他们， 加给他们什么呢？ 要使他们怀孕流产， 乳房枯干。
HOS|9|15|因他们在 吉甲 的一切恶事， 我在那里憎恶他们。 因他们所行的恶， 我必把他们赶出我的殿， 不再爱他们； 他们的领袖都是悖逆的。
HOS|9|16|以法莲 受击打， 其根枯干，不能结果， 即或生产， 我也要杀他们所生的爱子。
HOS|9|17|我的上帝必弃绝他们， 因为他们不听从他； 他们必飘流在列国中。
HOS|10|1|以色列 是茂盛的葡萄树， 结果繁多。 果子越多， 就越增添祭坛； 土地越肥美， 就越建造美丽的柱像。
HOS|10|2|他们心怀二意， 现今要定为有罪。 耶和华必拆毁他们的祭坛， 粉碎他们的柱像。
HOS|10|3|现在他们要说： “我们没有王； 因为我们不敬畏耶和华， 王又能为我们做什么呢？”
HOS|10|4|他们讲空话， 以假誓立约； 因此，惩罚如苦菜滋生 在田间的犁沟中。
HOS|10|5|撒玛利亚 的居民必因 伯．亚文 的牛犊惊恐； 它的百姓为它悲哀， 它的祭司为它战兢， 因为荣耀已经离开它。
HOS|10|6|人必将牛犊带到 亚述 ， 当作礼物献给大王。 以法莲 必蒙羞， 以色列 必因自己的计谋惭愧。
HOS|10|7|撒玛利亚 的王要灭亡， 如水面上的泡沫一般。
HOS|10|8|亚文 的丘坛， 以色列 犯罪的地方必毁坏， 荆棘和蒺藜必长在他们的祭坛上。 他们要向大山说：遮盖我们！ 向小山说：倒在我们身上！
HOS|10|9|以色列 啊， 你从 基比亚 的日子以来就时常犯罪， 他们仍停留在那里。 攻击罪孽之辈的战事岂不会临到 基比亚 吗？
HOS|10|10|我必随己意惩罚他们， 他们为双重的罪所缠； 万民必聚集攻击他们。
HOS|10|11|以法莲 是驯良的母牛犊，喜爱踹谷， 我要将轭套在它肥美的颈项上， 我要使 以法莲 被套住； 犹大 必耕田， 雅各 必耙地。
HOS|10|12|你们要为自己栽种公义， 收割慈爱。 你们要开垦荒地， 现今正是寻求耶和华的时候； 等他临到，公义必如雨降给你们。
HOS|10|13|你们耕种奸恶， 收割罪孽， 吃的是谎言的果实。 因你倚靠自己的行为， 仰赖你众多的勇士，
HOS|10|14|所以在你百姓中必掀起闹哄， 你一切的堡垒必被拆毁， 就如 沙勒幔 在争战的日子拆毁 伯．亚比勒 ， 将城中的母子一同摔死。
HOS|10|15|伯特利 啊，因你们的大恶， 你们必遭遇如此。 黎明来临， 以色列 的王必全然灭绝。
HOS|11|1|以色列 年幼的时候，我爱他， 就从 埃及 召我的儿子出来。
HOS|11|2|先知 越是呼唤他们， 他们越是远离 ， 向诸 巴力 献祭， 为雕刻的偶像烧香。
HOS|11|3|我曾教导 以法莲 行走， 我用膀臂 抱起他们， 他们却不知道是我医治他们。
HOS|11|4|我用慈绳爱索牵引他们； 我待他们如人松开牛两腮旁边的轭， 弯下身来喂养他们。
HOS|11|5|他们必不返回 埃及 地； 然而 亚述 人要作他们的王， 因他们不肯归向我。
HOS|11|6|刀剑必临到他们的城镇， 毁坏门闩，吞灭众人， 都因他们自己的计谋。
HOS|11|7|我的百姓偏要背离我， 他们虽向至高者呼求， 他却不抬举他们 。
HOS|11|8|以法莲 哪，我怎能舍弃你？ 以色列 啊，我怎能弃绝你？ 我怎能使你如 押玛 ？ 怎能使你如 洗扁 ？ 我回心转意， 我的怜悯燃了起来。
HOS|11|9|我必不发猛烈的怒气， 也不再毁灭 以法莲 。 因我是上帝，并非世人， 是你们中间的圣者； 我必不在怒中临到你们。
HOS|11|10|耶和华如狮子吼叫， 他的儿女必跟随他。 他一吼叫， 他们就从西方战兢而来。
HOS|11|11|他们必如雀鸟从 埃及 战兢而来， 又如鸽子从 亚述 地来到。 我必使他们住自己的房屋； 这是耶和华说的。
HOS|11|12|以法莲 用谎言围绕我， 以色列 家用诡计环绕我； 犹大 却仍与上帝同行 ， 向圣者忠心。
HOS|12|1|以法莲 以风为食物， 终日追逐东风， 增添虚谎和残暴， 与 亚述 立约， 也把油送到 埃及 。
HOS|12|2|耶和华指控 犹大 ， 要照 雅各 所行的惩罚他， 按他所做的报应他。
HOS|12|3|他在腹中抓住哥哥的脚跟， 壮年的时候与上帝角力，
HOS|12|4|他与天使角力，并且得胜。 他曾哀哭，恳求施恩。 在 伯特利 遇见耶和华， 耶和华在那里吩咐我们 ，
HOS|12|5|耶和华是万军之上帝， 耶和华是他可记念的名。
HOS|12|6|所以你当归向你的上帝， 谨守慈爱和公平， 常常等候你的上帝。
HOS|12|7|商人 手持诡诈的天平， 喜爱欺压。
HOS|12|8|以法莲 说： 我果然富有，得了财宝； 我所劳碌得来的一切 人必找不到我有什么可算为有罪的恶。
HOS|12|9|自从你出 埃及 地以来， 我就是耶和华－你的上帝； 我必使你再住帐棚， 如同节期的日子一样。
HOS|12|10|我已吩咐众先知， 又增加异象， 藉先知设比喻。
HOS|12|11|基列 没有罪孽吗？ 他们诚然是虚假的， 在 吉甲 献牛犊为祭； 他们的祭坛如同田间犁沟中的乱堆。
HOS|12|12|从前 雅各 逃到 亚兰 地， 以色列 为娶妻子工作， 为娶妻子而牧放。
HOS|12|13|后来耶和华藉先知领 以色列 从 埃及 上来， 也藉先知看顾他们。
HOS|12|14|然而 以法莲 大大惹动主怒， 他所流的血必归到他身上。 主必使他的羞辱归还给他。
HOS|13|1|从前 以法莲 说话，人都战兢， 他在 以色列 中居处高位； 但他因 巴力 犯罪就死了。
HOS|13|2|如今他们罪上加罪， 为自己铸造偶像， 凭自己的聪明用银子造偶像， 全都是匠人所制的。 论到它，有话说： 献祭的人都要亲吻牛犊。
HOS|13|3|因此，他们必如早晨的云雾， 又如速散的露水， 如被狂风吹离禾场的糠秕， 又如烟囱冒出的烟。
HOS|13|4|自从你出 埃及 地以来， 我就是耶和华－你的上帝； 除了我上帝以外，你不认识别的， 在我以外，并没有救主。
HOS|13|5|我曾在旷野， 就是那干旱之地认识你。
HOS|13|6|他们得到喂养，就饱足； 既得饱足，就心高气傲， 因而忘记了我。
HOS|13|7|因此我向他们如同狮子， 又如豹伏在道旁。
HOS|13|8|我如失去小熊的母熊，攻击他们， 撕裂他们的胸膛。 在那里我必如母狮吞吃他们， 如野兽撕开他们。
HOS|13|9|以色列 啊，你自取灭亡了 ， 因为我才是你的帮助。
HOS|13|10|现在，你的王在哪里呢？ 让他在你的各城中拯救你吧！ 你曾说“给我立君王和官长”， 那些治理你的又在哪里呢？
HOS|13|11|我在怒气中将王赐给你， 又在烈怒中将王废去。
HOS|13|12|以法莲 的罪孽被卷起来， 他的罪恶被收藏起来。
HOS|13|13|产妇的疼痛必临到他身上； 他是无智慧之子， 如同临盆时未出现的胎儿。
HOS|13|14|我必救赎他们脱离阴间， 救赎他们脱离死亡。 死亡啊，你的灾害在哪里？ 阴间哪，你的毁灭在哪里？ 怜悯必从我眼前消逝。
HOS|13|15|他在弟兄中虽然旺盛， 却有东风刮来， 就是耶和华的风从旷野上来。 他的泉源必干涸， 他的源头必枯竭， 这风必夺走他所积蓄的一切宝物。
HOS|13|16|撒玛利亚 要担当罪孽， 因为背叛自己的上帝。 他们必倒在刀下， 婴孩必被摔死， 孕妇必被剖开。
HOS|14|1|以色列 啊，你要归向耶和华－你的上帝， 你因自己的罪孽跌倒了。
HOS|14|2|当归向耶和华， 用言语向他说： “求你除尽罪孽，悦纳善行， 我们就用嘴唇的祭代替牛犊献上。
HOS|14|3|亚述 不能救我们， 我们不再骑马， 也不再对我们手所造的偶像说： ‘你是我们的上帝’； 孤儿在你那里得蒙怜悯。”
HOS|14|4|我必医治他们背道的病， 甘心爱他们， 因为我向他们所发的怒气已转消。
HOS|14|5|我必向 以色列 如甘露； 他必如百合花开放， 如 黎巴嫩 的树扎根。
HOS|14|6|他的嫩枝必延伸， 他的荣华如橄榄树， 香气如 黎巴嫩 的香柏树。
HOS|14|7|曾住在他荫下的必归回，使五谷生长 ， 他们要发旺如葡萄树， 他的名气 如 黎巴嫩 的酒。
HOS|14|8|以法莲 说： “我与偶像有何相干？” 我应允他，顾念他： 我如青翠的松树， 你的果实从我而来。
HOS|14|9|智慧人必明白这些事， 聪明人必知道这一切。 耶和华的道是正直的， 义人行在其中， 罪人却在其上跌倒。
JOEL|1|1|耶和华的话临到 毗土珥 的儿子 约珥 。
JOEL|1|2|老年人哪，当听这话； 这地所有的居民哪，要侧耳而听。 在你们的日子， 或你们祖先的日子， 曾发生过这样的事吗？
JOEL|1|3|你们要将这事传与子， 子传与孙， 孙传与后代。
JOEL|1|4|剪虫吃剩的，蝗虫来吃； 蝗虫吃剩的，蝻子来吃； 蝻子吃剩的，蚂蚱 来吃。
JOEL|1|5|醉酒的人哪，要清醒，要哭泣； 好酒的人哪，都要为甜酒哀号， 因为酒从你们的口中断绝了。
JOEL|1|6|有一队蝗虫 ，强盛且不可数， 上来侵犯我的地； 它的牙齿如狮子的牙齿， 如母狮的大牙。
JOEL|1|7|它毁坏我的葡萄树， 撕裂我的无花果树， 剥光又丢弃，使枝条露白。
JOEL|1|8|你要像童女腰束麻布， 为她年少时的丈夫哀号。
JOEL|1|9|耶和华的殿中断绝素祭和浇酒祭， 事奉耶和华的祭司都悲哀。
JOEL|1|10|田荒凉，地悲哀； 因为五谷毁坏， 新酒枯竭， 新的油也缺乏。
JOEL|1|11|农夫啊，要惭愧； 修整葡萄园的啊，你们要哀号； 因为大麦、小麦与田间的庄稼全都毁了。
JOEL|1|12|葡萄树枯干， 无花果树衰残， 石榴树、棕树、苹果树， 田野一切的树木都枯干； 众人的喜乐尽都消逝。
JOEL|1|13|祭司啊，当束上麻布痛哭； 事奉祭坛的啊，要哀号； 事奉我上帝的啊，你们要来，披上麻布过夜， 因为在你们上帝的殿中不再有素祭和浇酒祭了。
JOEL|1|14|你们要使禁食的日子分别为圣， 宣告严肃会， 召集长老和这地所有的居民 来到耶和华－你们上帝的殿， 向耶和华哀求。
JOEL|1|15|哀哉，这日子！ 因为耶和华的日子临近， 好像毁灭从全能者来到。
JOEL|1|16|粮食不是在我们眼前断绝了吗？ 欢喜快乐不是从我们上帝的殿中止息了吗？
JOEL|1|17|种子在土块下朽烂， 仓荒凉，廪破坏， 因为五谷枯干了。
JOEL|1|18|牲畜哀鸣， 牛群混乱，因无草场， 羊群也受苦。
JOEL|1|19|耶和华啊，我向你求告， 因为有火吞噬野地的草场， 火焰烧尽田野的树木。
JOEL|1|20|田野的走兽切慕你， 因为溪水干涸， 火吞噬了野地的草场。
JOEL|2|1|你们要在 锡安 吹角， 在我的圣山发出警报。 这地所有的居民要发颤， 因为耶和华的日子快到， 已经临近了。
JOEL|2|2|那是黑暗、阴森的日子， 是密云、乌黑的日子， 如同黎明笼罩山岭。 有一队蝗虫，又大又强， 自古以来没有像这样的， 以后直到万代也必没有。
JOEL|2|3|它们前面有火吞噬， 后面有火焰烧尽。 它们未到以前，地如 伊甸园 ， 过去以后，却成了荒凉的旷野， 没有一样能躲避它们。
JOEL|2|4|它们形状如马， 奔跑如战马。
JOEL|2|5|响声如战车在山顶上跳动， 如火焰吞噬碎秸， 好像强大的军队摆阵备战。
JOEL|2|6|在它们面前，万民伤恸， 脸都变色。
JOEL|2|7|它们如勇士奔跑， 如战士攀登城墙， 各行于自己的道路， 不乱队伍；
JOEL|2|8|它们并不彼此推挤， 各行于自己的大道， 冲过防御 ， 并不停止。
JOEL|2|9|它们蹦上城， 跳上墙， 爬上房屋， 从窗户进来，如同盗贼。
JOEL|2|10|在它们面前， 地动天摇， 日月昏暗， 星宿无光。
JOEL|2|11|耶和华在他的军旅前出声， 他的队伍庞大， 遵行他命令的强盛。 耶和华的日子大而可畏， 谁能当得起呢？
JOEL|2|12|然而你们现在要禁食，哭泣，哀号， 一心归向我。 这是耶和华说的。
JOEL|2|13|你们要撕裂心肠， 不要撕裂衣服。 归向耶和华－你们的上帝， 因为他有恩惠，有怜悯， 不轻易发怒， 有丰盛的慈爱， 并且会改变心意， 不降那灾难。
JOEL|2|14|谁知道他也许会回心转意，留下余福， 就是献给耶和华－你们上帝的素祭和浇酒祭。
JOEL|2|15|你们要在 锡安 吹角， 使禁食的日子分别为圣， 宣告严肃会。
JOEL|2|16|聚集百姓，使会众自洁； 召集老年人， 聚集孩童和在母怀吃奶的； 使新郎出内室， 新娘离开洞房。
JOEL|2|17|事奉耶和华的祭司 要在走廊和祭坛间哭泣，说： “耶和华啊，求你顾惜你的百姓， 不要使你的产业受羞辱， 在列国中成为笑柄。 为何让人在万民中说 ‘他们的上帝在哪里’呢？”
JOEL|2|18|耶和华为自己的地发热心， 怜悯他的百姓。
JOEL|2|19|耶和华应允他的百姓说： “看哪，我要赏赐你们五谷、新酒和新的油， 使你们饱足， 我必不再使你们受列国的羞辱。
JOEL|2|20|我要使北方来的队伍远离你们， 将他们赶到干旱荒芜之地： 前队赶入东海， 后队赶入西海； 臭气上升，恶臭腾空。 耶和华果然行了大事！
JOEL|2|21|“土地啊，不要惧怕， 要欢喜快乐， 因为耶和华行了大事。
JOEL|2|22|田野的走兽啊，不要惧怕， 因为旷野的草已生长， 树木结果， 无花果树、葡萄树也都效力 。
JOEL|2|23|“ 锡安 的民哪，你们要欢喜， 要因耶和华－你们的上帝快乐； 因他赏赐你们合宜的秋雨 ， 为你们降下甘霖， 秋雨和春雨，和先前一样。
JOEL|2|24|“禾场充满五谷， 池中漫溢新酒和新的油。
JOEL|2|25|我差遣到你们中间的大军队， 就是蝗虫、蝻子、蚂蚱、剪虫， 那些年间所吃的，我要补还给你们。
JOEL|2|26|“你们必吃得饱足， 赞美耶和华－你们上帝的名， 他为你们行了奇妙的事。 我的百姓不致羞愧，直到永远。
JOEL|2|27|你们必知道我是在 以色列 中， 又知道我是耶和华－你们的上帝，没有别的。 我的百姓不致羞愧，直到永远。”
JOEL|2|28|“以后，我要将我的灵浇灌凡有血肉之躯的。 你们的儿女要说预言， 你们的老人要做异梦， 你们的少年要见异象。
JOEL|2|29|在那些日子， 我要将我的灵浇灌我的仆人和婢女。
JOEL|2|30|“我要在天上地下显出奇事，有血，有火，有烟柱。
JOEL|2|31|太阳要变为黑暗，月亮要变为血，这都在耶和华大而可畏的日子未到以前。
JOEL|2|32|那时，凡求告耶和华名的就必得救；因为照耶和华所说的，在 锡安山 ，在 耶路撒冷 将有逃脱的人。凡耶和华所召的 ，都在余民之列。”
JOEL|3|1|“看哪，在那些日子，到那个时候，我使 犹大 和 耶路撒冷 被掳之人归回的时候，
JOEL|3|2|我要聚集万民，带他们下到 约沙法谷 去，在那里我要为我百姓，我产业 以色列 的缘故，向万民施行审判；因为他们把我的百姓分散到列国，瓜分了我的土地，
JOEL|3|3|为我的百姓抽签，以男孩换取妓女，为喝酒卖掉女孩。
JOEL|3|4|“ 推罗 、 西顿 和 非利士 四境的人哪，你们与我何干？你们要报复我吗？若要报复我，我必使报应速速归到你们头上。
JOEL|3|5|你们夺取我的金银，把我珍贵的宝物带入你们的庙宇 ，
JOEL|3|6|并将 犹大 人和 耶路撒冷 人卖给 希腊 人 ，使他们远离自己的疆土。
JOEL|3|7|看哪，我必激发他们离开你们把他们卖去的地方，又必使报应归到你们头上。
JOEL|3|8|我要将你们的儿女卖到 犹大 人手中，他们必转卖给远方的国家 示巴 人。这是耶和华说的。”
JOEL|3|9|当在列国中宣告： 预备打仗， 激发勇士， 使所有战士上前来。
JOEL|3|10|要将犁头打成刀剑， 镰刀打成戈矛； 弱者要说：“我是勇士。”
JOEL|3|11|四围的列国啊， 要速速前来， 一同聚集。 耶和华啊， 求你使你的勇士降临。
JOEL|3|12|列国都当兴起， 上到 约沙法谷 ； 因为我必坐在那里， 审判四围的列国。
JOEL|3|13|挥镰刀吧！因为庄稼熟了； 来踩踏吧！因为醡酒池满了。 酒池已经满溢， 因为他们的罪恶甚大。
JOEL|3|14|在 断定谷 有许多许多的人， 因为耶和华的日子临近 断定谷 了。
JOEL|3|15|日月昏暗， 星宿无光。
JOEL|3|16|耶和华必从 锡安 吼叫， 从 耶路撒冷 出声， 天地就震动。 耶和华却要作他百姓的避难所， 作 以色列 人的保障。
JOEL|3|17|你们就知道我是耶和华－你们的上帝， 我住在 锡安 －我的圣山。 耶路撒冷 必成为圣； 陌生人不再从其中经过。
JOEL|3|18|在那日，大山要滴甜酒， 小山要流奶， 犹大 的溪河都有水流出； 必有泉源从耶和华的殿中流出， 滋润 什亭谷 。
JOEL|3|19|埃及 必定荒凉， 以东 成为荒凉的旷野， 因为他们向 犹大 人行残暴， 又因他们在本地流无辜人的血。
JOEL|3|20|但 犹大 必存到永远， 耶路撒冷 必存到万代。
JOEL|3|21|我要免除 流人血的罪， 是先前未曾免除的， 耶和华居住在 锡安 。
AMOS|1|1|这是 犹大 王 乌西雅 在位与 约阿施 的儿子 以色列 王 耶罗波安 在位的时候，大地震前二年，从 提哥亚 来的牧人 阿摩司 所见的─他的话论到 以色列 。
AMOS|1|2|他说：“耶和华必从 锡安 吼叫， 从 耶路撒冷 出声； 牧人的草场哀伤， 迦密 的山顶枯干。”
AMOS|1|3|耶和华如此说： “ 大马士革 三番四次犯罪， 以铁的打谷机击打 基列 ， 我必不撤销对它的惩罚。
AMOS|1|4|我要降火在 哈薛 的王宫， 吞灭 便．哈达 的宫殿；
AMOS|1|5|我要折断 大马士革 的门闩， 剪除 亚文 平原的居民 和 伯．伊甸 的掌权者， 亚兰 人必被掳到 吉珥 。” 这是耶和华说的。
AMOS|1|6|耶和华如此说： “ 迦萨 三番四次犯罪， 掳掠全体百姓交给 以东 ， 我必不撤销对它的惩罚。
AMOS|1|7|我要降火在 迦萨 城内， 吞灭它的宫殿；
AMOS|1|8|我要剪除 亚实突 的居民 和 亚实基伦 的掌权者， 反手攻击 以革伦 ， 剩余的 非利士 人都必灭亡。” 这是主耶和华说的。
AMOS|1|9|耶和华如此说： “ 推罗 三番四次犯罪， 将全体百姓交给 以东 ， 不顾念弟兄的盟约， 我必不撤销对它的惩罚，
AMOS|1|10|我要降火在 推罗 城内， 吞灭它的宫殿。”
AMOS|1|11|耶和华如此说： “ 以东 三番四次犯罪， 怒气不停发作，永远怀着愤怒， 拿刀追赶兄弟，丝毫不存怜悯， 我必不撤销对它的惩罚。
AMOS|1|12|我要降火在 提幔 ， 吞灭 波斯拉 的宫殿。”
AMOS|1|13|耶和华如此说： “ 亚扪 人三番四次犯罪， 剖开 基列 的孕妇， 扩张自己的疆界， 我必不撤销对它的惩罚。
AMOS|1|14|我要在战争呐喊的日子， 在旋风狂吹时， 在 拉巴 城内放火， 吞灭它的宫殿；
AMOS|1|15|他们的君王和官长必一同被掳。” 这是耶和华说的。
AMOS|2|1|耶和华如此说： “ 摩押 三番四次犯罪， 把 以东 王的骸骨焚烧成灰， 我必不撤销对它的惩罚。
AMOS|2|2|我要降火在 摩押 ， 吞灭 加略 的宫殿， 摩押 必在闹哄、呐喊、吹角声中灭亡；
AMOS|2|3|我要剪除 摩押 的领袖， 把所有的官长和他一同杀戮。” 这是耶和华说的。
AMOS|2|4|耶和华如此说： “ 犹大 三番四次犯罪， 厌弃耶和华的训诲， 不遵守他的律例； 他们祖先所随从虚假的偶像 使他们走迷了， 我必不撤销对它的惩罚。
AMOS|2|5|我要降火在 犹大 ， 吞灭 耶路撒冷 的宫殿。”
AMOS|2|6|耶和华如此说： “ 以色列 三番四次犯罪， 为银子卖了义人， 为一双鞋卖了穷人， 我必不撤销对它的惩罚。
AMOS|2|7|他们把贫寒人的头践踏在地的尘土上 ， 又阻碍困苦人的道路。 父子与同一个女子行淫， 以致亵渎我的圣名。
AMOS|2|8|他们在各祭坛旁边， 躺卧在人所典当的衣服上， 又在他们上帝的殿里 喝受罚之人的酒。
AMOS|2|9|“我从他们面前除灭 亚摩利 人； 他虽高大如香柏树，强壮如橡树， 我却上灭其果，下绝其根。
AMOS|2|10|我曾将你们从 埃及 地领上来， 在旷野里引导你们四十年， 使你们得 亚摩利 人之地为业；
AMOS|2|11|我从你们子孙中兴起先知， 又从你们少年中兴起拿细耳人。 以色列 人哪，不是这样吗？” 这是耶和华说的。
AMOS|2|12|“你们却把酒给拿细耳人喝， 嘱咐先知说：‘不要说预言。’
AMOS|2|13|“看哪，我要把你们压下去， 如同装满禾捆的车压过一样。
AMOS|2|14|快跑的无从避难， 壮士无法使力， 勇士也不能自救；
AMOS|2|15|拿弓的站立不住， 腿快的不能逃脱， 骑马的也不能自救。
AMOS|2|16|到那日，勇士中最有胆量的， 必赤身逃跑。” 这是耶和华说的。
AMOS|3|1|以色列 人哪，当听耶和华责备你们的话，责备我从 埃及 地领上来的全家，说：
AMOS|3|2|“在地上万族中，我只认识你们； 因此，我必惩罚你们一切的罪孽。”
AMOS|3|3|二人若不同心， 岂能同行呢？
AMOS|3|4|狮子若无猎物， 岂会在林中咆哮呢？ 少壮狮子若无所得， 岂会从洞里吼叫呢？
AMOS|3|5|若未设圈套， 雀鸟岂能陷入地上的罗网呢？ 罗网若无所得， 岂会从地上翻起呢？
AMOS|3|6|城中若吹角， 百姓岂不战兢吗？ 灾祸若临到一城， 岂非耶和华所降的吗？
AMOS|3|7|主耶和华不会做任何事情， 除非先将奥秘指示他的仆人众先知。
AMOS|3|8|狮子吼叫，谁不惧怕呢？ 主耶和华既已说了，谁能不说预言呢？
AMOS|3|9|你们要在 亚实突 的宫殿 和 埃及 地的宫殿传扬，说： “要聚集在 撒玛利亚 的山上， 看城里有何等大的扰乱与欺压。”
AMOS|3|10|“他们以暴力抢夺， 堆积在自己的宫殿里， 却不懂得行正直的事。” 这是耶和华说的。
AMOS|3|11|所以主耶和华如此说： “敌人必来围攻这地， 削弱你的势力， 抢掠你的宫殿。”
AMOS|3|12|耶和华如此说：“牧人怎样从狮子口中抢回两条腿或耳朵的一小片，住 撒玛利亚 的 以色列 人得救也是如此，不过抢回床的一角和床榻的靠枕 而已。”
AMOS|3|13|主耶和华－万军之上帝说： “当听这话，警戒 雅各 家。
AMOS|3|14|我惩罚 以色列 罪孽的日子， 也要惩罚 伯特利 的祭坛； 祭坛的角必被砍下，坠落于地。
AMOS|3|15|我要拆毁过冬和避暑的房屋， 象牙的房屋必毁灭， 广厦豪宅都归无有。” 这是耶和华说的。
AMOS|4|1|“你们这些 撒玛利亚山 上的 巴珊 母牛啊， 当听这话！ 你们欺负贫寒人，压碎贫穷人， 对主人说：‘拿酒来，我们喝吧！’
AMOS|4|2|主耶和华指着自己的神圣起誓说： ‘看哪，日子将到，人必用钩子将你们钩去， 用鱼钩把你们中最后一个钩去。
AMOS|4|3|你们必从城墙的缺口 出去， 各人直往前行， 投向 哈门 。’” 这是耶和华说的。
AMOS|4|4|“ 以色列 人哪，任你们往 伯特利 去犯罪， 到 吉甲 增加罪过， 每早晨献上你们的祭物， 每三日纳你们的十一奉献；
AMOS|4|5|任你们献上有酵的感谢祭， 宣扬你们的甘心祭，使人听见， 因为这是你们所喜爱的。” 这是主耶和华说的。
AMOS|4|6|“我使你们在每一座城里牙齿干净， 使你们各处的粮食缺乏， 你们仍不归向我。” 这是耶和华说的。
AMOS|4|7|“在收割的前三个月， 我不降雨在你们那里， 我降雨在这城， 不降雨在那城； 这块地有雨， 那块无雨的地就必枯干。
AMOS|4|8|两三城的人挤到一个城去找水喝， 却喝不足， 你们仍不归向我。” 这是耶和华说的。
AMOS|4|9|“我以焚风 和霉烂攻击你们， 你们许多的菜园、葡萄园、 无花果树、橄榄树屡屡被剪虫 所吃， 你们仍不归向我。” 这是耶和华说的。
AMOS|4|10|“我降瘟疫在你们中间， 如在 埃及 的样子； 用刀杀戮你们的年轻人 和你们遭掳掠的马匹， 营中臭气扑鼻， 你们仍不归向我。” 这是耶和华说的。
AMOS|4|11|“我倾覆你们， 如同上帝从前倾覆 所多玛 、 蛾摩拉 一样； 你们好像从火中抢救出来的一根柴， 你们仍不归向我。” 这是耶和华说的。
AMOS|4|12|“因此， 以色列 啊，我要如此对待你； 因为我要这样对待你， 以色列 啊， 你当预备迎见你的上帝。”
AMOS|4|13|看哪，那创山，造风，将其心意指示人， 使晨光变幽暗，踩行在地之高处的， 他的名是耶和华－万军之上帝。
AMOS|5|1|以色列 家啊，听我为你们所作的哀歌：
AMOS|5|2|“ 以色列 民 跌倒，不得再起； 躺在地上，无人扶起。”
AMOS|5|3|主耶和华如此说： “ 以色列 家的城派出一千，只剩一百； 派出一百，只剩十个。”
AMOS|5|4|耶和华向 以色列 家如此说： “你们要寻求我，就必存活。
AMOS|5|5|不要往 伯特利 寻求， 不要进入 吉甲 ， 也不要过到 别是巴 ； 因为 吉甲 必被掳走， 伯特利 必归无有。”
AMOS|5|6|要寻求耶和华，就必存活， 免得他在 约瑟 家如火发出， 焚烧 伯特利 ，无人扑灭。
AMOS|5|7|你们这使公平变为茵蔯， 将公义丢弃于地的人哪！
AMOS|5|8|那造昴星和参星， 使死荫变为晨光， 使白昼变为黑夜， 召唤海水、 使其倾倒在地面上的， 耶和华是他的名。
AMOS|5|9|他快速摧毁强壮的人， 毁灭就临到堡垒。
AMOS|5|10|你们怨恨那在城门口断是非的， 憎恶那说正直话的。
AMOS|5|11|所以，因你们践踏贫寒人， 向他们勒索粮税； 你们虽建造石凿的房屋， 却不得住在其内； 虽栽植美好的葡萄园， 却不得喝其中所出的酒。
AMOS|5|12|我知道你们的罪过何其多， 你们的罪恶何其大； 你们迫害义人，收受贿赂， 在城门口屈枉贫穷人。
AMOS|5|13|所以智慧人在这样的时候必静默不言， 因为这是险恶的时候。
AMOS|5|14|你们要寻求良善， 不要寻求邪恶，就必存活。 这样，耶和华－万军之上帝 必照你们所说的与你们同在。
AMOS|5|15|要恨恶邪恶，喜爱良善， 在城门口秉公行义； 或者耶和华－万军之上帝 会施恩给 约瑟 的余民。
AMOS|5|16|因此，主耶和华－万军之上帝如此说： “在一切的广场上必有哀号的声音； 在各街市上必有人说： ‘哀哉！哀哉！’ 他们叫农夫来哭号， 叫善唱哀歌的来举哀；
AMOS|5|17|各葡萄园都有哀号的声音， 因为我必从你中间经过。” 这是耶和华说的。
AMOS|5|18|想望耶和华日子的人有祸了！ 为什么你们要耶和华的日子呢？ 那是黑暗没有光明的日子，
AMOS|5|19|好像人躲避狮子却遇见熊； 进房屋以手靠墙，却被蛇咬。
AMOS|5|20|耶和华的日子岂不是黑暗没有光明， 幽暗毫无光辉吗？
AMOS|5|21|“我厌恶你们的节期， 也不喜悦你们的严肃会。
AMOS|5|22|你们虽然向我献燔祭和素祭， 我却不悦纳， 也不看你们用肥畜献的平安祭。
AMOS|5|23|要使你们歌唱的声音远离我， 因为我不听你们琴瑟的乐曲。
AMOS|5|24|惟愿公平如大水滚滚， 公义如江河滔滔。
AMOS|5|25|“ 以色列 家啊，你们在旷野四十年，何尝将祭物和供物献给我呢？
AMOS|5|26|你们抬着你们的 撒古特 君王 ，和你们为自己所造之偶像 迦温 ，你们的神明之星。
AMOS|5|27|所以我要把你们掳到 大马士革 以外。”这是耶和华说的，他的名为万军之上帝。
AMOS|6|1|“那在 锡安 安逸， 在 撒玛利亚山 安稳， 为列国之首，具有名望， 且为 以色列 家所归向的，有祸了！
AMOS|6|2|你们要过到 甲尼 察看， 从那里往 哈马 大城去， 又下到 非利士 人的 迦特 ， 你们比这些国更好吗？ 或是他们的疆界比你们的疆界广大呢？
AMOS|6|3|你们以为降祸的日子尚远， 却使残暴的统治 临近。
AMOS|6|4|“那些躺卧在象牙床上，舒身在榻上的， 吃群中的羔羊和棚里的牛犊。
AMOS|6|5|他们以琴瑟逍遥歌唱， 为自己作曲 ，像 大卫 一样；
AMOS|6|6|以大碗喝酒，用上等油抹身， 却不为 约瑟 所受的苦难忧伤；
AMOS|6|7|所以，现在这些人必首先被掳， 逍遥的欢宴必消失。”
AMOS|6|8|主耶和华指着自己起誓说： “我憎恶 雅各 的骄傲，厌弃他的宫殿； 我必将城和其中一切所有的都交给敌人。” 这是耶和华－万军之上帝说的 。
AMOS|6|9|那时，若一房之内剩下十个人，也都必死。
AMOS|6|10|死人的叔伯要把尸首抬到屋外焚烧，就问房屋内间的人说：“你那里还有别人吗？”他说：“没有。”又说：“不要作声，不可提耶和华的名。”
AMOS|6|11|看哪，耶和华发命令， 把大房子拆成碎片， 小屋子裂为小块。
AMOS|6|12|马岂能在岩石上奔跑？ 人岂能在那里 用牛耕种呢？ 你们却使公平变为苦胆， 使公义的果子变为茵蔯。
AMOS|6|13|你们这些喜爱 罗．底巴 的，自夸说： “我们不是凭自己的力量攻占了 加宁 吗？”
AMOS|6|14|耶和华─万军之上帝说： “ 以色列 家，看哪，我必兴起一国攻击你们； 他们必欺压你们， 从 哈马口 直到 亚拉巴 的河。”
AMOS|7|1|主耶和华指示我一件事，在春天作物刚长出时，看哪，主 造了蝗虫；看哪，这是王收割后长出的春天作物。
AMOS|7|2|蝗虫吃尽那地青草的时候，我说： “主耶和华啊，求你赦免； 因为 雅各 弱小， 他怎能站立得住呢？”
AMOS|7|3|耶和华对这事改变心意， 耶和华说：“这灾可以免了。”
AMOS|7|4|主耶和华又指示我一件事，看哪，主耶和华命火施行审判，火就吞灭深渊，烧尽产业。
AMOS|7|5|我就说： “主耶和华啊，求你止息； 因为 雅各 弱小， 他怎能站立得住呢？”
AMOS|7|6|耶和华对这事改变心意， 主耶和华说：“这灾也可免了。”
AMOS|7|7|他又指示我一件事，看哪，主手拿铅垂线，站立在依铅垂线建好的墙边。
AMOS|7|8|耶和华对我说：“ 阿摩司 ，你看见什么？”我说：“铅垂线。”主说： “看哪，我要在我子民 以色列 中 吊起铅垂线， 不再宽恕他们。
AMOS|7|9|以撒 的丘坛必荒凉， 以色列 的圣所必荒废； 我要起来用刀攻击 耶罗波安 的家。”
AMOS|7|10|伯特利 的祭司 亚玛谢 派人到 以色列 王 耶罗波安 那里，说：“ 阿摩司 在 以色列 家中图谋背叛你，他所说的一切话，这地不能承担；
AMOS|7|11|因为 阿摩司 这样说： ‘ 耶罗波安 必被刀杀， 以色列 百姓必被掳， 离开本地。’”
AMOS|7|12|于是 亚玛谢 对 阿摩司 说：“你这先见哪，要逃到 犹大 地，在那里过活 ，在那里说预言；
AMOS|7|13|却不要在 伯特利 再说预言，因为这里有王的圣所，有王的宫殿。”
AMOS|7|14|阿摩司 对 亚玛谢 说：“我原不是先知，也不是先知的门徒；我是牧人，是修剪桑树的。
AMOS|7|15|耶和华带领我，叫我不再牧放羊群，对我说：‘你去向我子民 以色列 说预言。’
AMOS|7|16|“现在你要听耶和华的话。 你说：‘不要向 以色列 说预言， 也不要向 以撒 家传讲 。’
AMOS|7|17|所以耶和华如此说： ‘你的妻子要在城中作妓女， 你的儿女要倒在刀下； 你的地必有人用绳子量了瓜分， 你自己必死在不洁净之地； 以色列 百姓必被掳， 离开本地。’”
AMOS|8|1|主耶和华又指示我一件事，看哪，有一筐夏天的果子。
AMOS|8|2|他说：“ 阿摩司 ，你看见什么？”我说：“一筐夏天的果子。”耶和华对我说： “我子民 以色列 的结局 到了， 我必不再宽恕他们。
AMOS|8|3|那日，宫殿里的诗歌要变为哀号 ； 必有许多尸首抛在各处， 安静无声。” 这是主耶和华说的。
AMOS|8|4|你们这些践踏贫穷人、 使这地困苦人衰败的， 当听这话！
AMOS|8|5|你们说：“初一几时过去， 我们好卖粮； 安息日几时过去， 我们好摆开谷物； 我们要把伊法变小， 把舍客勒变大， 以诡诈的天平欺哄人，
AMOS|8|6|用银子买贫寒人， 以一双鞋换贫穷人， 把坏的谷物卖给人。”
AMOS|8|7|耶和华指着 雅各 的骄傲起誓说： “他们这一切的行为，我必永远不忘。
AMOS|8|8|地岂不因这事震动？ 其中的居民岂不悲哀吗？ 全地必如 尼罗河 涨起， 如 埃及 的 尼罗河 涌起退落。
AMOS|8|9|“到那日， 我要使太阳在正午落下， 使这地在白昼黑暗。” 这是主耶和华说的。
AMOS|8|10|“我要使你们的节期变为悲哀， 你们一切的歌曲变为哀歌； 我要使众人腰束麻布， 头上光秃； 我要使这悲哀如丧独子， 其结局如悲痛的日子。
AMOS|8|11|“看哪，日子将到， 我必命饥荒降在地上； 人饥饿非因无饼，干渴非因无水， 而是因不听耶和华的话。” 这是主耶和华说的。
AMOS|8|12|他们必飘流，从这海到那海， 从北边到东边，往来奔跑， 寻求耶和华的话， 却寻不着。
AMOS|8|13|“当那日，少年和美貌的少女 必因干渴而发昏。
AMOS|8|14|那些指着 撒玛利亚 的罪孽 起誓的，说： ‘ 但 哪，我们指着你那里的神明起誓’， 又说：‘我们指着通往 别是巴 的路起誓’， 这些人都必仆倒，永不再起。”
AMOS|9|1|我看见主站在祭坛旁，说： “你要击打柱顶，使门槛震动， 要剪除众人当中为首的， 他们中最后的 ，我必用刀杀戮； 无一人能逃避，无一人能逃脱。
AMOS|9|2|“虽然他们挖透阴间， 我的手必从那里拉出他们； 虽然他们爬到天上， 我必从那里拿下他们；
AMOS|9|3|虽然藏在 迦密山 顶， 我必在那里搜寻，擒拿他们； 虽然离开我眼前藏在海底， 我必在那里命令蛇咬他们；
AMOS|9|4|虽然被仇敌掳去， 我也必在那里命令刀剑杀戮他们； 我必定睛在他们身上， 降祸不降福。”
AMOS|9|5|万军的主耶和华触摸地，地就融化， 凡住在地上的都必悲哀； 全地必如 尼罗河 涨起， 如同 埃及 的 尼罗河 落下。
AMOS|9|6|那在天上建造楼阁、 在地上奠定穹苍、 召唤海水、 使其倾倒在地面上的， 耶和华是他的名。
AMOS|9|7|耶和华说：“ 以色列 人哪， 我岂不是看你们如 古实 人吗？ 我岂不是领 以色列 人出 埃及 地， 也领 非利士 人出 迦斐托 ， 领 亚兰 人出 吉珥 吗？
AMOS|9|8|看哪，主耶和华的眼目 察看这有罪的国度， 要把它从地面上灭绝， 却不将 雅各 家灭绝净尽。” 这是耶和华说的。
AMOS|9|9|“看哪，我发命令， 使 以色列 家在万国中飘流， 好像人用筛子筛谷， 连一粒也不落在地上。
AMOS|9|10|我子民中所有的罪人， 就是那些说 ‘灾祸必不靠近，必不追上我们’的， 都必死在刀下。”
AMOS|9|11|“在那日，我必重建 大卫 倒塌的帐幕， 修补其中的缺口； 我必建立那遭破坏的， 重新修造，如古时一般，
AMOS|9|12|使 以色列 人接管 以东 所剩余的 和所有称为我名下的国。 这是耶和华说的，他要行这事。
AMOS|9|13|“看哪，日子将到， 耕种的必接续收割的， 踹葡萄的必接续撒种的； 大山要滴下甜酒， 小山也被漫过。” 这是耶和华说的。
AMOS|9|14|“我要使 以色列 被掳的子民归回； 他们要重修荒废的城镇， 居住在其中； 栽植葡萄园，喝其中所出的酒， 修造果园，吃其中的果子。
AMOS|9|15|我要将他们栽植于本地， 他们必不再从我所赐给他们的地上被拔出。” 这是耶和华－你的上帝说的。
OBAD|1|1|俄巴底亚 所见的异象。 我们从耶和华那里得到消息， 有使者被差往列国去： “起来吧， 我们要起来与 以东 争战！” 主耶和华论 以东 如此说：
OBAD|1|2|看哪，我要使你在列国中为最小， 被人大大藐视。
OBAD|1|3|你狂傲的心欺骗了你， 你住在岩穴， 居所在高处， 心里说： “谁能把我拉下来到地上呢？”
OBAD|1|4|你虽如鹰高飞， 在星宿之间搭窝， 我必从那里拉你下来。 这是耶和华说的。
OBAD|1|5|盗贼若来到你那里， 小偷夜间来到， 岂不是只偷他们所需要的吗？ 摘葡萄的若来到你那里， 岂不留下几串吗？ 你竟全然灭绝！
OBAD|1|6|以扫 遭到搜查， 他隐藏的宝物竟被寻出！
OBAD|1|7|与你结盟的都驱赶你，直到边界， 与你和好的欺骗你，胜过你， 吃你饭的人设下圈套陷害你─ 他却毫无聪明 。
OBAD|1|8|到那日， 我岂不从 以东 除灭智慧人？ 从 以扫山 除灭聪明人？ 这是耶和华说的。
OBAD|1|9|提幔 哪， 你的勇士必惊惶， 以致 以扫山 的人都被杀戮剪除。
OBAD|1|10|因你向兄弟 雅各 施暴， 你必蒙羞， 永被剪除。
OBAD|1|11|当陌生人掳掠 雅各 的财物， 当外邦人进入他的城门， 为 耶路撒冷 抽签分取财物的日子， 你竟站在一旁，像与他们同伙。
OBAD|1|12|你兄弟遭难的日子， 你不该瞪着眼看； 犹大 人被灭的日子， 你不该幸灾乐祸； 他们遭难的日子， 你不该说狂傲的话。
OBAD|1|13|我子民遭灾的日子， 你不该进他们的城门； 他们遭灾的日子， 你不该瞪着眼看他们受苦； 他们遭灾的日子， 你不该伸手抢他们的财物。
OBAD|1|14|他们遭难的日子， 你不该站在岔路口 剪除他们逃脱的人， 你不该交出他们的幸存者。
OBAD|1|15|耶和华的日子临近万国； 你所做的，人也必向你照样做， 你的报应必归到自己头上。
OBAD|1|16|你们在我圣山怎样喝了苦杯， 万国必照样不停地喝， 且喝且吞， 他们就必归于无有。
OBAD|1|17|但在 锡安山 必有逃脱的人， 那山必成为圣； 雅各 家必得原有的产业 。
OBAD|1|18|雅各 家必成为大火， 约瑟 家成为火焰； 以扫 家必如碎秸， 遭燃烧，被吞灭， 以扫 家必无幸存者。 这是耶和华说的。
OBAD|1|19|他们必得 尼革夫 和 以扫山 ， 得 谢非拉 ， 非利士 人之地， 他们必得 以法莲 地和 撒玛利亚 地， 得 便雅悯 和 基列 ；
OBAD|1|20|被掳的 以色列 大军 必得 迦南 人的地，直到 撒勒法 ， 在 西法拉 被掳的 耶路撒冷 人 必得 尼革夫 的城镇。
OBAD|1|21|必有一些解救者 上到 锡安山 ，审判 以扫山 ， 国度就归耶和华了。
JONAH|1|1|耶和华的话临到 亚米太 的儿子 约拿 ，说：
JONAH|1|2|“起来，到 尼尼微 大城去，向其中的居民宣告，因为他们的恶已达到我面前。”
JONAH|1|3|约拿 却起身，逃往 他施 去躲避耶和华。他下到 约帕 ，遇见一条船要往 他施 去。 约拿 付了船费，就上船，与船上的人同往 他施 ，为要躲避耶和华。
JONAH|1|4|耶和华在海上刮起大风，海就狂风大作，船几乎破裂。
JONAH|1|5|水手都惧怕，各人哀求自己的神明。他们把船上的货物抛进海里，为要减轻载重。 约拿 却下到舱底，躺卧沉睡。
JONAH|1|6|船长到他那里，对他说：“你怎么还在沉睡呢？起来，求告你的神明，或者神明顾念我们，使我们不致灭亡。”
JONAH|1|7|船上的人彼此说：“来吧，我们来抽签，看看这灾难临到我们是因谁的缘故。”于是他们就抽签，抽出 约拿 来。
JONAH|1|8|他们对 约拿 说：“请你告诉我们，这灾难临到我们是因谁的缘故呢？你做什么行业？你从哪里来？你是哪一国的人？属哪一族？”
JONAH|1|9|他说：“我是 希伯来 人，我敬畏耶和华，天上的上帝，他创造了沧海和陆地。”
JONAH|1|10|那些人就大大惧怕，对他说：“你做的是什么事呢？”原来他们已经知道他在躲避耶和华，因为他告诉了他们。
JONAH|1|11|海浪越来越汹涌，他们就问他说：“我们当向你做什么，才能使海浪平静呢？”
JONAH|1|12|他对他们说：“你们把我抬起来，抛进海里，海就会平静了；我知道你们遭遇这大风浪是因我的缘故。”
JONAH|1|13|然而那些人竭力划桨，想要把船靠回陆地，却是不能；因风浪愈来愈大，扑向他们。
JONAH|1|14|于是他们求告耶和华说：“耶和华啊，求求你不要因这人的性命使我们灭亡，不要使流无辜人血的罪归给我们；因为你－耶和华随自己的旨意行事。”
JONAH|1|15|他们把 约拿 抬起来，抛进海里，海的狂浪就平息了。
JONAH|1|16|那些人就大大惧怕耶和华，向耶和华献祭许愿。
JONAH|1|17|耶和华安排一条大鱼吞下 约拿 ， 约拿 在鱼腹中三日三夜。
JONAH|2|1|约拿 在鱼腹中向耶和华－他的上帝祷告，
JONAH|2|2|说： “我在患难中求告耶和华， 他就应允我； 我从阴间的深处呼求， 你就俯听我的声音。
JONAH|2|3|你将我投下深渊， 直到海心； 大水环绕我， 你的波浪洪涛漫过我身。
JONAH|2|4|我说：‘我从你眼前被驱逐， 然而我仍要仰望你的圣殿。’
JONAH|2|5|众水环绕我，几乎淹没我； 深渊围住我； 海草缠绕我的头。
JONAH|2|6|我下沉到山的根基， 地的门闩将我永远关住。 耶和华－我的上帝啊， 你却将我的性命从地府里救出来。
JONAH|2|7|我心灵发昏时， 就想起耶和华。 我的祷告进入你的圣殿， 达到你面前。
JONAH|2|8|那信奉虚无神明 的人， 丢弃自己的慈爱；
JONAH|2|9|但我要以感谢的声音向你献祭。 我所许的愿，我必偿还。 救恩出于耶和华。”
JONAH|2|10|耶和华吩咐那鱼，鱼就把 约拿 吐在陆地上。
JONAH|3|1|耶和华的话第二次临到 约拿 ，说：
JONAH|3|2|“起来，到 尼尼微 大城去，把我告诉你的信息向其中的居民宣告。”
JONAH|3|3|约拿 就照耶和华的话起来，到 尼尼微 去。 尼尼微 是一座极大的城，约有三天的路程。
JONAH|3|4|约拿 进城，走了一天，宣告说：“再过四十天， 尼尼微 要倾覆了！”
JONAH|3|5|尼尼微 人就信服上帝，宣告禁食，从最大的到最小的都穿上麻衣。
JONAH|3|6|这消息传到 尼尼微 王那里，他就从宝座起来，脱下朝服，披上麻布，坐在灰中。
JONAH|3|7|他叫人通告 尼尼微 全城，说：“王和大臣有令，人、畜、牛、羊都不可尝任何东西，不可吃，也不可喝水。
JONAH|3|8|人与牲畜都要披上麻布，切切求告上帝。各人要回转离开恶道，离弃自己掌中的残暴。
JONAH|3|9|谁知道上帝也许会回心转意，不发烈怒，使我们不致灭亡。”
JONAH|3|10|上帝察看他们的行为，见他们离开恶道，上帝就改变心意，原先所说要降与他们的灾难，他不降了。
JONAH|4|1|这事令 约拿 大大不悦，甚至发怒。
JONAH|4|2|他就向耶和华祷告，说：“耶和华啊，这不就是我仍在本国的时候所说的吗？我知道你是有恩惠，有怜悯的上帝，不轻易发怒，有丰盛的慈爱，并且会改变心意，不降那灾难。我就是因为这样，才急速逃往 他施 去的呀！
JONAH|4|3|耶和华啊，现在求你取走我的性命吧！因为我死了比活着更好。”
JONAH|4|4|耶和华说：“你这样发怒，对吗？”
JONAH|4|5|约拿 出城，坐在城的东边，在那里为自己搭了一座棚。他坐在棚子的荫下，要看看城里会发生什么事。
JONAH|4|6|耶和华上帝安排了一棵蓖麻，使它生长高过 约拿 ，影子遮盖他的头，使他免受苦难； 约拿 因这棵蓖麻大大欢喜。
JONAH|4|7|次日黎明，上帝却安排一条虫来咬这蓖麻，以致枯干。
JONAH|4|8|太阳出来的时候，上帝安排炎热的东风，太阳曝晒 约拿 的头，使他发昏，他就为自己求死，说：“我死了比活着更好！”
JONAH|4|9|上帝对 约拿 说：“你因这棵蓖麻这样发怒，对吗？”他说：“我发怒以至于死，都是对的！”
JONAH|4|10|耶和华说：“这棵蓖麻你没有为它操劳，也不是你使它长大的；它一夜生长，一夜枯死，你尚且爱惜；
JONAH|4|11|何况这 尼尼微 大城，其中不能分辨左右手的就有十二万多人，还有许多牲畜，我岂能不爱惜呢？”
MIC|1|1|当 犹大 王 约坦 、 亚哈斯 、 希西家 在位的时候，耶和华的话临到 摩利沙 人 弥迦 ，他见到有关 撒玛利亚 和 耶路撒冷 的异象。
MIC|1|2|万民哪，你们都要听！ 地和其上所有的，要留心听！ 主耶和华要从他的圣殿 指证你们的不是。
MIC|1|3|看哪，耶和华从他的居所出来， 降临步行地之高处。
MIC|1|4|众山在他底下熔化， 诸谷崩裂， 如蜡熔在火中， 如水冲下山坡。
MIC|1|5|这都是因 雅各 的罪过， 因 以色列 家的罪恶。 雅各 的罪过在哪里呢？ 岂不是在 撒玛利亚 吗？ 犹大 的丘坛在哪里呢？ 岂不是在 耶路撒冷 吗？
MIC|1|6|因此，我必使 撒玛利亚 变为田野的废墟， 用以栽植葡萄； 我必把它的石头倒在山谷， 掀开它的地基。
MIC|1|7|城里一切雕刻的偶像必被打碎， 行淫的赏金全被火烧， 我要毁灭它的一切偶像； 因为从妓女的赏金积聚而来的， 它们仍归为妓女的赏金。
MIC|1|8|为此我要大声哀号， 赤身赤脚行走； 我要呼号如野狗， 哀鸣如鸵鸟。
MIC|1|9|因为 撒玛利亚 的创伤无法医治， 蔓延到 犹大 ， 到了我百姓的城门， 直达 耶路撒冷 。
MIC|1|10|不要在 迦特 宣扬 这事， 千万不要哭泣； 要在 伯．亚弗拉 翻滚于灰尘 中。
MIC|1|11|沙斐 的居民哪，要赤身羞愧地经过， 撒南 的居民不敢出门， 伯．以薛 哀哭，不再支持你们。
MIC|1|12|玛律 的居民心甚忧急，切望得着福气， 因为灾祸已从耶和华那里临到 耶路撒冷 的城门。
MIC|1|13|拉吉 的居民哪，要用快马 套车； 锡安 的罪由你而起， 以色列 的罪过在你那里显出。
MIC|1|14|因此，你要将送别礼送到 摩利设．迦特 ； 亚革悉 的众家族必用诡诈 待 以色列 诸王。
MIC|1|15|玛利沙 的居民哪， 我必使抢夺者来到你这里； 以色列 的贵族 必来到 亚杜兰 。
MIC|1|16|犹大 啊，为了你所喜爱的儿女， 你要剪发，剃光头， 要使你的头光秃，如同秃鹰， 因为他们被掳去离开你了。
MIC|2|1|祸哉，那些在床上图谋罪孽、筹划恶事的人！ 天一亮，他们因手中有能力就去行恶。
MIC|2|2|他们看上田地就占据， 贪图房屋便夺取； 他们欺压户主和他的家庭， 霸占人和他的产业。
MIC|2|3|所以耶和华如此说： 看哪，我筹划灾祸降与这家族； 这灾祸在你们颈项上无法解脱， 你们也不能昂首而行， 因为这是灾祸的时刻。
MIC|2|4|到那日，必有人为你们唱诗歌， 用悲哀的哀歌哀号，说： “我们全然败落， 我百姓的产业易主了！ 耶和华竟然使它离开我， 我们的田地为悖逆的人所瓜分了！”
MIC|2|5|因此，你必无人能在耶和华的会中 抽签拉绳 。
MIC|2|6|他们传讲说：“不可传讲； 人都不可传讲这些事， 羞辱不会临到我们。”
MIC|2|7|雅各 家啊，可这么说吗 ？ 耶和华没有耐心吗？ 这些事是他所行的吗？ 我的言语岂不是与行动正直的人有益吗？
MIC|2|8|然而，近来我的百姓兴起如仇敌。 你们剥去那些安然行路、不愿打仗之人身上的外衣，
MIC|2|9|把我百姓中的妇人从安乐家中赶出， 又将我的荣耀从她们孩子身上永远夺去。
MIC|2|10|起来，走吧！ 这里并非安歇之处； 因为不洁净带来毁坏， 且是大大的毁坏。
MIC|2|11|若有人心存虚假，用谎言说 ： “我向你们传讲可得清酒和烈酒 ”， 那人就必作这百姓的传讲者。
MIC|2|12|雅各 家啊，我定要聚集你们， 定要召集 以色列 的余民， 把他们安置在一处，如 波斯拉 的羊， 又如草场上的羊群， 人数众多，大大喧哗。
MIC|2|13|开路的在他们前面上去， 直闯过城门，从城门出去； 他们的王在前面行， 耶和华在他们的前头。
MIC|3|1|于是我说： 雅各 的领袖， 以色列 家的官长啊， 你们要听！ 你们岂不知道公平吗？
MIC|3|2|你们恶善好恶， 剥我百姓 身上的皮， 从他们的骨头上剔肉，
MIC|3|3|你们吃我百姓的肉， 剥他们的皮， 打断他们的骨头， 如切块 下锅， 如釜中的肉。
MIC|3|4|到了遭灾的时候，这些人要哀求耶和华， 他却不应允他们。 那时，因他们所行的恶， 他必转脸离开他们。
MIC|3|5|论到使我百姓走入歧途的先知， 他们牙齿有所嚼，就呼喊说：“平安！” 谁不给他们吃，就扬言攻击他， 耶和华如此说：
MIC|3|6|你们因此必遭遇黑夜，看不到异象； 遭遇幽暗，无法占卜。 太阳必向先知沉落， 白昼转为黑暗。
MIC|3|7|先见必抱愧， 占卜的必蒙羞， 他们全都捂着胡须， 因为上帝不应允他们。
MIC|3|8|至于我，我藉耶和华的灵， 满有能力、公平和勇气， 可向 雅各 述说他的过犯， 向 以色列 指出他的罪恶。
MIC|3|9|当听这话， 雅各 家的领袖， 以色列 家的官长啊！ 你们厌弃公平， 在一切事上屈枉正直；
MIC|3|10|以血建立 锡安 ， 以罪孽建造 耶路撒冷 。
MIC|3|11|城里的领袖为贿赂行审判， 祭司为酬劳施训诲， 先知为银钱行占卜； 他们却倚赖耶和华，说： “耶和华不是在我们中间吗？ 灾祸必不临到我们。”
MIC|3|12|因此，为你们的缘故， 锡安 要被耕种像一块田地， 耶路撒冷 要变为废墟， 这殿的山必如丛林的高处。
MIC|4|1|末后的日子， 耶和华殿的山必坚立， 超乎诸山，高举过于万岭； 万民都要流归这山。
MIC|4|2|必有许多民族前往，说： “来吧，我们登耶和华的山， 到 雅各 上帝的殿。 他必将他的道指教我们， 我们也要行他的路。” 因为教诲必出于 锡安 ， 耶和华的言语必出于 耶路撒冷 。
MIC|4|3|他必在许多民族中施行审判， 为远方强盛的国断定是非。 他们要将刀打成犁头， 把枪打成镰刀。 这国不举刀攻击那国， 他们也不再学习战事。
MIC|4|4|人人都要坐在自己的葡萄树 和无花果树下， 无人使他们惊吓； 这是万军之耶和华亲口说的。
MIC|4|5|万民都奉自己神明的名行事， 我们却要奉耶和华－我们上帝的名而行， 直到永永远远。
MIC|4|6|耶和华说：在那日， 我必聚集瘸腿的， 召集被赶逐的， 以及我所惩治的人。
MIC|4|7|我要使瘸腿的成为余民， 使被赶到远方的成为强盛之国。 耶和华要在 锡安山 作王治理他们， 从今直到永远。
MIC|4|8|你， 以得台 ， 锡安 的山冈啊， 先前的权柄必归给你， 耶路撒冷 的国权必将归还。
MIC|4|9|现在，你为何大声呼喊呢？ 你中间没有君王， 你的谋士灭绝， 以致疼痛抓住你， 如临产的妇人吗？
MIC|4|10|锡安 哪，你要疼痛生产， 仿佛临产的妇人； 因你必从城里出来，住在田野； 你要到 巴比伦 去， 在那里，你要蒙解救， 在那里，耶和华必救赎你 脱离仇敌的手掌。
MIC|4|11|现在，许多国家聚集攻击你，说： “让 锡安 被玷污！ 让我们亲眼看到！”
MIC|4|12|他们却不知道耶和华的意念， 也不明白他的筹算， 他聚集他们， 像把禾捆聚到禾场。
MIC|4|13|锡安 哪，起来踹谷吧！ 我必使你的角成为铁， 使你的蹄成为铜。 你必打碎许多民族， 将他们的财宝献给耶和华， 将他们的财富献给全地的主。
MIC|5|1|成群的民 哪，现在要聚集成队； 仇敌前来围攻我们， 要用杖击打 以色列 领袖的脸颊。
MIC|5|2|伯利恒 的 以法他 啊， 你在 犹大 诸城中虽小， 将来必有一位从你那里出来， 在 以色列 中为我作掌权者； 他的根源自亘古，从太初就有。
MIC|5|3|因此，耶和华要将 以色列 人交给敌人， 直到临产的妇人生下孩子； 那时，他其余的弟兄 必回到 以色列 人那里。
MIC|5|4|他必倚靠耶和华的大能， 倚靠耶和华－他上帝之名的威严， 站立并牧养， 使他们安然居住； 因为现在他必尊大， 直到地极。
MIC|5|5|这位就是和平 。 当 亚述 侵入我们领土， 践踏我们宫殿时， 我们就立七个牧者， 八个领袖攻击它。
MIC|5|6|他们要用刀剑毁坏 亚述 地 和 宁录 地的关口 。 当 亚述 侵入我们领土， 践踏我们边境时， 他必拯救我们。
MIC|5|7|雅各 的余民 必在许多民族中， 如从耶和华降下的露水， 又如甘霖降在草上； 他们不倚靠人， 也不仰赖世人。
MIC|5|8|雅各 的余民必在列国中， 在许多民族中， 如林间百兽中的狮子， 又如少壮狮子在羊群中； 他若经过就必践踏撕裂， 无人搭救。
MIC|5|9|愿你的手举起，高过敌人！ 愿你的仇敌都被剪除！
MIC|5|10|耶和华说：到那日， 我必从你中间剪除马匹， 毁坏战车；
MIC|5|11|除灭你国中的城镇， 拆毁你一切的堡垒；
MIC|5|12|除掉你手中的邪术， 你那里不再有占卜的人。
MIC|5|13|我必从你中间除灭雕刻的偶像和柱像， 你就不再跪拜自己手所造的；
MIC|5|14|我必从你中间拔除 亚舍拉 ， 毁灭你的城镇；
MIC|5|15|我必在怒气和愤怒中 报应那不听从我的列国。
MIC|6|1|当听耶和华说的话： 起来，向山岭争辩， 使冈陵听见你的声音。
MIC|6|2|山岭啊，要听耶和华的指控！ 大地永久的根基啊，要听！ 因耶和华控告他的百姓， 与 以色列 争辩。
MIC|6|3|“我的百姓啊，我向你做了什么呢？ 我在什么事上使你厌烦？ 你回答我吧！
MIC|6|4|我曾将你从 埃及 地领出来， 从为奴之家救赎你， 我差遣 摩西 、 亚伦 和 米利暗 在你前面带领。
MIC|6|5|我的百姓啊，当记念从前 摩押 王 巴勒 如何筹算， 比珥 的儿子 巴兰 如何回应他， 当记念从 什亭 到 吉甲 所发生的事， 好使你们明白耶和华公义的作为。”
MIC|6|6|“我朝见耶和华， 在至高上帝面前跪拜，当献上什么呢？ 难道献一岁的牛犊为燔祭来朝见他吗？
MIC|6|7|耶和华岂喜悦千千的公羊， 或是万万的油河吗？ 我岂可为自己的过犯献我的长子， 为自己的罪恶献我所亲生的吗？”
MIC|6|8|世人哪，耶和华已指示你何为善。 他向你所要的是什么呢？ 只要你行公义，好怜悯， 存谦卑的心与你的上帝同行。
MIC|6|9|耶和华向这城呼叫 ─看重你的名是真智慧 ─ 你们当听惩罚 和派定惩罚的人 。
MIC|6|10|恶人家中不是仍有不义之财 和惹人生气的变小了的伊法吗？
MIC|6|11|我若用不公道的天平 和袋中诡诈的法码， 岂可算为清白呢？
MIC|6|12|城里的有钱人遍行残暴， 其中的居民说谎话， 口中的舌头尽是诡诈。
MIC|6|13|因此，我也击打你，使你受伤 ， 因你的罪恶使你受惊骇。
MIC|6|14|你要吃，却吃不饱， 你的肚子仍是空空。 你必被挪去，不得逃脱； 如有逃脱的，我必交给刀剑。
MIC|6|15|你撒种，却不得收割； 踹橄榄，却不得油抹身； 有新酒，却不得酒喝。
MIC|6|16|因为你遵守 暗利 的规条， 行 亚哈 家一切所行的， 顺从他们的计谋； 因此，我必使你荒凉， 使你的居民遭人嗤笑， 你们也必担当我百姓的羞辱。
MIC|7|1|我有祸了！我好像夏日收割后的果子， 又如收成之后剩余的葡萄， 没有一挂可吃的， 也没有我心所渴想初熟的无花果。
MIC|7|2|地上的虔诚人灭尽了， 人世间已无正直的人； 他们都埋伏，为要流人的血， 用罗网猎取自己的弟兄。
MIC|7|3|他们双手善于作恶， 君王和审判官都索取贿赂； 位高的人吐出心中的欲望， 彼此勾结 。
MIC|7|4|他们当中最好的，不过像蒺藜； 最正直的，不过如荆棘篱笆。 你守候的日子，惩罚已经来到， 他们必扰乱不安。
MIC|7|5|不可倚赖邻舍， 不可信靠密友； 甚至对躺在你怀中的妻子 也要守住你的口。
MIC|7|6|因为儿子藐视父亲， 女儿抵挡母亲， 媳妇抗拒婆婆， 人的仇敌就是自己家里的人。
MIC|7|7|至于我，我要仰望耶和华， 等候那救我的上帝； 我的上帝必应允我。
MIC|7|8|我的仇敌啊，不要向我夸耀。 我虽跌倒，仍要起来； 虽坐在黑暗里，耶和华却作我的光。
MIC|7|9|我要承受耶和华的恼怒， 直到他为我辩护，为我伸冤， 因我得罪了他； 他要领我进入光明， 我必得见他的公义。
MIC|7|10|那时我的仇敌看见这事就羞愧， 他曾对我说：“耶和华－你的上帝在哪里？” 我必亲眼见他遭报， 现在，他必被践踏，如同街上的泥土。
MIC|7|11|你的城墙重修的日子到了！ 到那日，边界必扩展。
MIC|7|12|到那日，人必从 亚述 ， 从 埃及 的城镇， 从 埃及 到 大河 ， 从这海到那海， 从这山到那山， 都归到你这里。
MIC|7|13|然而，因居民的缘故， 为了他们行事的结果。 这地必然荒凉。
MIC|7|14|求你在 迦密 的树林中， 以你的杖牧放你独居的民， 你产业中的羊群； 愿他们像古时一样， 牧放在 巴珊 和 基列 。
MIC|7|15|我要显奇事给他们看， 好像出 埃及 地的时候一样。
MIC|7|16|列国看见，虽大有势力仍觉惭愧； 他们必用手捂口，掩耳不听。
MIC|7|17|他们要舔土如蛇， 又如地上爬行的动物， 战战兢兢离开他们的营寨； 他们必畏惧耶和华─我们的上帝， 也必因你而害怕。
MIC|7|18|有哪一个神明像你，赦免罪孽， 饶恕他产业中余民的罪过？ 他不永远怀怒，喜爱施恩。
MIC|7|19|他 必转回怜悯我们， 把我们的罪孽踏在脚下。 你必将他们 一切的罪投于深海。
MIC|7|20|你必按古时向我们列祖起誓的话， 以信实待 雅各 ， 向 亚伯拉罕 施慈爱。
NAH|1|1|论 尼尼微 的默示， 伊勒歌斯 人 那鸿 所见异象的书。
NAH|1|2|耶和华是忌邪 、报应的上帝。 耶和华施报应，大有愤怒； 耶和华向他的敌人报应， 向他的仇敌怀怒。
NAH|1|3|耶和华不轻易发怒，大有能力， 但耶和华万不以有罪的为无罪。 他的道路在旋风和暴风之中， 云彩为他脚下的尘土。
NAH|1|4|他斥责海，使海枯干， 使一切江河干涸。 巴珊 和 迦密 衰残， 黎巴嫩 的花草也衰残了。
NAH|1|5|大山因他震动， 小山也都融化； 大地在他面前突起， 世界和住在其间的也都如此。
NAH|1|6|他发愤恨，谁能立得住呢？ 他发烈怒，谁能当得起呢？ 他的愤怒如火倾泄而出， 磐石因他崩裂。
NAH|1|7|耶和华本为善， 在患难的日子为人的保障， 并且认识那些投靠他的人；
NAH|1|8|但他必以涨溢的洪水淹没其地方 ， 又驱逐仇敌进入黑暗。
NAH|1|9|你们筹划何种计谋攻击耶和华呢？ 他必终结一切， 仇敌 不会再度兴起。
NAH|1|10|你们像杂乱的荆棘， 像喝醉了的人， 又如枯干的碎秸，全然烧灭。
NAH|1|11|有一人从你那里出来， 图谋邪恶，设恶计攻击耶和华。
NAH|1|12|耶和华如此说： “他们虽然势力强大，人数众多， 也要被剪除，归于无有。 我虽曾使你受苦， 却不再使你受苦。
NAH|1|13|现在，我要从你身上折断他的轭， 解开捆绑你的绳索。”
NAH|1|14|耶和华已经发命令，指着你说： “你的名下必不再留后； 我要从你神明的庙中除灭雕刻的偶像和铸造的偶像， 我必因你的卑贱，为你预备坟墓。”
NAH|1|15|看哪，山上有报佳音、传平安之人的脚踪。 犹大 啊，守你的节期， 还你的愿吧！ 因为恶人不再侵犯你， 他已灭绝净尽了。
NAH|2|1|那打碎你的人 上到你面前。 要看守堡垒，把守道路， 要挺起腰来，大大使力。
NAH|2|2|耶和华复兴 雅各 的荣华， 像复兴 以色列 的荣华； 因为蹂躏者曾经蹂躏他们， 毁坏了他们的葡萄枝。
NAH|2|3|他勇士的盾牌是红的， 精兵都穿朱红衣服。 在预备打仗的日子， 战车上的铁闪烁如火 ， 柏木的枪杆也已举起 ；
NAH|2|4|战车在街上疾行， 在广场上来往奔驰， 形状如火把， 飞驰如闪电。
NAH|2|5|他 招聚他的贵族； 他们前行时绊跌， 速上城墙， 预备屏障。
NAH|2|6|河闸开放， 宫殿冲没。
NAH|2|7|这是命定之事： 王后赤身被掳 ， 宫女捶胸， 哀鸣如鸽子。
NAH|2|8|尼尼微 自古以来 如同聚水的池子； 现在居民都在逃跑 。 “站住！站住！” 却无人回转。
NAH|2|9|你们抢夺金子吧！ 你们抢夺银子吧！ 因为所积蓄的无穷， 华美的宝器无数。
NAH|2|10|荒芜，荒凉，全然荒废， 人心害怕，双膝颤抖， 腰部疼痛，脸都变色。
NAH|2|11|狮子的洞， 幼狮喂养之处在哪里呢？ 公狮、母狮、小狮出入， 无人使它们惊吓之地在哪里呢？
NAH|2|12|公狮撕碎的足够给幼狮吃， 又为母狮掐死猎物， 把猎物塞满它的洞穴， 把撕碎的装满它的窝。
NAH|2|13|看哪，我与你为敌，将它的战车 焚烧成烟，刀剑必吞灭你的少壮狮子；我必从地上除灭你的猎物，你使者的声音必不再听见。这是万军之耶和华说的。
NAH|3|1|祸哉！这流人血的城， 欺诈连连，抢夺充斥， 掳掠的事总不止息。
NAH|3|2|鞭声响亮，车轮轰轰， 马匹跳跃，战车奔腾；
NAH|3|3|骑兵争先，刀剑发光， 枪矛闪烁，被杀的甚多， 尸首成堆，尸骸无数， 人因尸骸而绊跌，
NAH|3|4|都因那美貌的妓女多有淫行， 惯行邪术， 藉淫行诱惑 列国， 用邪术诱惑万族。
NAH|3|5|看哪，我与你为敌， 掀开你的下摆，蒙在你脸上， 使列邦看见你的赤体， 使列国观看你的羞辱。 这是万军之耶和华说的。
NAH|3|6|我必将可憎污秽之物抛在你身上， 使你被藐视，为众人所观看。
NAH|3|7|凡看见你的，都必逃离你，说： “ 尼尼微 荒凉了！有谁为你悲伤呢？ 我何处找到安慰你的人呢？”
NAH|3|8|你能胜过 挪亚们 吗？ 它坐落在众河之间， 周围有水， 海 作它的城郭， 海 作它的城墙。
NAH|3|9|古实 和 埃及 是它的力量， 没有穷尽， 弗 人和 路比 人是它的帮手。
NAH|3|10|但它被流放，被人掳去， 它的婴孩也被摔碎在各街头； 人为它的贵族抽签， 它的权贵都被锁链锁住。
NAH|3|11|你也必喝醉，昏迷错乱， 并因仇敌的缘故寻求庇护。
NAH|3|12|你一切的堡垒必如无花果树上初熟的果子， 一经摇动，就落在想吃的人口中。
NAH|3|13|看哪，你中间的士兵是妇女， 你国中的关口向仇敌敞开， 你的门闩被火焚烧。
NAH|3|14|你要打水预备受困； 要加强防御， 取土踹泥， 做成砖模。
NAH|3|15|在那里，火要吞灭你， 刀必杀戮你， 如蝻子般吞灭你。 你人数增多如蝻子， 增多如蝗虫吧！
NAH|3|16|你增添商贾，多过天上的星宿； 如蝻子蜕皮飞去。
NAH|3|17|你的领袖多如蝗虫， 你的将军仿佛成群的蝗虫； 天凉时齐落在篱笆上， 太阳一出就飞去， 人不知道落在何处。
NAH|3|18|亚述 王啊， 你的牧人睡觉， 你的贵族躺卧 ， 你的百姓散在山间， 无人招聚。
NAH|3|19|你的损伤并未减轻， 你的伤痕极其重大。 凡听见这消息的人都因你拍掌。 有谁没有时常遭受你的暴行呢？
HAB|1|1|哈巴谷 先知所看见的默示。
HAB|1|2|耶和华啊，我呼求， 你不应允，要到几时呢？ 我向你呼喊“暴力！” 你还不拯救？
HAB|1|3|你为何使我看见罪孽？ 你为何坐视奸恶呢？ 毁灭和凶暴在我面前， 争执与纷争不断发生。
HAB|1|4|因此律法无效， 公理从未彰显。 因恶人围困义人， 所以公理遭受扭曲。
HAB|1|5|你们要向列国观看 ，注意看， 要惊奇，再惊奇！ 因为在你们的日子，有一件事发生 ， 尽管有人说了，你们还是不信。
HAB|1|6|看哪，我必兴起 迦勒底 人， 就是那残忍暴躁之民，通行遍地， 霸占不属自己的住处。
HAB|1|7|他威武可畏， 审判与威权都由他而出。
HAB|1|8|他的马比豹更快， 比晚上 的野狼更猛。 他的战马跳跃， 他的战马从远方而来 ； 他们飞跑，如鹰急速抓食，
HAB|1|9|都为施行残暴而来， 他们的脸面向东 ， 聚集俘虏，多如尘沙。
HAB|1|10|他讥诮列王， 嘲讽领袖， 嗤笑一切堡垒， 堆土攻取它。
HAB|1|11|那时，他如风猛然扫过， 他背叛，显为有罪； 他以自己的力量为神明。
HAB|1|12|耶和华－我的上帝，我的圣者啊， 你不是从亘古就有吗？ 我们必不致死。 耶和华啊，你派他为要行审判； 磐石啊，你立他为要惩治人。
HAB|1|13|你的眼目清洁， 不看邪恶，也不看奸恶， 为何你却看着人行诡诈呢？ 恶人吞灭比自己公义的人， 为何你保持沉默呢？
HAB|1|14|你为何使人如海中的鱼， 又如无人管辖的爬行动物呢？
HAB|1|15|他用钩子把他们全拉上来， 用罗网捕获他们， 拉渔网聚集他们。 因此，他欢喜快乐，
HAB|1|16|向罗网献祭， 向渔网烧香； 因为他藉此得丰盛的收获 与肥美的食物。
HAB|1|17|但他岂可因此屡屡倒空罗网 ， 时常杀戮列国的人，毫不顾惜呢？
HAB|2|1|我要站在我的了望台， 立在城楼 上观看， 看耶和华要对我说什么， 我可用什么话向他诉冤。
HAB|2|2|耶和华回答我，说： 将这默示清楚地写在看板上， 使人容易朗读 。
HAB|2|3|因为这默示有一定日期， 论及终局，绝不落空。 它虽然耽延，你要等候； 因为它必临到，不再迟延。
HAB|2|4|看哪，恶人自高自大，心不正直； 惟义人必因他的信得生 。
HAB|2|5|他因酒诡诈、 狂傲、不安于位； 他张开喉咙 ，好像阴间， 如死亡不能知足， 他聚集万国， 招聚万民全归自己。
HAB|2|6|这些人岂不都要提起诗歌和俗语，嘲讽他说： 祸哉！你增添不属自己的财物， 靠押金发财，要到几时呢？
HAB|2|7|咬伤你的 岂不忽然兴起， 扰害你的岂不突然崛起， 你就成为他们的掳物吗？
HAB|2|8|因你抢夺许多国家， 流人的血，向土地、城镇和全城的居民施行残暴， 各国残存之民都必抢夺你。
HAB|2|9|祸哉！那为本家积蓄不义之财、 在高处搭窝、指望得免灾祸的人！
HAB|2|10|你图谋剪除许多民族，犯了罪， 使自己的家蒙羞，自害己命。
HAB|2|11|墙里的石头要呼叫， 屋内的栋梁必应声。
HAB|2|12|祸哉！那以鲜血建城、 以罪孽造镇的人！
HAB|2|13|看哪，这不都是 出于万军之耶和华吗？ 万民劳碌得来的被火焚烧， 万族辛苦建造的，归于虚空。
HAB|2|14|全地都必认识耶和华的荣耀， 好像水充满海洋一般。
HAB|2|15|祸哉！那给邻舍酒喝，加上毒物 ， 使人喝醉，为要看见他们下体的人！
HAB|2|16|你满受羞辱，不得荣耀； 你也喝吧，显明你是未受割礼的 ！ 耶和华右手的杯必传到你那里， 你的荣耀就变为羞辱。
HAB|2|17|黎巴嫩 所受的残暴必淹没你， 野兽所遭遇的毁灭使你惊吓 ； 因你流人的血， 向土地、城镇和全城的居民施行残暴。
HAB|2|18|偶像有什么益处呢？ 制造者雕刻它， 铸成偶像，作虚假的教师； 制造者倚靠的是自己所做的哑巴偶像。
HAB|2|19|祸哉！那对木头说“醒起”， 对哑巴石头说“起来”的人！ 偶像岂能教导人呢？ 看哪，它以金银包裹，其中并无气息。
HAB|2|20|惟耶和华在他的圣殿中， 全地都当在他面前肃静。
HAB|3|1|哈巴谷 先知的祷告，调用流离歌。
HAB|3|2|耶和华啊，我听见你的名声； 耶和华啊，我惧怕你的作为。 求你在这些年间 复兴你的作为， 在这些年间将它显明出来 ； 在发怒的时候以怜悯为念。
HAB|3|3|上帝从 提幔 而来， 圣者从 巴兰山 临到； 他的荣光遮蔽诸天， 颂赞遍满全地。
HAB|3|4|他的辉煌如同日光， 从他手里发出光芒， 那里 隐藏他的能力。
HAB|3|5|在他前面有瘟疫流行， 在他脚下有热症发出。
HAB|3|6|他站立，震动 大地， 他观看，震动列国。 永久的山崩裂， 长存的岭塌陷， 他的作为与古时一样。
HAB|3|7|我见 古珊 的帐棚遭难， 米甸 地的幔子动摇。
HAB|3|8|耶和华啊，你岂是向江河发怒， 向江河生气， 向海洋发烈怒吗？ 你骑在马上， 坐在得胜的战车上，
HAB|3|9|你的弓全然显露 ， 箭是发誓的言语 ； 你以江河分开大地。
HAB|3|10|山岭见你，无不战抖； 大水泛滥而过， 深渊发声， 汹涌翻腾 。
HAB|3|11|因你的箭射出光芒， 你的枪闪出光耀， 日月都停在原处。
HAB|3|12|你发怒遍行大地， 以怒气责打列国，如打谷一般。
HAB|3|13|你出来拯救你的百姓， 拯救你的受膏者； 你打破恶人之家的头， 暴露其根基，直到颈项 。
HAB|3|14|你以其戈矛刺透他战士的头； 他们如旋风将我 刮散， 他们喜爱暗中吞吃困苦的人。
HAB|3|15|你骑马践踏海， 践踏汹涌的大水。
HAB|3|16|我听见这声音，身体战兢， 嘴唇发颤， 骨中朽烂， 在所立之处战兢 ； 但我安静等候 灾难之日临到那上来侵犯我们的民 。
HAB|3|17|虽然无花果树不发旺， 葡萄树不结果， 橄榄树也不收成， 田地不出粮食， 圈中绝了羊， 棚内也没有牛；
HAB|3|18|然而，我要因耶和华欢欣， 因救我的上帝喜乐。
HAB|3|19|主耶和华是我的力量， 他使我的脚快如母鹿， 又使我稳行在高处。 这歌交给圣咏团长，用丝弦的乐器。
ZEPH|1|1|当 亚们 的儿子 犹大 王 约西亚 在位的时候，耶和华的话临到 希西家 的玄孙， 亚玛利雅 的曾孙， 基大利 的孙子， 古示 的儿子 西番雅 。
ZEPH|1|2|耶和华说： “我必从地面上彻底除灭万物。
ZEPH|1|3|我必除灭人与牲畜， 除灭空中的鸟、海里的鱼、 绊脚石和恶人； 我必把人从地面上剪除， 这是耶和华说的。
ZEPH|1|4|我必伸手攻击 犹大 和 耶路撒冷 所有的居民； 从这地方剪除剩下的 巴力 、 事奉偶像之祭司的名字与祭司；
ZEPH|1|5|还有那些在屋顶拜天上万象的， 那些敬拜耶和华指着他起誓， 却又指着 米勒公 起誓的；
ZEPH|1|6|并那些转去不跟从耶和华， 不寻求耶和华，也不求问他的。”
ZEPH|1|7|在主耶和华面前要静默无声， 因为耶和华的日子快到了。 耶和华已经预备祭物， 将召来的人分别为圣。
ZEPH|1|8|“到了献祭给耶和华的日子， 我要惩罚领袖和王子， 及所有穿外邦衣服的人。
ZEPH|1|9|到那日，我必惩罚所有跳过门槛， 以残暴和诡诈塞满主人房屋的人。
ZEPH|1|10|“当那日，从 鱼门 必发出悲哀的声音， 从第二城区发出哀号的声音， 从山间发出破裂的大响声。 这是耶和华说的。
ZEPH|1|11|玛革提施 的居民哪，你们要哀号， 因为所有的商人 都灭亡了， 满载银子的人都被剪除。
ZEPH|1|12|那时，我必用灯巡查 耶路撒冷 ， 惩罚那些沉湎在酒渣上的人； 他们心里说： ‘耶和华必不降福，也不降祸。’
ZEPH|1|13|他们的财宝成为掠物， 房屋变为废墟。 他们建造房屋，却不得住在其内； 栽葡萄园，却不得喝其中所出的酒。”
ZEPH|1|14|耶和华的大日临近， 临近而且甚快； 那是耶和华日子的风声， 勇士必在那里痛痛地哭号。
ZEPH|1|15|那日是愤怒的日子， 急难困苦的日子， 荒废凄凉的日子， 黑暗幽冥的日子， 乌云密布的日子，
ZEPH|1|16|是吹角呐喊的日子， 要攻击坚固的城， 攻击高大的城楼。
ZEPH|1|17|我必使灾祸临到人身上， 使他们行走如同盲人， 因为他们得罪了耶和华； 他们的血必倒出如灰尘， 肉身抛弃如粪土。
ZEPH|1|18|当耶和华发怒的日子， 他们的金银不能救自己； 耶和华妒忌的火必烧灭全地， 要向地上所有的居民施行可怕的毁灭。
ZEPH|2|1|不知羞耻的国民哪， 趁命令尚未发出， 日子流逝如糠秕， 耶和华的烈怒尚未临到你们， 他发怒的日子未到以先， 你们应当聚集，聚集起来。
ZEPH|2|2|
ZEPH|2|3|世上遵守耶和华典章的谦卑人哪， 你们都当寻求耶和华， 寻求公义，寻求谦卑； 或许在耶和华发怒的日子得以隐藏。
ZEPH|2|4|迦萨 必遭遗弃 ， 亚实基伦 必然荒凉； 亚实突 人必在正午被赶出， 以革伦 也要连根拔除 。
ZEPH|2|5|祸哉，住沿海之地的 基利提 人！ 迦南 、 非利士 人之地啊，耶和华的话攻击你们： 我必毁灭你，以致无人居住。
ZEPH|2|6|沿海之地要变为草场， 牧人的住处 和羊群的圈。
ZEPH|2|7|这地必为 犹大 家的余民所得； 他们要在那里放牧， 晚上躺卧在 亚实基伦 的房屋中； 因为耶和华－他们的上帝必眷顾他们， 使被掳的人归回。
ZEPH|2|8|我听见 摩押 毁谤， 亚扪 人辱骂； 他们辱骂我的百姓， 自夸自大，侵犯他们的疆土。”
ZEPH|2|9|万军之耶和华－ 以色列 的上帝说： 因此，我指着我的永生起誓： 摩押 必如 所多玛 ， 亚扪 人必像 蛾摩拉 ， 都变为刺草、盐坑、永远荒废之地。 我百姓中剩余的必掳掠他们， 我国中的幸存者必得他们的地。
ZEPH|2|10|这事临到他们是因他们的骄傲， 他们自夸自大， 辱骂万军之耶和华的百姓。
ZEPH|2|11|耶和华必向他们显为可畏， 因他使地上的众神衰微； 列国的海岛各在自己的地方敬拜他。
ZEPH|2|12|你们 古实 人， 也是被我的刀所杀的。
ZEPH|2|13|耶和华要伸手攻击北方， 毁灭 亚述 ， 使 尼尼微 荒凉， 干旱如同旷野。
ZEPH|2|14|群畜，就是各类 的走兽必卧在其中， 鹈鹕和豪猪要宿在柱顶； 窗户有鸣叫的声音， 门槛毁坏 ， 他要毁坏香柏木板 。
ZEPH|2|15|这素来欢乐、安然居住的城， 心里说：“惟有我，除我以外再没有别的”， 现在竟然荒凉，成为野兽躺卧之处！ 凡经过的人都必摇着手嗤笑它。
ZEPH|3|1|祸哉，这欺压的城！ 悖逆，污秽，
ZEPH|3|2|不听从命令， 不领受训诲， 不倚靠耶和华， 不亲近它的上帝。
ZEPH|3|3|其中的领袖是咆哮的狮子， 审判官是晚上 的野狼， 不留一点到早晨。
ZEPH|3|4|它的先知是虚浮诡诈的人， 祭司亵渎圣所，强解律法。
ZEPH|3|5|耶和华在它中间行公义， 断不做非义的事， 每早晨显明他的公义，无日不然； 只是不义的人不知羞耻。
ZEPH|3|6|“我已经除灭列国， 使他们的城楼荒废。 我使他们街道荒凉， 无人经过； 他们的城镇毁坏， 没有人，没有居民。
ZEPH|3|7|我说：‘只要你敬畏我， 领受训诲； 其住处就不会照我原先所定的被剪除 。’ 然而，他们从早起来就在各样事上败坏自己。
ZEPH|3|8|“你们要等候我， 直到我兴起掳掠 的日子； 因为我已定意招聚列邦，聚集列国， 将我的恼怒，我一切的烈怒，都倾倒在它们身上。 我妒忌的火必烧灭全地。 这是耶和华说的。
ZEPH|3|9|“那时，我要改变万民， 使他们有清洁的嘴唇， 好求告耶和华的名， 同心合意事奉我。
ZEPH|3|10|那些向我祈求的， 我所分散的子民 ， 必从 古实河 的那一边， 献供物给我。
ZEPH|3|11|“当那日，你必不再因一切得罪我的事蒙羞， 因为那时我必从你中间除掉狂喜高傲的人， 在我的圣山上你也不再狂傲。
ZEPH|3|12|我却要在你中间留下困苦贫寒的百姓， 他们必投靠耶和华的名。
ZEPH|3|13|以色列 的余民必不行恶， 不说谎，口中没有诡诈的舌头； 他们吃喝躺卧， 无人使他们惊吓。”
ZEPH|3|14|锡安 哪，应当歌唱！ 以色列 啊，应当欢呼！ 耶路撒冷 啊，应当满心欢喜快乐！
ZEPH|3|15|耶和华已经免去对你的审判， 赶出你的仇敌。 以色列 的王－耶和华在你中间； 你必不再惧怕灾祸。
ZEPH|3|16|当那日，必有话对 耶路撒冷 说： “不要惧怕！ 锡安 哪，不要手软！
ZEPH|3|17|耶和华－你的上帝在你中间 大有能力，施行拯救。 他必因你欢欣喜乐， 他在爱中静默， 且因你而喜乐欢呼。
ZEPH|3|18|我要聚集那些因无节期而愁烦的人， 他们曾远离你， 是你的重担和羞辱 。
ZEPH|3|19|那时，看哪，我必对付所有苦待你的人， 拯救瘸腿的，召集被赶出的； 那些在全地受羞辱的， 我必使他们得称赞，享名声。
ZEPH|3|20|那时，我必领你们回来，召集你们； 我使你们被掳之人归回的时候， 我必使你们在地上的万民中享名声，得称赞； 这是耶和华说的。”
HAG|1|1|大流士 王第二年六月初一，耶和华的话藉 哈该 先知向 撒拉铁 的儿子 犹大 省长 所罗巴伯 和 约撒答 的儿子 约书亚 大祭司传讲，说：
HAG|1|2|“万军之耶和华如此说，这百姓说，建造耶和华殿的时候还没有到 。”
HAG|1|3|耶和华的话藉 哈该 先知传讲，说：
HAG|1|4|“这殿荒凉，你们自己还住天花板的房屋吗？
HAG|1|5|现在，万军之耶和华如此说，你们要省察自己的行为。
HAG|1|6|你们撒的种多，收的却少；你们吃，却不得饱；喝，却不得足；穿衣服，却不得暖；领工钱的，领了工钱却装入有破洞的袋中。
HAG|1|7|“万军之耶和华如此说，你们要省察自己的行为。
HAG|1|8|你们要上山取木料，建造这殿，我就因此喜乐，且得荣耀。这是耶和华说的。
HAG|1|9|你们盼望多得，看哪，所得的却少；你们收到家中，我就吹去。这是为什么呢？因为我的殿荒凉，你们各人却只为自己的房屋奔走。这是万军之耶和华说的。
HAG|1|10|所以，因你们的缘故 ，天不降甘露，地也不出土产。
HAG|1|11|我命令干旱临到土地、山冈、五谷、新酒、新油和地上的出产，也临到人和牲畜，以及一切人手劳碌得来的。”
HAG|1|12|那时， 撒拉铁 的儿子 所罗巴伯 、 约撒答 的儿子 约书亚 大祭司，和所有幸存的百姓都听从耶和华－他们上帝的话，就是 哈该 先知奉耶和华－他们上帝差遣所说的话；百姓在耶和华面前存敬畏的心。
HAG|1|13|耶和华的使者 哈该 奉耶和华差遣对百姓说：“我与你们同在。这是耶和华说的。”
HAG|1|14|耶和华激发 撒拉铁 的儿子 犹大 省长 所罗巴伯 、 约撒答 的儿子 约书亚 大祭司，和所有幸存百姓的心，他们就来为万军之耶和华－他们上帝的殿做工。
HAG|1|15|这是在 大流士 王第二年六月二十四日。
HAG|2|1|七月二十一日，耶和华的话藉 哈该 先知传讲，说：
HAG|2|2|“你要晓谕 撒拉铁 的儿子 犹大 省长 所罗巴伯 、 约撒答 的儿子 约书亚 大祭司，和所有幸存的百姓，说：
HAG|2|3|‘你们中间存留的，有谁见过这殿从前的荣耀呢？现在你们看如何？在你们眼中岂不是如同无有吗？
HAG|2|4|所罗巴伯 啊，现在，你当刚强！这是耶和华说的。 约撒答 的儿子 约书亚 大祭司啊，你当刚强！这是耶和华说的。这地的百姓啊，你们都当刚强做工，因为我与你们同在。这是万军之耶和华说的。
HAG|2|5|这是照着你们出 埃及 时我与你们立约的话。我的灵仍要住在你们中间，你们不必惧怕。
HAG|2|6|万军之耶和华如此说：过些时候，我必再一次震动天地、沧海与干地。
HAG|2|7|我必震动万国，万国的珍宝都必运来 ，我就使这殿充满荣耀。这是万军之耶和华说的。
HAG|2|8|银子是我的，金子也是我的。这是万军之耶和华说的。
HAG|2|9|这后来的殿的荣耀必大过先前的荣耀。这是万军之耶和华说的。在这地方我必赐平安。这是万军之耶和华说的。’”
HAG|2|10|大流士 王第二年九月二十四日，耶和华的话临到 哈该 先知，说：
HAG|2|11|“万军之耶和华如此说，你要向祭司请教律法，说：
HAG|2|12|‘看哪，若有人用衣服的边兜圣肉，这衣服的边接触了饼，或汤，或酒，或油，或别的食物，这些是否成为圣呢？’”祭司回答说：“不。”
HAG|2|13|哈该 又说：“若有人因摸尸体染了不洁净，然后接触任何东西，这东西就变为不洁净吗？”祭司回答说：“必不洁净。”
HAG|2|14|于是 哈该 说：“耶和华说，在我面前这民如此，这国也是如此；他们手里的各样工作都是如此；他们在那里所献的都不洁净。”
HAG|2|15|“现在，你们心里要想一想，从今日起，耶和华的殿还没有一块石头放在石头上的情况。
HAG|2|16|那时你们怎么了？ 有人来到二十斗的谷堆那里，却只得了十斗；有人来到酒池那里要取五十桶，却只得了二十桶。
HAG|2|17|我以焚风 、霉烂、冰雹攻击你们，和你们手上的各样工作，你们仍不归向我。这是耶和华说的。
HAG|2|18|你们心里要想一想，从今日起，就是从这九月二十四日起，从立耶和华殿根基的日子起，你们心里想一想：
HAG|2|19|仓里还有谷种吗？葡萄树、无花果树、石榴树、橄榄树虽没有结果子， 从今日起，我必赐福。”
HAG|2|20|这月二十四日，耶和华的话再次临到 哈该 ，说：
HAG|2|21|“你要告诉 犹大 省长 所罗巴伯 说，我必震动天地，
HAG|2|22|倾覆列国的宝座，除灭列邦列国的势力，并倾覆战车和坐在其上的。马和骑兵都必跌倒，各人被弟兄的刀所杀。
HAG|2|23|万军之耶和华说： 撒拉铁 的儿子我仆人 所罗巴伯 啊，这是耶和华说的，到那日，我必以你为印，因我拣选了你。这是万军之耶和华说的。”
ZECH|1|1|大流士 王第二年八月，耶和华的话临到 易多 的孙子， 比利家 的儿子 撒迦利亚 先知，说：
ZECH|1|2|“耶和华曾向你们祖先大发烈怒。
ZECH|1|3|你要对 以色列 人说，万军之耶和华如此说：你们要转向我，这是万军之耶和华说的，我就转向你们，这是万军之耶和华说的。
ZECH|1|4|不要效法你们的祖先。从前的先知呼叫他们说：‘万军之耶和华如此说，当回转离开你们的恶道恶行。’他们却不听，也不顺从我。这是耶和华说的。
ZECH|1|5|你们的祖先在哪里呢？那些先知能永远存活吗？
ZECH|1|6|然而我的言语和律例，就是我所吩咐我仆人众先知的，岂不临到你们的祖先吗？他们就回转，说：万军之耶和华定意按我们的所作所为对待我们，他也已经照样行了。”
ZECH|1|7|大流士 第二年十一月，就是细罢特月二十四日，耶和华的话临到 易多 的孙子， 比利家 的儿子 撒迦利亚 先知，说：
ZECH|1|8|“我夜间观看，看哪，有一人骑着红马，站在洼地的番石榴树中间。在他身后有红色、褐色和白色的马。”
ZECH|1|9|我说：“主啊，这是什么意思？”与我说话的天使说：“我要指示你这是什么意思。”
ZECH|1|10|那站在番石榴树中间的人回答说：“这是奉耶和华差遣，在遍地巡逻的。”
ZECH|1|11|他们对站在番石榴树中间耶和华的使者说：“我们在遍地巡逻，看哪，全地都安息平静。”
ZECH|1|12|于是，耶和华的使者说：“万军之耶和华啊，你恼恨 耶路撒冷 和 犹大 的城镇已经七十年了，你不施怜悯要到几时呢？”
ZECH|1|13|耶和华就用美善的话和安慰的话回答那与我说话的天使。
ZECH|1|14|与我说话的天使对我说：“你要宣告，万军之耶和华如此说：我为 耶路撒冷 而妒忌，为 锡安 大大妒忌。
ZECH|1|15|我非常恼怒那享安逸的列国，因我从前稍微恼怒，他们就越发加害。
ZECH|1|16|所以耶和华如此说：现在我回到 耶路撒冷 ，仍要施怜悯，我的殿要重建在其中，准绳必拉在 耶路撒冷 之上。这是万军之耶和华说的。
ZECH|1|17|你要再宣告，万军之耶和华如此说：我的城镇要再度繁荣发达。耶和华必再安慰 锡安 ，拣选 耶路撒冷 。”
ZECH|1|18|我举目观看，看哪，有四只角。
ZECH|1|19|我问那与我说话的天使：“这是什么意思？”他对我说：“这是击散 犹大 、 以色列 和 耶路撒冷 的角。”
ZECH|1|20|耶和华又把四个匠人指给我看。
ZECH|1|21|我问：“这些人来做什么呢？”他说：“那是击散 犹大 的角，使人不敢抬头；但这些匠人前来威吓列国，打掉列国的角，因为他们举起角来击散 犹大 地。”
ZECH|2|1|我举目观看，看哪，有一人手拿丈量的绳。
ZECH|2|2|我问：“你到哪里去？”他对我说：“要去丈量 耶路撒冷 ，看有多宽多长。”
ZECH|2|3|看哪，与我说话的天使出去 ，另有一位天使迎着他来，
ZECH|2|4|对他说：“你跑去告诉这个年轻人说， 耶路撒冷 必有人居住，如同无城墙的乡村，因为其中的人和牲畜很多。
ZECH|2|5|耶和华说：‘我要作 耶路撒冷 四围火的城墙，并要作城中的荣耀。’”
ZECH|2|6|耶和华说：“来，来！你们要从北方之地逃回；因我曾把你们分散到天的四方 。这是耶和华说的。”
ZECH|2|7|来！住 巴比伦 的 锡安 百姓啊，逃吧！
ZECH|2|8|万军之耶和华在显出荣耀之后，差遣我到掳掠你们的列国那里，他如此说：“碰你们的就是碰他自己 眼中的瞳人。
ZECH|2|9|看哪，我要挥手攻击他们，他们就必作自己奴仆的掳物。”你们就知道万军之耶和华差遣了我。
ZECH|2|10|耶和华说：“ 锡安 哪，应当欢乐歌唱，因为，看哪，我要来，要住在你中间。
ZECH|2|11|在那日，必有许多国家归附耶和华，作我的子民。我要住 在你中间。”你就知道万军之耶和华差遣我到你那里去。
ZECH|2|12|耶和华必收回 犹大 ，作为他圣地的产业，他必再度拣选 耶路撒冷 。
ZECH|2|13|凡血肉之躯都当在耶和华面前静默无声，因为他从他的圣所奋起了。
ZECH|3|1|天使 指给我看： 约书亚 大祭司站在耶和华的使者面前，撒但站在 约书亚 的右边控告他。
ZECH|3|2|耶和华向撒但说：“撒但哪，耶和华责备你！拣选 耶路撒冷 的耶和华责备你！这不是从火中抽出来的一根柴吗？”
ZECH|3|3|约书亚 穿着污秽的衣服，站在那使者面前。
ZECH|3|4|使者吩咐那些侍立在他面前的说：“脱去他污秽的衣服。”又对 约书亚 说：“你看，我使你的罪孽离开你，要给你穿上华美的衣服。”
ZECH|3|5|我说 ：“要将洁净的冠冕戴在他头上。”他们就把洁净的冠冕戴在他头上，给他穿上华美的衣服，耶和华的使者在旁边站立。
ZECH|3|6|耶和华的使者告诫 约书亚 说，
ZECH|3|7|万军之耶和华如此说：“你若遵行我的道，谨守我的命令，就可以管理我的家，看守我的院宇；我也要使你在这些侍立的人中间来往。
ZECH|3|8|约书亚 大祭司啊，你和坐在你面前的同伴都当听，因为他们是作预兆的：看哪，我必使我仆人 大卫 的苗裔 长出。
ZECH|3|9|看哪，这是我在 约书亚 面前所立的石头，这一块石头上有七眼。看哪，我要亲自雕刻这石头，并在一日之间除掉这地的罪孽。这是万军之耶和华说的。
ZECH|3|10|在那日，你们各人要请邻舍坐在葡萄树和无花果树下。这是万军之耶和华说的。”
ZECH|4|1|那与我说话的天使又来叫醒我，好像人睡觉时被唤醒一样。
ZECH|4|2|他问我：“你看见什么？”我说：“我看见了，看哪，有一个纯金的灯台，顶上有灯座，其上有七盏灯，每盏灯的上头有七根管子；
ZECH|4|3|旁边有两棵橄榄树，一棵在灯座的右边，一棵在灯座的左边。”
ZECH|4|4|我问与我说话的天使说：“主啊，这是什么意思？”
ZECH|4|5|与我说话的天使回答，对我说：“你不知道这是什么意思吗？”我说：“主啊，我不知道。”
ZECH|4|6|他回答我说：“这是耶和华指示 所罗巴伯 的话。万军之耶和华说：不是倚靠势力，不是倚靠才能，乃是倚靠我的灵方能成事 。
ZECH|4|7|大山哪，你算什么呢？在 所罗巴伯 面前，你必夷为平地。他安放顶上的那块石头，人就欢呼：‘愿恩惠、恩惠归与这殿！’”
ZECH|4|8|耶和华的话临到我，说：
ZECH|4|9|“ 所罗巴伯 的手立了这殿的根基，他的手也必完成这工，你就知道万军之耶和华差遣我到你们这里。
ZECH|4|10|谁藐视这日的事为小呢？他们见 所罗巴伯 手拿石垂线就欢喜。这七盏灯 是耶和华的眼睛，遍察全地。”
ZECH|4|11|我问天使说：“那么在灯台左右的这两棵橄榄树是什么意思呢？”
ZECH|4|12|我再次问他：“这两根橄榄树枝在两根流出金色油的金嘴旁边，是什么意思呢？”
ZECH|4|13|他对我说：“你不知道这是什么意思吗？”我说：“主啊，我不知道。”
ZECH|4|14|他说：“这是两位受膏者，侍立在全地之主的旁边。”
ZECH|5|1|我又举目观看，看哪，有一飞行的书卷。
ZECH|5|2|他问我：“你看见什么？”我回答：“我看见一飞行的书卷，长二十肘，宽十肘。”
ZECH|5|3|他对我说：“这就是向全地面发出的诅咒。凡偷窃的必按书卷这面的话除灭，凡起假誓的必按书卷那面的话除灭。
ZECH|5|4|万军之耶和华说：我要把这书卷送出去，进入偷窃者的家和指着我名起假誓者的家，停留在他家里，连房屋带木头和石头都毁灭了。”
ZECH|5|5|与我说话的天使前来，对我说：“你要举目观看，看那出现的是什么。”
ZECH|5|6|我问：“这是什么呢？”他说：“这出现的是量器 。”又说：“是他们的眼目，遍行全地 。”
ZECH|5|7|看哪，圆形的铅盖被抬起来，有一个妇人坐在量器中。
ZECH|5|8|天使说：“这是罪恶。”他就把妇人推进量器里，把铅盖压在量器的口上。
ZECH|5|9|于是我举目观看，看哪，有两个妇人前来，她们的翅膀中有风，翅膀如同鹳鸟的翅膀。她们把量器抬起来，悬在天地之间。
ZECH|5|10|我问那与我说话的天使：“她们要把量器抬到哪里去呢？”
ZECH|5|11|他对我说：“要抬到 示拿 地去，为它建造房屋；等预备妥当，就把它安放在自己的台座上。”
ZECH|6|1|我又举目观看，看哪，有四辆马车从两座山的中间出来；那两座山是铜山。
ZECH|6|2|第一辆车套着红马，第二辆车套着黑马，
ZECH|6|3|第三辆车套着白马，第四辆车套着带斑点的马，都是强壮的 。
ZECH|6|4|我就回应与我说话的天使说：“主啊，这是什么意思？”
ZECH|6|5|天使回答，对我说：“这是天的四风，是从全地之主面前出来的。”
ZECH|6|6|套着黑马的车往北方之地去，白马跟随在后；有斑点的马往南方之地去；
ZECH|6|7|那些壮马出来，急着要在地上巡逻。天使说：“你们只管在地上巡逻。”它们就在地上巡逻。
ZECH|6|8|他又呼叫我，告诉我说：“你看，往北方地去的已在北方之地使我放心。”
ZECH|6|9|耶和华的话临到我，说：
ZECH|6|10|“你要拿从 巴比伦 归来的被掳之人 黑玳 、 多比雅 、 耶大雅 所献的，当日就要进到 西番雅 的儿子 约西亚 的家里，
ZECH|6|11|拿这金银做冠冕，戴在 约撒答 的儿子 约书亚 大祭司的头上；
ZECH|6|12|对他说，万军之耶和华如此说：‘看哪，那名称为 大卫 苗裔的，要在本处生长，并要建造耶和华的殿。
ZECH|6|13|就是他，要建造耶和华的殿，他要承受尊荣，坐在位上掌王权；又有一位祭司坐在自己的位上，两职之间筹划和平。
ZECH|6|14|这冠冕要归 希连 、 多比雅 、 耶大雅 ，和 西番雅 的儿子 贤 ，放在耶和华的殿里作为纪念。’”
ZECH|6|15|远方的人要来建造耶和华的殿，你们因此就知道，万军之耶和华差遣我到你们这里来。你们若留意听从耶和华－你们上帝的话，这事必然成就。
ZECH|7|1|大流士 王第四年九月，就是基斯流月初四，耶和华的话临到 撒迦利亚 。
ZECH|7|2|那时 伯特利 人已经差遣 沙利色 和 利坚．米勒 ，并他们的人，去恳求耶和华的恩，
ZECH|7|3|问万军之耶和华殿中的祭司，又问先知：“我当如历年以来所行，在五月哭泣斋戒吗？”
ZECH|7|4|万军之耶和华的话临到我，说：
ZECH|7|5|“你要向这地全体百姓和祭司说：‘你们这七十年来，在五月、七月禁食悲哀，岂是真的向我禁食吗？
ZECH|7|6|你们吃喝，不是为自己吃，为自己喝吗？
ZECH|7|7|当 耶路撒冷 和四围的城镇有人居住，享繁荣， 尼革夫 和 谢非拉 也有人居住的时候，耶和华藉从前的先知所宣告的，你们不当听吗？’”
ZECH|7|8|耶和华的话临到 撒迦利亚 ，说：
ZECH|7|9|“万军之耶和华如此说：你们要按真正的公平来审判，彼此以慈爱怜悯相待。
ZECH|7|10|不可欺压寡妇、孤儿、寄居的和困苦的人。谁都不可心里谋害弟兄。
ZECH|7|11|他们却不留意；耸肩悖逆，耳朵发沉，不肯听从。
ZECH|7|12|他们的心坚硬如金刚石，不听律法和万军之耶和华藉着他的灵差遣从前先知所说的话。因此，万军之耶和华大发烈怒。
ZECH|7|13|万军之耶和华说：我曾呼唤他们，他们不听；将来他们呼求我，我也不听！
ZECH|7|14|我必以旋风将他们吹散到素不认识的万国中。他们离开以后，地就荒凉，无人来往经过；他们使美好之地荒凉了。”
ZECH|8|1|万军之耶和华的话临到我，说：
ZECH|8|2|“万军之耶和华如此说：我为 锡安 而妒忌，大大妒忌；我为了它妒忌而大发烈怒。
ZECH|8|3|耶和华如此说：我要回到 锡安 ，住在 耶路撒冷 中间。 耶路撒冷 必称为忠实的城，万军之耶和华的山必称为圣山。
ZECH|8|4|万军之耶和华如此说：将来必有年老的男女坐在 耶路撒冷 的广场上，各人因年纪老迈而手拿枴杖。
ZECH|8|5|城里的广场满有男孩女孩在玩耍。
ZECH|8|6|万军之耶和华如此说：在那些日子，即使这事在这余民眼中看为奇妙，难道在我眼中也看为奇妙吗？这是万军之耶和华说的。
ZECH|8|7|万军之耶和华如此说：看哪，我要从日出之地、从日落之地拯救我的子民。
ZECH|8|8|我要领他们来，使他们住在 耶路撒冷 中间。他们要作我的子民，我要作他们的上帝，都凭信实和公义。
ZECH|8|9|“万军之耶和华如此说：你们的手要坚强；这些日子，你们已听见先知的口，在万军之耶和华殿的根基立定、圣殿建造的日子所说的这些话。
ZECH|8|10|那些日子以前，人得不着工价，牲畜也无人雇用；且因敌人的缘故，出入不得平安；因我使人与人互相攻击。
ZECH|8|11|但如今，我对这余民必不像先前的日子。这是万军之耶和华说的。
ZECH|8|12|因为他们要平安撒种，葡萄树要结果子，土地必有出产，天也必降甘露。我要使这余民享受这一切。
ZECH|8|13|犹大 家和 以色列 家啊，你们从前在列国中怎样成为可诅咒的；照样，我要拯救你们，使你们得福 。不要惧怕，你们的手要坚强。
ZECH|8|14|“万军之耶和华如此说：你们祖先惹我发怒的时候，我怎样定意降祸，并不改变；万军之耶和华说，
ZECH|8|15|这些日子我也定意施恩给 耶路撒冷 和 犹大 家；你们不要惧怕。
ZECH|8|16|你们所当行的是这样：每个人要与邻舍说诚实话，在城门口要按真正的公平来审判，使人和睦。
ZECH|8|17|谁都不可心里谋害邻舍，也不可喜爱起假誓，因为这些事都为我所恨恶。这是耶和华说的。”
ZECH|8|18|万军之耶和华的话临到我，说：
ZECH|8|19|“万军之耶和华如此说：四月的禁食、五月的禁食、七月的禁食和十月的禁食，必成为 犹大 家的欢喜和快乐，以及美好的节期；所以你们要喜爱诚实与和平。
ZECH|8|20|“万军之耶和华如此说：将来还有众百姓和许多城镇的居民要来。
ZECH|8|21|这城的居民必到那城，说：‘我们快去恳求耶和华的恩，寻求万军之耶和华；我自己也要去。’
ZECH|8|22|必有许多民族和强盛的国家来到 耶路撒冷 寻求万军之耶和华，恳求耶和华的恩。
ZECH|8|23|万军之耶和华如此说：在那些日子，列国中说各种语言的人，必有十个人强拉住一个 犹大 人衣服的边，说：‘我们要与你们同去，因为我们听见上帝与你们同在了。’”
ZECH|9|1|耶和华的默示， 他的话临到 哈得拉 地、 大马士革 －因世人和 以色列 各支派的眼目都向着耶和华－
ZECH|9|2|和邻近的 哈马 ， 以及 推罗 和 西顿 。 因为它极有智慧，
ZECH|9|3|推罗 为自己建造坚固城 ， 堆起银子如尘沙， 纯金如街上的泥土。
ZECH|9|4|看哪，主必赶出它， 重创它海上的势力， 它必被火吞灭。
ZECH|9|5|亚实基伦 看见必惧怕， 迦萨 看见甚痛苦， 以革伦 因失了盼望而蒙羞； 迦萨 必不再有君王， 亚实基伦 也不再有人居住，
ZECH|9|6|混血的人要住在 亚实突 ； 我必除灭 非利士 人的骄傲。
ZECH|9|7|我要除去他口中带血之肉 和牙齿内可憎之物。 他必作余民归于我们的上帝， 在 犹大 像族长一样； 以革伦 必如 耶布斯 人。
ZECH|9|8|我要扎营在我的家， 敌军不得任意往来， 暴虐的人也不再经过， 因为我亲眼看顾。
ZECH|9|9|锡安 哪，应当大大喜乐； 耶路撒冷 啊，应当欢呼。 看哪，你的王来到你这里！ 他是公义的，并且施行拯救， 谦和地骑着驴， 骑着小驴，驴的驹子。
ZECH|9|10|我必除灭 以法莲 的战车 和 耶路撒冷 的战马； 战争的弓也必剪除。 他要向列国讲和平； 他的权柄必从这海管到那海， 从 大河 管到地极。
ZECH|9|11|锡安 哪，我因与你立约的血， 要从无水坑里释放你中间被囚的人。
ZECH|9|12|被囚而有指望的人哪，要转回堡垒； 我今日宣告，我必加倍补偿你。
ZECH|9|13|我为自己把 犹大 弯紧， 我使 以法莲 如满弓。 锡安 哪，我要唤起你的儿女， 希腊 啊，我要攻击你的儿女， 使你如勇士的刀。
ZECH|9|14|耶和华要显现在他们身上， 他的箭要射出如闪电。 主耶和华必吹角， 乘南方的旋风而行。
ZECH|9|15|万军之耶和华必保护他们； 他们要吞灭，要践踏弹弓的石头 ； 他们呐喊，狂饮 如喝酒， 如盛满的碗， 又如坛的四角。
ZECH|9|16|当那日，耶和华－他们的上帝 必看他的百姓如羊群，拯救他们； 因为他们如冠冕上的宝石， 在他的地上如旗帜高举 。
ZECH|9|17|他是何等善！ 他是何其美！ 五谷使少男强壮， 新酒使少女健美。
ZECH|10|1|春雨的季节，你们要向耶和华求雨。 耶和华发出雷电， 为众人降下大雨， 把田园的菜蔬赐给人。
ZECH|10|2|因为家中神像所言的是虚空， 占卜者所见的是虚假， 他们讲说假梦， 徒然安慰人。 所以众人如羊流离， 因无牧人就受欺压。
ZECH|10|3|我的怒气向牧人发作， 我必惩罚那为首的 ； 万军之耶和华眷顾他的羊群， 就是 犹大 家， 必使他们如战场上的骏马。
ZECH|10|4|房角石从他而出， 橛子从他而出， 战争的弓也从他而出， 每一个掌权的都从他而出。
ZECH|10|5|他们必如战场上的勇士， 践踏仇敌如街上的泥土。 他们必争战，因为耶和华与他们同在， 他们必使骑马的羞愧。
ZECH|10|6|我要坚固 犹大 家， 拯救 约瑟 家， 我要领他们归回，因我怜悯他们， 他们必像我未曾弃绝他们一样； 都因我是耶和华－他们的上帝， 我必应允他们。
ZECH|10|7|以法莲 人必如勇士， 他们心中畅快如同喝酒； 他们的儿女看见就欢喜， 他们的心必因耶和华喜乐。
ZECH|10|8|我要呼叫，聚集他们， 因我已经救赎他们。 他们的人数必增添， 如从前增添一样。
ZECH|10|9|我要将他们分散在列国中， 他们必在远方记得我； 他们与儿女都必存活， 他们要归回。
ZECH|10|10|我必使他们从 埃及 地归回， 从 亚述 召集他们， 领他们到 基列 地和 黎巴嫩 ； 这些还不够他们居住。
ZECH|10|11|耶和华 必经过苦海，击打海浪。 尼罗河 的深处全都枯干， 亚述 的骄傲必降卑， 埃及 的权杖必除去。
ZECH|10|12|我要使他们倚靠耶和华，得以坚固， 他们必奉他的名而行 ； 这是耶和华说的。
ZECH|11|1|黎巴嫩 哪，敞开你的门， 任火吞灭你的香柏树。
ZECH|11|2|哀号吧，松树！ 因为香柏树倾倒了，高大的树毁坏了。 哀号吧， 巴珊 的橡树！ 因为茂盛的树林倒下来了。
ZECH|11|3|听啊，有牧人在哀号， 因他们的荣华败落了； 听啊，有少壮狮子咆哮， 因 约旦河 旁的丛林荒废了。
ZECH|11|4|耶和华－我的上帝如此说：“你要牧养这群将宰的羊。
ZECH|11|5|买羊的宰了他们，却不认为自己有罪；卖他们的也说：‘耶和华是应当称颂的，因我富足了。’牧养他们的并不怜悯他们。
ZECH|11|6|我不再怜悯这地的居民。看哪，我要将这些人交在各人的邻舍和君王手中；他们必毁灭这地，我却不救任何一个脱离他们的手。这是耶和华说的。”
ZECH|11|7|于是，我牧养这群将宰的羊，就是羊群中最困苦的 ；我拿着两根杖，一根我称为“恩惠” ，一根称为“联合”。这样，我就牧养这群羊。
ZECH|11|8|一个月之内，我废除了三个牧人，因为我的心厌烦他们，他们的心也憎恶我。
ZECH|11|9|我就说：“我不牧养你们。要死的，由他死；灭亡的，由他灭亡；剩余的，由他们彼此吞食。”
ZECH|11|10|我拿起那根称为“恩惠”的杖，折断它，表明我废弃与万民所立的约。
ZECH|11|11|当日约就废了。因此，那些羊群中最困苦的 ，看着我，就知道这真是耶和华的话。
ZECH|11|12|我对他们说：“你们若看为美，就给我工价。不然，就罢了！”于是他们秤了三十块银钱作为我的工价。
ZECH|11|13|耶和华对我说：“把它丢给窑户。那是他们对我所估定的好价钱！”我就取这三十块银钱，在耶和华的殿中将它丢给窑户。
ZECH|11|14|我又折断第二根杖，就是称为“联合”的那根杖，表明我废弃 犹大 与 以色列 弟兄间的情谊。
ZECH|11|15|耶和华对我说：“你再把愚昧牧人所用的器具拿来，
ZECH|11|16|因为，看哪，我要在这地立一个牧人；他不看顾将亡的，不寻找分散的，不医治受伤的，也不牧养强壮的；却要吞吃肥羊的肉，撕裂它们的蹄。
ZECH|11|17|祸哉！无用的牧人丢弃羊群， 刀必临到他的膀臂和右眼上； 他的膀臂必全然枯干， 他的右眼也必昏暗失明。”
ZECH|12|1|耶和华的默示，他的话论到 以色列 。 铺张诸天、建立地基、造人里面之灵的耶和华说：
ZECH|12|2|“看哪，我要使 耶路撒冷 成为令四围列国百姓昏醉的杯； 耶路撒冷 被围困， 犹大 也一样受困 。
ZECH|12|3|在那日，我要使 耶路撒冷 成为万民的一块沉重石头，凡举起它的必受重伤；地上的万国都聚集攻击它。
ZECH|12|4|到那日，我必令一切的马匹惊惶，使骑马的癫狂。我必张开眼睛看顾 犹大 家，却使列国一切的马匹瞎眼。这是耶和华说的。
ZECH|12|5|犹大 的族长心里要说：‘ 耶路撒冷 的居民因倚靠万军之耶和华－他们的上帝，就成为我的力量 。’
ZECH|12|6|“那日，我必使 犹大 的族长如柴堆中的火盆，又如禾捆里的火把；他们必左右吞灭四围列国的百姓。 耶路撒冷 却仍屹立在本处，仍在 耶路撒冷 ！
ZECH|12|7|“耶和华要先拯救 犹大 的帐棚，免得 大卫 家的荣耀和 耶路撒冷 居民的荣耀胜过 犹大 。
ZECH|12|8|那日，耶和华必保护 耶路撒冷 的居民。他们中间软弱的在那日必如 大卫 ； 大卫 家必如上帝，如行在他们前面的耶和华的使者。
ZECH|12|9|那日，我必定意灭绝前来攻击 耶路撒冷 的万国。”
ZECH|12|10|“我要将那施恩与恳求的灵，浇灌 大卫 家和 耶路撒冷 的居民。他们必仰望我，就是他们所扎的那位。他们必为他悲伤，如丧独子，又为他哀哭，如丧长子。
ZECH|12|11|那日，在 耶路撒冷 必有大大的哀号，如 米吉多 平原上 哈达．临门 的哀号。
ZECH|12|12|这地必哀哭：一家一家地哭， 大卫 家的家族聚在一处，他们的妇女聚在一处； 拿单 家的家族聚在一处，他们的妇女聚在一处。
ZECH|12|13|利未 家的家族聚在一处，他们的妇女聚在一处； 示每 家的家族聚在一处，他们的妇女聚在一处。
ZECH|12|14|其余的各家，每一家的家族聚在一处，他们的妇女聚在一处。”
ZECH|13|1|“在那日，因罪恶与污秽的缘故，必有一泉源为 大卫 家和 耶路撒冷 的居民而开。”
ZECH|13|2|万军之耶和华说：“在那日，我要从地上除灭偶像的名，使它不再被记得；我也必使这地不再有先知，不再有污秽的灵。
ZECH|13|3|若还有人说预言，生他的父母必对他说：‘你不得存活，因为你假借耶和华的名说谎话。’生他的父母在他说预言时，要将他刺死。
ZECH|13|4|那日，凡作先知说预言的必因所论的异象羞愧，不再穿毛皮外袍哄骗人。
ZECH|13|5|他要说：‘我不是先知，我是耕地的；我从幼年就作人的奴仆。’
ZECH|13|6|有人对他说：‘你两手臂间是什么伤呢？’他说：‘这是我在亲友家中所受的伤。’”
ZECH|13|7|万军之耶和华说： 刀剑哪，兴起攻击我的牧人， 攻击我的同伴吧！ 要击打牧人，羊就分散了； 我必反手攻击那微小的。
ZECH|13|8|这全地的人， 三分之二将被剪除而死， 三分之一仍必存留。 这是耶和华说的。
ZECH|13|9|我要使这三分之一经过火， 熬炼他们，如熬炼银子； 试炼他们，如试炼金子。 他们要求告我的名， 我必应允他们。 我说：“这是我的子民。” 他们要说：“耶和华是我的上帝。”
ZECH|14|1|看哪，耶和华的日子临近了，你的财物必被抢掠，在你中间被瓜分。
ZECH|14|2|我要招聚万国与 耶路撒冷 争战；城必被攻取，房屋被抢夺，妇女被玷污，城中的一半被掳去；但其余的百姓不会从城中被剪除。
ZECH|14|3|那时，耶和华要出去与那些国家打仗，如同从前战争的日子打仗一样。
ZECH|14|4|那日，他的脚必站在 橄榄山 上，这山面向 耶路撒冷 的东边。 橄榄山 必从中间裂开，自东至西成为极大的谷；山的一半向北挪移，一半向南挪移。
ZECH|14|5|你们要从我的山谷中逃跑，因为山谷必延到 亚萨 。你们要逃跑，如在 犹大 王 乌西雅 年间逃避大地震一样 。耶和华－我的上帝必降临，所有的圣者与你 同来。
ZECH|14|6|在那日，必没有光，不会放晴，只有乌云 。
ZECH|14|7|耶和华所知道的那一日，没有白天，没有黑夜，到了晚上仍有亮光。
ZECH|14|8|在那日，必有活水从 耶路撒冷 出来，一半往东海流，一半往西海流；冬夏都是如此。
ZECH|14|9|耶和华要作全地的王。那日，耶和华必为独一无二，他的名也是独一无二。
ZECH|14|10|从 迦巴 直到 耶路撒冷 南方的 临门 ，全地要变为旷野。 耶路撒冷 要矗立于本处，从 便雅悯门 到 旧门 ，又到 角门 ，并从 哈楠业楼 ，直到王的酒池。
ZECH|14|11|人要住在其中，不再有诅咒； 耶路撒冷 必安然屹立。
ZECH|14|12|这是耶和华所降的灾殃，要攻击那些与 耶路撒冷 作战的万民；他们两脚站立时，肉要溃烂，眼在眶中溃烂，舌在口中也溃烂。
ZECH|14|13|那日，耶和华必使他们大大混乱。他们彼此用手揪住，用手互相攻击。
ZECH|14|14|犹大 也要在 耶路撒冷 打仗 。那时四围各国的财物，就是许许多多的金银和衣服，必被收聚。
ZECH|14|15|马匹、骡子、骆驼、驴和营中一切的牲畜所遭的灾殃与那灾殃一样。
ZECH|14|16|上来攻击 耶路撒冷 的列国中所有剩下的人，要年年上来敬拜大君王－万军之耶和华，并守住棚节。
ZECH|14|17|地上万族中，凡不上 耶路撒冷 敬拜大君王－万军之耶和华的，雨必不降在他们的地上。
ZECH|14|18|埃及 族若不上来，雨必不降在他们的地上；凡不上来守住棚节的列国，耶和华必用这灾攻击他们。
ZECH|14|19|这就是 埃及 的惩罚和那些不上来守住棚节之列国的惩罚。
ZECH|14|20|在那日，马的铃铛上要刻上“归耶和华为圣”。耶和华殿内的锅必如祭坛前的碗一样。
ZECH|14|21|耶路撒冷 和 犹大 一切的锅都必归万军之耶和华为圣。凡献祭的都必来取这锅，在其中煮肉。当那日，在万军之耶和华的殿中必不再有做买卖的人 。
MAL|1|1|耶和华的话，藉 玛拉基 传给 以色列 的默示。
MAL|1|2|耶和华说：“我曾爱你们。”你们却说：“你在何事上爱我们呢？”耶和华说：“ 以扫 不是 雅各 的哥哥吗？我却爱 雅各 ，
MAL|1|3|恶 以扫 ，使他的山岭荒凉，把他的地业交给旷野的野狗。”
MAL|1|4|以东 若说：“我们虽被毁坏，却要重建荒废之处。”万军之耶和华如此说：“任他们建造，我必拆毁；人必称他们为‘邪恶之境’，为‘耶和华永远恼怒之民’。”
MAL|1|5|你们必亲眼看见，你们要说：“耶和华在 以色列 疆界之外必尊为大！”
MAL|1|6|万军之耶和华对你们说：“儿子孝敬父亲，仆人敬畏主人；我既为父亲，孝敬我的在哪里呢？我既为主人，敬畏我的在哪里呢？你们这些藐视我名的祭司啊！”你们却说：“我们在何事上藐视你的名呢？”
MAL|1|7|“你们将不洁净的食物献在我的祭坛上，却说：‘我们在何事上使你不洁净呢？’你们说，耶和华的供桌是可藐视的。
MAL|1|8|你们将瞎眼的献为祭物，这不算为恶吗？将瘸腿的、有病的献上，这不算为恶吗？那么，请把这些献给你的省长，他岂会悦纳你 ，岂会抬举你呢？这是万军之耶和华说的。”
MAL|1|9|现在我劝你们要恳求上帝，好让他施恩给我们。这事既出于你们的手，他岂会抬举你们任何人呢？这是万军之耶和华说的。
MAL|1|10|万军之耶和华说：“甚愿你们中间有人把殿的门 关上，免得你们徒然在我坛上烧火。我不喜欢你们，也不从你们手中悦纳供物。”
MAL|1|11|万军之耶和华说：“从日出之地到日落之处，我的名在列国中必尊为大。在各处，人必奉我的名烧香，献洁净的供物，因为我的名在列国中必尊为大。
MAL|1|12|你们却亵渎我的名，说：‘主的供桌是不洁净的，供桌上的果子和食物是可藐视的。’
MAL|1|13|你们又说：‘看哪，这些事何等烦琐！’并嗤之以鼻 。这是万军之耶和华说的。你们把抢来的、瘸腿的、有病的拿来献上为祭，我岂能从你们手中悦纳它呢？这是耶和华说的。
MAL|1|14|行诡诈的人是可诅咒的！他的群畜中虽有公羊，他许了愿，却将有残疾的献给主。因我是大君王，我的名在列国中是可畏的。这是万军之耶和华说的。”
MAL|2|1|现在，众祭司啊，这诫命是给你们的。
MAL|2|2|万军之耶和华说：“你们若不听，不放在心上，不将荣耀归给我的名，我就使诅咒临到你们，使你们的福分变为诅咒；其实我已经诅咒了你们的福分，因你们不把诫命放在心上。
MAL|2|3|看哪，我要斥责你们的后裔，把粪抹在你们脸上，就是你们祭牲 的粪。人要把你们和粪一起抬出去，
MAL|2|4|你们就知道我颁这诫命给你们，使我与 利未 所立的约可以常存。这是万军之耶和华说的。
MAL|2|5|我曾与他立生命和平安的约。我将这两样赐给他，使他存敬畏的心；他就敬畏我，惧怕我的名。
MAL|2|6|真实的训诲在他口中，他的嘴唇中没有不义。他以平安和正直与我同行，使许多人回转离开罪孽。
MAL|2|7|祭司的嘴唇当守护知识，人也当从他口中寻求训诲，因为他是万军之耶和华的使者。
MAL|2|8|你们却偏离正道，使许多人在这训诲上绊跌。你们破坏了我与 利未 人所立的约。这是万军之耶和华说的。
MAL|2|9|所以我使你们被众百姓藐视，看为卑贱；因你们不遵守我的道，在律法上看人的情面 。”
MAL|2|10|我们岂不都有一位父吗？岂不是一位上帝创造了我们吗？为何互相行诡诈，亵渎了上帝与我们列祖所立的约呢？
MAL|2|11|犹大 行事诡诈，在 以色列 和 耶路撒冷 中行了可憎的事；因为 犹大 人亵渎耶和华所喜爱的圣殿，娶外邦神明的女子为妻。
MAL|2|12|凡做这事的，无论是清醒的 或回应的，即使献供物给万军之耶和华，耶和华也要将他从 雅各 的帐棚中剪除。
MAL|2|13|你们又再做这样的事，使哭泣和叹息的眼泪遮盖耶和华的祭坛，以致耶和华不再理会那供物，也不喜欢从你们的手中收纳。
MAL|2|14|你们还说：“这是为什么呢？”因为耶和华在你和你年轻时所娶的妻之间作证。她虽是你的配偶，你誓约 的妻，你却背弃她。
MAL|2|15|一个人如果还剩下一点灵性，他不会这么做。这人在寻找什么呢？上帝的后裔！ 当谨守你们的灵性，谁也不可背弃年轻时所娶的妻。
MAL|2|16|耶和华－ 以色列 的上帝说：“我恨恶休妻的事和衣服外面披上暴力的人。所以当谨守你们的心，不可行诡诈。这是万军之耶和华说的。”
MAL|2|17|你们用言语使耶和华厌烦，却说：“我们在何事上使他厌烦呢？”因为你们说：“凡行恶的，耶和华看为善，并且喜爱他们；”又说：“公平的上帝在哪里呢？”
MAL|3|1|万军之耶和华说：“看哪，我要差遣我的使者在我前面预备道路。你们所寻求的主必忽然来到他的殿；立约的使者，就是你们所仰慕的，看哪，快要来到。”
MAL|3|2|他来的日子，谁能当得起呢？他显现的时候，谁能立得住呢？因为他如炼金匠的火，如漂洗者的碱。
MAL|3|3|他必坐下如炼净银子的人，必洁净 利未 人，熬炼他们像金银一样；他们就凭公义献供物给耶和华。
MAL|3|4|那时， 犹大 和 耶路撒冷 所献的供物必蒙耶和华悦纳，仿佛古时之日、上古之年。
MAL|3|5|万军之耶和华说：“我必临近你们，施行审判。我必速速作见证，警戒那些行邪术的、犯奸淫的、起假誓的、剥削雇工工钱的、欺压孤儿寡妇的、屈枉寄居者的和不敬畏我的人。”
MAL|3|6|“我－耶和华是不改变的；所以， 雅各 的子孙啊，你们不致灭亡。
MAL|3|7|从你们祖先的日子以来，你们就偏离我的律例而不遵守。现在你们要转向我，我就转向你们。这是万军之耶和华说的。你们却说：‘我们如何转向呢？’
MAL|3|8|人岂可抢夺上帝呢？你们竟抢夺我！你们却说：‘我们在何事上抢夺你呢？’其实就是在你们当纳的十分之一奉献和当献的供物上。
MAL|3|9|因你们全国上下都抢夺我的供物，诅咒就临到你们身上。
MAL|3|10|你们要将当纳的十分之一全然送入仓库，使我家有粮，以此试试我，是否为你们敞开天上的窗户，倾福与你们，甚至无处可容。这是万军之耶和华说的。
MAL|3|11|我必为你们斥责蝗虫 ，不容它毁坏你们的土产。你们田间的葡萄树，果实未熟以先也不会掉落。这是万军之耶和华说的。
MAL|3|12|万国必称你们为有福的，因你们必成为喜乐之地。这是万军之耶和华说的。”
MAL|3|13|耶和华说：“你们用话顶撞我。”你们却说：“我们说了什么话顶撞你呢？”
MAL|3|14|你们说：“事奉上帝是枉然，我们遵守上帝所吩咐的，在万军之耶和华面前哀痛而行，有什么益处呢？
MAL|3|15|现在，我们称狂傲的人为有福，并且行恶的人得以建立；他们虽然试探上帝，却得以逃脱。”
MAL|3|16|那时，敬畏耶和华的人彼此谈论，耶和华侧耳而听，且有纪念册在他面前，记录那敬畏耶和华、思念他名的人。
MAL|3|17|万军之耶和华说：“在我所定的日子，他们必属我，是我宝贵的产业。我必怜悯他们，如同人怜悯那服侍他的儿子。
MAL|3|18|那时你们必再一次 看出义人和恶人，事奉上帝和不事奉上帝的人有何差别。”
MAL|4|1|万军之耶和华说：“看哪，那日临近，势如烧着的火炉，凡狂傲的和行恶的都如碎秸，在那日被烧尽，根与枝条无一存留。
MAL|4|2|但是，对你们敬畏我名的人，必有公义的太阳出现，其光线 有医治的能力。你们必出来跳跃如圈里的牛犊。
MAL|4|3|你们必践踏恶人；在我所定的日子，他们必成为你们脚掌下的灰尘。这是万军之耶和华说的。
MAL|4|4|“你们当记念我仆人 摩西 的律法，就是我在 何烈山 为 以色列 众人所吩咐他的律例典章。
MAL|4|5|“看哪，耶和华大而可畏之日未到以前，我要差遣 以利亚 先知到你们那里去。
MAL|4|6|他必使父亲的心转向儿女，儿女的心转向父亲，免得我来诅咒这地。”
MATT|1|1|亚伯拉罕 的后裔、 大卫 的子孙 耶稣基督的家谱：
MATT|1|2|亚伯拉罕 生 以撒 ， 以撒 生 雅各 ， 雅各 生 犹大 和他的兄弟，
MATT|1|3|犹大 从 她玛 氏生 法勒斯 和 谢拉 ， 法勒斯 生 希斯仑 ， 希斯仑 生 亚兰 ，
MATT|1|4|亚兰 生 亚米拿达 ， 亚米拿达 生 拿顺 ， 拿顺 生 撒门 ，
MATT|1|5|撒门 从 喇合 氏生 波阿斯 ， 波阿斯 从 路得 氏生 俄备得 ， 俄备得 生 耶西 ，
MATT|1|6|耶西 生 大卫 王。 大卫 从 乌利亚 的妻子生 所罗门 ，
MATT|1|7|所罗门 生 罗波安 ， 罗波安 生 亚比雅 ， 亚比雅 生 亚撒 ，
MATT|1|8|亚撒 生 约沙法 ， 约沙法 生 约兰 ， 约兰 生 乌西雅 ，
MATT|1|9|乌西雅 生 约坦 ， 约坦 生 亚哈斯 ， 亚哈斯 生 希西家 ，
MATT|1|10|希西家 生 玛拿西 ， 玛拿西 生 亚们 ， 亚们 生 约西亚 ，
MATT|1|11|百姓被迁到 巴比伦 的时候， 约西亚 生 耶哥尼雅 和他的兄弟。
MATT|1|12|迁到 巴比伦 之后， 耶哥尼雅 生 撒拉铁 ， 撒拉铁 生 所罗巴伯 ，
MATT|1|13|所罗巴伯 生 亚比玉 ， 亚比玉 生 以利亚敬 ， 以利亚敬 生 亚所 ，
MATT|1|14|亚所 生 撒督 ， 撒督 生 亚金 ， 亚金 生 以律 ，
MATT|1|15|以律 生 以利亚撒 ， 以利亚撒 生 马但 ， 马但 生 雅各 ，
MATT|1|16|雅各 生 约瑟 ，就是 马利亚 的丈夫；那称为基督的耶稣是从 马利亚 生的。
MATT|1|17|这样，从 亚伯拉罕 到 大卫 共有十四代，从 大卫 到迁至 巴比伦 的时候也有十四代，从迁至 巴比伦 的时候到基督又有十四代。
MATT|1|18|耶稣基督降生的事记在下面：他母亲 马利亚 已经许配给 约瑟 ，还没有迎娶， 马利亚 就从圣灵怀了孕。
MATT|1|19|她丈夫 约瑟 是个义人，不愿意当众羞辱她，想要暗地里把她休了。
MATT|1|20|正考虑这些事的时候，忽然主的使者在 约瑟 梦中向他显现，说：“ 大卫 的子孙 约瑟 ，不要怕，把你的妻子 马利亚 娶过来，因她所怀的孕是从圣灵来的。
MATT|1|21|她将要生一个儿子，你要给他起名叫耶稣，因他要将自己的百姓从罪恶里救出来。”
MATT|1|22|这整件事的发生，是要应验主藉先知所说的话：
MATT|1|23|“必有童女怀孕生子； 人要称他的名为 以马内利 。” （ 以马内利 翻出来就是“上帝与我们同在”。）
MATT|1|24|约瑟 醒来，就遵照主的使者的吩咐把妻子娶过来；
MATT|1|25|但是没有和她同房，直到她生了儿子 ，就给他起名叫耶稣。
MATT|2|1|在 希律 作王的时候，耶稣生在 犹太 的 伯利恒 。有几个博学之士 从东方来到 耶路撒冷 ，说：
MATT|2|2|“那生下来作 犹太 人之王的在哪里？我们在东方看见他的星，特来拜他。”
MATT|2|3|希律 王听见了，就心里不安； 耶路撒冷 全城的人也都不安。
MATT|2|4|他就召集了祭司长和民间的文士，问他们：“基督该生在哪里？”
MATT|2|5|他们说：“在 犹太 的 伯利恒 。因为有先知记着：
MATT|2|6|‘ 犹大 地的 伯利恒 啊， 你在 犹大 诸城中并不是最小的； 因为将来有一位统治者要从你那里出来， 牧养我 以色列 民。’”
MATT|2|7|于是， 希律 暗地里召了博学之士来，查问那星是什么时候出现的，
MATT|2|8|就派他们往 伯利恒 去，说：“你们去仔细寻访那小孩子，找到了就来报信，我也好去拜他。”
MATT|2|9|他们听了王的话就去了。忽然，在东方所看到的那颗星在前面引领他们，一直行到小孩子所在地方的上方就停住了。
MATT|2|10|他们看见那星，就非常欢喜；
MATT|2|11|进了房子，看见小孩子和他母亲 马利亚 ，就俯伏拜那小孩子，揭开宝盒，拿出黄金、乳香、没药，作为礼物献给他。
MATT|2|12|因为在梦中得到主的指示，不要回去见 希律 ，他们就从别的路回自己的家乡去了。
MATT|2|13|他们走后，忽然主的使者在 约瑟 梦中向他显现，说：“起来！带着小孩子和他母亲逃往 埃及 ，住在那里，等我的指示；因为 希律 要搜寻那小孩子来杀害他。”
MATT|2|14|约瑟 就起来，连夜带着小孩子和他母亲往 埃及 去，
MATT|2|15|住在那里，直到 希律 死了。这是要应验主藉先知所说的话：“我从 埃及 召我的儿子出来。”
MATT|2|16|希律 见自己被博学之士愚弄，极其愤怒，差人将 伯利恒 城里和四境所有的男孩，根据他向博学之士仔细查问到的时间，凡两岁以内的，都杀尽了。
MATT|2|17|这就应验了 耶利米 先知所说的话：
MATT|2|18|“在 拉玛 听见号啕大哭的声音， 是 拉结 哭她儿女； 她不肯受安慰， 因为他们都不在了。”
MATT|2|19|希律 死了以后，在 埃及 ，忽然主的使者在 约瑟 梦中向他显现，
MATT|2|20|说：“起来，带着小孩子和他母亲回 以色列 地去！因为要杀害这小孩子的人已经死了。”
MATT|2|21|约瑟 就起来，带着小孩子和他母亲进入 以色列 地去。
MATT|2|22|但是他因听见 亚基老 继承他父亲 希律 作了 犹太 王，怕到那里去；又在梦中得到主的指示，就往 加利利 境内去了。
MATT|2|23|他们到了一座城，名叫 拿撒勒 ，就住在那里。这是要应验先知所说的话：“他将称为 拿撒勒 人。”
MATT|3|1|在那些日子，施洗的 约翰 出来，在 犹太 的旷野宣讲：
MATT|3|2|“你们要悔改！因为天国近了。”
MATT|3|3|这人就是 以赛亚 先知所说的： “在旷野有声音呼喊着： 预备主的道， 修直他的路。”
MATT|3|4|这 约翰 身穿骆驼毛的衣服，腰束皮带，吃的是蝗虫和野蜜。
MATT|3|5|那时， 耶路撒冷 、全 犹太 和全 约旦河 地区的人，都到 约翰 那里去，
MATT|3|6|承认他们的罪，在 约旦河 里受他的洗。
MATT|3|7|约翰 看见许多法利赛人和撒都该人也来受洗，就对他们说：“毒蛇的孽种啊，谁指示你们逃避那将要来的愤怒呢？
MATT|3|8|你们要结出果子来，和悔改的心相称。
MATT|3|9|不要自己心里说：‘我们有 亚伯拉罕 为祖宗。’我告诉你们，上帝能从这些石头中给 亚伯拉罕 兴起子孙来。
MATT|3|10|现在斧子已经放在树根上，凡不结好果子的树就砍下来，丢在火里。
MATT|3|11|我是用水给你们施洗，叫你们悔改；但那在我以后来的，能力比我更大，我就是给他提鞋子也不配，他要用圣灵与火给你们施洗。
MATT|3|12|他手里拿着簸箕，要扬净他的谷物，把麦子收在仓里，把糠用不灭的火烧尽。”
MATT|3|13|当时，耶稣从 加利利 来到 约旦河 ，到了 约翰 那里，请 约翰 为他施洗。
MATT|3|14|约翰 想要阻止他，说：“我应该受你的洗，你怎么到我这里来呢？”
MATT|3|15|耶稣回答他：“暂且这样做吧，因为我们理当这样履行全部的义 。”于是 约翰 就依了他。
MATT|3|16|耶稣受了洗，随即从水里上来。天忽然为他 开了，他看见上帝的灵降下，仿佛鸽子落在他身上。
MATT|3|17|这时，天上有声音说：“这是我的爱子，我所喜爱的。”
MATT|4|1|当时，耶稣被圣灵引到旷野，受魔鬼的试探。
MATT|4|2|他禁食四十昼夜，后来就饿了。
MATT|4|3|那试探者进前来对他说：“你若是上帝的儿子，叫这些石头变成食物吧。”
MATT|4|4|耶稣却回答说：“经上记着： ‘人活着，不是单靠食物， 乃是靠上帝口里所出的一切话。’”
MATT|4|5|魔鬼就带他进了圣城，叫他站在圣殿顶上，
MATT|4|6|对他说：“你若是上帝的儿子，就跳下去！因为经上记着： ‘主要为你命令他的使者， 用手托住你， 免得你的脚碰在石头上。’”
MATT|4|7|耶稣对他说：“经上又记着：‘不可试探主—你的上帝。’”
MATT|4|8|魔鬼又带他上了一座很高的山，将世上的万国和万国的荣华都指给他看，
MATT|4|9|对他说：“你若俯伏拜我，我就把这一切赐给你。”
MATT|4|10|耶稣说：“撒但 ，退去！因为经上记着： ‘要拜主—你的上帝， 惟独事奉他。’”
MATT|4|11|于是，魔鬼离开了耶稣，立刻有天使来伺候他。
MATT|4|12|耶稣听见 约翰 下了监，就退到 加利利 去；
MATT|4|13|后来离开 拿撒勒 ，往 迦百农 去，住在那里。那地方靠海，在 西布伦 和 拿弗他利 地区。
MATT|4|14|这是要应验 以赛亚 先知所说的话：
MATT|4|15|“ 西布伦 ， 拿弗他利 ， 沿海的路， 约旦河 的东边， 外邦人的 加利利 —
MATT|4|16|那坐在黑暗里的百姓 看见了大光； 坐在死荫之地的人 有光照耀他们。”
MATT|4|17|从那时候，耶稣开始宣讲，说：“你们要悔改！因为天国近了。”
MATT|4|18|耶稣沿着 加利利 海边行走，看见两兄弟，就是那叫 彼得 的 西门 和他弟弟 安得烈 ，正往海里撒网；他们本是打鱼的。
MATT|4|19|耶稣对他们说：“来跟从我，我要叫你们得人如得鱼一样。”
MATT|4|20|他们立刻舍了网，跟从他。
MATT|4|21|耶稣从那里往前走，看见另外两兄弟，就是 西庇太 的儿子 雅各 和他弟弟 约翰 ，同他们的父亲 西庇太 在船上补网，耶稣就呼召他们。
MATT|4|22|他们立刻舍了船，辞别父亲，跟从了耶稣。
MATT|4|23|耶稣走遍 加利利 ，在各会堂里教导人，宣讲天国的福音，医治百姓各样的疾病。
MATT|4|24|他的名声传遍了 叙利亚 。那里的人把一切病人，就是有各样疾病和疼痛的、被鬼附的、癫痫的、瘫痪的，都带了来，耶稣就治好了他们。
MATT|4|25|当时，有一大群人从 加利利 、 低加坡里 、 耶路撒冷 、 犹太 、 约旦河 的东边，来跟从他。
MATT|5|1|耶稣看见这一群人，就上了山，坐下后，门徒到他跟前来，
MATT|5|2|他开口教导他们说：
MATT|5|3|“心灵贫穷的人有福了！ 因为天国是他们的。
MATT|5|4|哀恸的人有福了！ 因为他们必得安慰。
MATT|5|5|谦和的人有福了！ 因为他们必承受土地。
MATT|5|6|饥渴慕义的人有福了！ 因为他们必得饱足。
MATT|5|7|怜悯人的人有福了！ 因为他们必蒙怜悯。
MATT|5|8|清心的人有福了！ 因为他们必得见上帝。
MATT|5|9|缔造和平的人有福了！ 因为他们必称为上帝的儿子。
MATT|5|10|为义受迫害的人有福了！ 因为天国是他们的。
MATT|5|11|“人若因我辱骂你们，迫害你们，捏造各样坏话毁谤你们 ，你们就有福了！
MATT|5|12|要欢喜快乐，因为你们在天上的赏赐是很多的。在你们以前的先知，人也是这样迫害他们。”
MATT|5|13|“你们是地上的盐。盐若失了味，怎能叫它再咸呢？它不再有用，只好被丢在外面，任人践踏。
MATT|5|14|你们是世上的光。城造在山上是不能隐藏的。
MATT|5|15|人点灯，不放在斗底下，而是放在灯台上，就照亮一家的人。
MATT|5|16|你们的光也要这样照在人前，叫他们看见你们的好行为，把荣耀归给你们在天上的父。”
MATT|5|17|“不要以为我来是要废掉律法和先知。我来不是要废掉，而是要成全。
MATT|5|18|我实在告诉你们，就是到天地都废去，律法的一点一画也不能废去，直到一切都实现。
MATT|5|19|所以，无论谁废掉这诫命中最小的一条，又教导人也这样做，他在天国里要称为最小的。但无论谁遵行并如此教导人的，他在天国里要称为大。
MATT|5|20|我告诉你们，你们的义若不胜过文士和法利赛人的义，绝不能进天国。”
MATT|5|21|“你们听过有对古人说：‘不可杀人’；‘凡杀人的，必须受审判。’
MATT|5|22|但是我告诉你们：凡向弟兄动怒的，必须受审判；凡骂弟兄是废物的，必须受议会的审判；凡骂弟兄是白痴的，必须遭受地狱的火。
MATT|5|23|所以，你在祭坛上献祭物的时候，若想起有弟兄对你怀恨，
MATT|5|24|就要把祭物留在坛前，先去跟弟兄和好，然后来献祭物。
MATT|5|25|你同告你的冤家还在路上，就要赶快与他讲和，免得他把你送交给法官，法官交给警卫，你就下在监里了。
MATT|5|26|我实在告诉你，就是有一个大文钱 还没有还清，你也绝不能从那里出来。”
MATT|5|27|“你们听过有话说：‘不可奸淫。’
MATT|5|28|但是我告诉你们：凡看见妇女就动淫念的，这人心里已经与她犯奸淫了。
MATT|5|29|若是你的右眼使你跌倒，就把它挖出来，丢掉。宁可失去身体中的一部分，也不让整个身体被扔进地狱。
MATT|5|30|若是你的右手使你跌倒，就把它砍下来，丢掉。宁可失去身体中的一部分，也不让整个身体下地狱。”
MATT|5|31|“又有话说：‘无论谁休妻，都要给她休书。’
MATT|5|32|但是我告诉你们：凡休妻的，除非是因不贞的缘故，否则就是使她犯奸淫了；人若娶被休的妇人，也是犯奸淫了。”
MATT|5|33|“你们又听过有对古人说：‘不可背誓，所起的誓总要向主谨守。’
MATT|5|34|但是我告诉你们：什么誓都不可起。不可指着天起誓，因为天是上帝的宝座。
MATT|5|35|不可指着地起誓，因为地是他的脚凳；也不可指着 耶路撒冷 起誓，因为 耶路撒冷 是大君王的京城。
MATT|5|36|又不可指着你的头起誓，因为你不能使一根头发变黑变白。
MATT|5|37|你们的话，是，就说是；不是，就说不是。若再多说，就是出于那恶者。”
MATT|5|38|“你们听过有话说：‘以眼还眼，以牙还牙。’
MATT|5|39|但是我告诉你们：不要与恶人作对。有人打你的右脸，连另一边也转过去由他打。
MATT|5|40|有人想要告你，要拿你的里衣，连外衣也由他拿去。
MATT|5|41|有人强迫你走一里 路，你就跟他走二里。
MATT|5|42|有求你的，就给他；有向你借贷的，不可推辞。”
MATT|5|43|“你们听过有话说：‘要爱你的邻舍，恨你的仇敌。’
MATT|5|44|但是我告诉你们：要爱你们的仇敌，为那迫害你们的祷告。
MATT|5|45|这样，你们就可以作天父的儿女了。因为他叫太阳照好人，也照坏人；降雨给义人，也给不义的人。
MATT|5|46|你们若只爱那爱你们的人，有什么赏赐呢？就是税吏不也是这样做吗？
MATT|5|47|你们若只请你弟兄的安，有什么比别人强呢？就是外邦人不也是这样做吗？
MATT|5|48|所以，你们要完全，如同你们的天父是完全的。”
MATT|6|1|“你们要谨慎，不可故意在人面前表现虔诚，叫他们看见，若是这样，就不能得你们天父的赏赐了。
MATT|6|2|“所以，你施舍的时候，不可叫人在你前面吹号，像那假冒为善的人在会堂里和街道上所做的，故意要得人的称赞。我实在告诉你们，他们已经得了他们的赏赐。
MATT|6|3|你施舍的时候，不要让左手知道右手所做的，
MATT|6|4|好使你隐秘地施舍；你父在隐秘中察看，必然赏赐你。”
MATT|6|5|“你们祷告的时候，不可像那假冒为善的人，爱站在会堂里和十字路口祷告，故意让人看见。我实在告诉你们，他们已经得了他们的赏赐。
MATT|6|6|你祷告的时候，要进入内室，关上门，向那在隐秘中的父祷告；你父在隐秘中察看，必将赏赐你。
MATT|6|7|你们祷告，不可像外邦人那样重复一些空话，他们以为话多了必蒙垂听。
MATT|6|8|你们不可效法他们。因为在你们祈求以前，你们所需要的，你们的父早已知道了。”
MATT|6|9|“所以，你们要这样祷告： ‘我们在天上的父： 愿人都尊你的名为圣。
MATT|6|10|愿你的国降临； 愿你的旨意行在地上， 如同行在天上。
MATT|6|11|我们日用的饮食，今日赐给我们。
MATT|6|12|免我们的债， 如同我们免了人的债。
MATT|6|13|不叫我们陷入试探； 救我们脱离那恶者。 因为国度、权柄、荣耀，全是你的， 直到永远。阿们！ ’
MATT|6|14|“你们若饶恕人的过犯，你们的天父也必饶恕你们；
MATT|6|15|你们若不饶恕人 ，你们的天父也必不饶恕你们的过犯。”
MATT|6|16|“你们禁食的时候，不可像那假冒为善的人，脸上带着愁容；因为他们蓬头垢面，故意让人看出他们在禁食。我实在告诉你们，他们已经得了他们的赏赐。
MATT|6|17|你禁食的时候，要梳头洗脸，
MATT|6|18|不要让人看出你在禁食，只让你隐秘中的父看见；你父在隐秘中察看，必然赏赐你。”
MATT|6|19|“不要为自己在地上积蓄财宝；地上有虫子咬，能锈坏，也有贼挖洞来偷。
MATT|6|20|要在天上积蓄财宝；天上没有虫子咬，不会锈坏，也没有贼挖洞来偷。
MATT|6|21|因为你的财宝在哪里，你的心也在哪里。”
MATT|6|22|“眼睛是身体的灯。你的眼睛若明亮，全身就光明；
MATT|6|23|你的眼睛若昏花，全身就黑暗。你里面的光若黑暗了，那黑暗是何等大呢！”
MATT|6|24|“一个人不能服侍两个主；他不是恨这个爱那个，就是重这个轻那个。你们不能又服侍上帝，又服侍 玛门 。”
MATT|6|25|“所以，我告诉你们，不要为你们的生命忧虑吃什么喝什么 ，或为你们的身体忧虑穿什么。生命不胜于饮食吗？身体不胜于衣裳吗？
MATT|6|26|你们看一看那天上的飞鸟，也不种也不收，也不在仓里存粮，你们的天父尚且养活它们。你们不比飞鸟贵重得多吗？
MATT|6|27|你们哪一个能藉着忧虑使寿数多加一刻呢 ？
MATT|6|28|何必为衣裳忧虑呢？你们想一想野地里的百合花是怎么长起来的：它也不劳动也不纺线。
MATT|6|29|然而我告诉你们，就是 所罗门 极荣华的时候，他所穿戴的还不如这些花的一朵呢！
MATT|6|30|你们这小信的人哪！野地里的草今天还在，明天就丢在炉里，上帝还给它这样的妆饰，何况你们呢？
MATT|6|31|所以，不要忧虑，说：‘我们吃什么？喝什么？穿什么？’
MATT|6|32|这都是外邦人所求的。你们需要这一切东西，你们的天父都知道。
MATT|6|33|你们要先求上帝的国和他的义，这些东西都要加给你们了。
MATT|6|34|所以，不要为明天忧虑，因为明天自有明天的忧虑；一天的难处一天当就够了。”
MATT|7|1|“你们不要评断别人，免得你们被审判。
MATT|7|2|因为你们怎样评断别人，也必怎样被审判；你们用什么量器量给人，也必用什么量器量给你们。
MATT|7|3|为什么看见你弟兄眼中有刺，却不想自己眼中有梁木呢？
MATT|7|4|你自己眼中有梁木，怎能对你弟兄说‘让我去掉你眼中的刺’呢？
MATT|7|5|你这假冒为善的人！先去掉自己眼中的梁木，然后才能看得清楚，好去掉你弟兄眼中的刺。
MATT|7|6|不要把圣物给狗，也不要把你们的珍珠丢在猪面前，恐怕它们践踏了珍珠，转过来咬你们。”
MATT|7|7|“你们祈求，就给你们；寻找，就找到；叩门，就给你们开门。
MATT|7|8|因为凡祈求的，就得着；寻找的，就找到；叩门的，就给他开门。
MATT|7|9|你们中间谁有儿子求饼，反给他石头呢？
MATT|7|10|求鱼，反给他蛇呢？
MATT|7|11|你们虽然不好，尚且知道拿好东西给儿女，何况你们在天上的父，他岂不更要把好东西赐给求他的人吗？
MATT|7|12|所以，无论何事，你们想要人怎样待你们，你们也要怎样待人，因为这就是律法和先知的道理。”
MATT|7|13|“你们要进窄门。因为通往灭亡的门是宽的，路是大的，进去的人也多；
MATT|7|14|通往生命的门是窄的，路是小的，找到的人也少。”
MATT|7|15|“你们要防备假先知。他们到你们这里来，外面披着羊皮，里面却是残暴的狼。
MATT|7|16|岂能在荆棘上摘葡萄呢？岂能在蒺藜里摘无花果呢？凭着他们的果子，就可以认出他们来。
MATT|7|17|这样，凡好树都结好果子，而坏树结坏果子。
MATT|7|18|好树不能结坏果子，坏树也不能结好果子。
MATT|7|19|凡不结好果子的树就砍下来，丢在火里。
MATT|7|20|所以，凭着他们的果子就可以认出他们来。”
MATT|7|21|“不是每一个称呼我‘主啊，主啊’的人都能进天国；惟有遵行我天父旨意的人才能进去。
MATT|7|22|在那日必有许多人对我说：‘主啊，主啊，我们不是奉你的名传道，奉你的名赶鬼，奉你的名行许多异能吗？’
MATT|7|23|我要向他们宣告：‘我从来不认识你们，你们这些作恶的人，给我走开！’”
MATT|7|24|“所以，凡听了我这些话又去做的，好比一个聪明人把房子盖在磐石上。
MATT|7|25|风吹，雨打，水冲，撞击那房子，房子总不倒塌，因为根基立在磐石上。
MATT|7|26|凡听了我这些话而不去做的，好比一个无知的人把房子盖在沙土上。
MATT|7|27|风吹，雨打，水冲，撞击那房子，房子就倒塌了，并且倒塌得很厉害。”
MATT|7|28|耶稣讲完了这些话，众人对他的教导都感到惊奇，
MATT|7|29|因为他教导他们正像有权柄的人，不像他们的文士。
MATT|8|1|耶稣下了山，有一大群人跟着他。
MATT|8|2|这时，一个痲疯病人前来拜他，说：“主啊，你若肯，你能使我洁净。”
MATT|8|3|耶稣伸手摸他，说：“我肯，你洁净了吧！”他的痲疯病立刻就洁净了。
MATT|8|4|耶稣对他说：“你要注意，不可告诉任何人，只要去，让祭司为你检查，并献上 摩西 所吩咐的祭物，作为证据给众人看。”
MATT|8|5|耶稣进了 迦百农 ，有一个百夫长进前来，求他，
MATT|8|6|说：“主啊，我的僮仆瘫痪了，躺在家里，非常痛苦。”
MATT|8|7|耶稣说：“我去医治他。”
MATT|8|8|百夫长回答：“主啊，你到舍下来，我不敢当；只要你说一句话，我的僮仆就会痊愈。
MATT|8|9|因为我在人的权下，也有兵在我以下。我对这个说：‘去！’他就去；对那个说：‘来！’他就来；对我的仆人说：‘做这事！’他就去做。”
MATT|8|10|耶稣听了就很惊讶，对跟从的人说：“我实在告诉你们，这么大的信心，就是在 以色列 ，我也没有见过。
MATT|8|11|我又告诉你们，从东从西，将有许多人来，在天国里与 亚伯拉罕 、 以撒 、 雅各 一同坐席；
MATT|8|12|本国的子民反而被赶到外边黑暗里去，在那里要哀哭切齿了。”
MATT|8|13|耶稣对百夫长说：“你回去吧！照你的信心成全你了。”就在那时，他的僮仆好了。
MATT|8|14|耶稣到了 彼得 家里，见 彼得 的岳母正发烧躺着。
MATT|8|15|耶稣一摸她的手，烧就退了，于是她起来服事耶稣。
MATT|8|16|傍晚的时候，有人带着许多被鬼附的来到耶稣跟前，他只用一句话就把邪灵都赶出去，并且治好了一切有病的人。
MATT|8|17|这是要应验 以赛亚 先知所说的话： “他代替了我们的软弱， 担当了我们的疾病。”
MATT|8|18|耶稣见许多人围着他，就吩咐渡到对岸去。
MATT|8|19|有一个文士进前来对他说：“老师，你无论往哪里去，我都要跟从你。”
MATT|8|20|耶稣说：“狐狸有洞，天空的飞鸟有窝，人子却没有枕头的地方。”
MATT|8|21|又有一个门徒对耶稣说：“主啊，容许我先回去埋葬我的父亲。”
MATT|8|22|耶稣说：“让死人埋葬他们的死人。你跟从我吧！”
MATT|8|23|耶稣上了船，门徒跟着他。
MATT|8|24|海里忽然起了猛烈的风暴，以致船几乎被波浪淹没，耶稣却睡着了。
MATT|8|25|门徒去叫醒他，说：“主啊，救命啊，我们快没命啦！”
MATT|8|26|耶稣说：“你们这些小信的人哪，为什么胆怯呢？”于是他起来，斥责风和海，风和海就大大平静了。
MATT|8|27|众人惊讶地说：“这是怎样的一个人？连风和海都听从他。”
MATT|8|28|耶稣渡到对岸去，到 加大拉 人 的地区，有两个被鬼附的人从坟墓迎着他走来。他们极其凶猛，甚至没有人敢从那条路经过。
MATT|8|29|他们喊着说：“上帝的儿子，你为什么干扰我们？时候还没有到，你就上这里来叫我们受苦吗？”
MATT|8|30|离他们很远，有一大群猪正在吃食。
MATT|8|31|鬼就央求耶稣，说：“若要把我们赶出去，就打发我们进入猪群吧！”
MATT|8|32|耶稣对他们说：“去吧！”鬼就出来，进入猪群。一转眼，整群猪都闯下山崖，投进海里，淹死了。
MATT|8|33|放猪的就逃进城去，把这一切事和被鬼附的人所遭遇的都告诉众人。
MATT|8|34|全城的人都出来迎见耶稣，见了他以后，就央求他离开他们的地区。
MATT|9|1|耶稣上了船，渡过海，来到自己的城里。
MATT|9|2|有人用褥子抬着一个瘫子到耶稣跟前来。耶稣见他们的信心，就对瘫子说：“孩子，放心吧，你的罪赦了。”
MATT|9|3|这时，有几个文士心里说：“这个人说亵渎的话了。”
MATT|9|4|耶稣知道他们的心思，就说：“你们心里为什么怀着恶念呢？
MATT|9|5|说‘你的罪赦了’，或说‘你起来行走’，哪一样容易呢？
MATT|9|6|但要让你们知道，人子在地上有赦罪的权柄”，于是对瘫子说：“起来！拿你的褥子回家去吧。”
MATT|9|7|那人就起来，回家去了。
MATT|9|8|众人看见都畏惧，归荣耀给上帝，因为他把这样的权柄赐给人。
MATT|9|9|耶稣从那里往前走，看见一个人名叫 马太 ，在税关坐着，就对他说：“来跟从我！”他就起来跟从耶稣。
MATT|9|10|耶稣在屋里坐席的时候，有好些税吏和罪人来，与耶稣和他的门徒一同坐席。
MATT|9|11|法利赛人看见，就对耶稣的门徒说：“你们的老师为什么与税吏和罪人一同吃饭呢？”
MATT|9|12|耶稣听见，就说：“健康的人用不着医生；有病的人才用得着。
MATT|9|13|经上说：‘我喜爱怜悯，不喜爱祭祀。’这句话的意思，你们去揣摩。我不是来召义人，而是召罪人。”
MATT|9|14|那时， 约翰 的门徒来见耶稣，说：“我们和法利赛人常常 禁食，你的门徒却不禁食，这是为什么呢？”
MATT|9|15|耶稣对他们说：“新郎和宾客在一起的时候，宾客怎么能哀恸呢？但日子将到，新郎要被带走，那时候他们就要禁食了。
MATT|9|16|没有人把新布补在旧衣服上；因为所补上的会撕破那衣服，裂口就更大了。
MATT|9|17|也没有人把新酒装在旧皮袋里，若是这样，皮袋会胀破，酒就漏出来，皮袋也糟蹋了。相反地，把新酒装在新皮袋里，两样就都保全了。”
MATT|9|18|耶稣说这些话的时候，有一个会堂主管来，向他下跪，说：“我女儿刚死了，求你去按手在她身上，她就会活过来。”
MATT|9|19|耶稣就起来跟他去；门徒也跟了去。
MATT|9|20|这时，有一个女人，患了经血不止的病有十二年，来到耶稣背后，摸他的衣裳繸子；
MATT|9|21|因为她心里说：“我只要摸他的衣裳，就会痊愈。”
MATT|9|22|耶稣转过来，看见她，就说：“女儿，放心！你的信救了你。”从那时起，这女人就痊愈了。
MATT|9|23|耶稣到了会堂主管的家里，看见吹鼓手和乱哄哄的一群人，
MATT|9|24|就说：“退去吧！这女孩不是死了，而是睡着了。”他们就嘲笑他。
MATT|9|25|众人被赶出后，耶稣就进去，拉着女孩的手，女孩就起来了。
MATT|9|26|于是这消息传遍了那地方。
MATT|9|27|耶稣从那里往前走，有两个盲人跟着他，喊叫说：“ 大卫 之子，可怜我们吧！”
MATT|9|28|耶稣进了屋子，盲人就来到他跟前。耶稣说：“你们信我能做这事吗？”他们说：“主啊，我们信。”
MATT|9|29|耶稣就摸他们的眼睛，说：“照着你们的信心成全你们吧。”
MATT|9|30|他们的眼睛就开了。耶稣严严地叮嘱他们说：“要小心，不可让人知道。”
MATT|9|31|他们出去，竟把他的名声传遍了那地方。
MATT|9|32|他们出去的时候，有人把一个被鬼附的哑巴带到耶稣跟前来。
MATT|9|33|鬼被赶出去，哑巴就说出话来。众人都很惊讶，说：“在 以色列 ，从来没有见过这样的事。”
MATT|9|34|法利赛人却说：“他是靠着鬼王赶鬼的。”
MATT|9|35|耶稣走遍各城各乡，在他们的会堂里教导人，宣讲天国的福音，又医治各样的病症。
MATT|9|36|他看见一大群人，就怜悯他们；因为他们困苦无助，如同羊没有牧人一样。
MATT|9|37|于是他对门徒说：“要收的庄稼多，做工的人少。
MATT|9|38|所以，你们要求庄稼的主差遣做工的人出去收他的庄稼。”
MATT|10|1|耶稣叫了十二个门徒来，给他们权柄，能驱赶污灵和医治各样的疾病。
MATT|10|2|这十二使徒的名字如下：头一个叫 西门 （又称 彼得 ），还有他弟弟 安得烈 ， 西庇太 的儿子 雅各 和 雅各 的弟弟 约翰 ，
MATT|10|3|腓力 和 巴多罗买 ， 多马 和税吏 马太 ， 亚勒腓 的儿子 雅各 ，和 达太 ，
MATT|10|4|激进党的 西门 ，还有出卖耶稣的 加略 人 犹大 。
MATT|10|5|耶稣差遣这十二个人出去，吩咐他们说：“外邦人的路，你们不要走； 撒玛利亚 人的城，你们不要进；
MATT|10|6|宁可往 以色列 家迷失的羊那里去。
MATT|10|7|要边走边传，说‘天国近了’。
MATT|10|8|要医治病人，使死人复活，使痲疯病人洁净，把鬼赶出去。你们白白地得来，也要白白地给人。
MATT|10|9|腰袋里不要带金银铜钱；
MATT|10|10|途中不要带行囊，不要带两件内衣，也不要带鞋子和手杖，因为工人得饮食是应当的。
MATT|10|11|你们无论进哪一城、哪一村，要打听那里谁是合适的人，就住在他家，直住到离开的时候。
MATT|10|12|进他家时，要向那家请安。
MATT|10|13|那家若配得平安，你们所求的平安就临到那家；若不配得，你们所求的平安仍归你们。
MATT|10|14|凡不接待你们，不听你们话的人，你们离开那家，或是那城的时候，要跺掉你们脚上的尘土。
MATT|10|15|我实在告诉你们，在审判的日子， 所多玛 和 蛾摩拉 地方所受的，比那城还容易受呢！”
MATT|10|16|“看哪！我差你们出去，如同羊进入狼群，所以你们要机警如蛇，纯真如鸽。
MATT|10|17|你们要防备那些人，因为他们要把你们交给议会，也要在会堂里鞭打你们。
MATT|10|18|你们要为我的缘故被送到统治者和君王面前，对他们和外邦人作见证。
MATT|10|19|当人把你们交出时，不要担心怎样说话，或说什么话。到那时候，必赐给你们该说的话，
MATT|10|20|因为不是你们自己说的，而是你们父的灵在你们里面说的。
MATT|10|21|兄弟要把兄弟、父亲要把儿女置于死地；儿女要起来与父母为敌，害死他们。
MATT|10|22|而且你们要为我的名被众人憎恨。但坚忍到底的终必得救。
MATT|10|23|有人在这城迫害你们，就逃到另一城去。 我实在告诉你们， 以色列 的城镇，你们还没有走遍，人子就要来临。
MATT|10|24|“学生不高过老师，仆人不高过主人。
MATT|10|25|学生所遭遇的与老师一样，仆人所遭遇的与主人一样，也就够了。既然有人骂一家的主人是‘ 别西卜 ’ ，更何况他的家人呢？”
MATT|10|26|“所以，不要怕他们，因为掩盖的事没有不显露出来的，隐藏的事也没有不被知道的。
MATT|10|27|我在暗中告诉你们的，你们要在明处说出来；你们耳中所听的，要在屋顶上宣扬出来。
MATT|10|28|那杀人身体但不能灭人灵魂的，不要怕他们；惟有那能在地狱里毁灭身体和灵魂的，才要怕他。
MATT|10|29|两只麻雀不是卖一铜钱 吗？你们的父若不许，一只也不会掉在地上。
MATT|10|30|就是你们的头发也都数过了。
MATT|10|31|所以，不要惧怕，你们比许多的麻雀还贵重！”
MATT|10|32|“所以，凡在人面前认我的，我在我天上的父面前也必认他；
MATT|10|33|凡在人面前不认我的，我在我天上的父面前也必不认他。”
MATT|10|34|“你们不要以为我来是带给地上和平，我来并不是带来和平，而是刀剑。
MATT|10|35|因为我来是要叫 ‘人与父亲对立， 女儿与母亲对立， 媳妇与婆婆对立。
MATT|10|36|人的仇敌就是自己家里的人。’
MATT|10|37|爱父母胜过爱我的，不配作我的门徒；爱儿女胜过爱我的，不配作我的门徒。
MATT|10|38|不背自己的十字架跟从我的，不配作我的门徒。
MATT|10|39|得着性命的，要丧失性命；为我丧失性命的，要得着性命。”
MATT|10|40|“接纳你们的就是接纳我；接纳我的就是接纳差遣我来的那位。
MATT|10|41|把先知当作先知接纳的，必得先知的赏赐；把义人当作义人接纳的，必得义人的赏赐。
MATT|10|42|无论谁，只因门徒的名，就算把一杯凉水给这些小子中的一个喝，我实在告诉你们，他一定会得到赏赐。”
MATT|11|1|耶稣吩咐完了十二个门徒，就离开那里，往各城去传道，教导人。
MATT|11|2|约翰 在监狱里听见基督所做的事，就派他的门徒去，
MATT|11|3|问耶稣：“将要来的那位就是你吗？还是我们要等候另一位呢？”
MATT|11|4|耶稣回答他们：“你们去，把所听见、所看见的告诉 约翰 ：
MATT|11|5|就是盲人看见，瘸子行走，痲疯病人得洁净，聋子听见，死人复活，穷人听到福音。
MATT|11|6|凡不因我跌倒的有福了！”
MATT|11|7|他们一走，耶稣就对众人谈到 约翰 ，说：“你们从前到旷野去，是要看什么呢？看风吹动的芦苇吗？
MATT|11|8|你们出去到底是要看什么？看穿细软衣服的人吗？那穿细软衣服的人是在王宫里。
MATT|11|9|你们出去究竟是要看什么？是先知吗？是的，我告诉你们，他比先知大多了。
MATT|11|10|这个人就是经上所说的： ‘看哪，我要差遣我的使者在你面前， 他要在你前面为你预备道路。’
MATT|11|11|我实在告诉你们，凡女子所生的，没有一个比施洗 约翰 大；但在天国里，最小的比他还大。
MATT|11|12|从施洗 约翰 的日子到今天，天国受到强烈的攻击，强者夺取它 。
MATT|11|13|众先知和律法，直到 约翰 为止，都说了预言。
MATT|11|14|如果你们愿意接受，这人就是那要来的 以利亚 。
MATT|11|15|有耳的，就应当听！
MATT|11|16|“我该用什么来比这世代呢？这正像孩童坐在街市上向同伴呼喊：
MATT|11|17|‘我们为你们吹笛，你们不跳舞； 我们唱哀歌，你们不捶胸。’
MATT|11|18|约翰 来了，既不吃也不喝，人们就说他是被鬼附的；
MATT|11|19|人子来了，也吃也喝，他们又说这人贪食好酒，是税吏和罪人的朋友。而智慧是由它的果子来证实的 。”
MATT|11|20|那时，耶稣在一些城行了许多异能。因为城里的人不肯悔改，他就责备那些城说：
MATT|11|21|“ 哥拉汛 哪，你有祸了！ 伯赛大 啊，你有祸了！因为在你们中间所行的异能若行在 推罗 、 西顿 ，他们早已披麻蒙灰悔改了。
MATT|11|22|但我告诉你们，在审判的日子， 推罗 和 西顿 所受的，比你们还容易受呢！
MATT|11|23|迦百农 啊， 你以为要被举到天上吗？ 你要被推下阴间！ 因为在你那里所行的异能，若行在 所多玛 ，它还可以存留到今日。
MATT|11|24|但我告诉你们，在审判的日子， 所多玛 地方所受的，比你们还容易受呢！”
MATT|11|25|那时，耶稣说：“父啊，天地的主，我感谢你！因为你把这些事向聪明智慧的人隐藏起来，而向婴孩启示出来。
MATT|11|26|父啊，是的，因为你的美意本是如此。
MATT|11|27|一切都是我父交给我的；除了父，没有人知道子；除了子和子所愿意启示的人，没有人知道父。
MATT|11|28|凡劳苦担重担的人都到我这里来，我要使你们得安息。
MATT|11|29|我心里柔和谦卑，你们当负我的轭，向我学习；这样，你们的心灵就必得安息。
MATT|11|30|因为我的轭是容易的，我的担子是轻省的。”
MATT|12|1|那时，耶稣在安息日从麦田经过。他的门徒饿了，就摘麦穗来吃。
MATT|12|2|法利赛人看见，对耶稣说：“看哪，你的门徒在安息日做不合法的事了。”
MATT|12|3|耶稣对他们说：“ 大卫 和跟从他的人饥饿时所做的事，你们没有念过吗？
MATT|12|4|他怎么进了上帝的居所，吃了供饼呢？这饼是他和跟从他的人不可以吃的，惟独祭司才可以吃。
MATT|12|5|再者，律法上所记的，在安息日，祭司在圣殿里犯了安息日也不算有罪，你们没有念过吗？
MATT|12|6|但我告诉你们，比圣殿更大的在这里。
MATT|12|7|‘我喜爱怜悯，不喜爱祭祀。’你们若明白这话的意思，就不将无罪的当作有罪了。
MATT|12|8|因为人子是安息日的主。”
MATT|12|9|耶稣离开那地方，进了 犹太 人的会堂；
MATT|12|10|那里有个一只手萎缩了的人。有人为了要控告耶稣，就问他：“安息日治病合不合法？”
MATT|12|11|耶稣对他们说：“你们中间谁有一只羊在安息日掉在坑里，不抓住它，把它拉上来呢？
MATT|12|12|人比羊贵重得多了！所以，在安息日做善事是合法的。”
MATT|12|13|于是对那人说：“伸出手来！”他把手一伸，手就复原了，和另一只一样。
MATT|12|14|法利赛人出去，商议怎样除掉耶稣。
MATT|12|15|耶稣知道了，就离开那里，有一大群人跟着他。他把所有的病人都治好了，
MATT|12|16|又嘱咐他们不要把他宣扬出去。
MATT|12|17|这是要应验 以赛亚 先知所说的话：
MATT|12|18|“看哪，我所拣选的仆人， 我所亲爱，心所喜悦的； 我要将我的灵赐给他， 他必将公理传给外邦。
MATT|12|19|他不争吵，不喧嚷， 街上也没有人听见他的声音。
MATT|12|20|压伤的芦苇，他不折断， 将残的灯火，他不吹灭， 直到他使公理得胜。
MATT|12|21|外邦人都要仰望他的名。”
MATT|12|22|当时，有人把一个被鬼附，又盲又哑的人带到耶稣那里，耶稣医治他，那哑巴就能说话，又能看见。
MATT|12|23|众人都惊奇，说：“这不是 大卫 之子吗？”
MATT|12|24|但法利赛人听见，就说：“这个人赶鬼，无非是靠着鬼王 别西卜 罢了。”
MATT|12|25|耶稣知道他们的心思，就对他们说：“一国自相纷争，必定荒芜；一城一家自相纷争，必立不住。
MATT|12|26|若撒但赶出撒但，就是自相纷争，他的国怎能立得住呢？
MATT|12|27|我若靠着 别西卜 赶鬼，你们的子弟赶鬼又靠着谁呢？这样，他们要作你们的判官。
MATT|12|28|我若靠着上帝的灵赶鬼，那么，上帝的国就已临到你们了。
MATT|12|29|人怎能进壮士家里抢夺他的东西呢？除非先绑住那壮士，否则无法抢夺他的家。
MATT|12|30|不跟我一起的，就是反对我；不与我一起收聚的，就是在拆散。
MATT|12|31|所以我告诉你们，人一切的罪和亵渎的话都可得赦免，但是亵渎圣灵，总不得赦免。
MATT|12|32|凡说话干犯人子的，还可得赦免；但是说话干犯圣灵的，今世来世总不得赦免。”
MATT|12|33|“你们知道树好，果子也好；又知道树坏，果子也坏；因为看果子就可以知道树。
MATT|12|34|毒蛇的孽种啊，你们既是恶人，怎能说出好话来呢？因为心里所充满的，口里就说出来。
MATT|12|35|善人从他所存的善发出善来；恶人从他所存的恶发出恶来。
MATT|12|36|我告诉你们，凡是人所说的闲话，在审判的日子，要句句供出来；
MATT|12|37|因为要凭你的话定你为义，也要凭你的话定你有罪。”
MATT|12|38|当时，有几个文士和法利赛人对耶稣说：“老师，我们想请你显个神迹给我们看看。”
MATT|12|39|耶稣回答他们：“邪恶淫乱的世代求看神迹，除了先知 约拿 的神迹以外，再没有神迹给他们看了。
MATT|12|40|约拿 三日三夜在大鱼肚腹中，同样，人子也要三日三夜在地里面。
MATT|12|41|在审判的时候， 尼尼微 人要起来定这世代的罪，因为 尼尼微 人听了 约拿 所传的就悔改了。看哪，比 约拿 更大的在这里！
MATT|12|42|在审判的时候，南方的女王要起来定这世代的罪，因为她从地极而来，要听 所罗门 智慧的话。看哪，比 所罗门 更大的在这里！”
MATT|12|43|“污灵离了人身，走遍无水之地寻找安歇之处，却找不到。
MATT|12|44|于是他说：‘我要回到我原来的屋里去。’他到了，看见里面空着，打扫干净，修饰好了，
MATT|12|45|就去另带了七个比自己更恶的灵来，都进去住在那里。那人后来的景况比先前更坏了。这邪恶的世代也要如此。”
MATT|12|46|耶稣还在对众人说话的时候，不料，他母亲和他兄弟站在外边想要跟他说话。
MATT|12|47|有人告诉他：“看哪！你母亲和你兄弟站在外边，想要跟你说话。”
MATT|12|48|他却回答那对他说话的人，说：“谁是我的母亲？谁是我的兄弟？”
MATT|12|49|于是他伸手指着门徒，说：“看哪，我的母亲，我的兄弟！
MATT|12|50|凡遵行我天父旨意的人就是我的兄弟、姊妹和母亲。”
MATT|13|1|就在那天，耶稣从房子里出来，坐在海边。
MATT|13|2|有一大群人到他那里聚集，他只好上船坐下，众人都站在岸上。
MATT|13|3|他用比喻对他们讲了许多话。他说：“有一个撒种的出去撒种。
MATT|13|4|他撒的时候，有的落在路旁，飞鸟来把它们吃掉了。
MATT|13|5|有的落在土浅的石头地上，因为土不深，很快就长出苗来，
MATT|13|6|太阳出来一晒，因为没有根就枯干了。
MATT|13|7|有的落在荆棘里，荆棘长起来，把它挤住了。
MATT|13|8|又有的落在好土里，就结出果实，有一百倍的，有六十倍的，有三十倍的。
MATT|13|9|有耳的，就应当听！”
MATT|13|10|门徒进前来问耶稣：“对众人讲话，为什么用比喻呢？”
MATT|13|11|耶稣回答他们说：“因为天国的奥秘只让你们知道，不让他们知道。
MATT|13|12|凡有的，还要给他，让他有余；凡没有的，连他所有的也要夺去。
MATT|13|13|我之所以用比喻对他们讲，是因为 他们看却看不清， 听却听不见，也不明白。
MATT|13|14|在他们身上，正应验了 以赛亚 的预言： ‘你们听了又听，却不明白， 看了又看，却看不清。
MATT|13|15|因为这百姓的心麻木， 耳朵发沉， 眼睛闭着， 免得眼睛看见， 耳朵听见， 心里明白，回转过来， 我会医治他们。’
MATT|13|16|但你们的眼睛是有福的，因为看得见；你们的耳朵也是有福的，因为听得见。
MATT|13|17|我实在告诉你们，从前有许多先知和义人要看你们所看的，却没有看见；要听你们所听的，却没有听见。”
MATT|13|18|“所以，你们要听这撒种的比喻。
MATT|13|19|凡听见天国的道而不明白的，那恶者就来，把撒在他心里的夺了去；这就是撒在路旁的了。
MATT|13|20|撒在石头地上的，就是人听了道，立刻欢喜领受，
MATT|13|21|只因心里没有根，不过是暂时的，一旦为道遭受患难或迫害，立刻就跌倒。
MATT|13|22|撒在荆棘里的，就是人听了道，后来有世上的忧虑、钱财的迷惑把道挤住了，结不出果实。
MATT|13|23|撒在好土里的，就是人听了道，明白了，后来结了果实，有一百倍的，有六十倍的，有三十倍的。”
MATT|13|24|耶稣又设个比喻对他们说：“天国好比人撒好种在田里，
MATT|13|25|在人睡觉的时候，他的仇敌来，把杂草撒在麦子里就走了。
MATT|13|26|到长苗吐穗的时候，杂草也显出来。
MATT|13|27|地主的仆人进前来对他说：‘主人，你不是撒好种在田里吗？哪里来的杂草呢？’
MATT|13|28|主人回答他们：‘这是仇敌做的。’仆人对他说：‘你要我们去拔掉吗？’
MATT|13|29|主人说：‘不必，恐怕拔杂草，也把麦子连根拔出来。
MATT|13|30|让这两样一起长，等到收割。当收割的时候，我会对收割的人说，先把杂草拔出来，捆成捆，留着烧，把麦子收在我的仓里。’”
MATT|13|31|他又设个比喻对他们说：“天国好比一粒芥菜种，有人拿去种在田里。
MATT|13|32|它原比所有的种子都小，等到长起来，却比各样的菜都大，且成了树，以致天上的飞鸟来在它的枝上筑巢。”
MATT|13|33|他又对他们讲另一个比喻：“天国好比面酵，有妇人拿来放进三斗面里，直到全团都发起来。”
MATT|13|34|这都是耶稣用比喻对众人说的话，不用比喻，他就不对他们说什么。
MATT|13|35|这是要应验先知 所说的话： “我要开口说比喻， 说出从创世以来所隐藏的事。”
MATT|13|36|当时，耶稣离开众人，进了屋子。他的门徒进前来，说：“请把田间杂草的比喻讲给我们听。”
MATT|13|37|他回答：“那撒好种的就是人子，
MATT|13|38|田地就是世界，好种就是天国之子，杂草就是那恶者之子，
MATT|13|39|撒杂草的仇敌就是魔鬼，收割的时候就是世代的终结，收割的人就是天使。
MATT|13|40|正如把杂草拔出来用火焚烧，世代的终结也要如此。
MATT|13|41|人子要差遣他的使者，把一切使人跌倒的和作恶的从他国里挑出来，
MATT|13|42|丢在火炉里，在那里要哀哭切齿了。
MATT|13|43|那时，义人要在他们父的国里发出光来，像太阳一样。有耳的，就应当听！”
MATT|13|44|“天国好比宝贝藏在地里，人发现了就把它藏起来，欢欢喜喜地去变卖一切所有的，买这块地。
MATT|13|45|“天国又好比商人寻找好的珍珠，
MATT|13|46|发现一颗贵重的珍珠，就去变卖他一切所有的，买下这颗珍珠。”
MATT|13|47|“天国又好比网撒在海里，聚拢各种鱼类，
MATT|13|48|网一满，人们就把它拉上岸，坐下来，拣好的收在桶里，不好的丢掉。
MATT|13|49|世代的终结也要这样：天使要出来，把恶人从义人中分别出来，
MATT|13|50|丢在火炉里，在那里要哀哭切齿了。”
MATT|13|51|耶稣说：“这一切的话你们都明白了吗？”他们对他说：“明白了。”
MATT|13|52|他对他们说：“凡文士学习作天国的门徒，就像一个家的主人从他库里拿出新的和旧的东西来。”
MATT|13|53|耶稣说完了这些比喻，就离开那里，
MATT|13|54|来到自己的家乡，在会堂里教导人，以致他们都很惊奇，说：“这人哪来这样的智慧和异能呢？
MATT|13|55|这不是那木匠的儿子吗？他母亲不是叫 马利亚 吗？他兄弟们不是叫 雅各 、 约瑟 、 西门 、 犹大 吗？
MATT|13|56|他姊妹们不是都在我们这里吗？他这一切是从哪里来的呢？”
MATT|13|57|他们就厌弃他。耶稣对他们说：“先知除了在本乡和自己的家之外，没有不被尊敬的。”
MATT|13|58|耶稣因为他们不信，没有在那里行很多异能。
MATT|14|1|那时， 希律 分封王听见耶稣的名声，
MATT|14|2|就对臣仆说：“这是施洗的 约翰 从死人中复活，因此才有这些异能在他里面运行。”
MATT|14|3|原来， 希律 为他兄弟 腓力 的妻子 希罗底 的缘故，把 约翰 抓住绑了，关进监狱，
MATT|14|4|因为 约翰 曾对他说：“你占有这妇人是不合法的。”
MATT|14|5|希律 就想要杀他，可是怕民众，因为他们认为 约翰 是先知。
MATT|14|6|到了 希律 的生日， 希罗底 的女儿在众人面前跳舞，使 希律 欢喜，
MATT|14|7|于是 希律 发誓许诺随她所求的给她。
MATT|14|8|女儿被母亲指使，就说：“请把施洗 约翰 的头放在盘子里，拿来给我。”
MATT|14|9|王就忧愁，然而因他所发的誓，又因同席的人，就下令给她；
MATT|14|10|于是打发人去，在监狱里斩了 约翰 ，
MATT|14|11|把头放在盘子里，拿来给那女孩，她拿去给她母亲。
MATT|14|12|约翰 的门徒来，把尸体领去埋葬了，又去告诉耶稣。
MATT|14|13|耶稣听到了，就从那里上船，私下退到荒野的地方去。众人听到后，从各城来，步行跟随他。
MATT|14|14|耶稣出来，见有一大群人，就怜悯他们，治好了他们的病人。
MATT|14|15|傍晚的时候，门徒进前来，说：“这地方偏僻，而且时候已经晚了，请叫众人散去，他们好进村子，自己买些食物。”
MATT|14|16|耶稣对他们说：“不用他们去，你们给他们吃吧！”
MATT|14|17|门徒说：“我们这里只有五个饼、两条鱼。”
MATT|14|18|耶稣说：“拿过来给我。”
MATT|14|19|于是他吩咐众人坐在草地上，就拿着这五个饼和两条鱼，望着天祝福，擘开饼，递给门徒，门徒又递给众人。
MATT|14|20|他们都吃，并且吃饱了。门徒把剩下的碎屑收拾起来，装满了十二个篮子。
MATT|14|21|吃的人中，男的约有五千，还不算妇女和孩子。
MATT|14|22|耶稣随即催门徒上船，先渡到对岸，等他叫众人散去。
MATT|14|23|疏散了众人以后，他独自上山去祷告。到了晚上，只有他一人在那里。
MATT|14|24|那时船已离岸好几里 ，因风不顺，被浪颠簸。
MATT|14|25|天快亮的时候，耶稣在海面上走，往门徒那里去。
MATT|14|26|但门徒看见他在海面上走，就惊慌了，说：“是个鬼怪！”他们害怕得喊叫起来。
MATT|14|27|耶稣连忙对他们说：“放心！是我，不要怕！”
MATT|14|28|彼得 回答他说：“主啊，如果是你，请叫我从水面上走到你那里去。”
MATT|14|29|耶稣说：“你来吧！” 彼得 就从船上下去，在水面上走，往耶稣那里去；
MATT|14|30|只因见风很强 ，害怕起来，将要沉下去，就喊着说：“主啊，救我！”
MATT|14|31|耶稣立刻伸手拉住他，说：“你这小信的人哪，为什么疑惑呢？”
MATT|14|32|他们一上船，风就停了。
MATT|14|33|在船上的人都拜他，说：“你真是上帝的儿子。”
MATT|14|34|他们渡过了海，在 革尼撒勒 上岸。
MATT|14|35|那里的人认出耶稣，就打发人到整个周围地区去，把所有的病人带到他那里，
MATT|14|36|求耶稣让他们只摸一摸他的衣裳繸子，摸着的人就都好了。
MATT|15|1|那时，有法利赛人和文士从 耶路撒冷 来见耶稣，说：
MATT|15|2|“你的门徒为什么违反古人的传统？因为他们吃饭的时候不洗手。”
MATT|15|3|耶稣回答他们：“你们为什么因你们的传统而违反上帝的诫命呢？
MATT|15|4|上帝说：‘当孝敬父母’；又说：‘咒骂父母的，必须处死。’
MATT|15|5|你们倒说：‘无论谁对父母说：我所当供奉你的已经作了奉献，
MATT|15|6|就可以不孝敬他的父亲 。’这就是你们藉着传统，废了上帝的话。
MATT|15|7|假冒为善的人哪！ 以赛亚 指着你们所预言的说得好：
MATT|15|8|‘这百姓用嘴唇尊敬我， 他们的心却远离我。
MATT|15|9|他们把人的规条当作教义教导人； 他们拜我也是枉然。’”
MATT|15|10|耶稣叫了众人来，对他们说：“你们要听，也要明白。
MATT|15|11|从口里进去的不玷污人，从口里出来的才玷污人。”
MATT|15|12|当时，门徒进前来对他说：“法利赛人听见这话很反感，你知道吗？”
MATT|15|13|耶稣回答：“一切植物，若不是我天父栽植的，都要连根拔出来。
MATT|15|14|由他们吧！他们是瞎子作瞎子的向导 ；若是瞎子领瞎子，两个人都要掉在坑里。”
MATT|15|15|彼得 回应他说：“请将这比喻讲解给我们听。”
MATT|15|16|耶稣说：“连你们也还不明白吗？
MATT|15|17|难道你们不了解，凡进到口里的，是经过肚子，又排入厕所吗？
MATT|15|18|然而口里出来的是出于心里，这才玷污人。
MATT|15|19|因为出于心里的有种种恶念，如凶杀、奸淫、淫乱、偷盗、伪证、毁谤。
MATT|15|20|这些才玷污人。至于不洗手吃饭，那并不玷污人。”
MATT|15|21|耶稣离开那里，退到 推罗 、 西顿 境内。
MATT|15|22|有一个 迦南 妇人从那地方出来，喊着说：“主啊， 大卫 之子，可怜我！我女儿被鬼缠得很苦。”
MATT|15|23|耶稣却一言不答。门徒进前来，求他说：“这妇人在我们后头喊叫，请打发她走吧。”
MATT|15|24|耶稣回答：“我奉差遣只到 以色列 家迷失的羊那里去。”
MATT|15|25|那妇人来拜他，说：“主啊，帮帮我！”
MATT|15|26|他回答：“拿孩子的饼丢给小狗吃是不妥的。”
MATT|15|27|妇人说：“主啊，不错，可是小狗也吃它主人桌上掉下来的碎屑。”
MATT|15|28|于是耶稣回答她说：“妇人，你的信心很大！照你所要的成全你吧。”从那时起，她的女儿就好了。
MATT|15|29|耶稣离开那地方，来到靠近 加利利 的海边，就上山坐下。
MATT|15|30|有一大群人到他那里，带着瘸子、盲人、肢残的、聋哑的，和好些别的病人，都放在他脚前，他就治好了他们。
MATT|15|31|于是众人都惊讶，因为看见聋哑的说话，肢残的痊愈，瘸子行走，盲人看见，他们就归荣耀给 以色列 的上帝。
MATT|15|32|耶稣叫门徒来，说：“我怜悯这群人，因为他们同我在这里已经三天，没有吃的东西了。我不愿意叫他们饿着回去，恐怕他们在路上饿昏了。”
MATT|15|33|门徒说：“我们在这野地，哪里有这么多的饼让这许多人吃饱呢？”
MATT|15|34|耶稣对他们说：“你们有多少饼？”他们说：“有七个，还有几条小鱼。”
MATT|15|35|他就吩咐众人坐在地上，
MATT|15|36|拿着这七个饼和几条鱼，祝谢了，擘开，递给门徒；门徒又递给众人。
MATT|15|37|他们都吃，并且吃饱了，收拾剩下的碎屑，装满了七个筐子。
MATT|15|38|吃的人中，男的有四千，还不算妇女和孩子。
MATT|15|39|耶稣叫众人散去，就上船，来到 马加丹 境内。
MATT|16|1|法利赛人和撒都该人来试探耶稣，请他显个来自天上的神迹给他们看。
MATT|16|2|耶稣回答他们：“傍晚天发红，你们就说：‘明日天晴。’
MATT|16|3|早晨天色又红又暗，你们就说：‘今日有风雨。’你们知道分辨天上的气象，倒不能分辨这个时代的神迹 。
MATT|16|4|邪恶淫乱的世代求看神迹，除了 约拿 的神迹以外，再没有神迹给他们看了。”于是耶稣离开他们走了。
MATT|16|5|门徒渡到对岸，忘了带饼。
MATT|16|6|耶稣对他们说：“你们要谨慎，要防备法利赛人和撒都该人的酵。”
MATT|16|7|门徒彼此议论说：“这是因为我们没有带饼吧。”
MATT|16|8|耶稣知道了，就说：“你们这小信的人，为什么因为没有饼就彼此议论呢？
MATT|16|9|你们还不明白吗？不记得那五个饼分给五千人，你们收拾了多少篮子的碎屑吗？
MATT|16|10|也不记得那七个饼分给四千人，你们又收拾了多少筐子的碎屑吗？
MATT|16|11|我对你们说‘要防备法利赛人和撒都该人的酵’，这话不是指着饼说的，你们怎么不明白呢？”
MATT|16|12|门徒这才明白他所说的不是要他们防备饼的酵 ，而是要防备法利赛人和撒都该人的教训。
MATT|16|13|耶稣到了 凯撒利亚．腓立比 的境内，就问门徒：“人们说人子是谁？”
MATT|16|14|他们说：“有人说是施洗的 约翰 ；有人说是 以利亚 ；又有人说是 耶利米 或是先知中的一位。”
MATT|16|15|耶稣问他们：“你们说我是谁？”
MATT|16|16|西门．彼得 回答说：“你是基督，是永生上帝的儿子。”
MATT|16|17|耶稣回答他说：“ 约拿 的儿子 西门 ，你是有福的！因为这不是属血肉的启示你的，而是我在天上的父启示的。
MATT|16|18|我还告诉你，你是 彼得 ，我要把我的教会建造在这磐石上，阴间的权柄不能胜过它。
MATT|16|19|我要把天国的钥匙给你，凡你在地上所捆绑的，在天上也要捆绑；凡你在地上所释放的，在天上也要释放。”
MATT|16|20|当时，耶稣嘱咐门徒不可对任何人说他是基督。
MATT|16|21|从那时起，耶稣才向门徒明说，他必须上 耶路撒冷 去，受长老、祭司长和文士许多的苦，并且被杀，第三天复活。
MATT|16|22|彼得 就拉着他，责备他说：“主啊，千万不可如此！这事绝不可临到你身上。”
MATT|16|23|耶稣转过来，对 彼得 说：“撒但，退到我后边去！你是我的绊脚石，因为你不体会上帝的心意，而是体会人的意思。”
MATT|16|24|于是耶稣对门徒说：“若有人要跟从我，就当舍己，背起自己的十字架来跟从我。
MATT|16|25|因为凡要救自己生命的，要丧失生命；凡为我丧失生命的，要得着生命。
MATT|16|26|人若赚得全世界，赔上自己的生命，有什么益处呢？人还能拿什么换生命呢？
MATT|16|27|人子要在他父的荣耀里与他的众使者一起来临，那时候，他要照各人的行为报应各人。
MATT|16|28|我实在告诉你们，站在这里的，有人在没经历死亡以前，必定看见人子来到他的国里。”
MATT|17|1|过了六天，耶稣带着 彼得 、 雅各 和 雅各 的弟弟 约翰 ，领他们悄悄地上了高山。
MATT|17|2|他在他们面前变了形像，他的脸明亮如太阳，衣裳洁白如光。
MATT|17|3|忽然，有 摩西 和 以利亚 向他们显现，与耶稣说话。
MATT|17|4|彼得 回应，对耶稣说：“主啊，我们在这里真好！你若愿意，我就在这里搭三座棚，一座为你，一座为 摩西 ，一座为 以利亚 。”
MATT|17|5|说话之间，忽然有一朵明亮的云彩遮盖他们，又有声音从云彩里出来，说：“这是我的爱子，我所喜爱的。你们要听从他！”
MATT|17|6|门徒听见，就俯伏在地，极其害怕。
MATT|17|7|耶稣进前来，拍拍他们，说：“起来，不要害怕！”
MATT|17|8|他们举目，不见一人，只见耶稣独自一人。
MATT|17|9|下山的时候，耶稣嘱咐他们说：“人子还没有从死人中复活，你们不要把所看到的告诉人。”
MATT|17|10|门徒问耶稣：“那么，文士为什么说 以利亚 必须先来？”
MATT|17|11|耶稣回答：“ 以利亚 的确要来，并要复兴万事；
MATT|17|12|可是我告诉你们， 以利亚 已经来了，人不认识他，反倒任意待他。人子也将这样受他们的苦。”
MATT|17|13|门徒这才明白耶稣所说的是指施洗的 约翰 。
MATT|17|14|耶稣和门徒到了众人那里，有一个人来见耶稣，跪下，
MATT|17|15|说：“主啊，可怜我的儿子。他害癫痫病很苦，屡次跌进火里，屡次跌进水里。
MATT|17|16|我带他到你门徒那里，他们却不能医治他。”
MATT|17|17|耶稣回答：“唉！这又不信又悖谬的世代啊，我和你们在一起要到几时呢？我忍耐你们要到几时呢？把他带到我这里来！”
MATT|17|18|耶稣斥责那鬼，鬼就出来；从那时起，孩子就痊愈了。
MATT|17|19|门徒私下进前来问耶稣：“我们为什么不能赶出那鬼呢？”
MATT|17|20|耶稣对他们说：“是因你们的信心小。我实在告诉你们，你们若有信心像一粒芥菜种，就是对这座山说：‘你从这边移到那边’，它也会移过去，并且你们没有一件不能做的事了。 ”
MATT|17|21|
MATT|17|22|他们聚集在 加利利 的时候，耶稣对门徒说：“人子将要被交在人手里。
MATT|17|23|他们要杀害他，第三天他要复活。”门徒就非常忧愁。
MATT|17|24|他们到了 迦百农 ，收圣殿税 的人来见 彼得 ，说：“你们的老师不纳圣殿税吗？”
MATT|17|25|彼得 说：“纳。”他进了屋子，耶稣先对他说：“ 西门 ，你的意见如何？世上的君王向谁征收关税或丁税？是向自己的儿子呢？还是向外人呢？”
MATT|17|26|彼得 说：“是向外人。”耶稣对他说：“既然如此，儿子就可以免了。
MATT|17|27|但恐怕触犯他们，你往海边去钓鱼，把先钓上来的鱼拿起来，开了它的口，会发现一个司塔特 ，可以拿去给他们，作你我的税钱。”
MATT|18|1|当时，门徒前来问耶稣：“天国里谁是最大的？”
MATT|18|2|耶稣叫一个小孩子来，让他站在他们当中，
MATT|18|3|说：“我实在告诉你们，你们若不回转，变成像小孩子一样，绝不能进天国。
MATT|18|4|所以，凡自己谦卑像这小孩子的，他在天国里就是最大的。
MATT|18|5|凡为我的名接纳一个像这小孩子的，就是接纳我。”
MATT|18|6|“凡使这些信我的小子中的一个跌倒的，倒不如把大磨石拴在这人的颈项上，沉在深海里。
MATT|18|7|这世界有祸了，因为它使人跌倒；绊倒人的事是免不了的，但那绊倒人的有祸了！
MATT|18|8|如果你一只手或是一只脚使你跌倒，就把它砍下来扔掉。你缺一只手或是一只脚进入永生，比有两手两脚被扔进永火里还好。
MATT|18|9|如果你一只眼使你跌倒，就把它挖出来扔掉。你只有一只眼进入永生，比有两只眼被扔进地狱的火里还好。”
MATT|18|10|“你们要小心，不可轻看这些小子中的一个；我告诉你们，他们的天使在天上，常见我天父的面。
MATT|18|11|
MATT|18|12|“一个人若有一百只羊，其中一只走迷了路，你们的意见如何？他岂不留下这九十九只在山上，去找那只迷路的羊吗？
MATT|18|13|若是找到了，我实在告诉你们，他为这一只羊欢喜，比为那没有迷路的九十九只欢喜还大呢！
MATT|18|14|你们 在天上的父也是这样，不愿意失去这些小子中的一个。”
MATT|18|15|“若是你的弟兄得罪你 ，你要去，趁着只有他和你在一起的时候，指出他的错来。他若听你，你就赢得了你的弟兄；
MATT|18|16|他若不听，你就另外带一个或两个人同去，因为‘任何指控都要凭两个或三个证人的口述才能成立’。
MATT|18|17|他若是不听他们，就去告诉教会；若是不听教会，就把他看作外邦人和税吏。
MATT|18|18|“我实在告诉你们，凡你们在地上所捆绑的，在天上也要捆绑；凡你们在地上所释放的，在天上也要释放。
MATT|18|19|我又实在 告诉你们，若是你们中间有两个人在地上同心合意地求什么事，我在天上的父必为他们成全。
MATT|18|20|因为，哪里有两三个人奉我的名聚会，哪里就有我在他们中间。”
MATT|18|21|那时， 彼得 进前来，对耶稣说：“主啊，我弟兄得罪我，我当饶恕他几次呢？到七次够吗？”
MATT|18|22|耶稣说：“我告诉你，不是到七次，而是到七十个七次。
MATT|18|23|因为天国好像一个王要和他仆人算账。
MATT|18|24|他开始算的时候，有人带了一个欠一万他连得的仆人来。
MATT|18|25|因为他没有什么偿还之物，主人下令把他和他妻子儿女，以及一切所有的都卖了来偿还。
MATT|18|26|那仆人就俯伏向他叩头，说：‘宽容我吧，我都会还你的。’
MATT|18|27|那仆人的主人就动了慈心，把他释放了，并且免了他的债。
MATT|18|28|那仆人出来，遇见一个欠他一百个银币的同伴，就揪着他，扼住他的喉咙，说：‘把你所欠的还我！’
MATT|18|29|他的同伴就俯伏央求他，说：‘宽容我吧，我会还你的。’
MATT|18|30|他不肯，却把他下在监里，直到他还了所欠的债。
MATT|18|31|同伴们看见他所做的事就很悲愤，把这一切的事都告诉了主人。
MATT|18|32|于是主人叫了他来，对他说：‘你这恶奴才！你央求我，我就把你所欠的都免了；
MATT|18|33|你不应该怜悯你的同伴，像我怜悯你吗？’
MATT|18|34|主人就大怒，把他交给司刑的，直到他还清了所欠的债。
MATT|18|35|你们各人若不从心里饶恕你的弟兄，我天父也要这样待你们。”
MATT|19|1|耶稣说完了这些话，就离开 加利利 ，来到 犹太 的境内、 约旦河 的东边。
MATT|19|2|有一大群人跟着他，他就在那里治好了他们。
MATT|19|3|有些法利赛人来试探耶稣说：“无论什么缘故，人休妻都合法吗？”
MATT|19|4|耶稣回答：“那起初造人的，是造男造女，并且说：‘因此，人要离开父母，与妻子结合，二人成为一体。’这经文你们没有念过吗？
MATT|19|5|
MATT|19|6|既然如此，夫妻不再是两个人，而是一体的了。所以，上帝配合的，人不可分开。”
MATT|19|7|法利赛人说：“这样， 摩西 为什么吩咐给妻子休书就可以休她呢？”
MATT|19|8|耶稣说：“ 摩西 因为你们的心硬，所以准许你们休妻，但起初并不是这样。
MATT|19|9|我告诉你们，凡休妻另娶的，若不是为不贞的缘故，就是犯奸淫了。 ”
MATT|19|10|门徒对耶稣说：“丈夫和妻子的关系既是这样，倒不如不娶。”
MATT|19|11|耶稣对他们说：“这话不是人人都能领受的，惟独赐给谁，谁才能领受。
MATT|19|12|因为有人从母腹里就是不宜结婚的，也有因人为的缘故不宜结婚的，并有为天国的缘故自己不结婚的 。这话谁能领受，就领受吧。”
MATT|19|13|那时，有人带着小孩子来见耶稣，要他给他们按手祷告，门徒就责备那些人。
MATT|19|14|耶稣说：“让小孩子到我这里来，不要阻止他们，因为在天国的正是这样的人。”
MATT|19|15|耶稣给他们按手，然后离开那地方。
MATT|19|16|有一个人进前来问耶稣：“老师，我该做什么善事才能得永生？”
MATT|19|17|耶稣对他说：“你为什么问我关于善的事呢？只有一位是善良的。你若要进入永生，就该遵守诫命。”
MATT|19|18|他说：“哪些诫命？”耶稣说：“就是不可杀人；不可奸淫；不可偷盗；不可作假见证；
MATT|19|19|当孝敬父母；又当爱邻 如己。”
MATT|19|20|那青年说：“这一切我都遵守了，还缺少什么呢？”
MATT|19|21|耶稣说：“你若愿意作完全人，去变卖你所拥有的，分给穷人，就必有财宝在天上；然后来跟从我。”
MATT|19|22|那青年听见这话，就忧忧愁愁地走了，因为他的产业很多。
MATT|19|23|耶稣对门徒说：“我实在告诉你们，财主进天国是难的。
MATT|19|24|我再告诉你们，骆驼穿过针眼比财主进上帝的国还容易呢！”
MATT|19|25|门徒听见这话，就非常惊奇，说：“这样，谁能得救呢？”
MATT|19|26|耶稣看着他们，说：“在人这是不能，在上帝凡事都能。”
MATT|19|27|于是 彼得 回应，对他说：“看哪，我们已经撇下一切跟从你了，我们会得到什么呢？”
MATT|19|28|耶稣对他们说：“我实在告诉你们，你们这些跟从我的人，到了万物更新、人子坐在他荣耀宝座上的时候，你们也要坐在十二个宝座上，审判 以色列 十二个支派。
MATT|19|29|凡为我的名撇下房屋，或是兄弟、姊妹、父亲、母亲、 儿女、田地的，将得着百倍，并且承受永生。
MATT|19|30|然而，有许多在前的，将要在后；在后的，将要在前。”
MATT|20|1|“因为天国好比一家的主人清早去雇人进他的葡萄园做工。
MATT|20|2|他和工人讲定一天一个银币 ，就打发他们进葡萄园去。
MATT|20|3|约在上午九点钟出去，看见市场上还有闲站的人，
MATT|20|4|就对那些人说：‘你们也进葡萄园去，我会给你们合理的工钱。’
MATT|20|5|他们也进去了。约在正午和下午三点钟又出去，他也是这么做。
MATT|20|6|约在下午五点钟出去，他看见还有人站在那里，就问他们：‘你们为什么整天在这里闲站呢？’
MATT|20|7|他们说：‘因为没有人雇我们。’他说：‘你们也进葡萄园去。’
MATT|20|8|到了晚上，园主对工头说：‘叫工人都来，给他们工钱，从后来的起，到先来的为止。’
MATT|20|9|约在下午五点钟雇的人来了，各人领了一个银币。
MATT|20|10|那些最先雇的来了，以为可以多领，谁知也是各领一个银币。
MATT|20|11|他们领了工钱，就埋怨那家的主人说：
MATT|20|12|‘我们整天劳苦受热，那些后来的只做了一小时，你竟待他们和我们一样吗？’
MATT|20|13|主人回答其中的一人说：‘朋友，我没亏待你，你与我讲定的不是一个银币吗？
MATT|20|14|拿你的钱走吧！我乐意给那后来的和给你的一样，
MATT|20|15|难道我的东西不可随我的意思用吗？因为我作好人，你就眼红了吗？’
MATT|20|16|这样，那在后的，将要在前；在前的，将要在后了。”
MATT|20|17|耶稣上 耶路撒冷 去的时候，在路上把十二个门徒带到一边，对他们说：
MATT|20|18|“看哪，我们上 耶路撒冷 去，人子将被交给祭司长和文士；他们要定他死罪，
MATT|20|19|把他交给外邦人戏弄，鞭打，钉在十字架上；第三天他要复活。”
MATT|20|20|那时， 西庇太 儿子的母亲和她两个儿子上前来，向耶稣叩头，求他一件事。
MATT|20|21|耶稣问她：“你要什么呢？”她对耶稣说：“在你的国里，请让我这两个儿子一个坐在你右边，一个坐在你左边。”
MATT|20|22|耶稣回答：“你们不知道所求的是什么。我将要喝的杯，你们能喝吗？”他们对他说：“我们能。”
MATT|20|23|耶稣说：“我所喝的杯，你们要喝。可是坐在我的左右，不是我可以赐的，而是我父为谁预备就赐给谁。”
MATT|20|24|其余十个门徒听见，就对他们兄弟二人很生气。
MATT|20|25|耶稣叫了他们来，说：“你们知道，外邦人有君王作主治理他们，有大臣操权管辖他们。
MATT|20|26|但是在你们中间，不可这样。你们中间谁愿为大，就要作你们的用人；
MATT|20|27|谁愿为首，就要作你们的仆人。
MATT|20|28|正如人子来，不是要受人的服事，乃是要服事人，并且要舍命，作多人的赎价。”
MATT|20|29|他们出 耶利哥 的时候，有一大群人跟随耶稣。
MATT|20|30|有两个盲人坐在路旁，听说是耶稣经过，就喊着说：“主啊 ， 大卫 之子，可怜我们吧！”
MATT|20|31|众人责备他们，不许他们作声，他们却越发喊着说：“主啊 ， 大卫 之子，可怜我们吧！”
MATT|20|32|耶稣就站住，叫他们来，说：“你们要我为你们做什么？”
MATT|20|33|他们说：“主啊，让我们的眼睛能看见。”
MATT|20|34|耶稣动了慈心，摸了他们的眼睛，他们立刻看得见，就跟从耶稣。
MATT|21|1|耶稣和门徒快到 耶路撒冷 ，进了 橄榄山 的 伯法其 时，打发两个门徒，
MATT|21|2|对他们说：“你们往对面村子里去，会立刻看见一匹驴拴在那里，还有驴驹同在一处，解开它们，牵到我这里来。
MATT|21|3|若有人对你们说什么，你们就说：‘主要用它们。’那人会立刻让你们牵来。”
MATT|21|4|这事发生是要应验先知所说的话：
MATT|21|5|“要对 锡安 的儿女 说： 看哪，你的王来到你这里， 谦和地骑着驴， 骑着小驴—驴的驹子。”
MATT|21|6|门徒就照耶稣所吩咐的去做，
MATT|21|7|牵了驴和驴驹来，把他们的衣服搭在上面，耶稣就骑上。
MATT|21|8|许许多多的人把自己的衣服铺在路上，还有人砍下树枝来铺在路上。
MATT|21|9|前呼后拥的人群喊着说： “和散那 归于 大卫 之子！ 奉主名来的是应当称颂的！ 至高无上的，和散那！”
MATT|21|10|耶稣进了 耶路撒冷 ，全城都惊动了，说：“这是谁？”
MATT|21|11|众人说：“这是从 加利利 的 拿撒勒 来的先知耶稣。”
MATT|21|12|耶稣进了圣殿 ，赶出圣殿里所有在做买卖的人，推倒兑换银钱之人的桌子和卖鸽子之人的凳子，
MATT|21|13|对他们说：“经上记着： ‘我的殿要称为祷告的殿， 你们倒使它成为贼窝了。’”
MATT|21|14|在圣殿里有盲人和瘸子到耶稣跟前，他就治好了他们。
MATT|21|15|祭司长和文士看见耶稣所行的奇事，又见小孩子在圣殿里喊着说：“和散那归于 大卫 之子！”就很生气，
MATT|21|16|对他说：“这些人所喊的，你听到了吗？”耶稣对他们说：“听到了。经上说：‘你藉孩童和吃奶的口发出完全的赞美’，你们没有念过吗？”
MATT|21|17|于是他离开他们，出城到 伯大尼 去，在那里过夜。
MATT|21|18|早晨回城的时候，他饿了，
MATT|21|19|看见路旁有一棵无花果树，就走到跟前，在树上找不到什么，只有叶子，就对树说：“从今以后，你永不结果子！”那无花果树立刻枯干了。
MATT|21|20|门徒看见了，惊讶地说：“无花果树怎么立刻枯干了呢？”
MATT|21|21|耶稣回答他们：“我实在告诉你们，你们若有信心，不疑惑，不但能行我对无花果树所行的事，就是对这座山说：‘离开此地，投在海里！’也会实现。
MATT|21|22|你们祷告，无论求什么，只要信，就必得着。”
MATT|21|23|耶稣进了圣殿，正教导人的时候，祭司长和百姓的长老来问他：“你仗着什么权柄做这些事？给你这权柄的是谁呢？”
MATT|21|24|耶稣回答他们说：“我也要问你们一句话，你们若告诉我，我就告诉你们我仗着什么权柄做这些事。
MATT|21|25|约翰 的洗礼是从哪里来的？是从天上来的，还是从人间来的呢？”他们彼此商议说：“我们若说‘从天上来的’，他会对我们说：‘这样，你们为什么不信他呢？’
MATT|21|26|若说‘从人间来的’，我们又怕众人，因为大家都认为 约翰 是先知。”
MATT|21|27|于是他们回答耶稣：“我们不知道。”耶稣也对他们说：“我也不告诉你们，我仗着什么权柄做这些事。”
MATT|21|28|“有一件事，你们的意见如何？一个人有两个儿子。他来对大儿子说：‘孩子，今天到葡萄园里做工去。’
MATT|21|29|他回答：‘我不去’，以后自己懊悔，就去了。
MATT|21|30|他来对小儿子也是这样说。他回答：‘父亲大人，我去’，却不去。
MATT|21|31|这两个儿子是哪一个照着父亲的意愿做了呢？”他们说：“大儿子。”耶稣说：“我实在告诉你们，税吏和娼妓倒比你们先进上帝的国。
MATT|21|32|因为 约翰 到你们这里来指引你们走义路，你们却不信他，税吏和娼妓倒信了他。你们看见了以后，还是不悔悟去信他。”
MATT|21|33|“你们再听一个比喻：有一个家的主人开垦了一个葡萄园，四周围上篱笆，里面挖了一个榨酒池，盖了一座守望楼，租给园户，就出外远行去了。
MATT|21|34|收果子的时候快到了，他打发仆人到园户那里去收果子。
MATT|21|35|园户拿住仆人，打了一个，杀了一个，用石头打死了一个。
MATT|21|36|主人又打发别的仆人去，比先前更多；园户还是照样对待他们。
MATT|21|37|最后他打发自己的儿子到他们那里去，说：‘他们会尊敬我的儿子。’
MATT|21|38|可是，园户看见他儿子，彼此说：‘这是承受产业的。来，我们杀了他，占他的产业！’
MATT|21|39|于是他们拿住他，把他扔出葡萄园外，杀了。
MATT|21|40|葡萄园的主人来的时候，要怎样处置那些园户呢？”
MATT|21|41|他们说：“要狠狠地除灭那些恶人，将葡萄园转租给那些按时候交果子的园户。”
MATT|21|42|耶稣对他们说： “‘匠人所丢弃的石头 已作了房角的头块石头。 这是主所做的， 在我们眼中看为奇妙。’ 这段经文你们从来没有念过吗？
MATT|21|43|所以我告诉你们，上帝的国必从你们夺去，赐给那能结果子的民。
MATT|21|44|谁跌在这石头上，一定会跌得粉碎；这石头掉在谁的身上，就要把谁压得稀烂。 ”
MATT|21|45|祭司长和法利赛人听见他的比喻，就看出他是指着他们说的。
MATT|21|46|他们想要捉拿他，但是惧怕众人，因为众人认为他是先知。
MATT|22|1|耶稣又用比喻对他们说：
MATT|22|2|“天国好比一个王为他儿子摆设娶亲的宴席。
MATT|22|3|他打发仆人去，请那些被邀的人来赴宴，他们却不肯来。
MATT|22|4|王又打发别的仆人，说：‘你们去告诉那被邀的人，我的宴席已经预备好了，牛和肥畜已经宰了，各样都齐备，请你们来赴宴。’
MATT|22|5|那些人不理就走了，一个到自己田里去，一个做买卖去。
MATT|22|6|其余的抓住仆人，凌辱他们，把他们杀了。
MATT|22|7|王就大怒，发兵除灭那些凶手，烧毁他们的城。
MATT|22|8|于是王对仆人说：‘喜宴已经齐备，只是所邀的人不配。
MATT|22|9|所以你们要往岔路口上去，凡遇见的，都邀来赴宴。’
MATT|22|10|那些仆人就出去，到大路上，凡遇见的，不论善恶都招聚了来，宴席上就坐满了客人。
MATT|22|11|王进来见宾客，看到那里有一个没有穿礼服的，
MATT|22|12|就对他说：‘朋友，你到这里来怎么不穿礼服呢？’那人无言可答。
MATT|22|13|于是王对侍从说：‘捆起他的手脚，把他扔在外边的黑暗里；在那里他要哀哭切齿了。’
MATT|22|14|因为被召的人多，选上的人少。”
MATT|22|15|于是，法利赛人出去商议，怎样找话柄来陷害耶稣，
MATT|22|16|就打发他们的门徒同 希律 党人去见耶稣，说：“老师，我们知道你是诚实的，并且诚诚实实传上帝的道，无论谁你都一视同仁，因为你不看人的面子。
MATT|22|17|请告诉我们，你的意见如何？纳税给凯撒合不合法？”
MATT|22|18|耶稣看出他们的恶意，就说：“假冒为善的人哪，为什么试探我？
MATT|22|19|拿一个纳税的钱给我看！”他们就拿一个银币来给他。
MATT|22|20|耶稣问他们：“这像和这名号是谁的？”
MATT|22|21|他们说：“是凯撒的。”于是耶稣说：“这样，凯撒的归凯撒；上帝的归上帝。”
MATT|22|22|他们听了十分惊讶，就离开他走了。
MATT|22|23|那天，撒都该人来见耶稣。他们说没有复活这回事，于是问耶稣：
MATT|22|24|“老师， 摩西 说：‘某人若死了，没有孩子，他弟弟该娶他的妻子，为哥哥生子立后。’
MATT|22|25|从前，在我们这里有兄弟七人，第一个娶了妻，死了，没有孩子，撇下妻子给弟弟。
MATT|22|26|第二、第三，直到第七个，都是如此。
MATT|22|27|后来，那妇人也死了。
MATT|22|28|那么，在复活的时候，她是七个人中哪一个的妻子呢？因为他们都娶过她。”
MATT|22|29|耶稣回答他们说：“你们错了，因为不明白圣经，也不知道上帝的大能。
MATT|22|30|在复活的时候，人也不娶也不嫁，而是像天上的天使一样。
MATT|22|31|论到死人复活，上帝向你们所说的话，你们没有念过吗？
MATT|22|32|他说：‘我是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。’上帝不是死人的上帝，而是活人的上帝。”
MATT|22|33|众人听见这话，对他的教导非常惊讶。
MATT|22|34|法利赛人听见耶稣堵住了撒都该人的口，他们就聚集在一起。
MATT|22|35|其中有一个人是律法师 ，要试探耶稣，就问他：
MATT|22|36|“老师，律法上的诫命哪一条是最大的呢？”
MATT|22|37|耶稣对他说：“你要尽心、尽性、尽意爱主—你的上帝。
MATT|22|38|这是最大的，且是第一条诫命。
MATT|22|39|第二条也如此，就是要爱邻 如己。
MATT|22|40|这两条诫命是一切律法和先知书的总纲。”
MATT|22|41|法利赛人聚集的时候，耶稣问他们：
MATT|22|42|“论到基督，你们的意见如何？他是谁的后裔呢？”他们说：“是 大卫 的。”
MATT|22|43|耶稣说：“这样， 大卫 被圣灵感动，怎么还称他为主，说：
MATT|22|44|‘主对我主说： 你坐在我的右边， 等我把你的仇敌放在你脚下？’
MATT|22|45|大卫 既称他为主，他怎么又是 大卫 的后裔呢？”
MATT|22|46|没有一个人能回答一句话，从那日以后没有人敢再问他什么。
MATT|23|1|那时，耶稣对众人和门徒讲论，
MATT|23|2|说：“文士和法利赛人坐在 摩西 的位上，
MATT|23|3|所以凡他们所吩咐你们的，你们都要谨守遵行。但不要效法他们的行为，因为他们能说不能行。
MATT|23|4|他们把难挑的 重担捆起来，搁在人的肩上，但自己一个指头也不肯动。
MATT|23|5|他们所做的一切事都是要让人看见，所以把佩戴的经匣 加宽了，衣裳的繸子加长了，
MATT|23|6|喜爱宴席上的首座、会堂里的高位，
MATT|23|7|又喜欢人们在街市上向他们问安，称呼他们拉比 。
MATT|23|8|但你们不要接受拉比的称呼，因为只有一位是你们的老师；你们都是弟兄。
MATT|23|9|也不要称呼地上的人为父，因为只有一位是你们的父，就是在天上的父。
MATT|23|10|不要接受师傅的称呼，因为只有一位是你们的师傅，就是基督。
MATT|23|11|你们中间谁为大，谁就要作你们的用人。
MATT|23|12|凡自高的，必降为卑；自甘卑微的，必升为高。
MATT|23|13|“你们这假冒为善的文士和法利赛人有祸了！因为你们当着人的面把天国的门关了，自己不进去，要进去的人，你们也不容他们进去。
MATT|23|14|
MATT|23|15|“你们这假冒为善的文士和法利赛人有祸了！因为你们走遍海洋陆地，说服一个人入教，既入了教，却使他成为比你们加倍坏的地狱之子。
MATT|23|16|“你们这瞎眼的向导有祸了！你们说：‘凡指着圣所起誓的算不得什么；但是凡指着圣所中的金子起誓的，他就该谨守。’
MATT|23|17|你们这无知的瞎子啊，哪个更大呢？是金子，还是使金子成圣的圣所呢？
MATT|23|18|你们又说：‘凡指着祭坛起誓的算不得什么；但是凡指着坛上祭物起誓的，他就该谨守。’
MATT|23|19|你们这些瞎子啊，哪个更大呢？是祭物，还是使祭物成圣的坛呢？
MATT|23|20|所以，人指着祭坛起誓，就是指着坛和坛上一切所有的起誓；
MATT|23|21|人指着圣所起誓，就是指着圣所和那住在圣所里的起誓；
MATT|23|22|人指着天起誓，就是指着上帝的宝座和那坐在上面的起誓。
MATT|23|23|“你们这假冒为善的文士和法利赛人有祸了！因为你们将薄荷、大茴香、小茴香献上十分之一，那律法上更重要的事，就是公义、怜悯、信实，你们反倒不做；这原是你们该做的－至于那些奉献也不可废弃。
MATT|23|24|你们这瞎眼的向导，蠓虫你们就滤出来，骆驼你们倒吞下去。
MATT|23|25|“你们这假冒为善的文士和法利赛人有祸了！因为你们洗净杯盘的外面，里面却满了贪婪和放荡。
MATT|23|26|你这瞎眼的法利赛人，先洗净杯子 的里面，好使外面也干净了。
MATT|23|27|“你们这假冒为善的文士和法利赛人有祸了！因为你们好像粉饰了的坟墓，外面好看，里面却满了死人的骨头和一切的污秽。
MATT|23|28|你们也是如此，外面对人显出公义，里面却满了虚伪和不法的事。
MATT|23|29|“你们这假冒为善的文士和法利赛人有祸了！因为你们建造先知的坟，装修义人的墓，
MATT|23|30|说：‘若是我们在先祖的时代，必不和他们一同流先知的血。’
MATT|23|31|这样，你们就证明自己是杀害先知的人的子孙了。
MATT|23|32|你们去充满你们祖宗的恶贯吧！
MATT|23|33|你们这些蛇啊，毒蛇的孽种啊，怎能逃脱地狱的惩罚呢？
MATT|23|34|所以，我差遣先知、智慧人和文士到你们这里来，有的你们要杀害，要钉十字架；有的你们要在会堂里鞭打，从这城追逼到那城，
MATT|23|35|如此，地上所有义人流的血都归到你们身上，从义人 亚伯 的血起，直到你们在圣所和祭坛中间所杀的 巴拉加 的儿子 撒迦利亚 的血为止。
MATT|23|36|我实在告诉你们，这一切的罪都要归到这世代了。”
MATT|23|37|“ 耶路撒冷 啊， 耶路撒冷 啊，你常杀害先知，又用石头打死那奉差遣到你这里来的人。我多少次想聚集你的儿女，好像母鸡把小鸡聚集在翅膀底下，但是你们不愿意。
MATT|23|38|看吧，你们的家要被废弃成为荒芜。
MATT|23|39|我告诉你们，从今以后，你们绝不会再见到我，直到你们说：‘奉主名来的是应当称颂的！’”
MATT|24|1|耶稣出了圣殿，正离开的时候，门徒前来，把圣殿的建筑指给他看。
MATT|24|2|耶稣回应他们说：“你们不是看见这一切吗？我实在告诉你们，这里将没有一块石头会留在另一块石头上，而不被拆毁的。”
MATT|24|3|耶稣在 橄榄山 上坐着，门徒私下进前来问他：“请告诉我们，什么时候有这些事呢？你来临和世代的终结有什么预兆呢？”
MATT|24|4|耶稣回答他们：“你们要谨慎，免得有人迷惑你们。
MATT|24|5|因为将有好些人冒我的名来，说‘我是基督’，并且要迷惑许多人。
MATT|24|6|你们也将听见打仗和打仗的风声。注意，不要惊慌！因为这些事必须发生，但这还不是终结。
MATT|24|7|民要攻打民，国要攻打国，多处必有饥荒、地震。
MATT|24|8|这都是灾难 的起头。
MATT|24|9|那时，人要使你们陷在患难里，也要杀害你们；你们又要为我的名被万民憎恨。
MATT|24|10|那时，会有许多人跌倒，也会彼此陷害，彼此憎恨；
MATT|24|11|且有好些假先知起来，迷惑许多人。
MATT|24|12|因为不法的事增多，许多人的爱心渐渐冷淡了。
MATT|24|13|但坚忍到底的终必得救。
MATT|24|14|这天国的福音要传遍天下，对万民作见证，然后终结才来到。”
MATT|24|15|“当你们看见先知 但以理 所说的那‘施行毁灭的亵渎者’站在圣地（读这经的人要会意），
MATT|24|16|那时，在 犹太 的，应当逃到山上；
MATT|24|17|在屋顶上的，不要下来拿家里的东西；
MATT|24|18|在田里的，不要回去取衣裳。
MATT|24|19|在那些日子，怀孕的和奶孩子的就苦了。
MATT|24|20|你们要祈求，好让你们逃走的时候，不遇见冬天或安息日。
MATT|24|21|因为那时必有大灾难，自从世界的起头直到如今，从没有这样的灾难，将来也不会有。
MATT|24|22|若不减少那些日子，凡血肉之躯的，就没有一个能得救；可是为了选民，那些日子将减少。
MATT|24|23|那时，若有人对你们说：‘看哪，基督在这里！’或‘在那里！’你们不要信。
MATT|24|24|因为假基督和假先知将要起来，显大神迹、大奇事，如果可能，要把选民也迷惑了。
MATT|24|25|看哪，我已经预先告诉你们了。
MATT|24|26|若有人对你们说：‘看哪，基督在旷野里！’你们不要出去；或说：‘看哪，基督在内室中！’你们不要信。
MATT|24|27|好像闪电从东边发出，直照到西边，人子来临也要这样。
MATT|24|28|尸首在哪里，鹰也会聚在哪里。”
MATT|24|29|“那些日子的灾难一过去， 太阳要变黑， 月亮也不放光， 众星要从天上坠落， 天上的万象都要震动。
MATT|24|30|那时，人子的预兆要显在天上，地上的万族都要哀哭。他们要看见人子带着能力和大荣耀，驾着天上的云来临。
MATT|24|31|他要差遣天使，用大声的号筒，从四方，从天这边直到天那边，召集他的选民。”
MATT|24|32|“你们要从无花果树学习功课：当树枝发芽长叶的时候，你们就知道夏天近了。
MATT|24|33|同样，当你们看见这一切，就知道那时候近了，就在门口了。
MATT|24|34|我实在告诉你们，这世代还没有过去，这一切都要发生。
MATT|24|35|天地要废去，我的话却绝不废去。”
MATT|24|36|“但那日子，那时辰，没有人知道，连天上的天使也不知道，子也不知道，惟有父知道。
MATT|24|37|挪亚 的日子怎样，人子来临也要怎样。
MATT|24|38|在洪水以前的那些日子，人照常吃喝嫁娶，直到 挪亚 进方舟的那日，
MATT|24|39|不知不觉洪水来了，把他们全都冲去。人子来临也要这样。
MATT|24|40|那时，两个人在田里，一个被接去，一个被撇下。
MATT|24|41|两个女人推磨，一个被接去，一个被撇下。
MATT|24|42|所以，你们要警醒，因为不知道你们的主哪一天来到。
MATT|24|43|你们要知道，一家的主人若知道晚上什么时候有贼来，就必警醒，不让贼挖穿房屋。
MATT|24|44|所以，你们也要预备，因为在你们想不到的时候，人子就来了。”
MATT|24|45|“那么，谁是那忠心又精明的仆人，主人派他管理自己的家仆、按时分粮给他们的呢？
MATT|24|46|主人来到，看见仆人这样做，那仆人就有福了。
MATT|24|47|我实在告诉你们，主人要派他管理所有的财产。
MATT|24|48|如果那恶仆心里说：‘我的主人会来得迟’，
MATT|24|49|就动手打他的同伴，又和醉酒的人一同吃喝，
MATT|24|50|在想不到的日子，不知道的时候，那仆人的主人要来，
MATT|24|51|重重地惩罚他 ，定他和假冒为善的人同罪，在那里他要哀哭切齿了。”
MATT|25|1|“那时，天国好比十个童女拿着灯出去迎接新郎。
MATT|25|2|其中有五个是愚拙的，五个是聪明的。
MATT|25|3|愚拙的拿着灯，却没有带油；
MATT|25|4|聪明的拿着灯，又盛了油在器皿里。
MATT|25|5|新郎迟延的时候，她们都打盹，睡着了。
MATT|25|6|半夜有人喊：‘看，新郎来了，你们出来迎接他。’
MATT|25|7|那些童女就都起来挑亮她们的灯。
MATT|25|8|愚拙的对聪明的说：‘请分点油给我们，因为我们的灯要灭了。’
MATT|25|9|聪明的回答：‘恐怕不够你我用的；你们还是自己到卖油的那里去买吧。’
MATT|25|10|她们去买的时候，新郎到了。那预备好了的，与他进去共赴婚宴，门就关了。
MATT|25|11|其余的童女随后也来了，说：‘主啊，主啊，给我们开门！’
MATT|25|12|他却回答：‘我实在告诉你们，我不认识你们。’
MATT|25|13|所以，你们要警醒，因为那日子，那时辰，你们不知道。”
MATT|25|14|“天国又好比一个人要出外远行，就叫了仆人来，把他的家业交给他们。
MATT|25|15|他按着各人的才干，给他们银子：一个给了五千 ，一个给了二千 ，一个给了一千 ，就出外远行去了。
MATT|25|16|那领五千的立刻拿去做买卖，另外赚了五千。
MATT|25|17|那领二千的也照样另赚了二千。
MATT|25|18|但那领一千的去掘开地，把主人的银子埋藏了。
MATT|25|19|过了许久，那些仆人的主人来了，和他们算账。
MATT|25|20|那领五千的又带着另外的五千来，说：‘主啊，你交给我五千。请看，我又赚了五千。’
MATT|25|21|主人说：‘好，你这又善良又忠心的仆人，你在少许的事上忠心，我要派你管理许多的事，进来享受你主人的快乐吧！’
MATT|25|22|那领二千的也进前来，说：‘主啊，你交给我二千。请看，我又赚了二千。’
MATT|25|23|主人说：‘好，你这又善良又忠心的仆人，你在少许的事上忠心，我要派你管理许多的事，进来享受你主人的快乐吧！’
MATT|25|24|那领一千的也进前来，说：‘主啊，我知道你，你是个严厉的人：没有种的地方也要收割，没有播的地方也要收获，
MATT|25|25|我就害怕，去把你的一千银子埋藏在地里。请看，你的银子在这里。’
MATT|25|26|他的主人回答他说：‘你这又恶又懒的仆人，你既知道我没有种的地方也要收割，没有播的地方也要收获，
MATT|25|27|就该把我的银子放给兑换银钱的人，到我来的时候可以连本带利收回。
MATT|25|28|把他这一千夺过来，给那有一万 的。
MATT|25|29|因为凡有的，还要加给他，叫他有余；没有的，连他所有的也要夺过来。
MATT|25|30|把这无用的仆人丢在外面黑暗里，在那里他要哀哭切齿了。’”
MATT|25|31|“当人子在他荣耀里，同着众天使来临的时候，要坐在他荣耀的宝座上。
MATT|25|32|万民都要聚集在他面前。他要把他们分别出来，好像牧人分别绵羊、山羊一般，
MATT|25|33|把绵羊安置在右边，山羊在左边。
MATT|25|34|于是王要向他右边的说：‘你们这蒙我父赐福的，可来承受那创世以来为你们所预备的国。
MATT|25|35|因为我饿了，你们给我吃；渴了，你们给我喝；我流浪在外，你们留我住；
MATT|25|36|我赤身露体，你们给我穿；我病了，你们看顾我；我在监狱里，你们来看我。’
MATT|25|37|义人就回答：‘主啊，我们什么时候见你饿了，给你吃；渴了，给你喝？
MATT|25|38|什么时候见你流浪在外，留你住；或是赤身露体，给你穿？
MATT|25|39|又什么时候见你病了，或是在监狱里，来看你呢？’
MATT|25|40|王回答他们说：‘我实在告诉你们，这些事你们做在我弟兄中一个最小的身上，就是做在我身上了。’
MATT|25|41|“王又要向那左边的说：‘你们这被诅咒的人，离开我！进入那为魔鬼和他的使者所预备的永火里去！
MATT|25|42|因为我饿了，你们没有给我吃；渴了，你们没有给我喝；
MATT|25|43|我流浪在外，你们没有留我住；我赤身露体，你们没有给我穿；我病了，我在监狱里，你们没有来看顾我。’
MATT|25|44|他们也要回答：‘主啊，我们什么时候见你饿了，或渴了，或流浪在外，或赤身露体，或病了，或在监狱里，没有伺候你呢？’
MATT|25|45|王要回答：‘我实在告诉你们，这些事你们没有做在任何一个最小的弟兄身上，就是没有做在我身上了。’
MATT|25|46|这些人要往永刑里去；那些义人要往永生里去。”
MATT|26|1|耶稣说完了这一切的话，就对门徒说：
MATT|26|2|“你们知道，过两天是逾越节，人子将要被出卖，钉在十字架上。”
MATT|26|3|那时，祭司长和百姓的长老聚集在那称为 该亚法 的大祭司的院里。
MATT|26|4|大家商议要设计捉拿耶稣，把他杀掉。
MATT|26|5|可是他们说：“不可在过节的日子，恐怕百姓生乱。”
MATT|26|6|耶稣在 伯大尼 的痲疯病人 西门 家里，
MATT|26|7|有一个女人拿着一玉瓶极贵的香膏来，趁耶稣坐席的时候，浇在他的头上。
MATT|26|8|门徒看见就很不高兴，说：“何必这样浪费呢！
MATT|26|9|这香膏可以卖许多钱，周济穷人。”
MATT|26|10|耶稣看出他们的意思，就说：“为什么难为这女人呢？她在我身上做的是一件美事。
MATT|26|11|因为常有穷人和你们在一起，但是你们不常有我。
MATT|26|12|她把这香膏浇在我身上是为我安葬作准备的。
MATT|26|13|我实在告诉你们，普天之下，无论在什么地方传这福音，都要述说这女人所做的，来记念她。”
MATT|26|14|当时，十二使徒中有一个叫 加略 人 犹大 的，去见祭司长，
MATT|26|15|说：“我把他交给你们，你们愿意给我多少钱？”他们给了他三十块银钱。
MATT|26|16|从那时候起，他就找机会要把耶稣交给他们。
MATT|26|17|除酵节的第一天，门徒来问耶稣：“你要我们在哪里给你预备吃逾越节的宴席呢？”
MATT|26|18|耶稣说：“你们进城去，到某人那里，对他说：‘老师说：我的时候快到了，我要和我的门徒在你家里守逾越节。’”
MATT|26|19|门徒遵照耶稣所吩咐的去预备了逾越节的宴席。
MATT|26|20|到了晚上，耶稣和十二使徒坐席。
MATT|26|21|他们吃的时候，耶稣说：“我实在告诉你们，你们中间有一个人要出卖我。”
MATT|26|22|他们就非常忧愁，一个一个地问他：“主，该不是我吧？”
MATT|26|23|耶稣回答说：“同我蘸手在盘子里的，就是要出卖我的。
MATT|26|24|人子要去了，正如经上所写有关他的；但出卖人子的人有祸了！那人没有出生倒好。”
MATT|26|25|出卖耶稣的 犹大 回答他说：“拉比，该不是我吧？”耶稣说：“你自己说了。”
MATT|26|26|他们吃的时候，耶稣拿起饼来，祝福了，就擘开，递给门徒，说：“你们拿去，吃吧。这是我的身体。”
MATT|26|27|他又拿起杯来，祝谢了，递给他们，说：“你们都喝这个，
MATT|26|28|因为这是我立约的血，为许多人流出来，使罪得赦。
MATT|26|29|但我告诉你们，从今以后，我不再喝这葡萄汁，直到我在我父的国里与你们同喝新的那日子。”
MATT|26|30|他们唱了诗，就出来往 橄榄山 去。
MATT|26|31|那时，耶稣对他们说：“今夜，你们为我的缘故都要跌倒。因为经上记着： ‘我要击打牧人， 羊就分散了。’
MATT|26|32|但我复活以后，要在你们之前往 加利利 去。”
MATT|26|33|彼得 回答他说：“即使众人为你的缘故跌倒，我也绝不跌倒。”
MATT|26|34|耶稣说：“我实在告诉你，今夜鸡叫以前，你要三次不认我。”
MATT|26|35|彼得 说：“我就是必须和你同死，也绝不会不认你。”所有的门徒都是这样说。
MATT|26|36|耶稣和门徒来到一个地方，名叫 客西马尼 。他对他们说：“你们坐在这里，我到那边去祷告。”
MATT|26|37|于是他带着 彼得 和 西庇太 的两个儿子同去。他忧愁起来，极其难过，
MATT|26|38|就对他们说：“我心里非常忧伤，几乎要死；你们留在这里，和我一同警醒。”
MATT|26|39|他就稍往前走，俯伏在地，祷告说：“我父啊，如果可能，求你使这杯离开我。然而，不是照我所愿的，而是照你所愿的。”
MATT|26|40|他回到门徒那里，见他们睡着了，就对 彼得 说：“怎么样？你们不能同我警醒一小时吗？
MATT|26|41|总要警醒祷告，免得陷入试探。你们心灵固然愿意，肉体却软弱了。”
MATT|26|42|他第二次又去祷告说：“我父啊，这杯若不能离开我，必须我喝，就愿你的旨意成全。”
MATT|26|43|他又来，见他们睡着了，因为他们的眼睛困倦。
MATT|26|44|耶稣又离开他们，第三次去祷告，说的话跟先前一样。
MATT|26|45|然后他来到门徒那里，对他们说：“现在你们仍在睡觉安歇吗？看哪，时候到了，人子被出卖在罪人手里了。
MATT|26|46|起来，我们走吧！看哪，那出卖我的人快来了。”
MATT|26|47|耶稣还在说话的时候，十二使徒之一的 犹大 来了，还有一大群人带着刀棒，从祭司长和百姓的长老那里跟他同来。
MATT|26|48|那出卖耶稣的给了他们一个暗号，说：“我亲谁，谁就是。你们把他抓住。”
MATT|26|49|犹大 立刻进前来对耶稣说：“拉比，你好！”就跟他亲吻。
MATT|26|50|耶稣对他说：“朋友，你来要做的事，就做吧。 ”于是那些人上前，下手抓住耶稣。
MATT|26|51|忽然，有一个和耶稣一起的人伸手拔出刀来，把大祭司的仆人砍了一刀，削掉了他一只耳朵。
MATT|26|52|耶稣对他说：“收刀入鞘吧！凡动刀的，必死在刀下。
MATT|26|53|你想我不能求我父，现在为我差遣比十二营还多的天使来吗？
MATT|26|54|若是这样，经上所说事情必须如此发生的话怎么应验呢？”
MATT|26|55|就在那时，耶稣对众人说：“你们带着刀棒出来抓我，如同拿强盗吗？我天天坐在圣殿里教导人，你们并没有抓我。
MATT|26|56|但这整件事的发生，是要应验先知书上的话。”那时，门徒都离开他，逃走了。
MATT|26|57|抓耶稣的人把他带到大祭司 该亚法 那里去，文士和长老已经在那里聚集。
MATT|26|58|彼得 远远地跟着耶稣，直到大祭司的院子，进到里面，就和警卫同坐，要看结局怎样。
MATT|26|59|祭司长和全议会寻找假见证控告耶稣，要处死他。
MATT|26|60|虽然有好些人来作假见证，总找不到实据。最后有两个人前来，
MATT|26|61|说：“这个人曾说：‘我能拆毁上帝的殿，三日内又建造起来。’”
MATT|26|62|大祭司就站起来，对耶稣说：“这些人作证告你的事，你什么都不回答吗？”
MATT|26|63|耶稣却不言语。大祭司对他说：“我指着永生上帝命令你起誓告诉我们，你是不是基督—上帝的儿子？”
MATT|26|64|耶稣对他说：“你自己说了。然而，我告诉你们， 此后你们要看见人子 坐在权能者的右边， 驾着天上的云来临。”
MATT|26|65|大祭司就撕裂衣服，说：“他说了亵渎的话，我们何必再要证人呢？现在你们已经听见他这亵渎的话了。
MATT|26|66|你们的意见如何？”他们回答：“他该处死。”
MATT|26|67|他们就吐唾沫在他脸上，用拳头打他，也有打他耳光的，
MATT|26|68|说：“基督啊，向我们说预言吧！打你的是谁？”
MATT|26|69|彼得 在外面院子里坐着，有一个使女进前来，说：“你素来也是同那 加利利 人耶稣一起的。”
MATT|26|70|彼得 在众人面前却不承认，说：“我不知道你说的是什么！”
MATT|26|71|他出去，到了门口，又有一个使女看见他，就对那里的人说：“这个人是同 拿撒勒 人耶稣一起的。”
MATT|26|72|彼得 又不承认，起誓说：“我不认得那个人。”
MATT|26|73|过了不久，旁边站着的人前来，对 彼得 说：“你的确是他们一伙的，你的口音把你显露出来了。”
MATT|26|74|彼得 就赌咒发誓说：“我不认得那个人。”立刻鸡就叫了。
MATT|26|75|彼得 想起耶稣所说的话：“鸡叫以前，你要三次不认我。”他就出去痛哭。
MATT|27|1|到了早晨，众祭司长和百姓的长老商议要处死耶稣，
MATT|27|2|就把他绑着，解去，交给 彼拉多 总督。
MATT|27|3|这时，出卖耶稣的 犹大 看见耶稣已经定了罪，就后悔，把那三十块银钱拿回来给祭司长和长老，
MATT|27|4|说：“我出卖了无辜人的血有罪了。”他们说：“那跟我们有什么相干？你自己承当吧！”
MATT|27|5|犹大 就把那银钱丢在殿里，出去吊死了。
MATT|27|6|祭司长拾起银钱来，说：“这是血价，不可放在圣殿的银库里。”
MATT|27|7|他们商议，就用那银钱买了窑户的一块田，用来埋葬外乡人。
MATT|27|8|所以，那块田直到今日还叫做“血田”。
MATT|27|9|这就应验了先知 耶利米 所说的话：“他们用那三十块银钱，就是 以色列 人给那被估定的人所估定的价钱，
MATT|27|10|买了窑户的一块田；这是照着主所吩咐我的。”
MATT|27|11|耶稣站在总督面前，总督问他：“你是 犹太 人的王吗？”耶稣说：“是你说的。”
MATT|27|12|他被祭司长和长老控告的时候，什么都不回答。
MATT|27|13|彼拉多 就对他说：“他们作证告你这么多的事，你没有听见吗？”
MATT|27|14|耶稣仍不回答，连一句话也不说，以致总督觉得非常惊讶。
MATT|27|15|总督有一个常例，每逢这节期，随众人的意愿释放一个囚犯给他们。
MATT|27|16|当时有一个出名的囚犯叫 巴拉巴 。
MATT|27|17|众人聚集的时候， 彼拉多 就对他们说：“你们要我释放哪一个给你们？是 巴拉巴 呢？是称为基督的耶稣呢？”
MATT|27|18|总督原知道他们是因为嫉妒才把他解了来。
MATT|27|19|正坐堂的时候，他的夫人打发人来说：“这义人的事，你一点不可管，因为我今天在梦中因他受了许多的苦。”
MATT|27|20|祭司长和长老挑唆众人，要求释放 巴拉巴 ，除掉耶稣。
MATT|27|21|总督回答他们说：“这两个人，你们要我释放哪一个给你们呢？”他们说：“ 巴拉巴 。”
MATT|27|22|彼拉多 说：“这样，那称为基督的耶稣我怎么办他呢？”他们都说：“把他钉十字架！”
MATT|27|23|总督说：“为什么？他做了什么恶事呢？”他们更加喊着说：“把他钉十字架！”
MATT|27|24|彼拉多 见说也无济于事，反要生乱，就拿水在众人面前洗手，说：“流这人 的血，罪不在我，你们承当吧。”
MATT|27|25|众人都回答：“他的血归到我们和我们的子孙身上！”
MATT|27|26|于是 彼拉多 释放 巴拉巴 给他们，把耶稣鞭打后交给人钉十字架。
MATT|27|27|总督的兵把耶稣带进总督府，把全营的兵都聚集在耶稣那里。
MATT|27|28|他们脱了他的衣服，穿上一件朱红色的袍子，
MATT|27|29|用荆棘编了冠冕，戴在他头上，拿一根芦苇秆放在他右手里，跪在他面前，戏弄他，说：“万岁， 犹太 人的王！”
MATT|27|30|他们又向他吐唾沫，拿芦苇秆打他的头。
MATT|27|31|他们戏弄完了，就给他脱了袍子，又穿上他自己的衣服，带他出去，要钉十字架。
MATT|27|32|他们出去的时候，遇见一个 古利奈 人，名叫 西门 ，就强迫他同去，好背耶稣的十字架。
MATT|27|33|他们到了一个地方，名叫 各各他 ，就是“髑髅地”。
MATT|27|34|士兵拿苦胆调和的酒给耶稣喝。他尝了，不肯喝。
MATT|27|35|他们把他钉在十字架上，然后抽签分了他的衣服，
MATT|27|36|又坐在那里看守他。
MATT|27|37|他们在他头上方安了一个罪状牌，写着：“这是 犹太 人的王耶稣。”
MATT|27|38|当时，有两个强盗和他同钉十字架，一个在右边，一个在左边。
MATT|27|39|从那里经过的人讥笑他，摇着头，
MATT|27|40|说：“你这拆毁殿、三日又建造起来的，救救你自己吧！如果你是上帝的儿子，就从十字架上下来呀！”
MATT|27|41|众祭司长、文士和长老也同样嘲笑他，说：
MATT|27|42|“他救了别人，不能救自己。他是 以色列 的王，现在从十字架上下来，我们就信他。
MATT|27|43|他倚靠上帝，上帝若愿意，现在就来救他，因为他曾说‘我是上帝的儿子’。”
MATT|27|44|和他同钉的强盗也这样讥讽他。
MATT|27|45|从正午到下午三点钟，遍地都黑暗了。
MATT|27|46|约在下午三点钟，耶稣大声高呼，说：“以利！以利！拉马撒巴各大尼？”就是说：“我的上帝！我的上帝！为什么离弃我？”
MATT|27|47|站在那里的人，有的听见就说：“这个人呼叫 以利亚 呢！”
MATT|27|48|其中有一个人立刻跑去，拿海绵蘸满了醋，绑在芦苇秆上，送给他喝。
MATT|27|49|其余的人说：“且等着，看 以利亚 来不来救他。”
MATT|27|50|耶稣又大喊一声，气就断了。
MATT|27|51|忽然，殿的幔子从上到下裂为两半，地震动，磐石崩裂，
MATT|27|52|坟墓也开了，有许多已睡了的圣徒的身体也复活了。
MATT|27|53|耶稣复活以后，他们从坟墓里出来，进了圣城，向许多人显现。
MATT|27|54|百夫长和跟他一同看守耶稣的人看见地震和所经历的事，非常害怕，说：“他真是上帝的儿子！”
MATT|27|55|有好些妇女在那里，远远地观看，她们是从 加利利 跟随耶稣，来服事他的；
MATT|27|56|其中有 抹大拉 的 马利亚 ，又有 雅各 和 约瑟 的母亲 马利亚 ，并有 西庇太 两个儿子的母亲。
MATT|27|57|到了晚上，有一个财主，名叫 约瑟 ，是 亚利马太 来的，他也是耶稣的门徒。
MATT|27|58|这人去见 彼拉多 ，请求要耶稣的身体， 彼拉多 就吩咐给他。
MATT|27|59|约瑟 取了身体，用干净的细麻布裹好，
MATT|27|60|然后把他安放在自己的新墓穴里，就是他凿在岩石里的。他又把大石头滚到墓门口，然后离开。
MATT|27|61|有 抹大拉 的 马利亚 和另一个 马利亚 在那里，对着坟墓坐着。
MATT|27|62|次日，就是预备日的第二天，祭司长和法利赛人聚集来见 彼拉多 ，
MATT|27|63|说：“大人，我们记得那迷惑人的还活着的时候曾说：‘三天后我要复活。’
MATT|27|64|因此，请吩咐人将坟墓把守妥当，直到第三天，恐怕他的门徒来把他偷了去，就告诉百姓说：‘他从死人中复活了。’这样的话，那后来的迷惑就比先前的更厉害了。”
MATT|27|65|彼拉多 说：“你们有看守的兵，去吧！尽你们所能的把守妥当。”
MATT|27|66|他们就带着看守的兵同去，封了石头，将坟墓把守妥当。
MATT|28|1|安息日过后，七日的第一日，天快亮的时候， 抹大拉 的 马利亚 和另一个 马利亚 来看坟墓。
MATT|28|2|忽然，地大震动；因为有主的一个使者从天上下来，把石头滚开，坐在上面。
MATT|28|3|他的相貌如同闪电，衣服洁白如雪。
MATT|28|4|看守的人吓得浑身颤抖，甚至和死人一样。
MATT|28|5|天使回应妇女说：“不要害怕！我知道你们是寻找那钉十字架的耶稣。
MATT|28|6|他不在这里，照他所说的，他已经复活了。你们来！看看安放他的地方。
MATT|28|7|快去告诉他的门徒，说他已从死人中复活了，并且要比你们先到 加利利 去，在那里你们会看见他。看哪！我已经告诉你们了。”
MATT|28|8|妇女们急忙离开坟墓，又害怕，又大为欢喜，跑去告诉他的门徒。
MATT|28|9|忽然，耶稣迎上她们，说：“平安！”她们就上前抱住他的脚拜他。
MATT|28|10|耶稣对她们说：“不要害怕！你们去告诉我的弟兄，叫他们往 加利利 去，在那里会见到我。”
MATT|28|11|她们去的时候，看守的兵有几个进城去，把所发生的事都报告祭司长。
MATT|28|12|祭司长和长老聚集商议，就拿许多银钱给士兵，
MATT|28|13|说：“你们要这样说：‘夜间我们睡觉的时候，他的门徒来把他偷去了。’
MATT|28|14|若是这话被总督听见，有我们劝他，保你们无事。”
MATT|28|15|士兵收了银钱，就照所嘱咐他们的去做。这话就在 犹太 人中间流传，直到今日。
MATT|28|16|十一个门徒往 加利利 去，到了耶稣指定他们去的山上。
MATT|28|17|他们见了耶稣就拜他，然而还有人疑惑。
MATT|28|18|耶稣进前来，对他们说：“天上地下所有的权柄都赐给我了。
MATT|28|19|所以，你们要去，使万民作我的门徒，奉父、子、圣灵的名给他们施洗 ，
MATT|28|20|凡我所吩咐你们的，都教导他们遵守。看哪，我天天与你们同在，直到世代的终结。”
MARK|1|1|上帝的儿子 ，耶稣基督福音的起头。
MARK|1|2|正如 以赛亚 先知书上记着： “看哪，我要差遣我的使者在你面前， 他要为你预备道路。
MARK|1|3|在旷野有声音呼喊着： 预备主的道， 修直他的路。”
MARK|1|4|照这话，施洗 约翰 来到旷野 ，宣讲悔改的洗礼，使罪得赦。
MARK|1|5|犹太 全地和全 耶路撒冷 的人都出去，到 约翰 那里，承认他们的罪，在 约旦河 里受他的洗。
MARK|1|6|约翰 穿骆驼毛的衣服，腰束皮带，吃的是蝗虫和野蜜。
MARK|1|7|他宣讲，说：“有一位在我以后来的，能力比我更大，我就是弯腰给他解鞋带也不配。
MARK|1|8|我用水给你们施洗，他却要用圣灵给你们施洗。”
MARK|1|9|那时，耶稣从 加利利 的 拿撒勒 来，在 约旦河 里受了 约翰 的洗。
MARK|1|10|他从水里一上来，就看见天裂开了，圣灵仿佛鸽子降在他身上。
MARK|1|11|又有声音从天上来，说：“你是我的爱子，我喜爱你。”
MARK|1|12|圣灵立刻把耶稣催促到旷野里去。
MARK|1|13|他在旷野四十天，受撒但的试探，并与野兽同在一起，且有天使来伺候他。
MARK|1|14|约翰 下监以后，耶稣来到 加利利 ，宣讲上帝的福音，
MARK|1|15|说：“日期满了，上帝的国近了。你们要悔改，信福音！”
MARK|1|16|耶稣沿着 加利利 的海边走，看见 西门 和 西门 的弟弟 安得烈 在海上撒网；他们本是打鱼的。
MARK|1|17|耶稣对他们说：“来跟从我，我要叫你们得人如得鱼一样。”
MARK|1|18|他们立刻舍了网，跟从他。
MARK|1|19|耶稣稍往前走，又见 西庇太 的儿子 雅各 和他弟弟 约翰 在船上补网。
MARK|1|20|耶稣随即呼召他们，他们就把父亲 西庇太 和雇工留在船上，跟从了耶稣。
MARK|1|21|他们到了 迦百农 ，耶稣就在安息日进了会堂教导人。
MARK|1|22|他们对他的教导感到很惊奇，因为他教导他们正像有权柄的人，不像文士。
MARK|1|23|当时，会堂里有一个污灵附身的人，他在喊叫，
MARK|1|24|说：“ 拿撒勒 人耶稣，你为什么干扰我们？你来消灭我们吗？我知道你是谁，你是上帝的圣者。”
MARK|1|25|耶稣斥责他说：“不要作声，从这人身上出来吧！”
MARK|1|26|污灵使那人抽了一阵风，大声喊叫，就出来了。
MARK|1|27|众人都惊讶，以致彼此对问：“这是什么事？是个新的教导啊！他用权柄命令污灵，连污灵也听从了他。”
MARK|1|28|于是耶稣的名声立刻传遍了全 加利利 周围地区。
MARK|1|29|他们一出会堂，就同 雅各 和 约翰 进了 西门 和 安得烈 的家。
MARK|1|30|西门 的岳母正发烧躺着，就有人告诉耶稣。
MARK|1|31|耶稣进前拉着她的手，扶她起来，烧就退了，于是她服事他们。
MARK|1|32|傍晚日落的时候，有人带着一切害病的和被鬼附的，来到耶稣跟前。
MARK|1|33|全城的人都聚集在门前。
MARK|1|34|耶稣治好了许多害各样病的人，又赶出许多鬼，不许鬼说话，因为鬼认识他。
MARK|1|35|次日早晨，天未亮的时候，耶稣起来，到旷野地方去，在那里祷告。
MARK|1|36|西门 和同伴出去找他，
MARK|1|37|找到了就对他说：“众人都在找你！”
MARK|1|38|耶稣对他们说：“让我们往别处去，到邻近的乡村，我也好在那里传道，因为我是为这事出来的。”
MARK|1|39|于是他走遍全 加利利 ，在他们的会堂传道，并且赶鬼。
MARK|1|40|有一个痲疯病人来求耶稣，向他跪下 ，说：“你若肯，你能使我洁净。”
MARK|1|41|耶稣动了慈心，就伸手摸他，说：“我肯，你洁净了吧！”
MARK|1|42|痲疯病立刻离开他，他就洁净了。
MARK|1|43|耶稣严严地叮嘱他，立刻打发他走，
MARK|1|44|对他说：“你要注意，千万不可告诉任何人，只要去，让祭司为你检查，又因为你已经洁净，献上 摩西 所吩咐的祭物，作为证据给众人看。”
MARK|1|45|那人出去，倒说许多的话，把这件事传扬开了，使耶稣不能再公开进城，只好留在外边旷野地方，人从各处都到他跟前来。
MARK|2|1|过了些日子，耶稣又进了 迦百农 。人听说他在屋里，
MARK|2|2|于是许多人聚集，甚至连门前都没有空地；耶稣就对他们讲道。
MARK|2|3|有人带着一个瘫子来见耶稣，是由四个人抬来的；
MARK|2|4|因为人多，无法抬到耶稣跟前，就把他所在那房子的屋顶拆了，既拆通了，就把瘫子连所躺卧的褥子都缒下去。
MARK|2|5|耶稣见他们的信心，就对瘫子说：“孩子，你的罪赦了。”
MARK|2|6|有几个文士坐在那里，心里议论，说：
MARK|2|7|“这个人为什么这样说呢？他说亵渎的话了。除了上帝一位之外，谁能赦罪呢？”
MARK|2|8|耶稣心中立刻知道他们心里这样议论，就说：“你们心里为什么这样议论呢？
MARK|2|9|对瘫子说‘你的罪赦了’，或说‘起来！拿你的褥子行走’，哪一样容易呢？
MARK|2|10|但要让你们知道，人子在地上有赦罪的权柄。”就对瘫子说：
MARK|2|11|“我吩咐你，起来！拿你的褥子回家去吧。”
MARK|2|12|那人就起来，立刻拿着褥子，当着众人面前出去了，以致众人都惊奇，归荣耀给上帝，说：“我们从来没有见过这样的事！”
MARK|2|13|耶稣又到海边去，众人都到他跟前来，他就教导他们。
MARK|2|14|耶稣往前走，看见 亚勒腓 的儿子 利未 在税关坐着，就对他说：“来跟从我！”他就起来跟从耶稣。
MARK|2|15|耶稣在 利未 家里坐席的时候，有好些税吏和罪人与耶稣和他的门徒一同坐席，因为有很多人也跟随耶稣。
MARK|2|16|法利赛人中的文士 看见耶稣与罪人和税吏一同吃饭，就对他的门徒说：“他与税吏和罪人一同吃饭吗？”
MARK|2|17|耶稣听见，就对他们说：“健康的人用不着医生，有病的人才用得着。我不是来召义人，而是召罪人。”
MARK|2|18|那时， 约翰 的门徒和法利赛人都禁食。他们来问耶稣说：“ 约翰 的门徒和法利赛人的门徒禁食，你的门徒却不禁食，这是为什么呢？”
MARK|2|19|耶稣对他们说：“新郎和宾客在一起的时候，宾客怎么能禁食呢？只要新郎和他们在一起，他们不能禁食。
MARK|2|20|但日子将到，新郎要被带走，那日他们就要禁食了。
MARK|2|21|“没有人把新布缝在旧衣服上，若是这样，所补上的新布会撕破旧衣服，裂口就更大了。
MARK|2|22|也没有人把新酒装在旧皮袋里，若是这样，酒会胀破皮袋，酒和皮袋都糟蹋了 。相反地，新酒要装在新皮袋里 。”
MARK|2|23|有一个安息日，耶稣从麦田经过。他的门徒走路的时候，摘起麦穗来。
MARK|2|24|法利赛人对耶稣说：“看哪！他们为什么做安息日不合法的事呢？”
MARK|2|25|耶稣对他们说：“ 大卫 和跟从他的人饥饿需要食物时所做的事，你们没有念过吗？
MARK|2|26|他在 亚比亚他 作大祭司的时候，怎么进了上帝的居所，吃了供饼，又给跟从他的人吃呢？这饼除了祭司以外，人都不可以吃。”
MARK|2|27|他又对他们说：“安息日是为人设立的，人不是为安息日设立的。
MARK|2|28|所以，人子也是安息日的主。”
MARK|3|1|耶稣又进了会堂，在那里有一个人，他的一只手萎缩了。
MARK|3|2|众人为了要控告耶稣，就窥探他会不会在安息日医治那人。
MARK|3|3|耶稣对那手萎缩了的人说：“起来站在当中！”
MARK|3|4|他又问众人：“在安息日行善行恶，救命害命，哪样是合法的呢？”他们都不作声。
MARK|3|5|耶稣怒目环视他们，因他们的心刚硬而忧伤，就对那人说：“伸出手来！”他把手一伸，手就复原了。
MARK|3|6|法利赛人出去，立刻同 希律 一党的人商议怎样除掉耶稣。
MARK|3|7|耶稣和门徒退到海边去，有许多人从 加利利 跟随他。还有许多人听见他所做的事，就从 犹太 、 耶路撒冷 、 以土买 、 约旦河 的东边，以及 推罗 和 西顿 的附近地方来到他那里。
MARK|3|8|
MARK|3|9|因为人多，他吩咐门徒为他预备一只小船，免得众人拥挤他。
MARK|3|10|他治好了许多人，所以凡有疾病的，都挤着要摸他。
MARK|3|11|每当污灵看见他，就俯伏在他面前，喊着说：“你是上帝的儿子。”
MARK|3|12|耶稣再三嘱咐他们不要把他宣扬出去。
MARK|3|13|耶稣上了山，把自己所要的人召来，他们就来到他那里。
MARK|3|14|于是他设立十二个人，又称他们为使徒 ，要他们常和自己同在，也要差他们去传道，
MARK|3|15|并给他们权柄赶鬼。
MARK|3|16|他设立的十二个人 有 西门 －耶稣又给他起名叫 彼得 ，
MARK|3|17|还有 西庇太 的儿子 雅各 和 雅各 的弟弟 约翰 —耶稣又给他们起名叫 半尼其 ，就是雷的儿子—
MARK|3|18|又有 安得烈 、 腓力 、 巴多罗买 、 马太 、 多马 、 亚勒腓 的儿子 雅各 、 达太 和激进党的 西门 ，
MARK|3|19|还有出卖耶稣的 加略 人 犹大 。
MARK|3|20|耶稣进了屋子，众人又聚集，甚至他连饭也顾不得吃。
MARK|3|21|耶稣的家人听见，就出来要拉住他，因为他们说他癫狂了。
MARK|3|22|从 耶路撒冷 下来的文士说：“他是被 别西卜 附身的”，又说：“他是靠着鬼王赶鬼的。”
MARK|3|23|耶稣叫他们来，用比喻对他们说：“撒但怎能赶出撒但呢？
MARK|3|24|一国若自相纷争，那国就立不住；
MARK|3|25|一家若自相纷争，那家就立不住。
MARK|3|26|撒但若自相攻打纷争，他就立不住，必定灭亡。
MARK|3|27|没有人能进壮士家里，抢夺他的东西；除非先绑住那壮士，否则无法抢夺他的家。
MARK|3|28|我实在告诉你们，世人一切的罪和一切亵渎的话都可以得到赦免；
MARK|3|29|凡亵渎圣灵的，却永不得赦免，而要担当永远的罪。”
MARK|3|30|因为他们说：“他是被污灵附身的。”
MARK|3|31|那时，耶稣的母亲和他兄弟来，站在外边，打发人去叫他。
MARK|3|32|有许多人在耶稣周围坐着，他们就告诉他说：“看哪！你母亲、你兄弟和你姊妹 在外边找你。”
MARK|3|33|耶稣回答他们：“谁是我的母亲？谁是我的兄弟？”
MARK|3|34|就环视那周围坐着的人，说：“看哪，我的母亲，我的兄弟！
MARK|3|35|凡遵行上帝旨意的人就是我的兄弟姊妹和母亲。”
MARK|4|1|耶稣又在海边教导人。有一大群人到他那里聚集，他只好上船坐下。船在海里，众人都靠近海，站在岸上。
MARK|4|2|耶稣就用许多比喻教导他们。在教导的时候，他对他们说：
MARK|4|3|“你们听啊，有一个撒种的出去撒种。
MARK|4|4|他撒的时候，有的落在路旁，飞鸟来把它吃掉了。
MARK|4|5|有的落在土浅的石头地上，因为土不深，很快就长出苗来，
MARK|4|6|太阳出来一晒，因为没有根就枯干了。
MARK|4|7|有的落在荆棘里，荆棘长起来，把它挤住了，就结不出果实。
MARK|4|8|又有的落在好土里，就发芽长大，结出果实，有三十倍的，有六十倍的，有一百倍的。”
MARK|4|9|耶稣又说：“有耳可听的，就应当听！”
MARK|4|10|耶稣独自一人的时候，跟随他的人和十二使徒问他这些比喻的意思。
MARK|4|11|耶稣对他们说：“上帝国的奥秘只让你们知道，若是对外人讲，凡事就用比喻，
MARK|4|12|要 他们看了又看，却看不清， 听了又听，却不明白， 免得他们回转过来，获得赦免。”
MARK|4|13|耶稣又对他们说：“你们不明白这比喻吗？这样怎能明白一切的比喻呢？
MARK|4|14|撒种的人所撒的就是道。
MARK|4|15|那撒在路旁的种子，就是人听了道，撒但立刻来，把撒在他们心里的道夺了去。
MARK|4|16|那撒在石头地上的，就是人听了道，立刻欢喜领受，
MARK|4|17|因心里没有根，不过是暂时的，一旦为道遭受患难或迫害，立刻就跌倒。
MARK|4|18|还有那撒在荆棘里的，就是人听了道，
MARK|4|19|后来有世上的忧虑、钱财的迷惑，和别样的私欲进来，把道挤住了，结不出果实。
MARK|4|20|那撒在好土里的，就是人听了道，领受了，并且结了果实，有三十倍的，有六十倍的，有一百倍的。”
MARK|4|21|耶稣又对他们说：“人拿灯来，难道是要放在斗底下，床底下，而不放在灯台上吗？
MARK|4|22|因为掩藏的事没有不显出来的，隐瞒的事也没有不露出来的。
MARK|4|23|有耳可听的，就应当听！”
MARK|4|24|他又说：“你们要留心所听的。你们用什么量器来量，也将要用什么来量给你们，并且要多给你们。
MARK|4|25|因为有的，还要给他；没有的，连他所有的也要夺去。”
MARK|4|26|耶稣又说：“上帝的国如同人把种子撒在地上，
MARK|4|27|黑夜睡觉，白日起来，这种子就发芽生长，那人却不知道如何会这样。
MARK|4|28|土地自然而然地出产五谷，先发苗，后长穗，然后穗上结成饱满的谷子。
MARK|4|29|五谷熟了，就用镰刀去割，因为收成的时候到了。”
MARK|4|30|耶稣又说：“我们可用什么来比拟上帝的国呢？可用什么比喻来说明呢？
MARK|4|31|它像一粒芥菜种，种在地里的时候，虽比地上所有的种子都小，
MARK|4|32|但种下去以后，它长起来，比各样的菜都大，又长出大枝，以致天上的飞鸟可以在它的荫下筑巢。”
MARK|4|33|耶稣用许多这样的比喻，照他们所能听的，对他们讲道；
MARK|4|34|若不用比喻，他就不对他们讲，但私下没有人的时候，就把一切的道讲给门徒听。
MARK|4|35|那天晚上，耶稣对门徒说：“我们渡到对岸去吧。”
MARK|4|36|门徒离开众人，耶稣已在船上，他们就请他一同去；也有别的船和他同行。
MARK|4|37|忽然狂风大作，波浪打入船内，以致船灌满了水。
MARK|4|38|耶稣在船尾上，枕着枕头睡觉。门徒叫醒他，说：“老师！我们快没命了，你不管吗？”
MARK|4|39|耶稣醒了，斥责那风，向海说：“住了吧！静了吧！”风就止住，大大平静了。
MARK|4|40|耶稣对他们说：“为什么胆怯？你们还没有信心吗？”
MARK|4|41|他们就非常惧怕，彼此说：“这到底是谁？连风和海都听从他。”
MARK|5|1|他们渡到海的对岸，到 格拉森 人 的地区。
MARK|5|2|耶稣一下船，就有一个污灵附身的人从坟墓迎着他走来。
MARK|5|3|那人常住在坟墓里，没有人能捆住他，就是用铁链也不能；
MARK|5|4|因为人屡次用脚镣和铁链捆锁他，铁链被他挣断，脚镣也被他弄碎了，总没有人能制伏他。
MARK|5|5|他昼夜常在坟墓里和山中喊叫，又用石头打自己。
MARK|5|6|他远远看见耶稣，就跑过来拜他，
MARK|5|7|大声呼叫说：“至高上帝的儿子耶稣，你为什么干扰我？我指着上帝恳求你，不要叫我受苦！”
MARK|5|8|这是因耶稣曾吩咐他说：“污灵啊，从这人身上出来！”
MARK|5|9|耶稣问他：“你叫什么名字？”他说：“我名叫 群 ，因为我们数目众多。”
MARK|5|10|他就再三求耶稣不要叫他们离开那地方。
MARK|5|11|在山坡那里，有一大群猪正在吃食；
MARK|5|12|污灵就央求耶稣，说：“求你打发我们进入猪群，好附着它们。”
MARK|5|13|耶稣准了他们，污灵就出来，进入猪里，那群猪就闯下山崖，投进海里，淹死了。猪的数目约有二千。
MARK|5|14|放猪的逃跑了，去告诉城里和乡下的人。众人就来，要看发生了什么事。
MARK|5|15|他们来到耶稣那里，看见那被鬼附的人，就是曾被群鬼所附的，坐着，穿着衣服，神智清醒，他们就害怕。
MARK|5|16|看见这事的人把被鬼附的人所遇见的，和那群猪的事，都告诉了众人，
MARK|5|17|众人就央求耶稣离开他们的地区。
MARK|5|18|耶稣上船的时候，那曾被鬼附的人恳求要和耶稣在一起。
MARK|5|19|耶稣不许，却对他说：“你回家去，到你的亲友那里，将主为你所做多么大的事和他怎样怜悯你，都告诉他们。”
MARK|5|20|那人就走了，开始在 低加坡里 传扬耶稣为他做了多么大的事，众人就都惊讶。
MARK|5|21|耶稣又坐船 渡到对岸，有一大群人聚集到他身边；他正在海边。
MARK|5|22|有一个会堂主管，名叫 叶鲁 ，也来了，一见到耶稣，就俯伏在他脚前，
MARK|5|23|再三求他，说：“我的小女儿快要死了，求你去为她按手，使她痊愈，可以活下去。”
MARK|5|24|耶稣就和他同去。 有一大群人跟随他，拥挤着他。
MARK|5|25|有一个女人，患了经血不止的病有十二年，
MARK|5|26|在好多医生手里受了许多苦，又花尽了她所有的，一点也不见好，反而更重了。
MARK|5|27|她听见耶稣的事，就夹在众人中间，从后面来摸耶稣的衣裳，
MARK|5|28|因她想：“我只摸到他的衣裳，就会痊愈。”
MARK|5|29|于是她的流血立刻止住，她觉得身上的疾病好了。
MARK|5|30|耶稣顿时心里觉得有能力从自己身上出去，就在众人中间转过来，说：“谁摸我的衣裳？”
MARK|5|31|门徒对他说：“你看众人拥挤着你，还说‘谁摸我’呢？”
MARK|5|32|耶稣周围观看，要见做这事的女人。
MARK|5|33|那女人知道在自己身上所成的事，就恐惧战兢，来俯伏在耶稣跟前，将实情全告诉他。
MARK|5|34|耶稣对她说：“女儿，你的信救了你，平安地回去吧！你的疾病痊愈了。”
MARK|5|35|耶稣还在说话的时候，有人从会堂主管的家里来，说：“你的女儿死了，何必还劳驾老师呢？”
MARK|5|36|耶稣不理会他们所说的话，就对会堂主管说：“不要怕，只要信！”
MARK|5|37|于是他带着 彼得 、 雅各 和 雅各 的弟弟 约翰 同去，不许别人跟着他。
MARK|5|38|他们来到会堂主管的家里，耶稣看到一片吵闹，并有人大声哭泣哀号，
MARK|5|39|就进到里面，对他们说：“为什么大吵大哭呢？孩子不是死了，是睡着了。”
MARK|5|40|他们就嘲笑耶稣。耶稣把他们都赶出去，带着孩子的父母和跟随的人进了孩子所在的地方，
MARK|5|41|就拉着孩子的手，对她说：“大利大，古米！”翻出来就是说：“女孩，我吩咐你，起来！”
MARK|5|42|那女孩子立刻起来走动—她已经十二岁了；他们就非常惊奇。
MARK|5|43|耶稣切切地嘱咐他们，不要让人知道这事，又吩咐给她东西吃。
MARK|6|1|耶稣离开那里，来到自己的家乡；门徒也跟从他。
MARK|6|2|到了安息日，他在会堂里教导人。众人听见，就很惊奇，说：“这人哪来这本事呢？所赐给他的是什么智慧？他手所做的是何等的异能呢？
MARK|6|3|这不是那木匠吗？不是 马利亚 的儿子 雅各 、 约西 、 犹大 、 西门 的长兄吗？他姊妹们不也是在我们这里吗？”他们就厌弃他。
MARK|6|4|耶稣对他们说：“先知除了在本乡、本族和自己的家之外，没有不被尊敬的。”
MARK|6|5|耶稣在那里不能行什么异能，不过为几个病人按手，治好他们。
MARK|6|6|他也诧异他们不信。 耶稣走遍周围乡村教导人。
MARK|6|7|他叫了十二个使徒来，差遣他们两个两个地出去，也赐给他们权柄制伏污灵，
MARK|6|8|并且吩咐他们：途中不要带食物和行囊，腰袋里也不要带钱，除了手杖以外，什么都不要带；
MARK|6|9|只要穿鞋子，也不要穿两件内衣。
MARK|6|10|他又对他们说：“你们无论到何处，进哪家，就住在哪里，直到离开那地方。
MARK|6|11|若有什么地方的人不接待你们，不听你们，你们离开那里的时候，要跺掉你们脚上的尘土，证明他们的不是。”
MARK|6|12|使徒就出去传道，叫人悔改，
MARK|6|13|又赶出许多鬼，用油抹了许多病人，治好他们。
MARK|6|14|耶稣的名声传开了， 希律 王也听见。有人说：“施洗的 约翰 从死人中复活了，因此才有这些异能在他里面运行。”
MARK|6|15|但别人说：“他是 以利亚 。”又有人说：“是先知，正如先知中的一位。”
MARK|6|16|希律 听见却说：“是我所斩的 约翰 ，他复活了。”
MARK|6|17|原来， 希律 为他兄弟 腓力 的妻子 希罗底 的缘故，派人去抓了 约翰 ，把他绑了在监狱里，因为 希律 已经娶了那妇人。
MARK|6|18|约翰 曾对 希律 说：“你占有你兄弟的妻子是不合法的。”
MARK|6|19|于是 希罗底 怀恨他，想要杀他，只是不能。
MARK|6|20|因为 希律 怕 约翰 ，知道他是义人，是圣人，所以就保护他，虽然听了他的讲论十分困惑 ，仍然乐意听他。
MARK|6|21|有一天，恰巧是 希律 的生日， 希律 摆设宴席，请了大臣、千夫长和 加利利 的领袖。
MARK|6|22|他的女儿 希罗底 进来跳舞，使 希律 和同席的人都很高兴。王就对女孩说：“无论你要什么，向我求，我都会给你”；
MARK|6|23|又对她多次 起誓说：“无论你向我求什么，就是我国家的一半，我也会给你。”
MARK|6|24|她就出去对她母亲说：“我该求什么呢？”她母亲说：“施洗 约翰 的头。”
MARK|6|25|她就急忙进去见王，求他说：“我愿王立刻把施洗 约翰 的头放在盘子里给我。”
MARK|6|26|王就很忧愁，然而因他所发的誓，又因同席的人，不愿食言，
MARK|6|27|就立刻派一个卫兵，吩咐拿 约翰 的头来。卫兵就去，在监狱里斩了 约翰 ，
MARK|6|28|把头放在盘子里，拿来给那女孩，她就给她母亲。
MARK|6|29|约翰 的门徒听到了，就来把他的尸体领去，放在坟墓里。
MARK|6|30|使徒们聚集到耶稣那里，把一切所做的事、所传的道全告诉他。
MARK|6|31|他就说：“你们来，同我私下到荒野的地方去歇一歇。”这是因为来往的人多，他们连吃饭的时间也没有。
MARK|6|32|他们就坐船，私下往荒野的地方去。
MARK|6|33|众人看见他们走了，有许多认识他们的，就从各城步行，一同跑到那里，比他们先赶到了。
MARK|6|34|耶稣出来，见有一大群的人，就怜悯他们，因为他们如同羊没有牧人一般，于是开始教导他们许多事。
MARK|6|35|天已经很晚，门徒进前来，说：“这地方偏僻，而且天已经很晚了，
MARK|6|36|请叫众人散去，他们好往四面的乡镇村庄去，自己买些东西吃。”
MARK|6|37|耶稣回答他们说：“你们给他们吃吧！”门徒对他说：“我们要拿两百个银币去买饼给他们吃吗？”
MARK|6|38|耶稣说：“你们有多少饼？去看看。”他们知道后就说：“有五个，还有两条鱼。”
MARK|6|39|耶稣吩咐他们，叫众人一组一组地坐在青草地上。
MARK|6|40|众人就一群一群地坐下，有一百的，有五十的。
MARK|6|41|耶稣拿着这五个饼和两条鱼，望着天祝福，擘开饼，递给门徒，摆在众人面前，也把那两条鱼分给众人。
MARK|6|42|他们都吃，并且吃饱了。
MARK|6|43|门徒把饼和鱼的碎屑收拾起来，装满了十二个篮子。
MARK|6|44|吃饼的男人共有五千。
MARK|6|45|耶稣随即催门徒上船，先渡到对岸，到 伯赛大 去，等他叫众人散去。
MARK|6|46|他辞别了他们，就往山上去祷告。
MARK|6|47|到了晚上，船在海中，耶稣独自在岸上。
MARK|6|48|他看见门徒因风不顺，摇橹很苦。天快亮的时候，他在海面上走，往他们那里去，想要超过他们。
MARK|6|49|但门徒看见他在海面上走，以为是鬼怪，就喊叫起来；
MARK|6|50|因为他们都看见了他，甚为惊慌。耶稣连忙对他们说：“放心！是我，不要怕！”
MARK|6|51|于是他到他们那里，一上船，风就停了；他们心里十分惊奇。
MARK|6|52|这是因为他们不明白那分饼的事，心里还是愚顽。
MARK|6|53|他们渡过了海，在 革尼撒勒 靠岸，泊了船，
MARK|6|54|他们一下来，众人立刻认出是耶稣，
MARK|6|55|就跑遍那整个地区，听到他在哪里，就把有病的人用褥子抬到哪里。
MARK|6|56|耶稣所到的地方，或村中、或城里、或乡间，他们都把病人放在街市上，求耶稣让他们摸一摸他的衣裳繸子，摸着的人就都好了。
MARK|7|1|有法利赛人和几个从 耶路撒冷 来的文士聚集到耶稣那里。
MARK|7|2|他们曾看见他的门徒中有人用不洁净的手，就是没有洗的手吃饭。
MARK|7|3|法利赛人和所有的 犹太 人都拘守古人的传统，若不按规矩洗手就不吃饭；
MARK|7|4|从市场来，若不洗净也不吃饭；他们还拘守好些别的规矩，如洗杯、罐、铜器、床铺 等。
MARK|7|5|法利赛人和文士问他说：“你的门徒为什么不照古人的传统，竟然用不洁净的手吃饭呢？”
MARK|7|6|耶稣对他们说：“ 以赛亚 指着你们假冒为善的人所预言的说得好。如经上所记： ‘这百姓用嘴唇尊敬我， 他们的心却远离我。
MARK|7|7|他们把人的规条当作教义教导人； 他们拜我也是枉然。’
MARK|7|8|你们是离弃上帝的诫命，拘守人的传统。”
MARK|7|9|耶稣又说：“你们诚然是废弃上帝的诫命，为要守自己的传统。
MARK|7|10|摩西 说：‘当孝敬父母’；又说：‘咒骂父母的，必须处死。’
MARK|7|11|你们倒说：‘人若对父母说：我所当供奉你的已经作了各耳板’（各耳板就是奉献的意思），
MARK|7|12|你们就容许他不必再奉养父母。
MARK|7|13|这就是你们藉着继承传统，废了上帝的话。你们还做许多这样的事。”
MARK|7|14|耶稣又叫众人来，对他们说：“你们都要听我的话，也要明白。
MARK|7|15|从外面进去的不能玷污人，惟有从里面出来的才玷污人。 ”
MARK|7|16|
MARK|7|17|耶稣离开众人，进了屋子，门徒就问他这比喻的意思。
MARK|7|18|耶稣对他们说：“你们也是这样不明白吗？难道你们不了解，凡从外面进去的不能玷污人吗？
MARK|7|19|因为不是进入他的心，而是进入他的肚子，又排入厕所。”（这是说，各样的食物都是洁净的。）
MARK|7|20|耶稣又说：“从人里面出来的，那才玷污人；
MARK|7|21|因为从人心里发出种种恶念，如淫乱、偷盗、凶杀、
MARK|7|22|奸淫、贪婪、邪恶、诡诈、淫荡、嫉妒、毁谤、骄傲、狂妄。
MARK|7|23|这一切的恶都是从里面出来，且能玷污人。”
MARK|7|24|耶稣从那里起身，往 推罗 境内去，进了一家，他不愿意人知道，却隐藏不住。
MARK|7|25|立刻有一个妇人，她的小女儿被污灵附着，一听见耶稣的事，就来俯伏在他脚前。
MARK|7|26|这妇人是 希腊 人，属 叙利亚 的 腓尼基 族。她求耶稣从她女儿身上赶出那鬼。
MARK|7|27|耶稣对她说：“让孩子们先吃饱，拿孩子的饼丢给小狗吃是不妥的。”
MARK|7|28|妇人回答：“主啊，桌子底下的小狗也吃小孩子的碎屑呀！”
MARK|7|29|耶稣对她说：“凭着这句话，你回去吧，鬼已经离开你的女儿了。”
MARK|7|30|她就回家去，见小孩子躺在床上，鬼已经出去了。
MARK|7|31|耶稣又离开了 推罗 地区，经过 西顿 ，就从 低加坡里 境内来到 加利利海 。
MARK|7|32|有人带着一个耳聋舌结的人来见耶稣，求他为他按手。
MARK|7|33|耶稣领他离开众人，到一边去，就用指头探他的耳朵，吐唾沫抹他的舌头，
MARK|7|34|望天叹息，对他说：“以法大！”就是说“开了吧！”
MARK|7|35|他的耳朵立刻 开了，舌结也解了，他说话也清楚了。
MARK|7|36|耶稣嘱咐他们不要告诉人；但他越嘱咐，他们越发传扬。
MARK|7|37|众人分外惊奇，说：“他所做的事样样都好，他甚至使聋子听见，哑巴说话。”
MARK|8|1|那时，又有一大群人聚集，没有什么吃的。耶稣叫门徒来，说：
MARK|8|2|“我怜悯这群人，因为他们同我在这里已经三天，没有吃的东西了。
MARK|8|3|我若叫他们饿着回家，他们会在路上饿昏，因为其中有从远处来的。”
MARK|8|4|门徒回答：“在这野地，从哪里能得饼使这些人吃饱呢？”
MARK|8|5|耶稣问他们：“你们有多少饼？”他们说：“七个。”
MARK|8|6|他吩咐众人坐在地上，就拿着这七个饼祝谢了，擘开，递给门徒，叫他们摆开，门徒就摆在众人面前。
MARK|8|7|他们还有几条小鱼；耶稣祝谢了，就吩咐也摆在众人面前。
MARK|8|8|他们都吃，并且吃饱了，收拾剩下的碎屑，有七筐子。
MARK|8|9|人数约有四千。耶稣打发他们走了，
MARK|8|10|随即同门徒上船，来到 大玛努他 境内。
MARK|8|11|法利赛人出来盘问耶稣，要求他从天上显个神迹给他们看，想要试探他。
MARK|8|12|耶稣心里深深叹息，说：“这世代为什么求神迹呢？我实在告诉你们，没有神迹给这世代看。”
MARK|8|13|他就离开他们，又上船往海的对岸去了。
MARK|8|14|门徒忘了带饼，在船上除了一个饼，没有别的食物。
MARK|8|15|耶稣嘱咐他们说：“你们要谨慎，要防备法利赛人的酵和 希律 的酵。”
MARK|8|16|他们彼此议论说：“这是因为我们没有饼吧。”
MARK|8|17|耶稣知道了，就说：“你们为什么因为没有饼就议论呢？你们还不领悟，还不明白吗？你们的心还是愚顽吗？
MARK|8|18|你们有眼睛，看不见吗？有耳朵，听不到吗？也不记得吗？
MARK|8|19|我擘开那五个饼分给五千人，你们收拾的碎屑装满了多少个篮子呢？”他们说：“十二个。”
MARK|8|20|“又擘开那七个饼分给四千人，你们收拾的碎屑装满了多少个筐子呢？”他们说：“七个。”
MARK|8|21|耶稣说：“你们还不明白吗？”
MARK|8|22|他们来到 伯赛大 ，有人带一个盲人来，求耶稣摸他。
MARK|8|23|耶稣拉着盲人的手，领他到村外，就吐唾沫在他眼睛上，为他按手，问他：“你看见什么？”
MARK|8|24|他抬头一看，说：“我看见人，他们好像树木，并且行走。”
MARK|8|25|随后耶稣又按手在他眼睛上，他定睛一看，就复原了，样样都看得清楚了。
MARK|8|26|耶稣打发他回家，说：“连这村子你也不要进去。”
MARK|8|27|耶稣和门徒出去，往 凯撒利亚．腓立比 附近的村庄去。在路上，他问门徒：“人们说我是谁？”
MARK|8|28|他们对他说：“是施洗的 约翰 ；有人说是 以利亚 ；又有人说是先知中的一位。”
MARK|8|29|他又问他们：“你们说我是谁？” 彼得 回答他：“你是基督。”
MARK|8|30|于是耶稣切切地嘱咐他们不可对任何人说起他。
MARK|8|31|从此，他教导他们说：“人子必须受许多的苦，被长老、祭司长和文士弃绝，并且被杀，三天后复活。”
MARK|8|32|耶稣明白地说了这话， 彼得 就拉着他，责备他。
MARK|8|33|耶稣转过来看着门徒，斥责 彼得 说：“撒但，退到我后边去！因为你不体会上帝的心意，而是体会人的意思。”
MARK|8|34|于是他叫众人和门徒来，对他们说：“若有人要跟从我，就当舍己，背起自己的十字架来跟从我。
MARK|8|35|因为凡要救自己生命的，必丧失生命；凡为我和福音丧失生命的，必救自己的生命。
MARK|8|36|人就是赚得全世界，赔上自己的生命，有什么益处呢？
MARK|8|37|人还能拿什么换生命呢？
MARK|8|38|凡在这淫乱罪恶的世代，把我和我的道当作可耻的，人子在他父的荣耀里与圣天使一同来临的时候，也要把那人当作可耻的。”
MARK|9|1|耶稣又对他们说：“我实在告诉你们，站在这里的，有人在没经历死亡以前，必定看见上帝的国带着能力临到。”
MARK|9|2|过了六天，耶稣带着 彼得 、 雅各 、 约翰 ，领他们悄悄地上了高山。他在他们面前变了形像，
MARK|9|3|衣服放光，极其洁白，地上漂布的人没有一个能漂得那样白。
MARK|9|4|有 以利亚 和 摩西 向他们显现，并且与耶稣说话。
MARK|9|5|彼得 对耶稣说：“拉比 ，我们在这里真好！我们来搭三座棚，一座为你，一座为 摩西 ，一座为 以利亚 。”
MARK|9|6|彼得 不知道说什么才好，因为他们很害怕。
MARK|9|7|有一朵云彩来遮盖他们，又有声音从云彩里出来，说：“这是我的爱子，你们要听从他！”
MARK|9|8|门徒连忙向周围观看，不再看见任何人，只见耶稣同他们在一起。
MARK|9|9|下山的时候，耶稣嘱咐他们说：“人子还没有从死人中复活，你们不要把所看到的告诉人。”
MARK|9|10|门徒将这话存记在心，彼此议论“从死人中复活”是什么意思。
MARK|9|11|他们就问耶稣：“文士为什么说 以利亚 必须先来？”
MARK|9|12|耶稣说：“ 以利亚 的确先来复兴万事。经上不是指着人子说，他要受许多的苦和被人轻慢吗？
MARK|9|13|我告诉你们， 以利亚 已经来了，他们任意待他，正如经上指着他说的。”
MARK|9|14|他们到了门徒那里，看见有一大群人围着他们，又有文士和他们辩论。
MARK|9|15|众人一见耶稣，都很惊奇，就跑上去向他问安。
MARK|9|16|耶稣问他们：“你们和他们辩论什么？”
MARK|9|17|众人中的一个回答：“老师，我带了我的儿子到你这里来，他被哑巴的灵附着。
MARK|9|18|无论在哪里，那灵拿住他，把他摔倒，他就口吐白沫，牙关紧锁，身体僵硬。我请过你的门徒把那灵赶出去，他们却不能。”
MARK|9|19|耶稣回答：“唉！这不信的世代啊，我和你们在一起要到几时呢？我忍耐你们要到几时呢？把他带到我这里！”
MARK|9|20|他们就带了他来。那灵一见耶稣，就使他重重地抽风，倒在地上，翻来覆去，口吐白沫。
MARK|9|21|耶稣问他父亲：“他得这病有多久了呢？”父亲说：“从小的时候。
MARK|9|22|那灵屡次把他扔在火里、水里，要治死他。你若能做什么，求你怜悯我们，帮助我们。”
MARK|9|23|耶稣对他说：“‘你若能’，在信的人，凡事都能。”
MARK|9|24|孩子的父亲立刻喊着说：“我信；求你帮助我的不信！”
MARK|9|25|耶稣看见众人都跑上来，就斥责那污灵说：“你这聋哑的灵，我命令你从他里头出来，再不要进去！”
MARK|9|26|那灵大喊一声，使孩子猛烈地抽了一阵风，就出来了。孩子好像死了一般，以致众人多半说：“他死了。”
MARK|9|27|但耶稣拉着他的手，扶他起来，他就站起来了。
MARK|9|28|耶稣进了屋子，门徒就私下问他：“我们为什么不能赶出那灵呢？”
MARK|9|29|耶稣对他们说：“非用祷告 ，这一类的邪灵总赶不出来。”
MARK|9|30|他们离开那地方，经过 加利利 ；耶稣不愿意人知道，
MARK|9|31|因为他正教导门徒说：“人子将要被交在人手里，他们要杀害他；被杀以后，三天后他要复活。”
MARK|9|32|门徒却不明白这话，又不敢问他。
MARK|9|33|他们来到 迦百农 。耶稣在屋里问门徒说：“你们在路上议论的是什么？”
MARK|9|34|门徒不作声，因为他们在路上彼此争论谁最大。
MARK|9|35|耶稣坐下，叫十二个使徒来，说：“若有人愿意为首，他要作众人之后，作众人的用人。”
MARK|9|36|于是耶稣领一个小孩过来，让他站在门徒当中，又抱起他来，对他们说：
MARK|9|37|“凡为我的名接纳一个像这小孩子的，就是接纳我；凡接纳我的，不是接纳我，而是接纳那差我来的。”
MARK|9|38|约翰 对耶稣说：“老师，我们看见一个人奉你的名赶鬼，我们就阻止他，因为他不跟从我们。”
MARK|9|39|耶稣说：“不要阻止他，因为没有人奉我的名行异能，反倒轻易毁谤我。
MARK|9|40|不抵挡我们的，就是帮助我们的。
MARK|9|41|凡因你们是属基督，给你们一杯水喝的，我实在告诉你们，他一定会得到赏赐。”
MARK|9|42|“凡使这些信我的小子 中的一个跌倒的，倒不如把大磨石拴在这人的颈项上，扔在海里。
MARK|9|43|如果你一只手使你跌倒，就把它砍下来；你缺一只手进入永生，比有两只手落到地狱，入那不灭的火里去还好。
MARK|9|44|
MARK|9|45|如果你一只脚使你跌倒，就把它砍下来；你瘸腿进入永生，比有两只脚被扔进地狱里还好。
MARK|9|46|
MARK|9|47|如果你一只眼使你跌倒，就去掉它；你只有一只眼进入上帝的国，比有两只眼被扔进地狱里还好。
MARK|9|48|在那里，虫是不死的，火是不灭的。
MARK|9|49|因为每个人必被火像盐一般腌起来。
MARK|9|50|盐本是好的，若失了咸味，你们怎能用它调味呢？你们中间要有盐，彼此和睦。”
MARK|10|1|耶稣从那里起身，来到 犹太 的境内， 约旦河 的东边。众人又聚集到他那里，他又照常教导他们。
MARK|10|2|有法利赛人来问他说：“男人休妻合不合法？”意思是要试探他。
MARK|10|3|耶稣回答他们说：“ 摩西 吩咐你们的是什么？”
MARK|10|4|他们说：“ 摩西 准许写了休书就可以休妻。”
MARK|10|5|耶稣对他们说：“ 摩西 因为你们的心硬，所以写这诫命给你们。
MARK|10|6|但从起初创造的时候，上帝造人是造男造女。
MARK|10|7|因此，人要离开他的父母，与妻子结合 ，
MARK|10|8|二人成为一体。既然如此，夫妻不再是两个人，而是一体的了。
MARK|10|9|所以，上帝配合的，人不可分开。”
MARK|10|10|他们到了屋里，门徒又问他这事。
MARK|10|11|耶稣对他们说：“凡休妻另娶的，就是犯奸淫，辜负他的妻子；
MARK|10|12|妻子若离弃丈夫另嫁，也是犯奸淫了。”
MARK|10|13|有人带着小孩子来见耶稣，要他摸他们，门徒就责备那些人。
MARK|10|14|耶稣看见就很生气，对门徒说：“让小孩到我这里来，不要阻止他们，因为在上帝国的正是这样的人。
MARK|10|15|我实在告诉你们，凡要接受上帝国的，若不像小孩子，绝不能进去。”
MARK|10|16|于是他抱着小孩子，给他们按手，为他们祝福。
MARK|10|17|耶稣刚上路的时候，有一个人跑来，跪在他面前，问他：“善良的老师，我该做什么事才能承受永生？”
MARK|10|18|耶稣对他说：“你为什么称我是善良的？除了上帝一位之外，再没有善良的。
MARK|10|19|诫命你是知道的：‘不可杀人；不可奸淫；不可偷盗；不可作假见证；不可亏负人；当孝敬父母。’”
MARK|10|20|他对耶稣说：“老师，这一切我从小都遵守了。”
MARK|10|21|耶稣看着他，就爱他，对他说：“你还缺少一件：去变卖你所有的，分给穷人，就必有财宝在天上；然后来跟从我。”
MARK|10|22|他听见这话，脸就变了色，忧忧愁愁地走了，因为他的产业很多。
MARK|10|23|耶稣看了看周围，对门徒说：“有钱财的人进上帝的国是何等的难哪！”
MARK|10|24|门徒对他的话非常惊奇。耶稣又对他们说：“孩子们， 要进上帝的国是何等的难哪！
MARK|10|25|骆驼穿过针眼比财主进上帝的国还容易呢！”
MARK|10|26|门徒就更为惊讶，彼此对问：“这样，谁能得救呢？”
MARK|10|27|耶稣看着他们，说：“在人不能，在上帝却不然，因为在上帝凡事都能。”
MARK|10|28|彼得 就对他说：“看哪，我们已经撇下一切跟从你了。”
MARK|10|29|耶稣说：“我实在告诉你们，凡为我和福音撇下房屋，或是兄弟、姊妹、父亲、母亲、儿女、田地，
MARK|10|30|没有不在今世得百倍的，就是房屋、兄弟、姊妹、母亲、儿女、田地，并且要受迫害，在来世得永生。
MARK|10|31|然而，有许多在前的，将要在后；在后的，将要在前。”
MARK|10|32|他们行路上 耶路撒冷 去。耶稣在前头走，他们很惊讶，跟从的人也害怕。耶稣又叫十二使徒来，把自己将要遭遇的事告诉他们，
MARK|10|33|说：“看哪，我们上 耶路撒冷 去，人子将被交给祭司长和文士；他们要定他死罪，又交给外邦人。
MARK|10|34|他们要戏弄他，向他吐唾沫，鞭打他，杀害他；三天后，他要复活。”
MARK|10|35|西庇太 的儿子 雅各 和 约翰 进前来，对耶稣说：“老师，我们无论求你什么，愿你为我们做。”
MARK|10|36|耶稣对他们说：“要我为你们做什么？”
MARK|10|37|他们对他说：“在你的荣耀里，请赐我们一个坐在你右边，一个坐在你左边。”
MARK|10|38|耶稣对他们说：“你们不知道所求的是什么。我所喝的杯，你们能喝吗？我所受的洗，你们能受吗？”
MARK|10|39|他们对他说：“我们能。”耶稣对他们说：“我所喝的杯，你们要喝；我所受的洗，你们也要受。
MARK|10|40|可是坐在我的左右，不是我可以赐的，而是为谁预备就赐给谁。”
MARK|10|41|其余十个门徒听见，就对 雅各 和 约翰 很生气。
MARK|10|42|耶稣叫了他们来，对他们说：“你们知道，外邦人有君王作主治理他们，有大臣操权管辖他们。
MARK|10|43|但是在你们中间，不可这样。你们中间谁愿为大，就要作你们的用人；
MARK|10|44|在你们中间谁愿为首，就要作众人的仆人。
MARK|10|45|因为人子来，并不是要受人的服事，乃是要服事人，并且要舍命作多人的赎价。”
MARK|10|46|他们到了 耶利哥 。耶稣同门徒并许多人离开 耶利哥 的时候，有一个讨饭的盲人，是 底买 的儿子 巴底买 ，坐在路旁。
MARK|10|47|他听见是 拿撒勒 的耶稣，就喊了起来，说：“ 大卫 之子耶稣啊，可怜我吧！”
MARK|10|48|有许多人责备他，不许他作声，他却越发喊着：“ 大卫 之子啊，可怜我吧！”
MARK|10|49|耶稣就站住，说：“叫他过来。”他们就叫那盲人，对他说：“放心，起来！他在叫你啦。”
MARK|10|50|盲人就丢下衣服，跳起来，走到耶稣那里。
MARK|10|51|耶稣回答他说：“你要我为你做什么？”盲人对他说：“拉波尼 ，我要能看见。”
MARK|10|52|耶稣对他说：“你去吧！你的信救了你。”盲人立刻看得见，就在路上跟随耶稣。
MARK|11|1|耶稣和门徒快到 耶路撒冷 ，来到 伯法其 和 伯大尼 ，在 橄榄山 那里。耶稣打发两个门徒，
MARK|11|2|对他们说：“你们往对面村子里去，一进去的时候会看见一匹驴驹拴在那里，是从来没有人骑过的，把它解开，牵来。
MARK|11|3|若有人对你们说：‘为什么做这事？’你们就说：‘主要用它，但会立刻把它牵回到这里来。’”
MARK|11|4|他们去了，看见一匹驴驹拴在门外街道上，就把它解开。
MARK|11|5|在那里站着的人，有几个说：“你们解开驴驹做什么？”
MARK|11|6|门徒照着耶稣的话说，那些人就任凭他们牵去了。
MARK|11|7|他们把驴驹牵到耶稣那里，把自己的衣服搭在上面，耶稣就骑上。
MARK|11|8|有许多人把衣服铺在路上，还有人把田间的树枝砍下来铺上。
MARK|11|9|前呼后拥的人都喊着说： “和散那 ！ 奉主名来的是应当称颂的！
MARK|11|10|那将要来的我祖 大卫 之国是应当称颂的！ 至高无上的，和散那！”
MARK|11|11|耶稣到了 耶路撒冷 ，进入圣殿，看了周围的一切。天色已晚，他就和十二使徒出城，往 伯大尼 去。
MARK|11|12|第二天，他们从 伯大尼 出来，耶稣饿了。
MARK|11|13|他远远地看见一棵无花果树，树上有叶子，就过去，看是不是在树上可以找到什么。他到了树下，竟找不到什么，只有叶子，因为不是无花果的季节。
MARK|11|14|耶稣就对树说：“从今以后，永没有人吃你的果子。”他的门徒都听到了。
MARK|11|15|他们来到 耶路撒冷 。耶稣一进圣殿，就赶出在圣殿里做买卖的人，推倒兑换银钱之人的桌子和卖鸽子之人的凳子；
MARK|11|16|也不许人拿着器具从圣殿里经过。
MARK|11|17|他教导他们说：“经上不是记着： ‘我的殿要称为万国祷告的殿吗？ 你们倒使它成为贼窝了。’”
MARK|11|18|祭司长和文士听见这话，就想法子要除掉耶稣，却又怕他，因为众人都对他的教导感到惊奇。
MARK|11|19|每天晚上，他们 都到城外去。
MARK|11|20|早晨，他们从那里经过，看见无花果树连根都枯干了。
MARK|11|21|彼得 想起耶稣的话来，就对他说：“拉比，你看！你所诅咒的无花果树已经枯干了。”
MARK|11|22|耶稣回答：“你们对上帝要有信心。
MARK|11|23|我实在告诉你们，无论何人对这座山说：‘离开此地，投在海里！’他心里若不疑惑，只信所说的必成，就为他实现。
MARK|11|24|所以我告诉你们，凡你们祷告祈求的，无论是什么，只要信你们已经得着了，就为你们实现。
MARK|11|25|你们站着祷告的时候，若想起有人得罪你们，就该饶恕他，好让你们在天上的父也饶恕你们的过犯。 ”
MARK|11|26|
MARK|11|27|他们又来到 耶路撒冷 。耶稣在圣殿里行走的时候，祭司长、文士和长老进前来，
MARK|11|28|问他说：“你仗着什么权柄做这些事？给你权柄做这些事的是谁呢？”
MARK|11|29|耶稣对他们说：“我要问你们一句话，你们回答我，我就告诉你们我仗着什么权柄做这些事。
MARK|11|30|约翰 的洗礼是从天上来的，还是从人间来的呢？你们回答我吧。”
MARK|11|31|他们彼此商议说：“我们若说‘从天上来的’，他会说：‘这样，你们为什么不信他呢？’
MARK|11|32|但若说‘从人间来的’，却又怕众人，因为大家认为 约翰 确是先知。”
MARK|11|33|于是他们回答耶稣：“我们不知道。”耶稣说：“我也不告诉你们，我仗着什么权柄做这些事。”
MARK|12|1|耶稣就用比喻对他们说：“有人开垦了一个葡萄园，四周围上篱笆，挖了一个榨酒池，盖了一座守望楼，租给园户，就出外远行去了。
MARK|12|2|到了时候，他打发一个仆人到园户那里，要向他们收葡萄园的果子。
MARK|12|3|他们拿住他，打了他，叫他空手回去。
MARK|12|4|园主再打发一个仆人到他们那里。他们打伤他的头，并且侮辱他。
MARK|12|5|园主又打发一个仆人去，他们就杀了他。以后又打发好些仆人去，有的被他们打了，有的被他们杀了。
MARK|12|6|园主还有一位，是他的爱子，最后又打发他去，说：‘他们会尊敬我的儿子。’
MARK|12|7|那些园户却彼此说：‘这是承受产业的。来，我们杀了他，产业就归我们了！’
MARK|12|8|于是他们拿住他，杀了他，把他扔出葡萄园。
MARK|12|9|这样，葡萄园主要怎么做呢？他要来除灭那些园户，将葡萄园转给别人。
MARK|12|10|‘匠人所丢弃的石头 已作了房角的头块石头。 这是主所做的， 在我们眼中看为奇妙。’ 这经文你们没有念过吗？”
MARK|12|11|
MARK|12|12|他们看出这比喻是指着他们说的，就想要捉拿他，但是惧怕众人，于是离开他走了。
MARK|12|13|后来，他们打发几个法利赛人和 希律 党人到耶稣那里，要用他自己的话陷害他。
MARK|12|14|他们来了，就对他说：“老师，我们知道你是诚实的，无论谁你都一视同仁；因为你不看人的面子，而是诚诚实实传上帝的道。纳税给凯撒合不合法？
MARK|12|15|我们该不该纳？”耶稣知道他们的虚伪，就对他们说：“你们为什么试探我？拿一个银币来给我看。”
MARK|12|16|他们就拿了来。耶稣问他们：“这像和这名号是谁的？”他们对他说：“是凯撒的。”
MARK|12|17|耶稣对他们说：“凯撒的归凯撒；上帝的归上帝。”他们对他非常惊讶。
MARK|12|18|撒都该人来见耶稣。他们说没有复活这回事，于是问耶稣：
MARK|12|19|“老师， 摩西 为我们写下这话：‘某人的哥哥若死了，撇下妻子，没有孩子，他该娶哥哥的妻子，为哥哥生子立后。’
MARK|12|20|那么，有兄弟七人，第一个娶了妻，死了，没有留下孩子。
MARK|12|21|第二个娶了她，也死了，没有留下孩子。第三个也是这样。
MARK|12|22|那七个人都没有留下孩子。最后，那妇人也死了。
MARK|12|23|在复活的时候， 她是哪一个的妻子呢？因为他们七个人都娶过她。”
MARK|12|24|耶稣说：“你们错了，不正是因为不明白圣经，也不知道上帝的大能吗？
MARK|12|25|当人从死人中复活后，也不娶也不嫁，而是像天上的天使一样。
MARK|12|26|论到死人复活，你们没有念过 摩西 书中《荆棘篇》上所记载的吗？上帝对 摩西 说：‘我是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。’
MARK|12|27|上帝不是死人的上帝，而是活人的上帝。你们是大错了。”
MARK|12|28|有一个文士来，听见他们的辩论，知道耶稣回答得好，就问他说：“诫命中哪一条是第一呢？”
MARK|12|29|耶稣回答：“第一是：‘ 以色列 啊，你要听，主—我们的上帝是独一的主。
MARK|12|30|你要尽心、尽性、尽意、尽力爱主—你的上帝。’
MARK|12|31|第二是：‘要爱邻 如己。’再没有比这两条诫命更大的了。”
MARK|12|32|那文士对耶稣说：“好，老师，你说得对，上帝是一位，除了他以外，再没有别的了；
MARK|12|33|并且尽心、尽智、尽力爱他，又爱邻如己，要比一切燔祭和祭祀好得多。”
MARK|12|34|耶稣见他回答得有智慧，就对他说：“你离上帝的国不远了。”从此以后，没有人敢再问他什么。
MARK|12|35|耶稣在圣殿里教导人，问他们说：“文士怎么说基督是 大卫 的后裔呢？
MARK|12|36|大卫 被圣灵感动，说： ‘主对我主说： 你坐在我的右边， 等我把你的仇敌放在你脚下 。’
MARK|12|37|大卫 亲自称他为主，他怎么又是 大卫 的后裔呢？”一大群的人都喜欢听他。
MARK|12|38|他在教导的时候，说：“你们要防备文士。他们好穿长袍走来走去，喜欢人们在街市上向他们问安，
MARK|12|39|又喜爱会堂里的高位，宴席上的首座。
MARK|12|40|他们侵吞寡妇的家产，假意作很长的祷告。这些人要受更重的惩罚！”
MARK|12|41|耶稣面向圣殿银库坐着，看众人怎样把钱投入银库。有好些财主投了许多钱。
MARK|12|42|有一个穷寡妇来，投了两个小文钱 ，就是一个大文钱 。
MARK|12|43|耶稣叫门徒来，对他们说：“我实在告诉你们，这穷寡妇投入银库里的比众人所投的更多。
MARK|12|44|因为，众人都是拿有余的捐献，但这寡妇，虽然自己不足，却把她一生所有的全都投进去了。”
MARK|13|1|耶稣从圣殿里出来的时候，有一个门徒对他说：“老师，请看，这是多么了不起的石头！多么了不起的建筑！”
MARK|13|2|耶稣对他说：“你看见这些宏伟的建筑吗？这里将没有一块石头会留在另一块石头上而不被拆毁的。”
MARK|13|3|耶稣在 橄榄山 上，面向圣殿坐着； 彼得 、 雅各 、 约翰 和 安得烈 私下问他说：
MARK|13|4|“请告诉我们，什么时候有这些事呢？这一切事将成的时候有什么预兆呢？”
MARK|13|5|耶稣说：“你们要谨慎，免得有人迷惑你们。
MARK|13|6|将有好些人冒我的名来，说‘我是基督’，并且要迷惑许多人。
MARK|13|7|当你们听见打仗和打仗的风声，不要惊慌；这些事必须发生，但这还不是终结。
MARK|13|8|民要攻打民，国要攻打国，多处必有地震、饥荒。这都是灾难 的起头。
MARK|13|9|但你们自己要谨慎；因为有人要把你们交给议会，并且你们在会堂里要受鞭打，又为我的缘故站在统治者和君王面前，对他们作见证。
MARK|13|10|然而，福音必须先传给万民。
MARK|13|11|有人把你们解送去受审的时候，不要事先担心说什么；到那时候，赐给你们什么话，你们就说什么；因为说话的不是你们，而是圣灵。
MARK|13|12|兄弟要把兄弟、父亲要把儿女置于死地；儿女要起来与父母为敌，害死他们；
MARK|13|13|而且你们要为我的名被众人憎恨。但坚忍到底的终必得救。”
MARK|13|14|“当你们看见那‘施行毁灭的亵渎者’站在不当站的地方（读这经的人要会意），那时，在 犹太 的，应当逃到山上；
MARK|13|15|在屋顶上的，不要下来，也不要进家里去拿东西；
MARK|13|16|在田里的，不要回去取衣裳。
MARK|13|17|在那些日子，怀孕的和奶孩子的就苦了。
MARK|13|18|你们要祈求，叫这事不在冬天发生。
MARK|13|19|因为，在那些日子必有灾难，自从上帝创造万物直到如今，从没有这样的灾难，将来也不会有。
MARK|13|20|若不是主减少那些日子，凡血肉之躯的，就没有一个能得救；但是为了他所拣选的选民，他将那些日子减少了。
MARK|13|21|那时，若有人对你们说：‘看哪，基督在这里！看哪，在那里！’你们不要信。
MARK|13|22|因为假基督和假先知将要起来，显神迹奇事，如果可能，连选民也迷惑了。
MARK|13|23|你们要谨慎！凡事我都预先告诉你们了。”
MARK|13|24|“在那些日子、那灾难以后， 太阳要变黑，月亮也不放光，
MARK|13|25|众星要从天上坠落， 天上的万象都要震动。
MARK|13|26|那时，他们要看见人子带着大能力和荣耀驾云来临。
MARK|13|27|他要差遣天使，从四方，从地极直到天边，召集他的选民。”
MARK|13|28|“你们要从无花果树学习功课：当树枝发芽长叶的时候，你们就知道夏天近了。
MARK|13|29|同样，当你们看见这些事发生，就知道那时候近了，就在门口了。
MARK|13|30|我实在告诉你们，这世代还没有过去，这一切都要发生。
MARK|13|31|天地要废去，我的话却绝不废去。”
MARK|13|32|“但那日子，那时辰，没有人知道，连天上的天使也不知道，子也不知道，惟有父知道。
MARK|13|33|你们要谨慎，要警醒 ，因为你们不知道那时刻几时来到。
MARK|13|34|这事正如一个人离家远行，授权给仆人们，分派各人的工作，又吩咐看门的警醒。
MARK|13|35|所以，你们要警醒，因为你们不知道这家的主人什么时候来，是晚上，或半夜，或鸡叫时，或早晨，
MARK|13|36|免得他忽然来到，看见你们睡着了。
MARK|13|37|我对你们所说的话，也是对众人说的：要警醒！”
MARK|14|1|过两天是逾越节，又是除酵节，祭司长和文士在想法子怎样设计捉拿耶稣，把他杀掉。
MARK|14|2|他们说：“不可在过节的日子，恐怕百姓生乱。”
MARK|14|3|耶稣在 伯大尼 痲疯病人 西门 家里坐席的时候，有一个女人拿着一玉瓶极贵的纯哪哒 香膏来，打破玉瓶，把膏浇在耶稣的头上。
MARK|14|4|有几个人心中很不高兴，说：“何必这样浪费香膏呢？
MARK|14|5|这香膏可以卖三百多个银币周济穷人。”他们就对那女人生气。
MARK|14|6|耶稣说：“由她吧！为什么难为她呢？她在我身上做的是一件美事。
MARK|14|7|因为常有穷人和你们在一起，要向他们行善，随时都可以，但是你们不常有我。
MARK|14|8|她所做的是尽她所能的；她是为了我的安葬，把香膏预先浇在我身上。
MARK|14|9|我实在告诉你们，普天之下，无论在什么地方传这福音，都要述说这女人所做的，来记念她。”
MARK|14|10|十二使徒中有一个 加略 人 犹大 ，去见祭司长，要把耶稣交给他们。
MARK|14|11|他们听见就很高兴，又应许给他银子；他就想怎样找机会把耶稣交给他们。
MARK|14|12|除酵节的第一天，就是宰逾越节羔羊的那一天，门徒对耶稣说：“你要我们到哪里去预备你吃逾越节的宴席呢？”
MARK|14|13|耶稣就打发两个门徒，对他们说：“你们进城去，会有人拿着一罐水迎面而来，你们就跟着他。
MARK|14|14|无论他进哪一家，你们就对那家的主人说：‘老师问：我的客房在哪里？我和我的门徒要在那里吃逾越节的宴席。’
MARK|14|15|他会带你们看一间摆设齐全、准备妥当的楼上大厅，你们就在那里为我们预备。”
MARK|14|16|门徒出去，进了城，所看到的正如耶稣所说的。他们就预备了逾越节的宴席。
MARK|14|17|到了晚上，耶稣和十二使徒都来了。
MARK|14|18|他们坐席，正吃的时候，耶稣说：“我实在告诉你们，你们中间有一个与我同吃的人要出卖我了。”
MARK|14|19|他们就忧愁起来，一个个地问他：“不是我吧？”
MARK|14|20|耶稣对他们说：“是十二人中的一个，就是同我蘸饼在盘子里的那个人。
MARK|14|21|人子要去了，正如经上所写有关他的；但出卖人子的人有祸了！那人没有出生倒好。”
MARK|14|22|他们吃的时候，耶稣拿起饼来，祝福了，就擘开，递给他们，说：“你们拿去，这是我的身体。”
MARK|14|23|他又拿起杯来，祝谢了，递给他们；他们都喝了。
MARK|14|24|耶稣对他们说：“这是我立约的血，为许多人流出来的。
MARK|14|25|我实在告诉你们，我不再喝这葡萄汁，直到我在上帝的国里喝新的那日子。”
MARK|14|26|他们唱了诗，就出来往 橄榄山 去。
MARK|14|27|耶稣对他们说：“你们都要跌倒，因为经上记着： ‘我要击打牧人， 羊就分散了。’，　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　　
MARK|14|28|但我复活以后，要在你们之前往 加利利 去。”
MARK|14|29|彼得 说：“虽然众人跌倒，但我不会。”
MARK|14|30|耶稣对他说：“我实在告诉你，今天夜里，鸡叫两遍 以前，你要三次不认我。”
MARK|14|31|彼得 却极力地说：“我就是必须和你同死，也绝不会不认你。”所有的门徒 都是这样说。
MARK|14|32|他们来到一个地方，名叫 客西马尼 。耶稣对门徒说：“你们坐在这里，我去祷告。”
MARK|14|33|于是他带着 彼得 、 雅各 和 约翰 同去。他惊恐起来，极其难过，
MARK|14|34|对他们说：“我心里非常忧伤，几乎要死；你们留在这里，要警醒。”
MARK|14|35|他就稍往前走，俯伏在地，祷告说，如果可能，就叫那时候离开他。
MARK|14|36|他说：“阿爸，父啊！在你凡事都能；求你将这杯撤去。然而，不是照我所愿的，而是照你所愿的。”
MARK|14|37|耶稣回来，见他们睡着了，就对 彼得 说：“ 西门 ，你睡着了吗？不能警醒一小时吗？
MARK|14|38|总要警醒祷告，免得陷入试探。你们心灵固然愿意，肉体却软弱了。”
MARK|14|39|耶稣又去祷告，说的话跟先前一样。
MARK|14|40|他又来，见他们睡着了，因为他们的眼睛很困倦；他们也不知道怎么回答他。
MARK|14|41|他第三次来对他们说：“现在你们仍在睡觉安歇吗？够了，时候到了。看哪，人子被出卖在罪人手里了。
MARK|14|42|起来，我们走吧！看哪，那出卖我的人快来了。”
MARK|14|43|耶稣还在说话的时候，忽然十二使徒之一的 犹大 来了，还有一群人带着刀棒，从祭司长、文士和长老那里跟他同来。
MARK|14|44|那出卖耶稣的人曾给他们一个暗号，说：“我亲谁，谁就是。你们把他抓住，稳妥地带走。”
MARK|14|45|犹大 来了，随即到耶稣跟前，说：“拉比”，就跟他亲吻。
MARK|14|46|他们就下手抓住他。
MARK|14|47|旁边站着的人，有一个拔出刀来，把大祭司的仆人砍了一刀，削掉了他一只耳朵。
MARK|14|48|耶稣回应他们说：“你们带着刀棒出来拿我，如同拿强盗吗？
MARK|14|49|我天天教导人，同你们在殿里，你们并没有抓我。但这是要应验经上的话。”
MARK|14|50|门徒都离开他，逃走了。
MARK|14|51|有一个青年光着身子，只披一块麻布，跟随耶稣，众人就抓住他。
MARK|14|52|他却丢下麻布，赤身逃走了。
MARK|14|53|他们把耶稣带到大祭司那里，又有众祭司长、长老和文士都来一同聚集。
MARK|14|54|彼得 远远地跟着耶稣，直到进了大祭司的院子，和警卫一同坐在火边取暖。
MARK|14|55|祭司长和全议会寻找见证控告耶稣，要处死他，却找不到实据。
MARK|14|56|因为有好些人作假见证告他，他们的见证又各不相符。
MARK|14|57|又有几个人站起来，作假见证告他说：
MARK|14|58|“我们听见他说：‘我要拆毁这人手所造的殿，三日内另造一座不是人手所造的。’”
MARK|14|59|就是这样，他们的见证还是不相符。
MARK|14|60|大祭司起来站在中间，问耶稣说：“这些人作证告你的事，你什么都不回答吗？”
MARK|14|61|耶稣却不言语，一句也不回答。大祭司又问他：“你是不是基督，那当称颂者的儿子？”
MARK|14|62|耶稣说：“我是。 你们要看见人子 坐在那权能者的右边， 驾着天上的云来临。”
MARK|14|63|大祭司就撕裂衣服，说：“我们何必再要证人呢？
MARK|14|64|你们已经听见他这亵渎的话了。你们的决定如何？”他们都判定他该处死。
MARK|14|65|于是有人开始向他吐唾沫，又蒙着他的脸，用拳头打他，对他说：“你说预言吧！”警卫把他拉过来，打他耳光。
MARK|14|66|彼得 在下边院子里，大祭司的一个使女来了，
MARK|14|67|见 彼得 取暖，就看着他，说：“你素来也是同 拿撒勒 人耶稣一起的。”
MARK|14|68|彼得 却不承认，说：“我不知道，也不明白你说的是什么！”于是他出来，到了前院，鸡就叫了 。
MARK|14|69|那使女看见他，又对旁边站着的人说：“这个人也是他们一伙的。”
MARK|14|70|彼得 又不承认。过了不久，旁边站着的人又对 彼得 说：“你真是他们一伙的，因为你也是 加利利 人。”
MARK|14|71|彼得 就赌咒发誓说：“我不认得你们说的这个人。”
MARK|14|72|立刻，鸡叫了第二遍。 彼得 想起耶稣对他所说的话：“鸡叫两遍以前，你要三次不认我。”他就忍不住哭了。
MARK|15|1|一到早晨，众祭司长、长老、文士，和全议会的人大家商议，就把耶稣绑着，解去，交给 彼拉多 。
MARK|15|2|彼拉多 问他：“你是 犹太 人的王吗？”耶稣回答：“是你说的。”
MARK|15|3|祭司长们告他许多的事。
MARK|15|4|彼拉多 又问他：“你看，他们告你这么多的事，你什么都不回答吗？”
MARK|15|5|耶稣仍不回答，以致 彼拉多 觉得惊讶。
MARK|15|6|每逢这节期， 彼拉多 照众人所求的，释放一个囚犯给他们。
MARK|15|7|有一个人名叫 巴拉巴 ，和作乱的人监禁在一起。他们作乱的时候曾杀过人。
MARK|15|8|众人上去求 彼拉多 照常例给他们办理。
MARK|15|9|彼拉多 说：“你们要我释放 犹太 人的王给你们吗？”
MARK|15|10|他原知道祭司长们是因嫉妒才把耶稣解了来。
MARK|15|11|但是祭司长们煽动众人，宁可要他释放 巴拉巴 给他们。
MARK|15|12|彼拉多 又说：“那么，你们称为 犹太 人的王的 ，要 我怎么办他呢？”
MARK|15|13|他们又再喊着：“把他钉十字架！”
MARK|15|14|彼拉多 说：“为什么？他做了什么恶事呢？”他们更加喊着：“把他钉十字架！”
MARK|15|15|彼拉多 要讨好众人，就释放 巴拉巴 给他们，把耶稣鞭打后交给人钉十字架。
MARK|15|16|士兵把耶稣带进总督府的庭院里，叫齐了全营的兵。
MARK|15|17|他们给他穿上紫袍，又用荆棘编了冠冕给他戴上，
MARK|15|18|然后向他致敬，说：“万岁， 犹太 人的王！”
MARK|15|19|他们又拿一根芦苇秆打他的头，向他吐唾沫，屈膝拜他。
MARK|15|20|他们戏弄完了，就给他脱了紫袍，又穿上他自己的衣服，带他出去，要把他钉十字架。
MARK|15|21|有一个 古利奈 人 西门 ，就是 亚历山大 和 鲁孚 的父亲，从乡下来，经过那地方，他们就强迫他同去，好背耶稣的十字架。
MARK|15|22|他们带耶稣到了一个地方叫 各各他 （翻出来就是“髑髅地”），
MARK|15|23|拿没药调和的酒给耶稣，他却不受。
MARK|15|24|于是他们把他钉在十字架上，抽签分他的衣服，看谁得什么。
MARK|15|25|他们把他钉十字架的时候是上午九点钟。
MARK|15|26|罪状牌上写的是：“ 犹太 人的王。”
MARK|15|27|他们又把两个强盗和他同钉十字架，一个在右边，一个在左边。
MARK|15|28|
MARK|15|29|从那里经过的人讥笑他，摇着头，说：“哼！你这拆毁殿、三日又建造起来的，
MARK|15|30|救救你自己，从十字架上下来呀！”
MARK|15|31|众祭司长和文士也这样嘲笑他，彼此说：“他救了别人，不能救自己。
MARK|15|32|以色列 的王基督，现在从十字架上下来，好让我们看见就信了呀！”那和他同钉的人也讥讽他。
MARK|15|33|到了正午，全地都黑暗了，直到下午三点钟。
MARK|15|34|下午三点钟的时候，耶稣大声呼喊：“以罗伊！以罗伊！拉马撒巴各大尼？”（翻出来就是：我的上帝！我的上帝！为什么离弃我？）
MARK|15|35|旁边站着的人，有的听见就说：“看哪，他叫 以利亚 呢！”
MARK|15|36|有一个人跑去，把海绵蘸满了醋，绑在芦苇秆上，送给他喝，说：“且等着，看 以利亚 会不会来把他放下来。”
MARK|15|37|耶稣大喊一声，气就断了。
MARK|15|38|殿的幔子从上到下裂为两半。
MARK|15|39|对面站着的百夫长看见耶稣这样断气 ，就说：“这人真是上帝的儿子！”
MARK|15|40|还有些妇女远远地观看，其中有 抹大拉 的 马利亚 ，又有小 雅各 和 约西 的母亲 马利亚 ，并有 撒罗米 ，
MARK|15|41|就是耶稣在 加利利 的时候，跟随他、服事他的那些人，还有同耶稣上 耶路撒冷 的好些妇女。
MARK|15|42|到了晚上，因为这是预备日，就是安息日的前一日，
MARK|15|43|有 亚利马太 的 约瑟 前来，他是尊贵的议员，也是盼望着上帝国的，他放胆进去见 彼拉多 ，请求要耶稣的身体。
MARK|15|44|彼拉多 诧异耶稣已经死了，就叫百夫长来，问他耶稣是不是死了很久；
MARK|15|45|既从百夫长得知实情，就把耶稣的身体赐给 约瑟 。
MARK|15|46|约瑟 买了细麻布，把耶稣取下来，用细麻布裹好，安放在岩石中凿出来的墓穴里，又滚来一块石头挡住墓门。
MARK|15|47|抹大拉 的 马利亚 和 约西 的母亲 马利亚 都看见安放他的地方。
MARK|16|1|过了安息日， 抹大拉 的 马利亚 、 雅各 的母亲 马利亚 ，和 撒罗米 ，买了香料，要去膏耶稣的身体。
MARK|16|2|七日的第一日清早，太阳出来后，她们来到坟墓那里，
MARK|16|3|彼此说：“谁要替我们把石头从墓门滚开呢？”
MARK|16|4|她们抬头一看，看见石头已经滚开了，原来那石头很大。
MARK|16|5|她们进了坟墓，看见一个年轻人坐在右边，穿着白袍，就很惊奇。
MARK|16|6|那年轻人对她们说：“不要惊慌！你们寻找那钉十字架的 拿撒勒 人耶稣，他已经复活了，不在这里。来看安放他的地方。
MARK|16|7|你们去，对他的门徒和 彼得 说：‘他要比你们先到 加利利 去，在那里你们会看见他，正如他从前所告诉你们的。’”
MARK|16|8|于是她们出来，从坟墓那里逃走，又发抖又惊讶，什么也没有告诉人，因为她们害怕。 〔
MARK|16|9|凡耶稣所吩咐的，她们简洁地告诉 彼得 和他周围的人。这些事以后，耶稣亲自藉着他的门徒，从东到西，把那神圣、不朽、永远拯救的福音传出去。阿们！〕 〔 在七日的第一日清早，耶稣复活了，先向 抹大拉 的 马利亚 显现；耶稣曾从她身上赶出七个鬼。
MARK|16|10|她去告诉那向来跟随耶稣的人；那时他们正哀恸哭泣。
MARK|16|11|他们听见耶稣活了，被 马利亚 看见，可是不信。〕 〔
MARK|16|12|这些事以后，门徒中有两个人往乡下去；正走着的时候，耶稣以另一种形像向他们显现。
MARK|16|13|他们去告诉其余的门徒，那些门徒还是不信。〕 〔
MARK|16|14|后来十一使徒坐席的时候，耶稣向他们显现，责备他们不信，心里刚硬，因为他们不信那些在他复活以后看见他的人。
MARK|16|15|他又对他们说：“你们往普天下去，传福音给万民 听。
MARK|16|16|信而受洗的必然得救，不信的必被定罪。
MARK|16|17|信的人将有神迹随着他们：就是奉我的名赶鬼；说新方言；
MARK|16|18|手 能拿蛇；若喝了什么毒物，也不会受害；手按病人，病人就好了。”〕 〔
MARK|16|19|主耶稣 和他们说完了话以后，被接到天上，坐在上帝的右边。
MARK|16|20|门徒出去，到处传福音。主和他们同工，藉着伴随的神迹证实所传的道。 〕
LUKE|1|1|提阿非罗 大人哪，有好些人提笔作书，述说在我们中间所实现的事，是照传道的人从起初亲眼看见又传给我们的。这些事我从起头都详细考察了，我也想按着次序写给你，
LUKE|1|2|
LUKE|1|3|
LUKE|1|4|要让你知道所学的道都是确实的。
LUKE|1|5|在 希律 作 犹太 王的时候， 亚比雅 班里有一个祭司，名叫 撒迦利亚 ；他妻子是 亚伦 的后代，名叫 伊利莎白 。
LUKE|1|6|他们两人在上帝面前都是义人，遵行主的一切诫命和条例，没有可指责的。
LUKE|1|7|只是他们没有孩子，因为 伊利莎白 不生育，两个人又年纪老迈了。
LUKE|1|8|撒迦利亚 按班次在上帝面前执行祭司的职务，
LUKE|1|9|照祭司的规矩抽签，进到主的殿里烧香。
LUKE|1|10|烧香的时候，众百姓在外面祷告。
LUKE|1|11|有主的一个使者站在香坛的右边，向他显现。
LUKE|1|12|撒迦利亚 看见，就惊慌害怕。
LUKE|1|13|天使对他说：“ 撒迦利亚 ，不要害怕，因为你的祈祷已经被听见了。你的妻子 伊利莎白 要给你生一个儿子，你要给他起名叫 约翰 。
LUKE|1|14|你必欢喜快乐；有许多人因他出世也必喜乐。
LUKE|1|15|他在主面前将要为大，淡酒烈酒都不喝，从母腹里就被圣灵充满。
LUKE|1|16|他要使许多 以色列 人回转，归于主—他们的上帝。
LUKE|1|17|他将有 以利亚 的精神和能力，走在主的前面，叫父亲的心转向儿女，叫悖逆的人转向义人的智慧，又为主预备迎接他的百姓。”
LUKE|1|18|撒迦利亚 对天使说：“我怎么能知道这事呢？我已经老了，我的妻子也年纪老迈了。”
LUKE|1|19|天使回答他说：“我是站在上帝面前的 加百列 ，奉差遣来对你说话，把这好信息报给你。
LUKE|1|20|到了时候，这些话必然应验；只因你不信我的话，你会成为哑巴，不能说话，直到这些事实现的日子。”
LUKE|1|21|百姓等候 撒迦利亚 ，诧异他在圣所里迟延那么久。
LUKE|1|22|到他出来，却不能和他们说话，他们就知道他在圣所里见了异象；他直向他们打手势，因为他成了哑巴。
LUKE|1|23|他供职的日子一满，就回家去了。
LUKE|1|24|这些日子以后，他的妻子 伊利莎白 就怀孕，隐藏了五个月；
LUKE|1|25|她说：“主在眷顾我的日子，这样看顾我，要除掉我在人前的羞耻。”
LUKE|1|26|到了第六个月，天使 加百列 奉上帝的差遣往 加利利 的一座城去，这城名叫 拿撒勒 ，
LUKE|1|27|到一个童女那里，她已经许配 大卫 家的一个人，名叫 约瑟 ；童女的名字叫 马利亚 。
LUKE|1|28|天使进去，对她说：“蒙大恩的女子，你好，主和你同在！”
LUKE|1|29|马利亚 因这话就很惊慌，又反覆思考这样问候是什么意思。
LUKE|1|30|天使对她说： “ 马利亚 ，不要怕，你在上帝面前已经蒙恩了。
LUKE|1|31|你要怀孕生子，要给他起名叫耶稣。
LUKE|1|32|他将要为大，称为至高者的儿子； 主上帝要把他祖先 大卫 的王位给他。
LUKE|1|33|他要作 雅各 家的王，直到永远； 他的国没有穷尽。”
LUKE|1|34|马利亚 对天使说：“我没有出嫁，怎么会有这事呢？”
LUKE|1|35|天使回答她说： “圣灵要临到你身上； 至高者的能力要庇荫你， 因此，那要出生的圣者要称为上帝的儿子 。
LUKE|1|36|况且，你的亲戚 伊利莎白 ，就是那素来称为不生育的，在年老的时候也怀了男胎，现在怀孕六个月了。
LUKE|1|37|因为，出于上帝的话，没有一句不带能力的。”
LUKE|1|38|马利亚 说：“我是主的使女，愿意照你的话实现在我身上。”于是天使离开她去了。
LUKE|1|39|在那些日子， 马利亚 起身，急忙前往山区，来到 犹大 的一座城，
LUKE|1|40|进了 撒迦利亚 的家，向 伊利莎白 问安。
LUKE|1|41|伊利莎白 一听到 马利亚 问安，所怀的胎就在腹里跳动。 伊利莎白 被圣灵充满，
LUKE|1|42|高声喊着说： “你在妇女中是有福的！ 你所怀的胎也是有福的！
LUKE|1|43|我主的母亲到我这里来，为何这事临到我呢？
LUKE|1|44|因为你问安的声音一入我耳，我腹里的胎就欢喜跳动。
LUKE|1|45|这相信的女子是有福的！因为主对她所说的话都要应验。”
LUKE|1|46|马利亚 说： “我心尊主为大；
LUKE|1|47|我灵以上帝我的救主为乐；
LUKE|1|48|因为他顾念他使女的卑微； 从今以后，万代要称我有福。
LUKE|1|49|因为那有权能的为我做了大事； 他的名是圣的。
LUKE|1|50|他怜悯敬畏他的人， 直到世世代代。
LUKE|1|51|他用膀臂施展大能； 他赶散心里妄想的狂傲人。
LUKE|1|52|他叫有权柄的失位， 叫卑贱的升高。
LUKE|1|53|他叫饥饿的饱餐美食， 叫富足的空手回去。
LUKE|1|54|他扶助了他的仆人 以色列 ，不忘记施怜悯，
LUKE|1|55|正如他对我们的列祖说过， ‘怜悯 亚伯拉罕 和他的后裔，直到永远。’”
LUKE|1|56|马利亚 和 伊利莎白 同住，约有三个月，然后回家去了。
LUKE|1|57|伊利莎白 的产期到了，生了一个儿子。
LUKE|1|58|邻里亲属听见主向她大施怜悯，就和她一同欢乐。
LUKE|1|59|到了第八日，他们来给孩子行割礼，并要照他父亲的名字叫他 撒迦利亚 。
LUKE|1|60|他母亲回应说：“不！要叫他 约翰 。”
LUKE|1|61|他们对她说：“你亲族中没有叫这名字的。”
LUKE|1|62|他们就向他父亲打手势，问他这孩子要叫什么名字。
LUKE|1|63|他要了一块写字的板，写上：“他的名字是 约翰 。”他们就都惊讶。
LUKE|1|64|撒迦利亚 的口立刻开了，舌头也松了，就开始说话称颂上帝。
LUKE|1|65|周围居住的人都惧怕；这一切的事就传遍了 犹太 山区。
LUKE|1|66|凡听见的人都把这事放在心里，他们说：“这个孩子将来会怎么样呢？”因为有主的手与他同在。
LUKE|1|67|他父亲 撒迦利亚 被圣灵充满，就预言说：
LUKE|1|68|“主— 以色列 的上帝是应当称颂的！ 因他眷顾他的百姓，为他们施行救赎，
LUKE|1|69|在他仆人 大卫 家中， 为我们兴起了拯救的角，
LUKE|1|70|正如主藉着古时候圣先知的口所说的，
LUKE|1|71|‘他拯救我们脱离仇敌， 脱离一切恨我们之人的手。
LUKE|1|72|他向我们列祖施怜悯， 记得他的圣约，
LUKE|1|73|就是他对我们祖宗 亚伯拉罕 所起的誓，
LUKE|1|74|叫我们既从仇敌手中被救出来， 就可以终身在他面前， 无所惧怕地用圣洁和公义事奉他。
LUKE|1|75|
LUKE|1|76|孩子啊，你要称为至高者的先知； 因为你要走在主的前面，为他预备道路，
LUKE|1|77|叫他的百姓因罪得赦， 认识救恩；
LUKE|1|78|因我们上帝怜悯的心肠， 叫清晨的日光从高天临到我们，
LUKE|1|79|要照亮坐在黑暗中死荫里的人， 把我们的脚引到和平的路上。’”
LUKE|1|80|这孩子渐渐长大，心灵坚强，住在旷野，直到他在 以色列 人面前公开出现的日子。
LUKE|2|1|在那些日子，凯撒 奥古斯都 降旨，叫全国人民都登记户籍。
LUKE|2|2|这第一次登记户籍是在 居里扭 作 叙利亚 总督的时候行的。
LUKE|2|3|众人各归各城，办理登记。
LUKE|2|4|约瑟 也从 加利利 的 拿撒勒城 上 犹太 去，到了 大卫 的城名叫 伯利恒 ，因为他是 大卫 家族的人，
LUKE|2|5|要和他所聘之妻 马利亚 一同登记户籍。那时 马利亚 已经怀孕。
LUKE|2|6|他们在那里的时候， 马利亚 的产期到了，
LUKE|2|7|就生了头胎的儿子，用布包起来，放在马槽里，因为客店里没有地方。
LUKE|2|8|在 伯利恒 的野外有牧羊人，夜间值班看守羊群。
LUKE|2|9|有主的一个使者站在他们旁边，主的荣光四面照着他们，牧羊人就很惧怕。
LUKE|2|10|那天使对他们说：“不要惧怕！看哪！因为我报给你们大喜的信息，是关乎万民的：
LUKE|2|11|因今天在 大卫 的城里，为你们生了救主，就是主基督。
LUKE|2|12|你们要看见一个婴孩，包着布，卧在马槽里，那就是给你们的记号。”
LUKE|2|13|忽然，有一大队天兵同那天使赞美上帝说：
LUKE|2|14|“在至高之处荣耀归与上帝！ 在地上平安归与他所喜悦的人！”
LUKE|2|15|众天使离开他们，升天去了。牧羊人彼此说：“我们往 伯利恒 去，看看所成的事，就是主所告诉我们的。”
LUKE|2|16|他们急忙去了，找到 马利亚 和 约瑟 ，还有那婴孩卧在马槽里。
LUKE|2|17|他们看见，就把天使论这孩子的话传开了。
LUKE|2|18|听见的人都诧异牧羊人对他们所说的话。
LUKE|2|19|马利亚 却把这一切的事存在心里，反覆思考。
LUKE|2|20|牧羊人回去了，因所听见所看见的一切事，正如天使向他们所说的，就归荣耀于上帝，赞美他。
LUKE|2|21|满了八天，他们就给孩子行割礼，又给他起名叫耶稣；这是他还没有在母腹里成胎以前天使所起的名。
LUKE|2|22|按 摩西 律法满了洁净的日子，他们就带着孩子上 耶路撒冷 去，要把他献给主。
LUKE|2|23|正如主的律法上所记：“凡头生的男子必归主为圣”；
LUKE|2|24|又要照主的律法上所说，用一对斑鸠，或用两只雏鸽献祭。
LUKE|2|25|那时，在 耶路撒冷 有一个人，名叫 西面 ；这人又公义又虔诚，素常盼望 以色列 的安慰者来到，又有圣灵在他身上。
LUKE|2|26|他得了圣灵的启示，知道自己未死以前必看见主所立的基督。
LUKE|2|27|他受了圣灵的感动，进入圣殿，正遇见耶稣的父母抱着孩子进来，要照律法的规矩而行。
LUKE|2|28|西面 就把他抱过来，称颂上帝说：
LUKE|2|29|“主啊，如今可以照你的话， 容你的仆人安然去世；
LUKE|2|30|因为我的眼睛已经看见你的救恩，
LUKE|2|31|就是你在万民面前所预备的：
LUKE|2|32|是启示外邦人的光， 是你民 以色列 的荣耀。”
LUKE|2|33|孩子的父母因论耶稣的这些话就惊讶。
LUKE|2|34|西面 给他们祝福，又对孩子的母亲 马利亚 说：“这孩子被立，是要叫 以色列 中许多人跌倒，许多人兴起；又要成为毁谤的对象，
LUKE|2|35|叫许多人心里的意念显露出来；你自己的心也要被剑刺透。”
LUKE|2|36|又有位女先知，名叫 亚拿 ，是 亚设 支派 法内力 的女儿，年纪已经老迈，从童女出嫁，同丈夫住了七年，
LUKE|2|37|就寡居了，现在已经八十四岁 。她不离开圣殿，禁食祈求，昼夜事奉上帝。
LUKE|2|38|正当那时，她进前来感谢上帝，对一切盼望 耶路撒冷 得救赎的人讲论这孩子的事。
LUKE|2|39|约瑟 和 马利亚 照主的律法办完了一切的事，就回 加利利 ，到自己的城 拿撒勒 去了。
LUKE|2|40|孩子渐渐长大，强健起来，充满智慧，又有上帝的恩典在他身上。
LUKE|2|41|每年逾越节，他父母都上 耶路撒冷 去。
LUKE|2|42|当他十二岁的时候，他们按着过节的规矩上去。
LUKE|2|43|守满了节期，他们回去，孩童耶稣仍旧在 耶路撒冷 。他的父母并不知道，
LUKE|2|44|以为他在同行的人中间，走了一天的路程才在亲属和熟悉的人中找他，
LUKE|2|45|既找不着，就回 耶路撒冷 去找他。
LUKE|2|46|过了三天，他们发现他在圣殿里，坐在教师中间，一面听，一面问。
LUKE|2|47|凡听见他的人都对他的聪明和应对感到惊奇。
LUKE|2|48|他父母看见就很惊奇。他母亲对他说：“我儿啊，为什么对我们这样做呢？看哪，你父亲和我很焦急，到处找你！”
LUKE|2|49|耶稣对他们说：“为什么找我呢？难道你们不知道我应当在我父的家里吗？ ”
LUKE|2|50|他所说的这话，他们不明白。
LUKE|2|51|他就同他们下去，回到 拿撒勒 ，并且顺从他们。他母亲把这一切的事都存在心里。
LUKE|2|52|耶稣的智慧和身量 ，并上帝和人喜爱他的心，都一齐增长。
LUKE|3|1|凯撒 提庇留 在位第十五年， 本丢．彼拉多 作 犹太 总督， 希律 作 加利利 分封的王，他兄弟 腓力 作 以土利亚 和 特拉可尼 地区分封的王， 吕撒聂 作 亚比利尼 分封的王，
LUKE|3|2|亚那 和 该亚法 作大祭司。那时， 撒迦利亚 的儿子 约翰 在旷野里，上帝的话临到他。
LUKE|3|3|他就走遍 约旦河 一带地方，宣讲悔改的洗礼，使罪得赦。
LUKE|3|4|正如 以赛亚 先知书上所记的话： “在旷野有声音呼喊着： 预备主的道， 修直他的路！
LUKE|3|5|一切山洼都要填满； 大小山冈都要削平！ 弯弯曲曲的地方要改为笔直； 高高低低的道路要改为平坦！
LUKE|3|6|凡血肉之躯的，都要看见上帝的救恩！”
LUKE|3|7|约翰 对那出来要受他洗的众人说：“毒蛇的孽种啊，谁指示你们逃避那将要来的愤怒呢？
LUKE|3|8|你们要结出果子来，和悔改的心相称。不要自己心里说：‘我们有 亚伯拉罕 为祖宗。’我告诉你们，上帝能从这些石头中给 亚伯拉罕 兴起子孙来。
LUKE|3|9|现在斧子已经放在树根上，凡不结好果子的树就砍下来，丢在火里。”
LUKE|3|10|众人问他：“这样，我们该做什么呢？”
LUKE|3|11|约翰 回答：“有两件衣裳的，就分给那没有的；有食物的，也该这样做。”
LUKE|3|12|也有税吏来要受洗，对他说：“老师，我们该做什么呢？”
LUKE|3|13|约翰 对他们说：“除了规定的数目，不要多收。”
LUKE|3|14|也有士兵问他说：“我们该做什么呢？” 约翰 说：“不要勒索任何人，也不要敲诈人；自己有粮饷就该知足。”
LUKE|3|15|百姓期待基督的来临；他们心里猜测，或许 约翰 是基督。
LUKE|3|16|约翰 对众人说：“我是用水给你们施洗，但有一位能力比我更大的要来，我就是给他解鞋带也不配。他要用圣灵与火给你们施洗。
LUKE|3|17|他手里拿着簸箕，要扬净他的谷物，把麦子收在仓里，把糠用不灭的火烧尽。”
LUKE|3|18|约翰 又用许多别的话劝百姓，向他们传福音。
LUKE|3|19|希律 分封王，因他兄弟之妻 希罗底 的缘故，并因他所做的一切恶事，受了 约翰 的责备。
LUKE|3|20|希律 在一切事上又添了这一件，就是把 约翰 收在监里。
LUKE|3|21|众百姓都受了洗，耶稣也受了洗。他正祷告的时候，天开了，
LUKE|3|22|圣灵降在他身上，形状仿佛鸽子；又有声音从天上来，说：“你是我的爱子，我喜爱你。”
LUKE|3|23|耶稣开始传道，年纪约有三十岁。依人看来，他是 约瑟 的儿子， 约瑟 是 希里 的儿子，
LUKE|3|24|希里 是 玛塔 的儿子， 玛塔 是 利未 的儿子， 利未 是 麦基 的儿子， 麦基 是 雅拿 的儿子， 雅拿 是 约瑟 的儿子，
LUKE|3|25|约瑟 是 玛他提亚 的儿子， 玛他提亚 是 亚摩斯 的儿子， 亚摩斯 是 拿鸿 的儿子， 拿鸿 是 以斯利 的儿子， 以斯利 是 拿该 的儿子，
LUKE|3|26|拿该 是 玛押 的儿子， 玛押 是 玛他提亚 的儿子， 玛他提亚 是 西美 的儿子， 西美 是 约瑟 的儿子， 约瑟 是 犹大 的儿子， 犹大 是 约亚拿 的儿子，
LUKE|3|27|约亚拿 是 利撒 的儿子， 利撒 是 所罗巴伯 的儿子， 所罗巴伯 是 撒拉铁 的儿子， 撒拉铁 是 尼利 的儿子， 尼利 是 麦基 的儿子，
LUKE|3|28|麦基 是 亚底 的儿子， 亚底 是 哥桑 的儿子， 哥桑 是 以摩当 的儿子， 以摩当 是 珥 的儿子， 珥 是 约细 的儿子，
LUKE|3|29|约细 是 以利以谢 的儿子， 以利以谢 是 约令 的儿子， 约令 是 玛塔 的儿子， 玛塔 是 利未 的儿子，
LUKE|3|30|利未 是 西缅 的儿子， 西缅 是 犹大 的儿子， 犹大 是 约瑟 的儿子， 约瑟 是 约南 的儿子， 约南 是 以利亚敬 的儿子，
LUKE|3|31|以利亚敬 是 米利亚 的儿子， 米利亚 是 买南 的儿子， 买南 是 玛达他 的儿子， 玛达他 是 拿单 的儿子， 拿单 是 大卫 的儿子，
LUKE|3|32|大卫 是 耶西 的儿子， 耶西 是 俄备得 的儿子， 俄备得 是 波阿斯 的儿子， 波阿斯 是 沙拉 的儿子， 沙拉 是 拿顺 的儿子 ，
LUKE|3|33|拿顺 是 亚米拿达 的儿子， 亚米拿达 是 亚民 的儿子， 亚民 是 亚尼 的儿子， 亚尼 是 希斯仑 的儿子 ， 希斯仑 是 法勒斯 的儿子， 法勒斯 是 犹大 的儿子，
LUKE|3|34|犹大 是 雅各 的儿子， 雅各 是 以撒 的儿子， 以撒 是 亚伯拉罕 的儿子， 亚伯拉罕 是 他拉 的儿子， 他拉 是 拿鹤 的儿子，
LUKE|3|35|拿鹤 是 西鹿 的儿子， 西鹿 是 拉吴 的儿子， 拉吴 是 法勒 的儿子， 法勒 是 希伯 的儿子， 希伯 是 沙拉 的儿子，
LUKE|3|36|沙拉 是 该南 的儿子， 该南 是 亚法撒 的儿子， 亚法撒 是 闪 的儿子， 闪 是 挪亚 的儿子， 挪亚 是 拉麦 的儿子，
LUKE|3|37|拉麦 是 玛土撒拉 的儿子， 玛土撒拉 是 以诺 的儿子， 以诺 是 雅列 的儿子， 雅列 是 玛勒列 的儿子， 玛勒列 是 该南 的儿子， 该南 是 以挪士 的儿子，
LUKE|3|38|以挪士 是 塞特 的儿子， 塞特 是 亚当 的儿子， 亚当 是上帝的儿子。
LUKE|4|1|耶稣满有圣灵，从 约旦河 回来，圣灵把他引到旷野，
LUKE|4|2|四十天受魔鬼的试探。在那些日子，他没有吃什么，日子满了，他饿了。
LUKE|4|3|魔鬼对他说：“你若是上帝的儿子，叫这块石头变成食物吧。”
LUKE|4|4|耶稣回答：“经上记着： ‘人活着，不是单靠食物。 ’”
LUKE|4|5|魔鬼又领他上了高山，霎时间把天下万国都指给他看，
LUKE|4|6|对他说：“这一切权柄和荣华我都要给你，因为这原是交给我的，我愿意给谁就给谁。
LUKE|4|7|你若在我面前下拜，这一切都归你。”
LUKE|4|8|耶稣回答他说：“经上记着： ‘要拜主—你的上帝， 惟独事奉他。’”
LUKE|4|9|魔鬼又领他到 耶路撒冷 去，叫他站在圣殿顶上，对他说：“你若是上帝的儿子，从这里跳下去！
LUKE|4|10|因为经上记着： ‘主要为你命令他的使者保护你；
LUKE|4|11|他们要用手托住你， 免得你的脚碰在石头上。’”
LUKE|4|12|耶稣回答他说：“经上说：‘不可试探主—你的上帝。’”
LUKE|4|13|魔鬼用完了各样的试探，就离开耶稣，再等时机。
LUKE|4|14|耶稣带着圣灵的能力回到 加利利 ，他的名声传遍了四方。
LUKE|4|15|他在各会堂里教导人，众人都称赞他。
LUKE|4|16|耶稣来到 拿撒勒 ，就是他长大的地方。在安息日，照他素常的规矩进了会堂，站起来要念圣经。
LUKE|4|17|有人把 以赛亚 先知的书交给他，他就打开，找到一处写着：
LUKE|4|18|“主的灵在我身上， 因为他用膏膏我， 叫我传福音给贫穷的人； 差遣我宣告： 被掳的得释放， 失明的得看见， 受压迫的得自由，
LUKE|4|19|宣告上帝悦纳人的禧年。”
LUKE|4|20|于是他把书卷起来，交还给管理人，就坐下。会堂里的人都定睛看他。
LUKE|4|21|耶稣对他们说：“你们听见的这段经文，今天已经应验了。”
LUKE|4|22|众人都称赞他，并对他口中所出的恩言感到惊讶；他们说：“这不是 约瑟 的儿子吗？”
LUKE|4|23|耶稣对他们说：“你们一定会用这俗语向我说：‘医生，你医治自己吧！我们听见你在 迦百农 所做的事，也该在你自己的家乡做吧。’”
LUKE|4|24|他又说：“我实在告诉你们，没有先知在自己家乡被人接纳的。
LUKE|4|25|我对你们说实话，在 以利亚 的时候，天闭塞了三年六个月，遍地有大饥荒，那时， 以色列 中有许多寡妇，
LUKE|4|26|以利亚 并没有奉差往她们中任何一个人那里去，只奉差往 西顿 的 撒勒法 一个寡妇那里去。
LUKE|4|27|在 以利沙 先知的时候， 以色列 中有许多痲疯病人，但除了 叙利亚 的 乃缦 ，没有一个得洁净的。”
LUKE|4|28|会堂里的人听见这些话，都怒气填胸，
LUKE|4|29|就起来赶他出城。他们的城造在山上；他们带他到山崖，要把他推下去。
LUKE|4|30|他却从他们中间穿过去，走了。
LUKE|4|31|耶稣下到 迦百农 ，就是 加利利 的一座城，在安息日教导众人。
LUKE|4|32|他们对他的教导感到很惊奇，因为他的话里有权柄。
LUKE|4|33|在会堂里有一个人，被污鬼的灵附着，大声喊叫说：
LUKE|4|34|“唉！ 拿撒勒 人耶稣，你为什么干扰我们？你来消灭我们吗？我知道你是谁，你是上帝的圣者。”
LUKE|4|35|耶稣斥责他说：“不要作声，从这人身上出来吧！”鬼把那人摔倒在众人中间，就出来了，却没有伤害他。
LUKE|4|36|众人都惊讶，彼此对问：“这是什么道理呢？因为他用权柄能力命令污灵，污灵就出来。”
LUKE|4|37|于是耶稣的名声传遍了周围各地。
LUKE|4|38|耶稣出了会堂，进了 西门 的家。 西门 的岳母在发高烧，有些人为她求耶稣。
LUKE|4|39|耶稣站在她旁边，斥责那高烧，烧就退了。她立刻起来服事他们。
LUKE|4|40|日落的时候，凡有病人的，不论害什么病，都带到耶稣那里。耶稣给他们每一个人按手，治好他们。
LUKE|4|41|又有鬼从好些人身上出来，喊着说：“你是上帝的儿子！”耶稣斥责他们，不许他们说话，因为他们知道他是基督。
LUKE|4|42|天亮的时候，耶稣出来，走到荒野的地方。众人去找他，到了他那里，要留住他，不让他离开他们。
LUKE|4|43|但耶稣对他们说：“我也必须在别的城传上帝国的福音，因我奉差原是为此。”
LUKE|4|44|于是耶稣在 犹太 的各会堂传道。
LUKE|5|1|耶稣站在 革尼撒勒 湖边，众人拥挤他，要听上帝的道。
LUKE|5|2|他见有两只船靠在湖边，打鱼的人却离开船，洗网去了。
LUKE|5|3|有一只船是 西门 的，耶稣就上去，请他把船撑开，稍微离岸，就坐下，在船上教导众人。
LUKE|5|4|他讲完了，对 西门 说：“把船开到水深的地方下网打鱼。”
LUKE|5|5|西门 说：“老师，我们整夜劳累，并没有打着什么。但依从你的话，我就下网。”
LUKE|5|6|他们下了网，圈住许多鱼，网险些裂开，
LUKE|5|7|就招手叫另一只船上的同伴来帮助。他们就来，把鱼装满了两只船，船甚至要沉下去。
LUKE|5|8|西门．彼得 看见，就俯伏在耶稣膝前，说：“主啊，离开我，我是个罪人。”
LUKE|5|9|他和一切跟他一起的人对打到了这一网的鱼都很惊讶。
LUKE|5|10|他的伙伴 西庇太 的儿子 雅各 、 约翰 ，也是这样。耶稣对 西门 说：“不要怕！从今以后，你要得人了。”
LUKE|5|11|他们把两只船靠了岸，就撇下所有的，跟从了耶稣。
LUKE|5|12|有一回，耶稣在一个城里，有人满身长了痲疯，看见他，就俯伏在地，求他说：“主啊，你若肯，你能使我洁净。”
LUKE|5|13|耶稣伸手摸他，说：“我肯，你洁净了吧！”痲疯病立刻离开了他。
LUKE|5|14|耶稣吩咐他：“你不可告诉任何人，只要去，把自己给祭司察看，又因为你已经洁净，要照 摩西 所吩咐的献上祭物，作为证据给众人看。”
LUKE|5|15|但耶稣的名声越发传扬出去。有一大群人聚集来听道，也希望耶稣医治他们的病。
LUKE|5|16|耶稣却退到旷野去祷告。
LUKE|5|17|有一天，耶稣教导人，有法利赛人和律法教师在旁边坐着；他们是从 加利利 各乡村、 犹太 和 耶路撒冷 来的。主的能力与耶稣同在，使他能治好病人。
LUKE|5|18|这时，有些人用褥子抬着一个瘫子，要把他抬进去放在耶稣面前，
LUKE|5|19|却因人多，找不出法子抬进去，就上了房顶，从瓦间把他连褥子缒到当中，在耶稣面前。
LUKE|5|20|耶稣见他们的信心，就说：“朋友，你的罪赦了。”
LUKE|5|21|文士和法利赛人就开始议论说：“这个人是谁，竟说亵渎的话？除了上帝一位之外，谁能赦罪呢？”
LUKE|5|22|耶稣知道他们所议论的，就回答他们说：“你们心里为什么议论呢？
LUKE|5|23|说‘你的罪赦了’，或说‘你起来行走’，哪一样容易呢？
LUKE|5|24|但要让你们知道，人子在地上有赦罪的权柄。”他就对瘫子说：“我吩咐你，起来！拿你的褥子回家去吧。”
LUKE|5|25|那人当着众人面前立刻起来，拿了他所躺卧的褥子回家去，归荣耀给上帝。
LUKE|5|26|众人都惊奇，也归荣耀给上帝，并且满心惧怕，说：“我们今日看见不寻常的事了！”
LUKE|5|27|这些事以后，耶稣出去，看见一个税吏，名叫 利未 ，在税关坐着，就对他说：“来跟从我！”
LUKE|5|28|他就撇下所有的，起来跟从耶稣。
LUKE|5|29|利未 在自己家里为耶稣大摆宴席，有一大群税吏和别的人与他们一同坐席。
LUKE|5|30|法利赛人和文士就向耶稣的门徒发怨言说：“你们为什么跟税吏和罪人一同吃喝呢？”
LUKE|5|31|耶稣回答他们：“健康的人用不着医生；有病的人才用得着。
LUKE|5|32|我不是来召义人悔改，而是召罪人悔改。”
LUKE|5|33|他们对耶稣说：“ 约翰 的门徒常常禁食祈祷，法利赛人的门徒也是这样，惟独跟你在一起的又吃又喝。”
LUKE|5|34|耶稣对他们说：“新郎和宾客在一起的时候，你们怎么能叫宾客禁食呢？
LUKE|5|35|但日子将到，新郎要被带走，那些日子他们就要禁食了。”
LUKE|5|36|耶稣又讲一个比喻，对他们说：“没有人把新衣服撕下一块来补在旧衣服上，若是这样，会把新的撕裂了，并且所撕下来的那块新的和旧的也不相称。
LUKE|5|37|也没有人把新酒装在旧皮袋里；若是这样，新酒会胀破皮袋，酒就漏出来，皮袋也糟蹋了。
LUKE|5|38|相反地，新酒必须装在新皮袋里。
LUKE|5|39|没有人喝了陈酒又想喝新的；他总说陈的好。”
LUKE|6|1|有一个安息日 ，耶稣从麦田经过。他的门徒摘了麦穗，用手搓着吃。
LUKE|6|2|有几个法利赛人说：“你们为什么做安息日不合法的事呢？”
LUKE|6|3|耶稣回答他们：“ 大卫 和跟从他的人饥饿时所做的事，你们没有念过吗？
LUKE|6|4|他怎么进了上帝的居所，拿供饼吃，又给跟从的人吃呢？这饼惟独祭司可以吃，别人都不可以吃。”
LUKE|6|5|他又对他们说：“人子是安息日的主。”
LUKE|6|6|又有一个安息日，耶稣进了会堂教导人，在那里有一个人，他的右手萎缩了。
LUKE|6|7|文士和法利赛人窥探耶稣会不会在安息日治病，为要找把柄告他。
LUKE|6|8|耶稣却知道他们的意念，就对那萎缩了手的人说：“起来，站在当中！”那人就起来，站着。
LUKE|6|9|耶稣对他们说：“我问你们，在安息日行善行恶，救命害命，哪样是合法的呢？”
LUKE|6|10|他就环视众人，对那人说：“伸出手来！”他照着做，他的手就复原了。
LUKE|6|11|他们怒气填胸，彼此商议怎样对付耶稣。
LUKE|6|12|在那些日子，耶稣出去，上山祈祷，整夜向上帝祷告。
LUKE|6|13|到了天亮，他叫门徒来，就从他们中间挑选十二个人，称他们为使徒。
LUKE|6|14|这十二个人有 西门 （耶稣又给他起名叫 彼得 ），还有他弟弟 安得烈 ，又有 雅各 和 约翰 ， 腓力 和 巴多罗买 ，
LUKE|6|15|马太 和 多马 ， 亚勒腓 的儿子 雅各 和激进党的 西门 ，
LUKE|6|16|雅各 的儿子 犹大 和后来成为出卖者的 加略 人 犹大 。
LUKE|6|17|耶稣和他们下了山，站在一块平地上；在一起的有许多门徒，又有许多百姓从全 犹太 和 耶路撒冷 ，并 推罗 、 西顿 的海边来，
LUKE|6|18|都要听他讲道，又希望耶稣医治他们的病；还有被污灵缠磨的，也得了医治。
LUKE|6|19|众人都想要摸他，因为有能力从他身上发出来，治好了他们。
LUKE|6|20|耶稣举目看着门徒，说： “贫穷的人有福了！ 因为上帝的国是你们的。
LUKE|6|21|现在饥饿的人有福了！ 因为你们将得饱足。 现在哭泣的人有福了！ 因为你们将要欢笑。
LUKE|6|22|人为人子的缘故憎恨你们，拒绝你们，辱骂你们，把你们当恶人除掉你们的名，你们就有福了！
LUKE|6|23|在那日，你们要欢欣雀跃，因为你们在天上的赏赐是很多的；他们的祖宗也是这样待先知的。
LUKE|6|24|但你们富足的人有祸了！ 因为你们已经受过安慰。
LUKE|6|25|你们现在饱足的人有祸了！ 因为你们将要饥饿。 你们现在欢笑的人有祸了！ 因为你们将要哀恸哭泣。
LUKE|6|26|人都说你们好的时候，你们有祸了！因为他们的祖宗也是这样待假先知的。”
LUKE|6|27|“可是我告诉你们这些听的人，要爱你们的仇敌！要善待恨你们的人！
LUKE|6|28|要祝福诅咒你们的人！要为凌辱你们的人祷告！
LUKE|6|29|有人打你的脸，连另一边也由他打。有人拿你的外衣，连内衣也由他拿去。
LUKE|6|30|凡求你的，就给他；有人拿走你的东西，不要讨回来。
LUKE|6|31|“你们想要人怎样待你们，你们也要怎样待人。
LUKE|6|32|你们若只爱那爱你们的人，有什么可感谢的呢？就是罪人也爱那爱他们的人。
LUKE|6|33|你们若善待那善待你们的人，有什么可感谢的呢？就是罪人也是这样做。
LUKE|6|34|你们若借给人，希望从他收回，有什么可感谢的呢？就是罪人也借给罪人，再如数收回。
LUKE|6|35|你们倒要爱仇敌，要善待他们，并要借给人不指望偿还，你们的赏赐就很多了，你们必作至高者的儿子，因为他恩待那忘恩的和作恶的。
LUKE|6|36|你们要仁慈，像你们的父是仁慈的。”
LUKE|6|37|“你们不要评断别人，就不被审判；你们不要定人的罪，就不被定罪；你们要饶恕人，就必蒙饶恕。
LUKE|6|38|你们要给人，就必有给你们的，并且用十足的升斗，连摇带按，上尖下流地倒在你们怀里；因为你们用什么量器量给人，也必用什么量器量给你们。”
LUKE|6|39|耶稣又用比喻对他们说：“瞎子岂能领瞎子，两个人不是都要掉在坑里吗？
LUKE|6|40|学生不高过老师，凡学成了的会和老师一样。
LUKE|6|41|为什么看见你弟兄眼中有刺，却不想自己眼中有梁木呢？
LUKE|6|42|你不见自己眼中有梁木，怎能对你弟兄说：‘让我去掉你眼中的刺’呢？你这假冒为善的人！先去掉自己眼中的梁木，然后才能看得清楚，好去掉你弟兄眼中的刺。”
LUKE|6|43|“没有好树结坏果子，也没有坏树结好果子。
LUKE|6|44|每一种树木可以从其果子看出来。人不是从荆棘上摘无花果的，也不是从蒺藜里摘葡萄的。
LUKE|6|45|善人从他心里所存的善发出善来，恶人从他所存的恶发出恶来；因为心里所充满的，口里就说出来。”
LUKE|6|46|“你们为什么称呼我‘主啊，主啊’，却不照我的话做呢？
LUKE|6|47|凡到我这里来，听了我的话又去做的，我要告诉你们他像什么人：
LUKE|6|48|他像一个人盖房子，把地挖深，将根基立在磐石上，到发大水的时候，水冲那房子，房子总不动摇，因为盖造得好。
LUKE|6|49|但听了不去做的，就像一个人在土地上盖房子，没有根基，水一冲，立刻倒塌了，并且那房子损坏得很厉害。”
LUKE|7|1|耶稣对百姓讲完了这一切的话，就进了 迦百农 。
LUKE|7|2|有一个百夫长所器重的仆人害病，快要死了。
LUKE|7|3|百夫长风闻耶稣的事，就托 犹太 人的几个长老去求耶稣来救他的仆人。
LUKE|7|4|他们到了耶稣那里，切切地求他说：“你为他做这事是他配得的；
LUKE|7|5|因为他爱我们的民族，为我们建造会堂。”
LUKE|7|6|耶稣就和他们同去。离那家不远，百夫长托几个朋友去见耶稣，对他说：“主啊，不必劳驾，因你到舍下来，我不敢当。
LUKE|7|7|我也自以为不配去见你，只要你说一句话，就会让我的僮仆得痊愈。
LUKE|7|8|因为我被派在人的权下，也有兵在我之下。我对这个说：‘去！’他就去；对那个说：‘来！’他就来；对我的仆人说：‘做这事！’他就去做。”
LUKE|7|9|耶稣听到这些话，就很惊讶，转身对跟随的众人说：“我告诉你们，这么大的信心，就是在 以色列 ，我也没有见过。”
LUKE|7|10|那差来的人回到百夫长家里，发现仆人已经好了。
LUKE|7|11|过了不久 ，耶稣往一座城去，这城名叫 拿因 ，他的门徒和一大群人与他同行。
LUKE|7|12|当他走近城门时，有一个死人被抬出来。这人是他母亲独生的儿子，而他母亲又是寡妇。城里的许多人与她一同送殡。
LUKE|7|13|主看见那寡妇就怜悯她，对她说：“不要哭。”
LUKE|7|14|于是耶稣进前来，按着杠，抬的人就站住了。耶稣说：“年轻人，我吩咐你，起来！”
LUKE|7|15|那死人就坐了起来，开始说话，耶稣就把他交给他的母亲。
LUKE|7|16|众人都惊奇，归荣耀给上帝，说：“有大先知在我们当中兴起了！”又说：“上帝眷顾了他的百姓！”
LUKE|7|17|关于耶稣的这事就传遍了 犹太 和周围地区。
LUKE|7|18|约翰 的门徒把这些事都告诉 约翰 。于是 约翰 叫了两个门徒来，
LUKE|7|19|差他们到主 那里去，说：“将要来的那位就是你吗？还是我们要等候别人呢？”
LUKE|7|20|那两个人来到耶稣那里，说：“施洗的 约翰 差我们来问你：‘将要来的那位就是你吗？还是我们要等候别人呢？’”
LUKE|7|21|就在那时，耶稣治好了许多患疾病的，得瘟疫的，被邪灵附身的，又开恩使好些盲人能看见。
LUKE|7|22|耶稣回答他们：“你们去，把所看见、所听见的告诉 约翰 ：就是盲人看见，瘸子行走，痲疯病人得洁净，聋子听见，死人复活，穷人听到福音。
LUKE|7|23|凡不因我跌倒的有福了！”
LUKE|7|24|约翰 所差来的人一走，耶稣就对众人谈到 约翰 ，说：“你们从前到旷野去，是要看什么呢？被吹动的芦苇吗？
LUKE|7|25|你们出去到底是要看什么？穿细软衣服的人吗？看哪，那穿华丽衣服、宴乐度日的人是在王宫里。
LUKE|7|26|你们出去究竟是要看什么？是先知吗？是的，我告诉你们，他比先知大多了。
LUKE|7|27|这个人就是经上所说的： ‘看哪，我要差遣我的使者在你面前， 他要在你前面为你预备道路。’
LUKE|7|28|我告诉你们，凡女子所生的，没有比 约翰 大的；但在上帝国里，最小的比他还大。”
LUKE|7|29|众百姓和税吏已受过 约翰 的洗，听见这话，就以上帝为义；
LUKE|7|30|但法利赛人和律法师没有受过 约翰 的洗，竟废弃了上帝为他们所定的旨意。
LUKE|7|31|主又说：“这样，我该用什么来比这世代的人呢？他们好像什么呢？
LUKE|7|32|这正像孩童坐在街市上，彼此喊叫： ‘我们为你们吹笛，你们不跳舞； 我们唱哀歌，你们不啼哭。’
LUKE|7|33|施洗的 约翰 来，不吃饼，不喝酒，你们说他是被鬼附的。
LUKE|7|34|人子来，也吃也喝，你们又说这人贪食好酒，是税吏和罪人的朋友。
LUKE|7|35|而智慧是由所有智慧的人来证实的。”
LUKE|7|36|有一个法利赛人请耶稣和他吃饭，耶稣就到那法利赛人家里去坐席。
LUKE|7|37|那城里有一个女人，是个罪人，知道耶稣在法利赛人家里坐席，就拿着盛满香膏的玉瓶，
LUKE|7|38|站在耶稣背后，挨着他的脚哭，眼泪滴湿了耶稣的脚，就用自己的头发擦干，又用嘴连连亲他的脚，把香膏抹上。
LUKE|7|39|请耶稣的法利赛人看见这事，心里说：“这人若是先知，一定知道摸他的是谁，是个怎样的女人；她是个罪人哪！”
LUKE|7|40|耶稣回应他说：“ 西门 ，我有话要对你说。” 西门 说：“老师，请说。”
LUKE|7|41|耶稣说：“有两个人欠了某一个债主的钱，一个欠五百个银币，一个欠五十个银币。
LUKE|7|42|因为他们无力偿还，债主就开恩赦免了他们两个人的债。那么，这两个人哪一个更爱他呢？”
LUKE|7|43|西门 回答：“我想是那多得赦免的人。”耶稣对他说：“你的判断不错。”
LUKE|7|44|于是他转过来向着那女人，对 西门 说：“你看见这女人吗？我进了你的家，你没有给我水洗脚，但这女人用眼泪滴湿了我的脚，又用头发擦干。
LUKE|7|45|你没有亲我，但这女人从我进来就不住地亲我的脚。
LUKE|7|46|你没有用油抹我的头，但这女人用香膏抹我的脚。
LUKE|7|47|所以我告诉你，她许多的罪都赦免了，因为她爱的多；而那少得赦免的，爱的就少。”
LUKE|7|48|于是耶稣对那女人说：“你的罪都赦免了。”
LUKE|7|49|同席的人心里说：“这是什么人，竟赦免人的罪呢？”
LUKE|7|50|耶稣对那女人说：“你的信救了你，平安地回去吧！”
LUKE|8|1|过了不久，耶稣周游各城各乡传道，宣讲上帝国的福音。和他同去的有十二个使徒，
LUKE|8|2|还有曾被邪灵所附，被疾病所缠，而已经治好的几个妇女，其中有称为 抹大拉 的 马利亚 ，曾有七个鬼从她身上赶出来，
LUKE|8|3|又有 希律 的管家 苦撒 的妻子 约亚拿 ，和 苏撒拿 以及好些别的妇女，她们都是用自己的财物供给耶稣和使徒。
LUKE|8|4|当一大群人聚集，又有人从各城里出来见耶稣的时候，耶稣用比喻说：
LUKE|8|5|“有一个撒种的出去撒种。他撒的时候，有的落在路旁，被人践踏，天上的飞鸟又来把它吃掉了。
LUKE|8|6|有的落在磐石上，一出来就枯干了，因为得不着滋润。
LUKE|8|7|有的落在荆棘里，荆棘跟它一同生长，把它挤住了。
LUKE|8|8|又有的落在好土里，生长起来，结实百倍。”耶稣说完这些话，大声说：“有耳可听的，就应当听！”
LUKE|8|9|门徒问耶稣这比喻是什么意思。
LUKE|8|10|他说：“上帝国的奥秘只让你们知道，至于别人，就用比喻，要 他们看也看不见， 听也不明白。”
LUKE|8|11|“这比喻是这样的：种子就是上帝的道。
LUKE|8|12|那些在路旁的，就是人听了道，随后魔鬼来，从他们心里把道夺去，以免他们信了得救。
LUKE|8|13|那些在磐石上的，就是人听道，欢喜领受，但没有根，不过暂时相信，等到碰上试炼就退后了。
LUKE|8|14|那落在荆棘里的，就是人听了道，走开以后，被今生的忧虑、钱财、宴乐挤住了，结不出成熟的子粒来。
LUKE|8|15|那落在好土里的，就是人听了道，并用纯真善良的心持守它，耐心等候结果实。”
LUKE|8|16|“没有人点灯用器皿盖上，或放在床底下，而是放在灯台上，让进来的人看见亮光。
LUKE|8|17|因为掩藏的事没有不显出来的，隐瞒的事也没有不露出来被人知道的。
LUKE|8|18|所以，你们应当小心怎样听。因为凡有的，还要给他；凡没有的，连他自以为有的也要夺去。”
LUKE|8|19|耶稣的母亲和他兄弟来看他，因为人多，不能到他跟前。
LUKE|8|20|有人告诉他说：“你母亲和你兄弟站在外边，要见你。”
LUKE|8|21|耶稣回答他们：“听了上帝的道而遵行的人，就是我的母亲，我的兄弟了。”
LUKE|8|22|有一天，耶稣和门徒上了船，他对门徒说：“我们渡到湖的对岸去吧。”他们就开了船。
LUKE|8|23|船行的时候，耶稣睡着了。湖上忽然起了狂风，船将灌满了水，很危险。
LUKE|8|24|门徒去叫醒他，说：“老师！老师！我们快没命啦！”耶稣醒了，斥责那狂风大浪，风浪就止住，平静了。
LUKE|8|25|耶稣对他们说：“你们的信心在哪里呢？”他们又惧怕又惊讶，彼此说：“这到底是谁？他吩咐风和水，连风和水都听从他。”
LUKE|8|26|他们到了 格拉森 人的地区，就在 加利利 的对面。
LUKE|8|27|耶稣上了岸，就有城里一个被鬼附的人迎着他走来。这个人好久不穿衣服，不住在屋子里，而住在坟墓里。
LUKE|8|28|他看见耶稣，就喊叫着俯伏在他面前，大声说：“至高上帝的儿子耶稣，你为什么干扰我？我求你，不要叫我受苦！”
LUKE|8|29|这是因耶稣曾吩咐污灵从这人身上出来。原来这污灵屡次抓住他；他常被人看守，又被铁链和脚镣捆锁，他竟把锁链挣断，被鬼赶到旷野去。
LUKE|8|30|耶稣问他：“你的名字叫什么？”他说：“ 群 ”；这是因为附着他的鬼多。
LUKE|8|31|鬼就央求耶稣不要命令他们到无底坑里去。
LUKE|8|32|那里有一大群猪正在山坡上吃食，鬼央求耶稣准他们进入猪里；耶稣准了他们。
LUKE|8|33|于是鬼从那人出来，进入猪里，那群猪就闯下山崖，投进湖里，淹死了。
LUKE|8|34|放猪的看见这事就逃跑了，去告诉城里和乡下的人。
LUKE|8|35|众人出来，要看发生了什么事；到了耶稣那里，发现那人坐在耶稣脚前，鬼已离开了他，穿着衣服，神智清醒，他们就害怕。
LUKE|8|36|看见这事的人把被鬼附的人怎么得医治的事告诉他们。
LUKE|8|37|格拉森 周围地区的人，因为害怕得很，都求耶稣离开他们；耶稣就上船回去了。
LUKE|8|38|鬼已从身上出去的那人恳求要和耶稣在一起，耶稣却打发他回去，说：
LUKE|8|39|“你回家去，传讲上帝为你做了多么大的事。”他就走遍全城，传扬耶稣为他做了多么大的事。
LUKE|8|40|耶稣回来的时候，众人迎接他，因为他们都等候着他。
LUKE|8|41|有一个会堂主管，名叫 叶鲁 ，来俯伏在耶稣脚前，求耶稣到他家里去，
LUKE|8|42|因为他有一个独生女，约十二岁，快要死了。 耶稣去的时候，众人簇拥着他。
LUKE|8|43|有一个女人，患了经血不止的病有十二年，在医生手里花尽了一生所有的 ，但没有人能治好她。
LUKE|8|44|她来到耶稣背后，摸他的衣裳繸子，经血立刻止住了。
LUKE|8|45|耶稣说：“摸我的是谁？”众人都不承认。 彼得 说：“老师，众人拥拥挤挤紧靠着你。”
LUKE|8|46|耶稣说：“有人摸了我，因为我觉得有能力从我身上出去。”
LUKE|8|47|那女人知道瞒不住了，就战战兢兢地俯伏在耶稣跟前，把摸他的缘故和怎样立刻痊愈的事，当着众人都说出来。
LUKE|8|48|耶稣对她说：“女儿，你的信救了你。平安地回去吧！”
LUKE|8|49|耶稣还在说话的时候，有人从会堂主管的家里来，说：“你的女儿死了，不要劳驾老师了。”
LUKE|8|50|耶稣听见就对他说：“不要怕，只要信！她必得痊愈。”
LUKE|8|51|耶稣到了他的家，除了 彼得 、 约翰 、 雅各 ，和女儿的父母，不许别人同他进去。
LUKE|8|52|众人都在为这女孩哀哭捶胸。耶稣说：“不要哭，她不是死了，是睡着了。”
LUKE|8|53|他们知道她已经死了，就嘲笑耶稣。
LUKE|8|54|耶稣拉着她的手，呼叫着：“孩子，起来吧！”
LUKE|8|55|她的灵魂就回来了，她立刻起来。耶稣吩咐给她东西吃。
LUKE|8|56|她的父母非常惊奇；耶稣吩咐他们不要把所发生的事告诉任何人。
LUKE|9|1|耶稣叫齐了十二使徒，给他们能力和权柄制伏一切的鬼，医治疾病，
LUKE|9|2|又差遣他们宣讲上帝的国，医治病人，
LUKE|9|3|对他们说：“途中什么都不要带；不要带手杖和行囊，不要带食物和银钱，也不要带两件内衣 。
LUKE|9|4|你们无论进哪一家，就住在哪里，也从那里离开。
LUKE|9|5|凡不接待你们的，你们离开那城的时候，要跺掉你们脚上的尘土，证明他们的不是。”
LUKE|9|6|于是使徒出去，走遍各乡传福音，到处治病。
LUKE|9|7|希律 分封王听见耶稣所做的一切事，就困惑起来，因为有人说：“ 约翰 从死人中复活了。”
LUKE|9|8|又有人说：“ 以利亚 显现了。”还有人说：“古时的一个先知又活了。”
LUKE|9|9|希律 说：“ 约翰 我已经斩了，但这是什么人？关于他，我竟听到这样的事！”于是 希律 想要见他。
LUKE|9|10|使徒们回来，把所做的事告诉耶稣，耶稣就私下带他们离开那里，往一座叫 伯赛大 的城去。
LUKE|9|11|众人知道了，就跟着他去；耶稣接待他们，对他们讲论上帝国的事，治好那些需要医治的人。
LUKE|9|12|太阳快要下山，十二使徒进前来对他说：“请叫众人散去，他们好往四面村庄乡镇里去借宿和找吃的，因为我们这里地方偏僻。”
LUKE|9|13|耶稣对他们说：“你们给他们吃吧！”他们说：“我们不过有五个饼、两条鱼，若不去为这许多人买食物就不够。”
LUKE|9|14|那时，男人约有五千。耶稣对门徒说：“叫他们分组坐下，每组大约五十个人。”
LUKE|9|15|门徒就这样做了，叫众人都坐下。
LUKE|9|16|耶稣拿着这五个饼和两条鱼，望着天祝福，擘开，递给门徒，摆在众人面前。
LUKE|9|17|所有的人都吃，并且吃饱了。他们把剩下的碎屑收拾起来，装满了十二个篮子。
LUKE|9|18|耶稣独自祷告的时候，门徒也同他在那里。耶稣问他们：“众人说我是谁？”
LUKE|9|19|他们回答：“是施洗的 约翰 ；有人说是 以利亚 ；还有人说是古时的一个先知又活了。”
LUKE|9|20|耶稣问他们：“你们说我是谁？” 彼得 回答：“是上帝所立的基督。”
LUKE|9|21|耶稣切切吩咐他们，命令他们不可把这事告诉任何人；
LUKE|9|22|又说：“人子必须受许多的苦，被长老、祭司长和文士弃绝，并且被杀，第三天复活。”
LUKE|9|23|耶稣又对众人说：“若有人要跟从我，就当舍己，天天背起自己的十字架来跟从我。
LUKE|9|24|因为凡要救自己生命的，必丧失生命；凡为我丧失生命的，他必救自己的生命。
LUKE|9|25|人就是赚得全世界，却丧失了自己，或赔上自己，有什么益处呢？
LUKE|9|26|凡把我和我的道当作可耻的，人子在自己的荣耀里，和天父与圣天使的荣耀里来临的时候，也要把那人当作可耻的。
LUKE|9|27|我实在告诉你们，站在这里的，有人在没经历死亡以前，必定看见上帝的国。”
LUKE|9|28|说了这些话以后约有八天，耶稣带着 彼得 、 约翰 、 雅各 上山去祷告。
LUKE|9|29|正祷告的时候，他的面貌改变了，衣服洁白放光。
LUKE|9|30|忽然有 摩西 和 以利亚 两个人同耶稣说话；
LUKE|9|31|他们在荣光里显现，谈论耶稣去世的事，就是他在 耶路撒冷 将要完成的事。
LUKE|9|32|彼得 和他的同伴都打盹，但一清醒，就看见耶稣的荣光和与他一起站着的那两个人。
LUKE|9|33|二人正要和耶稣分离的时候， 彼得 对耶稣说：“老师，我们在这里真好！我们来搭三座棚，一座为你，一座为 摩西 ，一座为 以利亚 。”他却不知道自己在说些什么。
LUKE|9|34|说这些话的时候，有一朵云彩来遮盖他们；他们一进入云彩就很惧怕。
LUKE|9|35|有声音从云彩里出来，说：“这是我的儿子，我所拣选的 。你们要听从他！”
LUKE|9|36|声音停止后，只见耶稣独自一人。当那些日子，门徒保持沉默，不把所看见的事告诉任何人。
LUKE|9|37|第二天，他们下了山，有一大群人来迎见耶稣。
LUKE|9|38|其中有一人喊着说：“老师！求你看看我的儿子，因为他是我的独子。
LUKE|9|39|他被灵拿住就突然喊叫，那灵又使他抽风，口吐白沫，并且重重地伤害他，不轻易放过他。
LUKE|9|40|我求过你的门徒把那灵赶出去，他们却不能。”
LUKE|9|41|耶稣回答：“唉！这又不信又悖谬的世代啊，我和你们在一起，忍耐你们，要到几时呢？把你的儿子带到这里来！”
LUKE|9|42|他正来的时候，那鬼把他摔倒，使他重重地抽风。耶稣斥责那污灵，把孩子治好了，交给他父亲。
LUKE|9|43|众人都诧异上帝的大能 。 众人正惊讶于耶稣所做的一切事的时候，耶稣对门徒说：
LUKE|9|44|“你们要把这些话听进去，因为人子将要被交在人手里。”
LUKE|9|45|门徒却不明白这话，其中的意思对他们隐藏着，使他们不能明白，他们也不敢问这话的意思。
LUKE|9|46|门徒互相议论，他们中间谁最大。
LUKE|9|47|耶稣看出他们心中的议论，就领一个小孩子来，叫他站在自己旁边，
LUKE|9|48|对他们说：“凡为我的名接纳这小孩子的，就是接纳我；凡接纳我的，就是接纳那差我来的。你们中间最小的，他就是最大的。”
LUKE|9|49|约翰 回应说：“老师，我们看见一个人奉你的名赶鬼，我们就阻止他，因为他不与我们一同跟从你。”
LUKE|9|50|耶稣对他说：“不要阻止他，因为不抵挡你们的，就是帮助你们的。”
LUKE|9|51|耶稣被接上升的日子将到，他决定面向 耶路撒冷 走去。
LUKE|9|52|他打发使者在他前头走；他们进了 撒玛利亚 的一个村庄，要为他作准备。
LUKE|9|53|那里的人不接待他，因为他面向着 耶路撒冷 去。
LUKE|9|54|他的门徒 雅各 和 约翰 看见了，就说：“主啊！你要我们吩咐火从天上降下来，烧灭他们 吗？”
LUKE|9|55|耶稣转身责备两个门徒。
LUKE|9|56|于是他们就往别的村庄去了。
LUKE|9|57|他们在路上走的时候，有一个人对耶稣说：“你无论往哪里去，我都要跟从你。”
LUKE|9|58|耶稣对他说：“狐狸有洞，天空的飞鸟有窝，人子却没有枕头的地方。”
LUKE|9|59|他又对另一个人说：“来跟从我！”那人说：“主啊 ，容许我先回去埋葬我的父亲。”
LUKE|9|60|耶稣对他说：“让死人埋葬他们的死人，你只管去传讲上帝的国。”
LUKE|9|61|又有一人说：“主啊，我要跟从你，但容许我先去辞别我家里的人。”
LUKE|9|62|耶稣对他说：“手扶着犁向后看的人，不配进上帝的国。”
LUKE|10|1|这些事以后，主另外指定七十二个人 ，差遣他们两个两个地在他前面，往自己所要到的各城各地去。
LUKE|10|2|他对他们说：“要收的庄稼多，做工的人少。所以，你们要求庄稼的主差遣做工的人出去收他的庄稼。
LUKE|10|3|你们去吧！看！我差你们出去，如同羔羊进入狼群。
LUKE|10|4|不要带钱囊，不要带行囊，不要带鞋子；在路上也不要向人问安。
LUKE|10|5|无论进哪一家，先要说：‘愿这一家平安。’
LUKE|10|6|那里若有当得平安的人，你们所求的平安就必临到那家，不然，将归还你们。
LUKE|10|7|你们要住在那家，吃喝他们所供给的，因为工人得工钱是应当的；不要从这家搬到那家。
LUKE|10|8|无论进哪一城，人若接待你们，给你们摆上什么食物，你们就吃什么。
LUKE|10|9|要医治那城里的病人，对他们说：‘上帝的国临近你们了。’
LUKE|10|10|无论进哪一城，人若不接待你们，你们就到大街上去，说：
LUKE|10|11|‘就是你们城里的尘土粘在我们的脚上，我们也当着你们擦去。但是，你们该知道上帝的国临近了。’
LUKE|10|12|我告诉你们，在那日子， 所多玛 所受的，比那城还容易受呢！”
LUKE|10|13|“ 哥拉汛 哪，你有祸了！ 伯赛大 啊，你有祸了！因为在你们中间所行的异能，若行在 推罗 、 西顿 ，他们早已披麻蒙灰，坐在地上悔改了。
LUKE|10|14|在审判的时候， 推罗 和 西顿 所受的，比你们还容易受呢！
LUKE|10|15|迦百农 啊， 你以为要被举到天上吗？ 你要被推下阴间！”
LUKE|10|16|耶稣又对门徒说：“听从你们的就是听从我；弃绝你们的就是弃绝我；弃绝我的就是弃绝差遣我来的那位。”
LUKE|10|17|那七十二个人欢欢喜喜地回来，说：“主啊，因你的名，就是鬼也服了我们。”
LUKE|10|18|耶稣对他们说：“我看见撒但从天上坠落，像闪电一样。
LUKE|10|19|我已经给你们权柄可以践踏蛇和蝎子，又胜过仇敌一切的能力，绝没有什么能害你们。
LUKE|10|20|然而，不要因灵服了你们就欢喜，而要因你们的名记录在天上欢喜。”
LUKE|10|21|正当那时，耶稣被圣灵感动而欢喜快乐，说：“父啊，天地的主，我感谢你！因为你把这些事向聪明智慧的人隐藏起来，而向婴孩启示出来。父啊，是的，因为你的美意本是如此。
LUKE|10|22|一切都是我父交给我的。除了父，没有人知道子是谁；除了子和子所愿意启示的人，没有人知道父是谁。”
LUKE|10|23|耶稣转身私下对门徒说：“看见你们所看见的，那眼睛有福了。
LUKE|10|24|我告诉你们，从前有许多先知和君王要看你们所看的，却没有看见，要听你们所听的，却没有听见。”
LUKE|10|25|有一个律法师起来试探耶稣，说：“老师！我该做什么才可以承受永生？”
LUKE|10|26|耶稣对他说：“律法上写的是什么？你是怎样念的呢？”
LUKE|10|27|他回答说：“你要尽心、尽性、尽力、尽意爱主—你的上帝，又要爱邻 如己。”
LUKE|10|28|耶稣对他说：“你回答得正确，你这样做就会得永生。”
LUKE|10|29|那人要证明自己有理，就对耶稣说：“谁是我的邻舍呢？”
LUKE|10|30|耶稣回答：“有一个人从 耶路撒冷 下 耶利哥 去，落在强盗手中。他们剥去他的衣裳，把他打个半死，丢下他走了。
LUKE|10|31|偶然有一个祭司从那条路下来，看见他就从另一边过去了。
LUKE|10|32|又有一个 利未 人来到那里，看见他，也照样从另一边过去了。
LUKE|10|33|可是，有一个 撒玛利亚 人路过那里，看见他就动了慈心，
LUKE|10|34|上前用油和酒倒在他的伤处，包裹好了，扶他骑上自己的牲口，带他到旅店里去，照应他。
LUKE|10|35|第二天，他拿出两个银币来，交给店主，说：‘请你照应他，额外的费用，我回来时会还你。’
LUKE|10|36|你想，这三个人哪一个是落在强盗手中那人的邻舍呢？”
LUKE|10|37|他说：“是怜悯他的。”耶稣对他说：“你去，照样做吧！”
LUKE|10|38|他们继续前行，耶稣进了一个村庄。有一个女人，名叫 马大 ，接他到自己家里。
LUKE|10|39|她有一个妹妹，名叫 马利亚 ，在主的脚前坐着听他的道。
LUKE|10|40|马大 伺候的事多，心里忙乱，进前来，说：“主啊，我的妹妹留下我一个人伺候，你不在意吗？请吩咐她来帮助我。”
LUKE|10|41|主回答说：“ 马大 ， 马大 ，你为许多的事操心烦恼，
LUKE|10|42|但是不可少的只有一件 。 马利亚 已经选择了那上好的福分，是没有人能从她夺去的。”
LUKE|11|1|耶稣在一个地方祷告。祷告完了，有个门徒对他说：“主啊，求你教导我们祷告，像 约翰 教导他的门徒一样。”
LUKE|11|2|耶稣对他们说：“你们祷告的时候，要说： ‘父啊， 愿人都尊你的名为圣； 愿你的国降临；
LUKE|11|3|我们日用的饮食，天天赐给我们。
LUKE|11|4|赦免我们的罪， 因为我们也赦免凡亏欠我们的人。 不叫我们陷入试探。 ’”
LUKE|11|5|耶稣又对他们说：“你们中间谁有一个朋友半夜到他那里去，对他说：‘朋友！请借给我三个饼；
LUKE|11|6|因为我有一个朋友旅途中来到我这里，我没有东西招待他。’
LUKE|11|7|那人在里面回答：‘不要打扰我，门已经关了，孩子们也同我在床上了，我不能起来给你。’
LUKE|11|8|我告诉你们，虽不因他是朋友起来给他，也会因他不顾面子地直求，起来照他所需要的给他。
LUKE|11|9|我又告诉你们，祈求，就给你们；寻找，就找到；叩门，就给你们开门。
LUKE|11|10|因为凡祈求的，就得着；寻找的，就找到；叩门的，就给他开门。
LUKE|11|11|你们中间作父亲的，谁有儿子 求鱼，反拿蛇当鱼给他呢？
LUKE|11|12|求鸡蛋，反给他蝎子呢？
LUKE|11|13|你们虽然不好，尚且知道拿好东西给儿女，何况 天父，他岂不更要把圣灵赐给求他的人吗？”
LUKE|11|14|耶稣赶出一个使人成为哑巴的鬼 ，鬼出去了，哑巴就说出话来；众人都很惊讶。
LUKE|11|15|其中却有人说：“他是靠着鬼王 别西卜 赶鬼。”
LUKE|11|16|又有人试探耶稣，要他显个来自天上的神迹。
LUKE|11|17|他知道他们的意念，就对他们说：“一国自相纷争，必定荒芜；一家自相纷争，就必败落。
LUKE|11|18|撒但若自相纷争，他的国怎能立得住呢？因为你们说我是靠着 别西卜 赶鬼。
LUKE|11|19|我若靠着 别西卜 赶鬼，你们的子弟赶鬼又靠着谁呢？这样，他们要作你们的判官。
LUKE|11|20|我若靠着上帝的能力赶鬼，那么，上帝的国就已临到你们了。
LUKE|11|21|壮士全副武装，看守自己的住宅，他所有的都很安全；
LUKE|11|22|但有一个比他更强的来攻击他，并且战胜了他，就夺去他所倚靠的盔甲兵器，又分了他的掠物。
LUKE|11|23|不跟我一起的，就是反对我；不与我一起收聚的，就是在拆散。”
LUKE|11|24|“污灵离了人身，走遍无水之地寻找安歇之处，却找不到。就说：‘我要回到我原来的屋里去。’
LUKE|11|25|他到了，看见里面打扫干净，修饰好了，
LUKE|11|26|就去另带了七个比自己更恶的灵来，都进去住在那里。那人后来的景况比先前更坏了。”
LUKE|11|27|耶稣正说这些话的时候，众人中间有一个女人高声对他说：“怀你胎乳养你的有福了！”
LUKE|11|28|耶稣却说：“更有福的是听上帝的道而遵守的人！”
LUKE|11|29|当众人越来越拥挤的时候，耶稣说：“这世代是一个邪恶的世代。他们求看神迹，除了 约拿 的神迹以外，再没有神迹给他们看了。
LUKE|11|30|约拿 怎样为 尼尼微 人成了神迹，人子也要照样为这世代的人成为神迹。
LUKE|11|31|在审判的时候，南方的女王要起来定这世代的人的罪，因为她从地极而来，要听 所罗门 智慧的话。看哪，比 所罗门 更大的在这里！
LUKE|11|32|在审判的时候， 尼尼微 人要起来定这世代的罪，因为 尼尼微 人听了 约拿 所传的就悔改了。看哪，比 约拿 更大的在这里！”
LUKE|11|33|“没有人点灯放在地窖里，或是斗底下 ，总是放在灯台上，让进来的人看见亮光。
LUKE|11|34|你的眼睛就是身体的灯。当你的眼睛明亮，全身就光明，当眼睛昏花，全身就黑暗。
LUKE|11|35|所以，你要注意，免得你里面的光暗了。
LUKE|11|36|若是你全身光明，毫无黑暗，就必全然光明，如同灯的明光照亮你。”
LUKE|11|37|耶稣正说话的时候，有一个法利赛人请他吃饭，耶稣就进去坐席。
LUKE|11|38|这法利赛人看见耶稣饭前不先洗手就很诧异。
LUKE|11|39|主对他说：“如今你们法利赛人洗净杯盘的外面，你们里面却满了贪婪和邪恶。
LUKE|11|40|无知的人哪！造外面的，不也造了里面吗？
LUKE|11|41|只要把杯盘里面的施舍给人，对你们来说一切就都洁净了。
LUKE|11|42|“但是你们法利赛人有祸了！因为你们将薄荷、芸香，和各样蔬菜献上十分之一，疏忽了公义和爱上帝的事；这原是你们该做的—至于其他也不可忽略。
LUKE|11|43|你们法利赛人有祸了！因为你们喜爱会堂里的高位，又喜欢人们在街市上向你们问安。
LUKE|11|44|你们有祸了！因为你们如同不显露的坟墓，走在上面的人并不知道。”
LUKE|11|45|律法师中有一个回答耶稣，说：“老师，你这样说也把我们侮辱了。”
LUKE|11|46|耶稣说：“你们律法师也有祸了！因为你们把难挑的担子放在别人身上，自己却不肯动一个指头去减轻这些担子。
LUKE|11|47|你们有祸了！因为你们建造先知的坟墓，那些先知正是你们的祖宗所杀的。
LUKE|11|48|可见你们祖宗所做的事，你们是证人，你们也赞同，因为他们杀了先知，你们建造先知的坟墓。
LUKE|11|49|所以，上帝的智慧也曾说：‘我要差遣先知和使徒到他们那里去，有的他们要残杀，有的他们要迫害’，
LUKE|11|50|为使创世以来所流众先知的血的罪都归在这世代的人身上，
LUKE|11|51|就是从 亚伯 的血起，直到被杀在祭坛和圣所中间的 撒迦利亚 的血为止。是的，我告诉你们，这都要向这世代的人追讨。
LUKE|11|52|你们律法师有祸了！因为你们把知识的钥匙夺了去，自己不进去，要进去的人，你们也阻挡他们。”
LUKE|11|53|耶稣从那里出来，文士和法利赛人就开始极力地催逼他，盘问他许多事，
LUKE|11|54|伺机要抓他的话柄。
LUKE|12|1|这时，有几万人聚集，甚至彼此践踏。耶稣就先对门徒说：“你们要防备法利赛人的酵，就是假冒为善。
LUKE|12|2|掩盖的事没有不显露出来的，隐藏的事也没有不被人知道的。
LUKE|12|3|因此，你们在暗中所说的，将要在明处被人听见；在密室附耳所说的，将要在屋顶上被人宣扬。”
LUKE|12|4|“我的朋友，我对你们说，那最多只能杀人身体而不能再做什么的，不要怕他们。
LUKE|12|5|我提醒你们该怕的是谁：该怕那杀了以后又有权柄把人扔在地狱里的。是的，我告诉你们，正要怕他。
LUKE|12|6|五只麻雀不是卖二铜钱 吗？但在上帝面前，一只也不被忘记；
LUKE|12|7|就是你们的头发也都数过了。不要惧怕，你们比许多的麻雀还贵重！”
LUKE|12|8|“我又告诉你们，凡在人面前认我的，人子在上帝的使者面前也必认他；
LUKE|12|9|在人面前不认我的，人子在上帝的使者面前也必不认他。
LUKE|12|10|凡说话干犯人子的，还可得赦免；但是亵渎圣灵的，总不得赦免。
LUKE|12|11|有人带你们到会堂、官长和掌权的人面前，不要担心怎么答辩，说什么话；
LUKE|12|12|因为就在那时候，圣灵要指教你们该说的话。”
LUKE|12|13|人群中有一个人对耶稣说：“老师！请你吩咐我的兄弟和我分家产。”
LUKE|12|14|耶稣对他说：“你这个人！谁立我作你们的判官，或给你们分家产的呢？”
LUKE|12|15|于是他对他们说：“你们要谨慎自守，躲避一切的贪心，因为人的生命不在于家道丰富。”
LUKE|12|16|然后他用比喻对他们说：“有一个财主，田地出产丰富。
LUKE|12|17|他自己心里想：‘我的出产没有地方储藏，怎么办呢？’
LUKE|12|18|就说：‘我要这么办：要把我的仓库拆了，另盖更大的，在那里好储藏我一切的粮食和财物，
LUKE|12|19|然后要对我自己说：你这个人哪，你有许多财物积存，可供多年享用，只管安安逸逸吃喝快乐吧！’
LUKE|12|20|上帝却对他说：‘无知的人哪！今夜就要你的性命，你所预备的要归谁呢？’
LUKE|12|21|凡为自己积财，在上帝面前却不富足的，也是这样。”
LUKE|12|22|耶稣又对门徒说：“所以，我告诉你们，不要为生命忧虑吃什么，为身体忧虑穿什么。
LUKE|12|23|因为生命胜于饮食，身体胜于衣裳。
LUKE|12|24|你们想一想乌鸦：它们既不种也不收，既没有仓又没有库，上帝尚且养活它们。你们比飞鸟要贵重得多呢！
LUKE|12|25|你们哪一个能藉着忧虑使寿数多加一刻呢 ？
LUKE|12|26|这最小的事你们尚且不能做，何必忧虑其余的事呢？
LUKE|12|27|你们想一想百合花是怎么长起来的：它也不劳动，也不纺线。然而我告诉你们，就是 所罗门 极荣华的时候，他所穿戴的还不如这些花的一朵呢！
LUKE|12|28|你们这小信的人哪！野地里的草今天还在，明天就丢在炉里，上帝还给它这样的妆饰，何况你们呢？
LUKE|12|29|你们不要求吃什么，喝什么，也不要挂虑。
LUKE|12|30|这都是世上的外邦人所求的；你们需要这些东西，你们的父都知道。
LUKE|12|31|你们只要求他的国，这些东西就必加给你们了。
LUKE|12|32|你们这小群，不要惧怕，因为你们的父乐意把国赐给你们。
LUKE|12|33|你们要变卖财产周济人，为自己预备永不坏的钱囊和用不尽的财宝在天上，就是贼不能近，虫不能蛀的地方。
LUKE|12|34|因为你们的财宝在哪里，你们的心也在哪里。”
LUKE|12|35|“你们要束紧腰带，灯也要点着，
LUKE|12|36|好像仆人等候自己的主人从婚宴上回来。他来叩门，就立刻给他开门。
LUKE|12|37|主人来了，看见仆人警醒，那些仆人就有福了。我实在告诉你们，主人会叫他们坐席，自己束上腰带，前来伺候他们。
LUKE|12|38|他或是半夜来，或是天亮之前来，看见仆人这样，那些仆人就有福了。
LUKE|12|39|你们要知道，一家的主人若知道贼什么时候来，就 不容贼挖穿房屋。
LUKE|12|40|你们也要预备，因为在你们想不到的时候，人子就来了。”
LUKE|12|41|彼得 说：“主啊，这比喻是对我们说的呢？还是也对众人呢？”
LUKE|12|42|主说：“那么，谁是那忠心又精明的管家，主人要派他管理自己的家仆，按时定量分粮给他们的呢？
LUKE|12|43|主人来到，看见仆人这样做，那仆人就有福了。
LUKE|12|44|我实在告诉你们，主人要派他管理所有的财产。
LUKE|12|45|如果那仆人心里说‘我的主人会来得迟’，就动手打僮仆和使女，并且吃喝醉酒，
LUKE|12|46|在想不到的日子，不知道的时候，那仆人的主人要来，重重地惩罚他 ，定他和不忠心的人同罪。
LUKE|12|47|仆人知道主人的意思，却没预备，又未顺他的意思做，那仆人要多受责打；
LUKE|12|48|至于那不知道而做了当受责打的事的，要少受责打。多给谁，就向谁多取；多托谁，就向谁多要。”
LUKE|12|49|“我来是要把火丢在地上，假如已经烧起来，不也是我所希望的吗？
LUKE|12|50|我有当受的洗还没有受，在这事完成之前，我是多么地焦急！
LUKE|12|51|你们以为我来是要使地上太平吗？不！我告诉你们，是使人纷争。
LUKE|12|52|从今以后，一家五个人将要纷争，三个和两个相争，两个和三个相争：
LUKE|12|53|父亲和儿子相争， 儿子和父亲相争； 母亲和女儿相争， 女儿和母亲相争； 婆婆和媳妇相争， 媳妇和婆婆相争。”
LUKE|12|54|耶稣又对众人说：“你们看见西边起了云彩，就说：‘要下大雨了’，果然就有；
LUKE|12|55|起了南风，你们就说：‘要燥热了’，也就有了。
LUKE|12|56|假冒为善的人哪，你们知道分辨天地的气象，怎么不知道分辨这是什么时代呢？”
LUKE|12|57|“你们又为何不自己判断什么是合理的呢？
LUKE|12|58|你同告你的冤家去见官，还在路上，要尽力跟他和解，免得他拉你到法官面前，法官把你交给法警，法警把你下在监里。
LUKE|12|59|我告诉你，就是最后一小文钱 还没有还清，你也绝不能从那里出来。”
LUKE|13|1|正当那时，有些在场的人把 彼拉多 使 加利利 人的血搀杂在他们祭物中的事，告诉耶稣。
LUKE|13|2|耶稣对他们说：“你们以为这些 加利利 人比其他的 加利利 人更有罪，所以受这害吗？
LUKE|13|3|我告诉你们，不是的！你们若不悔改，都同样要灭亡！
LUKE|13|4|从前 西罗亚 楼倒塌，压死了十八个人，你们以为那些人比一切住在 耶路撒冷 的人更有罪吗？
LUKE|13|5|我告诉你们，不是的！你们若不悔改，都照样要灭亡！”
LUKE|13|6|于是，耶稣用比喻说：“有一个人在葡萄园里栽了一棵无花果树。他前来在树上找果子，却找不到，
LUKE|13|7|就对园丁说：‘看哪，我这三年来到这棵无花果树前找果子，竟找不到。把它砍了吧，何必白占土地呢？’
LUKE|13|8|园丁回答：‘主啊，今年且留着，等我在树周围掘开土，加上肥料，
LUKE|13|9|以后若结果子便罢，不然再把它砍了。’”
LUKE|13|10|安息日，耶稣在一个会堂里教导人。
LUKE|13|11|有一个女人被灵附身，病了十八年，腰弯得一点都直不起来。
LUKE|13|12|耶稣看见，就叫她过来，对她说：“妇人，你的病好了！”
LUKE|13|13|于是用双手按着她，她立刻直起腰来，就归荣耀给上帝。
LUKE|13|14|会堂的主管因为耶稣在安息日治病，就很生气，对众人说：“有六天应当做工，那六天之内可以来求医，在安息日却不可。”
LUKE|13|15|主回答他：“假冒为善的人哪，难道你们各人在安息日不解开槽上的牛和驴，牵去喝水吗？
LUKE|13|16|何况她本是 亚伯拉罕 的后裔，被撒但捆绑了十八年，不该在安息日这天解开她的绑吗？”
LUKE|13|17|耶稣说这些话，他的敌人都惭愧了；所有的人因他所做一切荣耀的事都很欢喜。
LUKE|13|18|耶稣说：“上帝的国像什么？我拿什么来比拟呢？
LUKE|13|19|它好比一粒芥菜种，有人拿去种在园子里，长大成树，天上的飞鸟在它的枝上筑巢。”
LUKE|13|20|他又说：“我拿什么来比拟上帝的国呢？
LUKE|13|21|它好比面酵，有妇人拿来放进三斗面里，直到全团都发起来。”
LUKE|13|22|耶稣往 耶路撒冷 去，在所经过的各城各乡教导人。
LUKE|13|23|有一个人问他：“主啊，得救的人很少吧？” 耶稣对众人说：
LUKE|13|24|“你们要努力进窄门。我告诉你们，将来有许多人想要进去，却不能。
LUKE|13|25|等到一家之主起来关了门，你们才站在外面敲门，说：‘主啊，给我们开门！’他要回答你们说：‘我不认识你们，不知道你们是哪里来的。’
LUKE|13|26|那时，你们要说：‘我们在你面前吃过喝过，你也在我们的街上教导过人。’
LUKE|13|27|他要对你们说：‘我 告诉你们，我不知道你们是哪里来的。你们这一切不义的人，给我走开！’
LUKE|13|28|你们要看见 亚伯拉罕 、 以撒 、 雅各 和众先知都在上帝的国里，你们却被赶到外面，在那里要哀哭切齿了。
LUKE|13|29|从东从西，从南从北，将有人来，在上帝的国里坐席。
LUKE|13|30|看吧，在后的，将要在前；在前的，将要在后。”
LUKE|13|31|就在那时，有几个法利赛人来对耶稣说：“离开这里到别处去吧，因为 希律 想要杀你。”
LUKE|13|32|耶稣对他们说：“你们去告诉那个狐狸：‘你看吧，今天明天我赶鬼治病，第三天我的事就成了。’
LUKE|13|33|虽然这样，今天明天后天我必须向前走，因为先知是不可能在 耶路撒冷 之外被害的。
LUKE|13|34|耶路撒冷 啊， 耶路撒冷 啊，你常杀害先知，又用石头打死那奉差遣到你这里来的人。我多少次想聚集你的儿女，好像母鸡把小鸡聚集在翅膀底下，可是你们不愿意。
LUKE|13|35|看吧，你们的家要被废弃。我告诉你们，你们绝不会再见到我，直到你们说：‘奉主名来的是应当称颂的！’”
LUKE|14|1|安息日，耶稣到一个法利赛人的领袖家里去吃饭，他们就窥探他。
LUKE|14|2|这时在他面前有一个患水肿病的人。
LUKE|14|3|耶稣回答律法师和法利赛人，说：“安息日治病合不合法？”
LUKE|14|4|他们却不说话。耶稣扶着那人，治好了他，叫他走了。
LUKE|14|5|耶稣对他们说：“你们中间谁有儿子 或有牛在安息日掉在井里，不立刻拉他上来呢？”
LUKE|14|6|他们对这些事不能反驳。
LUKE|14|7|耶稣见所请的客人选择首位，就用比喻对他们说：
LUKE|14|8|“你被人请去赴婚宴，不要坐在首位上，恐怕主人请了比你尊贵的客人，
LUKE|14|9|请了你和他的那人前来，对你说：‘请让座给这一位吧。’你就羞羞惭惭地退到末位去了。
LUKE|14|10|你被请的时候，去坐在末位上，好让主人来对你说：‘朋友，请上座。’那时，你在同席的人面前就有光彩了。
LUKE|14|11|因为凡自高的，必降为卑；自甘卑微的，必升为高。”
LUKE|14|12|耶稣又对请他的人说：“你准备午饭或晚餐，不要请你的朋友、弟兄、亲属和富足的邻舍，免得他们回请你，你就得了报答。
LUKE|14|13|你摆设宴席，倒要请那贫穷的、残疾的、瘸腿的、失明的，
LUKE|14|14|你就有福了！因为他们没有什么可报答你。到义人复活的时候，你要得到报答。”
LUKE|14|15|同席的有一人听见这些话，就对耶稣说：“在上帝国里吃饭的有福了！”
LUKE|14|16|耶稣对他说：“有人摆设大宴席，请了许多客人。
LUKE|14|17|到了坐席的时候，他打发仆人去对所请的人说：‘请来吧！样样都已齐备了。’
LUKE|14|18|众人异口同声地推辞。头一个对他说：‘我买了一块地，必须去看看。请你准我辞了。’
LUKE|14|19|另一个说：‘我买了五对牛，要去试一试。请你准我辞了。’
LUKE|14|20|又有一个说：‘我才娶了妻子，所以不能去。’
LUKE|14|21|那仆人回来，把这些事都告诉了主人。这家的主人就发怒，对仆人说：‘快出去，到城里大街小巷，领那贫穷的、残疾的、失明的、瘸腿的来。’
LUKE|14|22|仆人说：‘主啊，你所吩咐的已经办了，还有空位。’
LUKE|14|23|主人对仆人说：‘你出去，到大街小巷强拉人进来，坐满我的屋子。
LUKE|14|24|我告诉你们，先前所请的人没有一个可以尝到我的宴席。’”
LUKE|14|25|有一大群人和耶稣同行。他转过来对他们说：
LUKE|14|26|“无论什么人到我这里来，若不爱我胜过爱 自己的父母、妻子、儿女、兄弟、姊妹，甚至自己的性命，就不能作我的门徒。
LUKE|14|27|凡不背着自己的十字架来跟从我的，也不能作我的门徒。
LUKE|14|28|你们哪一个要盖一座楼，不先坐下来计算费用，看能不能盖成？
LUKE|14|29|免得安了地基，不能盖成，看见的人都笑话他，说：
LUKE|14|30|‘这个人开了工，却不能完工。’
LUKE|14|31|或是一个王出去和别的王打仗，岂不先坐下来酌量，他能不能用一万兵去抵抗那领二万兵来攻打他的吗？
LUKE|14|32|若是不能，他就趁敌人还远的时候，派使者去谈和平的条件。
LUKE|14|33|这样，你们无论什么人，若不撇下一切所有的，就不能作我的门徒。”
LUKE|14|34|“盐本是好的；盐若失了味，怎能叫它再咸呢？
LUKE|14|35|或用在田里，或堆在粪里，都不合适，只好丢在外面。有耳可听的，就应当听！”
LUKE|15|1|许多税吏和罪人都挨近耶稣，要听他讲道。
LUKE|15|2|法利赛人和文士私下议论说：“这个人接纳罪人，又同他们吃饭。”
LUKE|15|3|耶稣就用比喻对他们说：
LUKE|15|4|“你们中间谁有一百只羊，失去其中的一只，不把这九十九只留在旷野，去找那失去的羊，直到找着呢？
LUKE|15|5|找到了，他就欢欢喜喜地把羊扛在肩上。
LUKE|15|6|他回到家里，请朋友和邻舍来，对他们说：‘你们和我一同欢喜吧，我失去的羊已经找到了！’
LUKE|15|7|我告诉你们，一个罪人悔改，在天上也要这样为他欢喜，比为九十九个不用悔改的义人欢喜还大呢！”
LUKE|15|8|“同样，哪一个妇人有十块钱 ，若失落一块，不点上灯，打扫屋子，细细地找，直到找着呢？
LUKE|15|9|找到了，她就请朋友和邻舍来，对她们说：‘你们和我一同欢喜吧，我失落的那块钱已经找到了！’
LUKE|15|10|我告诉你们，一个罪人悔改，上帝的使者也是这样为他欢喜。”
LUKE|15|11|耶稣又说：“一个人有两个儿子。
LUKE|15|12|小儿子对父亲说：‘父亲，请你把我应得的家业分给我。’他父亲就把财产分给他们。
LUKE|15|13|过了不多几天，小儿子把他一切所有的都收拾起来，往远方去了。在那里，他任意放荡，浪费钱财。
LUKE|15|14|他耗尽了一切所有的，又恰逢那地方有大饥荒，就穷困起来。
LUKE|15|15|于是他去投靠当地的一个居民，那人打发他到田里去放猪。
LUKE|15|16|他恨不得拿猪所吃的豆荚充饥，也没有人给他什么吃的。
LUKE|15|17|他醒悟过来，就说：‘我父亲有多少雇工，粮食有余，我倒在这里饿死吗？
LUKE|15|18|我要起来，到我父亲那里去，对他说：父亲！我得罪了天，又得罪了你，
LUKE|15|19|从今以后，我不配称为你的儿子，把我当作一个雇工吧。’
LUKE|15|20|于是他起来，往他父亲那里去。相离还远，他父亲看见，就动了慈心，跑去拥抱着他，连连亲他。
LUKE|15|21|儿子对他说：‘父亲！我得罪了天，又得罪了你，从今以后，我不配称为你的儿子。’
LUKE|15|22|父亲却吩咐仆人：‘快把那上好的袍子拿出来给他穿，把戒指戴在他指头上，把鞋穿在他脚上，
LUKE|15|23|把那肥牛犊牵来宰了，我们来吃喝庆祝；
LUKE|15|24|因为我这个儿子是死而复活，失而复得的。’他们就开始庆祝。
LUKE|15|25|“那时，大儿子正在田里。他回来，离家不远时，听见奏乐跳舞的声音，
LUKE|15|26|就叫一个僮仆来，问是什么事。
LUKE|15|27|僮仆对他说：‘你弟弟回来了，你父亲因为他无灾无病地回来，把肥牛犊宰了。’
LUKE|15|28|大儿子就生气，不肯进去，他父亲出来劝他。
LUKE|15|29|他对父亲说：‘你看，我服侍你这么多年，从来没有违背过你的命令，而你从来没有给我一只小山羊，叫我和朋友们一同快乐。
LUKE|15|30|但你这个儿子和娼妓吃光了你的财产，他一回来，你倒为他宰了肥牛犊。’
LUKE|15|31|父亲对他说：‘儿啊！你常和我同在，我所有的一切都是你的；
LUKE|15|32|可是你这个弟弟是死而复活，失而复得的，所以我们理当欢喜庆祝。’”
LUKE|16|1|耶稣又对门徒说：“某财主有一个管家，有人向主人告管家浪费他的财物。
LUKE|16|2|主人叫他来，对他说：‘我听到了，你做的是什么事？把你所经管的交代清楚，你不能再作我的管家了。’
LUKE|16|3|那管家心里说：‘主人辞我，不用我再作管家，我将来做什么呢？锄地嘛，没有力气；讨饭嘛，怕羞。
LUKE|16|4|我知道怎么做，好叫人们在我不作管家之后，接我到他们家里去。’
LUKE|16|5|于是他把欠他主人债的，一个一个地叫了来，问头一个说：‘你欠我主人多少？’
LUKE|16|6|他说：‘一百篓 油。’管家对他说：‘拿你的账，快坐下，写五十。’
LUKE|16|7|他问另一个说：‘你欠多少？’他说：‘一百石麦子。’管家对他说：‘拿你的账，写八十。’
LUKE|16|8|主人就夸奖这不义的管家做事精明，因为今世之子应付自己的世代比光明之子更加精明。
LUKE|16|9|我又告诉你们，要藉着那不义的钱财结交朋友，到了钱财无用的时候，他们可以接你们到永远的住处 去。
LUKE|16|10|人在最小的事上忠心，在大事上也忠心；在最小的事上不义，在大事上也不义。
LUKE|16|11|若是你们在不义的钱财上不忠心，谁还把那真实的钱财托付你们呢？
LUKE|16|12|如果你们在别人的东西上不忠心，谁还把你们自己的东西给你们呢？
LUKE|16|13|一个仆人不能服侍两个主；他不是恨这个爱那个，就是重这个轻那个。你们不能又服侍上帝，又服侍 玛门 。”
LUKE|16|14|法利赛人是贪爱钱财的；他们听见这一切话，就嘲笑耶稣。
LUKE|16|15|耶稣对他们说：“你们是在人面前自称为义的，你们的心，上帝却知道；因为人以为尊贵的，是上帝看为可憎恶的。
LUKE|16|16|律法和先知到 约翰 为止，从此上帝国的福音传开了，人人努力要进去。
LUKE|16|17|天地废去比律法的一点一画落空还要容易。
LUKE|16|18|凡休妻另娶的，就是犯奸淫；娶被丈夫休了的妇人的，也是犯奸淫。”
LUKE|16|19|“有一个财主穿着紫色袍和细麻布衣服，天天奢华宴乐。
LUKE|16|20|又有一个讨饭的，名叫 拉撒路 ，浑身长疮，被人放在财主门口，
LUKE|16|21|想得财主桌子上掉下来的碎食充饥，甚至还有狗来舔他的疮。
LUKE|16|22|后来那讨饭的死了，被天使带去放在 亚伯拉罕 的怀里。财主也死了，并且埋葬了。
LUKE|16|23|他在阴间受苦，举目远远地望见 亚伯拉罕 ，又望见 拉撒路 在他怀里，
LUKE|16|24|他就喊着说：‘我祖 亚伯拉罕 哪，可怜我吧！请打发 拉撒路 来，用指头尖蘸点水，凉凉我的舌头，因为我在这火焰里，极其痛苦。’
LUKE|16|25|亚伯拉罕 说：‘孩子啊，你该回想你生前享过福， 拉撒路 也同样受过苦，如今他在这里得安慰，你却受痛苦。
LUKE|16|26|除此之外，在你们和我们之间，有深渊隔开，以致人要从这边过到你们那边是不可能的；要从那边过到这边也是不可能的。’
LUKE|16|27|财主说：‘我祖啊，既然这样，求你打发 拉撒路 到我父家去，
LUKE|16|28|因为我还有五个兄弟，他可以警告他们，免得他们也来到这痛苦的地方。’
LUKE|16|29|亚伯拉罕 说：‘他们有 摩西 和先知的话可以听从。’
LUKE|16|30|他说：‘不！我祖 亚伯拉罕 哪，假如有一个人从死人中到他们那里去，他们一定会悔改。’
LUKE|16|31|亚伯拉罕 对他说：‘如果他们不听从 摩西 和先知的话，就是有人从死人中复活，他们也不会信服的。’”
LUKE|17|1|耶稣又对门徒说：“绊倒人的事是免不了的，但那绊倒人的有祸了！
LUKE|17|2|人若把这些小子中的一个绊倒的，还不如把磨石拴在他的颈项上，丢在海里。
LUKE|17|3|你们要谨慎！若是你的弟兄犯罪，就劝戒他；他若懊悔，就饶恕他。
LUKE|17|4|如果他一天七次得罪你，又七次回头，说：‘我懊悔了’，你总要饶恕他。”
LUKE|17|5|使徒对主说：“请加增我们的信心。”
LUKE|17|6|主说：“你们若有信心像一粒芥菜种，就是对这棵桑树说：‘你要连根拔起，栽在海里’，它也会听从你们。”
LUKE|17|7|“你们当中谁有仆人耕地或是放羊，从田里回来，就对他说‘你快来坐下吃饭’呢？
LUKE|17|8|他岂不对仆人说‘你给我预备晚饭，束上带子伺候我，等我吃喝完了，你才可以吃喝’吗？
LUKE|17|9|仆人照所吩咐的去做，主人还谢谢他吗？
LUKE|17|10|这样，你们做完了一切所吩咐的，要说：‘我们是无用的仆人，所做的本是我们该做的。’”
LUKE|17|11|耶稣往 耶路撒冷 去，经过 撒玛利亚 和 加利利 中间的地区。
LUKE|17|12|他进入一个村子，有十个痲疯病人迎面而来，远远地站着，
LUKE|17|13|高声说：“耶稣，老师啊，可怜我们吧！”
LUKE|17|14|耶稣看见，就对他们说：“你们去，把身体给祭司检查。”他们正去的时候就洁净了。
LUKE|17|15|其中有一个见自己已经好了，就回来大声归荣耀给上帝，
LUKE|17|16|又俯伏在耶稣脚前感谢他。这人是 撒玛利亚 人。
LUKE|17|17|耶稣回答说：“洁净了的不是十个人吗？那九个在哪里呢？
LUKE|17|18|除了这外族人，再没有别人回来归荣耀给上帝吗？”
LUKE|17|19|于是他对那人说：“起来，走吧，你的信救了你！”
LUKE|17|20|法利赛人问：“上帝的国几时来到？”耶稣回答：“上帝的国来到，不是眼睛看得见的。
LUKE|17|21|人也不能说：‘看哪，在这里！’或说：‘在那里！’因为上帝的国就在你们心里 。”
LUKE|17|22|他又对门徒说：“那些日子将到，你们渴望能看见人子的一个日子，却看不见。
LUKE|17|23|有人要对你们说：‘看哪，在那里！’或说：‘看哪，在这里！’你们不要出去，也不要追随他们。
LUKE|17|24|好像闪电从天这边一闪直照到天那边，人子在他的日子 也要这样。
LUKE|17|25|可是他必须先受许多苦，又被这世代所弃绝。
LUKE|17|26|挪亚 的日子怎样，人子的日子也要怎样。
LUKE|17|27|那时，人又吃又喝，又娶又嫁，直到 挪亚 进方舟的那日，洪水就来，把他们全都灭了。
LUKE|17|28|同样，就像在 罗得 的日子，人又吃又喝，又买又卖，又耕种又建造，
LUKE|17|29|到 罗得 离开 所多玛 的那日，有火与硫磺从天上降下来，把他们全都灭了。
LUKE|17|30|人子显现的日子也要这样。
LUKE|17|31|在那日，人在屋顶上，东西在屋里，不要下来拿；人在田里，也不要回家。
LUKE|17|32|你们想想 罗得 的妻子吧！
LUKE|17|33|凡想保全性命的，要丧失性命；凡丧失性命的，要保存性命。
LUKE|17|34|我告诉你们，在那一夜，两个人在一张床上，一个被接去，一个被撇下。
LUKE|17|35|两个女人一同推磨，一个被接去，一个被撇下。 ”
LUKE|17|36|
LUKE|17|37|门徒回答他说：“主啊，在哪里呢？”耶稣对他们说：“尸首在哪里，鹰也会聚在哪里。”
LUKE|18|1|耶稣对门徒讲了一个比喻，为了要他们常常祷告，不可灰心。
LUKE|18|2|他说：“某城有一个官，不惧怕上帝，也不尊重人。
LUKE|18|3|那城里有个寡妇，常到他那里，说：‘我有一个冤家，求你给我伸冤。’
LUKE|18|4|他很久不受理，后来心里说：‘我虽不惧怕上帝，也不尊重人，
LUKE|18|5|只因这寡妇烦扰我，我就给她伸冤吧，免得她常来纠缠我。’”
LUKE|18|6|主说：“你们听这不义的官所说的话。
LUKE|18|7|上帝的选民昼夜呼吁他，他岂会延迟不给他们伸冤吗？
LUKE|18|8|我告诉你们，他很快就要给他们伸冤。然而，人子来的时候，能在世上找到这样的信德吗？”
LUKE|18|9|耶稣向那些自以为义而藐视别人的人讲了这比喻：
LUKE|18|10|“有两个人上圣殿去祷告，一个是法利赛人，一个是税吏。
LUKE|18|11|法利赛人独自站着，自言自语地祷告说：‘上帝啊，我感谢你，我不像别人勒索、不义、奸淫，也不像这个税吏。
LUKE|18|12|我每周禁食两次，凡我所得的都献上十分之一。’
LUKE|18|13|那税吏远远地站着，连举目望天也不敢，只捶着胸，说：‘上帝啊，开恩可怜我这个罪人！’
LUKE|18|14|我告诉你们，这人回家去比那人倒算为义了。因为凡自高的，必降为卑；自甘卑微的，必升为高。”
LUKE|18|15|有人甚至连婴孩也带来见耶稣，要他摸他们，门徒看见就责备那些人。
LUKE|18|16|耶稣却叫他们来，说：“让小孩子到我这里来，不要阻止他们，因为在上帝国的正是这样的人。
LUKE|18|17|我实在告诉你们，凡要接受上帝国的，若不像小孩子，绝不能进去。”
LUKE|18|18|有一个官问耶稣说：“善良的老师，我该做什么事才能承受永生？”
LUKE|18|19|耶稣对他说：“你为什么称我是善良的？除了上帝一位之外，再没有善良的。
LUKE|18|20|诫命你是知道的：‘不可奸淫；不可杀人；不可偷盗；不可作假见证；当孝敬父母。’”
LUKE|18|21|那人说：“这一切我从小都遵守了。”
LUKE|18|22|耶稣听见了，就对他说：“你还缺少一件：要变卖你一切所有的，分给穷人，就必有财宝在天上；你还要来跟从我。”
LUKE|18|23|他听见这些话，就很忧愁，因为他很富有。
LUKE|18|24|耶稣见他变得很忧愁 ，就说：“有钱财的人进上帝的国是何等的难哪！
LUKE|18|25|骆驼穿过针眼比财主进上帝的国还容易呢！”
LUKE|18|26|听见的人说：“这样，谁能得救呢？”
LUKE|18|27|耶稣说：“在人所不能的事，在上帝都能。”
LUKE|18|28|彼得 说：“看哪，我们已经撇下自己所有的跟从你了。”
LUKE|18|29|耶稣对他们说：“我实在告诉你们，凡是为上帝的国撇下房屋，或是妻子、兄弟、父母、儿女的，
LUKE|18|30|没有不在今世得更多倍，而在来世得永生的。”
LUKE|18|31|耶稣把十二使徒带到一边，对他们说：“看哪，我们上 耶路撒冷 去，先知所写的一切事都要成就在人子身上。
LUKE|18|32|他将被交给外邦人；他们要戏弄他，凌辱他，向他吐唾沫，
LUKE|18|33|并要鞭打他，杀害他；第三天他要复活。”
LUKE|18|34|这些事门徒一点也不明白，这话的意思对他们是隐藏的；他们不知道所说的是什么。
LUKE|18|35|耶稣将近 耶利哥 的时候，有一个盲人坐在路旁讨饭。
LUKE|18|36|他听见许多人经过，就问是什么事。
LUKE|18|37|他们告诉他，是 拿撒勒 人耶稣经过。
LUKE|18|38|他就呼叫说：“ 大卫 之子耶稣啊，可怜我吧！”
LUKE|18|39|在前头走的人就责备他，不许他作声，他却越发喊叫：“ 大卫 之子啊，可怜我吧！”
LUKE|18|40|耶稣就站住，吩咐把他领过来，他到了跟前，就问他：
LUKE|18|41|“你要我为你做什么？”他说：“主啊，我要能看见。”
LUKE|18|42|耶稣对他说：“你看见吧！你的信救了你。”
LUKE|18|43|那盲人立刻看得见了，就跟随耶稣，一路归荣耀给上帝。众人看见这事，也都赞美上帝。
LUKE|19|1|耶稣进了 耶利哥 ，要从那里经过。
LUKE|19|2|有一个人名叫 撒该 ，作税吏长，是个财主。
LUKE|19|3|他要看看耶稣是怎样的人，只因人多，他的身材又矮，所以看不见。
LUKE|19|4|于是他跑到前头，爬上桑树，要看耶稣，因为耶稣要从那里经过。
LUKE|19|5|耶稣到了那里，抬头一看，对他说：“ 撒该 ，快下来！今天我必须住在你家里。”
LUKE|19|6|他就急忙下来，欢欢喜喜地接待耶稣。
LUKE|19|7|众人看见，都私下议论说：“他竟然到罪人家里去住宿。”
LUKE|19|8|撒该 站着对主说：“主啊，我把所有的一半给穷人；我若勒索了谁，就还他四倍。”
LUKE|19|9|耶稣对他说：“今天救恩到了这家，因为他也是 亚伯拉罕 的子孙。
LUKE|19|10|人子来是要寻找和拯救失丧的人。”
LUKE|19|11|众人正听见这些话的时候，耶稣因为将近 耶路撒冷 ，又因他们以为上帝的国快要显现，就接着讲了一个比喻，
LUKE|19|12|说：“有一个贵族往远方去，为要取得王位，然后回来。
LUKE|19|13|他叫了自己的十个仆人来，交给他们十锭银子，说：‘你们去做生意，直到我回来。’
LUKE|19|14|他本国的百姓却恨他，打发使者随后去，说：‘我们不愿意这个人作我们的王。’
LUKE|19|15|他得了王位回来，就吩咐叫那领了银子的仆人来，要知道他们做生意赚了多少。
LUKE|19|16|头一个上来，说：‘主啊，你的一锭银子已经赚了十锭。’
LUKE|19|17|主人对他说：‘好，我善良的仆人，你既在最小的事上忠心，你有权柄管十座城。’
LUKE|19|18|第二个来，说：‘主啊，你的一锭银子已经赚了五锭。’
LUKE|19|19|主人也对这个说：‘你管五座城。’
LUKE|19|20|又有一个来说：‘主啊！看哪，你的一锭银子在这里，我把它包在手巾里存着。
LUKE|19|21|我向来怕你，因为你是严厉的人：没有放的，也要去拿；没有种的，也要去收。’
LUKE|19|22|主人对他说：‘你这恶仆，我要凭你的话定你的罪。你既知道我是严厉的人，没有放的也去拿，没有种的也去收，
LUKE|19|23|为什么不把我的银子存在银行，等我来的时候，连本带利都取回来呢？’
LUKE|19|24|于是他对那些站在旁边的人说：‘把他这一锭夺过来，给那有十锭的。’
LUKE|19|25|他们对他说：‘主啊，他已经有十锭了。’
LUKE|19|26|主人说：‘我告诉你们，凡有的，还要给他；没有的，连他所有的也要夺过来。
LUKE|19|27|至于我那些仇敌，不要我作他们王的，把他们拉来，在我面前杀了！’”
LUKE|19|28|耶稣说完了这些话，就走在前面，上 耶路撒冷 去。
LUKE|19|29|快到 伯法其 和 伯大尼 ，在名叫 橄榄山 的地方，他打发两个门徒，
LUKE|19|30|说：“你们往对面村子里去，进去的时候会看见一匹驴驹拴在那里，是从来没有人骑过的，把它解开，牵来。
LUKE|19|31|若有人问为什么解开它，你们就这样说：‘主要用它。’”
LUKE|19|32|被打发的人去了，所遇见的正如耶稣对他们所说的。
LUKE|19|33|他们解开驴驹的时候，主人问他们：“为什么解开驴驹？”
LUKE|19|34|他们说：“主要用它。”
LUKE|19|35|他们把驴驹牵到耶稣那里，把自己的衣服搭在上面，扶耶稣骑上。
LUKE|19|36|他前进的时候，众人把衣服铺在路上。
LUKE|19|37|他将近 耶路撒冷 ，正下 橄榄山 的时候，一大群门徒因所见过的一切异能，都欢呼起来，大声赞美上帝，
LUKE|19|38|说： “奉主名来的王 是应当称颂的！ 在天上有和平； 在至高之处有荣光。”
LUKE|19|39|人群中有几个法利赛人对耶稣说：“老师，责备你的门徒吧！”
LUKE|19|40|耶稣回答：“我告诉你们，若是这些人闭口不说，石头也要呼叫起来。”
LUKE|19|41|耶稣快到 耶路撒冷 ，看见那城，就为它哀哭，
LUKE|19|42|说：“但愿你在这日子知道有关你平安的事，不过这事现在是隐藏的，你的眼睛看不出来。
LUKE|19|43|因为日子将到，你的仇敌要筑起土垒包围你，四面困住你，
LUKE|19|44|并要消灭你和你里头的儿女，连一块石头也不留在另一块石头上，因为你不知道你蒙眷顾的时候。”
LUKE|19|45|耶稣一进圣殿就赶出在里面做买卖的人，
LUKE|19|46|对他们说：“经上说： ‘我的殿是祷告的殿， 你们倒使它成为贼窝了。’”
LUKE|19|47|耶稣天天在圣殿里教导人。祭司长、文士和百姓的领袖都想杀他，
LUKE|19|48|但找不出方法来，因为百姓都侧耳听他。
LUKE|20|1|有一天，耶稣在圣殿里教导百姓，宣讲福音的时候，祭司长、文士和长老上前来，
LUKE|20|2|问他说：“你告诉我们，你仗着什么权柄做这些事？给你这权柄的是谁呢？”
LUKE|20|3|耶稣回答他们：“我也要问你们一句话，你们告诉我。
LUKE|20|4|约翰 的洗礼是从天上来的，还是从人间来的呢？”
LUKE|20|5|他们彼此商量说：“我们若说‘从天上来的’，他会说‘这样，你们为什么不信他呢？’
LUKE|20|6|我们若说‘从人间来的’，所有的百姓都会用石头打死我们，因为他们信 约翰 是先知。”
LUKE|20|7|于是他们回答：“我们不知道是从哪里来的。”
LUKE|20|8|耶稣对他们说：“我也不告诉你们，我仗着什么权柄做这些事。”
LUKE|20|9|耶稣用这个比喻对百姓说：“有人开垦了一个葡萄园，租给园户，就出外远行，去了许久。
LUKE|20|10|到了时候，他打发一个仆人到园户那里去，叫他们把园中当纳的果子交给他；园户竟打了他，叫他空手回去。
LUKE|20|11|园主又打发另一个仆人去，他们也打了他，并且侮辱他，叫他空手回去。
LUKE|20|12|园主又打发第三个仆人去，他们也打伤了他，把他推出去了。
LUKE|20|13|葡萄园主说：‘我要怎么做呢？我要打发我的爱子去，或许他们会尊敬他。’
LUKE|20|14|可是，园户看见他，彼此说：‘这是承受产业的。我们杀了他，产业就归我们了！’
LUKE|20|15|于是他们把他扔出葡萄园外，杀了。这样，葡萄园主要怎么处置他们呢？
LUKE|20|16|他要来除灭那些园户，将葡萄园转给别人。”听见的人说：“绝对不可！”
LUKE|20|17|耶稣看着他们，说：“那么，经上记着： ‘匠人所丢弃的石头 已作了房角的头块石头。’ 这是什么意思呢？
LUKE|20|18|凡跌在那石头上的，一定会跌得粉碎；那石头掉在谁的身上，就要把谁压得稀烂。”
LUKE|20|19|文士和祭司长看出这比喻是指着他们说的，当时就想要下手拿他，只是惧怕百姓。
LUKE|20|20|于是他们窥探耶稣，打发奸细装作好人，要在他的话上抓把柄，好把他交给总督处置。
LUKE|20|21|奸细就问耶稣：“老师，我们知道你所讲所教的都很正确，也不看人的面子，而是诚诚实实传上帝的道。
LUKE|20|22|我们纳税给凯撒合不合法？”
LUKE|20|23|耶稣看出他们的诡诈，就对他们说：
LUKE|20|24|“拿一个银币来给我看。这像和这名号是谁的？”他们说：“是凯撒的。”
LUKE|20|25|耶稣对他们说：“这样，凯撒的归凯撒，上帝的归上帝。”
LUKE|20|26|他们无法当着百姓在他的话上抓到把柄，又因他的对答而惊讶，就闭口不言了。
LUKE|20|27|有些撒都该人来见耶稣。他们说没有复活这回事，于是问耶稣：
LUKE|20|28|“老师， 摩西 为我们写下这话：‘某人的哥哥若死了，有妻无子，他该娶哥哥的妻子，为哥哥生子立后。’
LUKE|20|29|那么，有兄弟七人，第一个娶了妻，没有孩子死了。
LUKE|20|30|第二个、
LUKE|20|31|第三个也娶过她；同样地，七个人都娶过她，没有留下孩子就死了。
LUKE|20|32|后来，那妇人也死了。
LUKE|20|33|那么，在复活的时候，那妇人是哪一个的妻子呢？因为他们七个人都娶过她。”
LUKE|20|34|耶稣对他们说：“这世代的人有娶有嫁，
LUKE|20|35|惟有配得那要来的世代和从死人中复活的人不娶也不嫁。
LUKE|20|36|因为他们不能再死，和天使一样；既然是复活的人，他们就是上帝的儿子。
LUKE|20|37|至于死人复活， 摩西 在《荆棘篇》上就指明了，他称主是 亚伯拉罕 的上帝， 以撒 的上帝， 雅各 的上帝。
LUKE|20|38|上帝不是死人的上帝，而是活人的上帝，因为对他来说，人都是活的。”
LUKE|20|39|有几个文士说：“老师，你说得好。”
LUKE|20|40|以后，他们不敢再问他什么了。
LUKE|20|41|耶稣对他们说：“人们怎么说基督是 大卫 的后裔呢？
LUKE|20|42|《诗篇》 上 大卫 自己说： “主对我主说： ‘你坐在我的右边，
LUKE|20|43|等我使你的仇敌作你的脚凳。’
LUKE|20|44|大卫 既称他为主，他怎么又是 大卫 的后裔呢？”
LUKE|20|45|众百姓听的时候，耶稣对他的门徒说：
LUKE|20|46|“你们要防备文士。他们好穿长袍走来走去，喜欢人们在街市上向他们问安，又喜爱会堂里的高位，宴席上的首座。
LUKE|20|47|他们侵吞寡妇的家产，假意作很长的祷告。这些人要受更重的惩罚！”
LUKE|21|1|耶稣抬头观看，见财主把捐项投入圣殿银库，
LUKE|21|2|又见一个穷寡妇投了两个小文钱 ，
LUKE|21|3|就说：“我实在告诉你们，这穷寡妇所投的比众人更多。
LUKE|21|4|因为众人都是拿有余的捐献，但这寡妇，虽然自己不足，却把一生所有的都投进去了。”
LUKE|21|5|有人谈论圣殿是用美石和供物装饰的，耶稣就说：
LUKE|21|6|“你们所看见的这一切，日子将到，没有一块石头会留在另一块石头上而不被拆毁的。”
LUKE|21|7|他们问他：“老师，什么时候有这些事呢？这些事将临到的时候有什么预兆呢？”
LUKE|21|8|耶稣说：“你们要谨慎，不要受迷惑，因为将有好些人冒我的名来，说‘我是基督’，又说‘时候近了’，你们不要跟从他们！
LUKE|21|9|当你们听见打仗和动乱的事，不要惊惶；因为这些事必须先发生，但终结不会立刻就到。”
LUKE|21|10|于是耶稣对他们说：“民要攻打民，国要攻打国，
LUKE|21|11|将有大地震，多处必有饥荒、瘟疫，又有可怕的异象和大神迹从天上显现。
LUKE|21|12|但这一切的事以前，有人要下手拿你们，迫害你们，把你们交给会堂，并且关在监里，又为我名的缘故拉你们到君王和统治者面前。
LUKE|21|13|但这些事终必成为你们作见证的机会。
LUKE|21|14|所以，你们要立定心意，不要预先考虑怎样申辩；
LUKE|21|15|因为我必赐你们口才和智慧，是你们一切敌人所敌不住、驳不倒的。
LUKE|21|16|连你们的父母、兄弟、亲族、朋友也要把你们交给官府；你们中间也将有被他们害死的。
LUKE|21|17|你们要为我的名被众人憎恨。
LUKE|21|18|然而，你们连一根头发也不会损失。
LUKE|21|19|你们凭着坚忍，就必保全性命。”
LUKE|21|20|“当你们看见 耶路撒冷 被兵围困，就可知道它成为荒芜的日子近了。
LUKE|21|21|那时，在 犹太 的，应当逃到山上；在城里的，应当出来；在乡下的，不要进城。
LUKE|21|22|因为这是报应的日子，要使经上所写的都得应验。
LUKE|21|23|在那些日子，怀孕的和奶孩子的就苦了。因为将有大灾难降在这地方，也有愤怒临到这百姓。
LUKE|21|24|他们要倒在刀下，又被掳到各国去。 耶路撒冷 要被外邦人践踏，直到外邦人的日子满了。”
LUKE|21|25|“日月星辰要显出预兆，地上的邦国也有困苦，因海中波浪的响声而惶惶不安。
LUKE|21|26|人想到那要临到世界的事，就都吓得魂不附体，因为天上的万象都要震动。
LUKE|21|27|那时，他们要看见人子带着能力和大荣耀驾云来临。
LUKE|21|28|一有这些事，你们就当挺身昂首，因为你们得救赎的日子近了。”
LUKE|21|29|耶稣对他们讲了一个比喻说：“你们看无花果树和各样的树，
LUKE|21|30|树叶一长出来，你们看了自然就知道夏天近了。
LUKE|21|31|同样，当你们看见这些事发生，就知道上帝的国近了。
LUKE|21|32|我实在告诉你们，这世代还没有过去，一切都要发生。
LUKE|21|33|天地要废去，我的话却绝不废去。”
LUKE|21|34|“你们要谨慎，免得被贪食、醉酒和今生的忧虑压住你们的心，那日子就忽然临到你们，
LUKE|21|35|如同罗网一样，因为那日子要临到所有居住在地面上的人。
LUKE|21|36|你们要时时警醒，常常祈求，使你们能逃避这一切要来的事，得以站立在人子面前。”
LUKE|21|37|耶稣每日在圣殿里教导人，每夜出城到 橄榄山 住宿。
LUKE|21|38|众百姓清早上圣殿，到耶稣那里听他讲道。
LUKE|22|1|除酵节，又叫逾越节，近了。
LUKE|22|2|祭司长和文士在想法子怎样杀害耶稣，因他们惧怕百姓。
LUKE|22|3|这时，撒但入了那称为 加略 人 犹大 的心。他本是十二使徒里的一个。
LUKE|22|4|他去跟祭司长和守殿官商量怎样把耶稣交给他们。
LUKE|22|5|他们很高兴，就约定给他银子。
LUKE|22|6|他应允了，就找机会，要趁众人不在跟前的时候把耶稣交给他们。
LUKE|22|7|除酵节到了，这一天必须宰逾越节的羔羊。
LUKE|22|8|耶稣打发 彼得 和 约翰 ，说：“你们去为我们预备逾越节的宴席，好让我们吃。”
LUKE|22|9|他们问他：“你要我们在哪里预备？”
LUKE|22|10|耶稣对他们说：“你们进了城，会有人拿着一罐水迎面而来，你们就跟着他，到他所进的房子里去，
LUKE|22|11|对那家的主人说：‘老师问：客房在哪里？我和我的门徒要在那里吃逾越节的宴席。’
LUKE|22|12|他会带你们看一间摆设齐全的楼上大厅，你们就在那里预备。”
LUKE|22|13|他们去了，所看到的正如耶稣所说的。他们就预备了逾越节的宴席。
LUKE|22|14|时候到了，耶稣坐席，使徒们也和他同坐。
LUKE|22|15|耶稣对他们说：“我非常渴望在受害以前和你们吃这逾越节的宴席。
LUKE|22|16|我告诉你们，我不再吃这宴席，直到它实现在上帝的国里。”
LUKE|22|17|耶稣接过杯来，祝谢了，说：“你们拿这杯，大家分着喝。
LUKE|22|18|我告诉你们，从今以后，我不再喝这葡萄汁，直等上帝的国来到。”
LUKE|22|19|他又拿起饼来，祝谢了，就擘开，递给他们，说：“这是我的身体，为你们舍的，你们要如此行，为的是记念我。”
LUKE|22|20|饭后他照样拿起杯来，说：“这杯是用我的血所立的新约，为你们流出来的。
LUKE|22|21|但是，看哪，那出卖我的人的手跟我一同在桌子上。
LUKE|22|22|人子固然要照所预定的离去，但那出卖人子的人有祸了！”
LUKE|22|23|于是他们开始互相追问他们中间哪一个会做这事。
LUKE|22|24|门徒中间也起了争论：他们中哪一个可算为大。
LUKE|22|25|耶稣对他们说：“外邦人有君王为主治理他们，那掌权管他们的称为恩主。
LUKE|22|26|但你们不可这样。你们中间最大的，倒要成为最小的；为领袖的，倒要像服事人的。
LUKE|22|27|是谁为大？是坐席的还是服事人的呢？不是坐席的大吗？然而，我在你们中间是如同服事人的。
LUKE|22|28|“我在试炼之中，常和我同在的就是你们。
LUKE|22|29|我把国赐给你们，正如我父赐给我一样，
LUKE|22|30|使你们在我的国里坐在我的席上吃喝，并且坐在宝座上审判 以色列 十二个支派。”
LUKE|22|31|主又说：“ 西门 ， 西门 ！撒但要得着你们，好筛你们像筛麦子一样；
LUKE|22|32|但我已经为你祈求，使你不至于失了信心。你回头以后，要坚固你的弟兄。”
LUKE|22|33|彼得 对他说：“主啊，我已准备好要同你坐牢，与你同死。”
LUKE|22|34|耶稣说：“ 彼得 ，我告诉你，今日鸡还没有叫，你要三次说不认得我。”
LUKE|22|35|耶稣又对他们说：“我差你们出去的时候，没有钱囊，没有行囊，没有鞋子，你们缺少什么没有？”他们说：“没有。”
LUKE|22|36|耶稣对他们说：“但如今，有钱囊的要带着，有行囊的也一样；没有刀的要卖衣服买刀。
LUKE|22|37|我告诉你们，经上写着说：‘他被列在罪犯之中。’这话必须应验在我身上，因为那关于我的事必然成就。”
LUKE|22|38|他们说：“主啊，请看！这里有两把刀。”耶稣对他们说：“够了。”
LUKE|22|39|耶稣出来，照常往 橄榄山 去，门徒也跟随他。
LUKE|22|40|到了那地方，他就对他们说：“你们要祷告，免得陷入试探。”
LUKE|22|41|于是他离开他们约有一块石头扔出去那么远，跪下祷告，
LUKE|22|42|说：“父啊！你若愿意，求你将这杯撤去；然而，不是照我的意愿，而是要成全你的旨意。” 〔
LUKE|22|43|有一位天使从天上显现，加添他的力量。
LUKE|22|44|耶稣非常痛苦焦虑，祷告更加恳切，汗如大血点滴在地上。 〕
LUKE|22|45|祷告完了，他起来，到门徒那里，见他们因为忧愁都睡着了，
LUKE|22|46|就对他们说：“你们为什么睡觉呢？起来祷告，免得陷入试探！”
LUKE|22|47|耶稣还在说话的时候，来了一群人。十二使徒之一名叫 犹大 的，走在前头，接近耶稣，要亲他。
LUKE|22|48|耶稣对他说：“ 犹大 ，你用亲吻来出卖人子吗？”
LUKE|22|49|左右的人见了要发生的事，就说：“主啊，我们拿刀砍好不好？”
LUKE|22|50|其中有一个人把大祭司的仆人砍了一刀，削掉了他的右耳。
LUKE|22|51|耶稣回答说：“算了，住手吧！”就摸那人的耳朵，把他治好了。
LUKE|22|52|耶稣对那些来抓他的祭司长、守殿官和长老说：“你们带着刀棒出来，如同对付强盗吗？
LUKE|22|53|我天天同你们在圣殿里，你们不下手抓我。现在却是你们的时候，黑暗掌权了。”
LUKE|22|54|他们拿住耶稣，把他带走，进入大祭司的住宅。 彼得 远远地跟着。
LUKE|22|55|他们在院子中间生了火，一同坐着， 彼得 也坐在他们当中。
LUKE|22|56|有一个使女看见 彼得 面向火光坐着，就定睛看他，说：“这个人素来也是同那人一起的。”
LUKE|22|57|彼得 却不承认，说：“你这个女人，我不认得他！”
LUKE|22|58|过了一会儿，又有一个人看见他，说：“你也是他们一伙的。” 彼得 说：“你这个人，我不是！”
LUKE|22|59|约过了一小时，又有一个人坚持说：“他实在是同那人一起的，因为他也是 加利利 人。”
LUKE|22|60|彼得 说：“你这个人，我不知道你在说什么！”正说话之间，鸡就叫了。
LUKE|22|61|主转过身来看 彼得 ， 彼得 就想起主对他所说的话：“今日鸡叫以前，你要三次不认我。”
LUKE|22|62|他就出去痛哭。
LUKE|22|63|看守耶稣的人戏弄他，打他，
LUKE|22|64|又蒙着他的眼，问他：“你说预言吧！打你的是谁？”
LUKE|22|65|他们还用许多别的话辱骂他。
LUKE|22|66|天一亮，民间的众长老、祭司长和文士都聚集，把耶稣带到他们的议会里，
LUKE|22|67|说：“如果你是基督，就告诉我们。”耶稣对他们说：“我若告诉你们，你们也不信；
LUKE|22|68|我若问你们，你们也不回答。
LUKE|22|69|从今以后，人子要坐在权能者上帝的右边。”
LUKE|22|70|他们都说：“那么，你是上帝的儿子了？”耶稣对他们说：“你们说我是。”
LUKE|22|71|他们说：“我们何必再要见证呢？他亲口所说的，我们都亲耳听见了。”
LUKE|23|1|众人都起来，把耶稣解到 彼拉多 面前。
LUKE|23|2|他们开始控告他说：“我们见这人煽惑我们的国民，禁止我们纳税给凯撒，并说自己是基督，是王。”
LUKE|23|3|彼拉多 问耶稣：“你是 犹太 人的王吗？”耶稣回答：“是你说的。”
LUKE|23|4|彼拉多 对祭司长们和众人说：“我查不出这人有什么罪来。”
LUKE|23|5|但他们越发竭力地说：“他煽动百姓，在 犹太 全地传道，从 加利利 起，直到这里了。”
LUKE|23|6|彼拉多 一听见，就问：“这人是 加利利 人吗？”
LUKE|23|7|既知道耶稣属 希律 所管， 彼拉多 就把他送到 希律 那里去。那时 希律 正在 耶路撒冷 。
LUKE|23|8|希律 看见耶稣就非常高兴；因为听见过他的事，早就想要见他，并且指望看他行些神迹，
LUKE|23|9|于是问他许多的话，耶稣却一言不答。
LUKE|23|10|那些祭司长和文士都站着，竭力控告他。
LUKE|23|11|希律 和他的士兵就藐视耶稣，戏弄他，给他穿上华丽的衣服，把他送回 彼拉多 那里去。
LUKE|23|12|从前 希律 和 彼拉多 彼此有仇，在那一天竟成了朋友。
LUKE|23|13|彼拉多 传齐了众祭司长、官长和百姓，
LUKE|23|14|对他们说：“你们解这人到我这里，说他是煽惑百姓的。看哪，我也曾在你们面前审问他，并没有查出这人犯过你们控告他的任何罪；
LUKE|23|15|就是 希律 也是如此，所以把他送回来。可见他没有做什么该死的事。
LUKE|23|16|所以，我要责打他，把他释放。”
LUKE|23|17|
LUKE|23|18|众人却一齐喊着说：“除掉这个人！释放 巴拉巴 给我们！”
LUKE|23|19|这 巴拉巴 是因在城里作乱和杀人而下在监里的。
LUKE|23|20|彼拉多 愿意释放耶稣，就再次向他们讲话。
LUKE|23|21|无奈他们喊着说：“把他钉十字架！把他钉十字架！”
LUKE|23|22|彼拉多 第三次对他们说：“为什么呢？这人做了什么恶事呢？我并没有查出他有什么该死的罪来。所以，我要责打他，把他释放。”
LUKE|23|23|他们大声催逼 彼拉多 ，要求他把耶稣钉十字架；他们的声音终于得胜。
LUKE|23|24|彼拉多 这才照他们的要求定案；
LUKE|23|25|又把他们所要求的那因作乱和杀人而下在监里的人释放了，而把耶稣交给他们，随他们的意思处置。
LUKE|23|26|他们把耶稣带去的时候，有一个 古利奈 人 西门 从乡下来，他们就拿住他，把十字架搁在他身上，叫他背着跟在耶稣后面。
LUKE|23|27|有许多百姓跟随耶稣，其中有好些妇女为他号啕痛哭。
LUKE|23|28|耶稣转身对她们说：“ 耶路撒冷 的女子，不要为我哭，要为你们自己和你们的儿女哭。
LUKE|23|29|因为日子将到，人要说：‘不生育的、未曾怀孕的，和未曾哺乳孩子的有福了！’
LUKE|23|30|那时，人要向大山说： ‘倒在我们身上！’ 向小山说： ‘遮盖我们！’
LUKE|23|31|他们若在树木青绿的时候做这些事，那么在枯干的时候将会怎么样呢？”
LUKE|23|32|另外有两个犯人也被带来和耶稣一同处死。
LUKE|23|33|到了一个地方，名叫髑髅地，他们就在那里把耶稣钉在十字架上，又钉了两个犯人：一个在右边，一个在左边。 〔
LUKE|23|34|这时，耶稣说：“父啊！赦免他们，因为他们所做的，他们不知道。” 〕士兵就抽签分他的衣服。
LUKE|23|35|百姓站在那里观看。官长也嘲笑他，说：“他救了别人，他若是基督，是上帝所拣选的，救救他自己吧！”
LUKE|23|36|士兵也戏弄他，上前拿醋送给他喝，
LUKE|23|37|说：“你若是 犹太 人的王，救救你自己吧！”
LUKE|23|38|在耶稣上方有一个牌子写着：“这是 犹太 人的王。”
LUKE|23|39|同钉的犯人中有一个讥笑他，说：“你不是基督吗？救救你自己和我们吧！”
LUKE|23|40|另一个就应声责备他，说：“你是一样受刑的，还不怕上帝吗？
LUKE|23|41|我们是应得的，因为我们是自作自受，但这个人没有做过一件不对的事。”
LUKE|23|42|他对耶稣说：“耶稣啊，你进入你国的时候，求你记念我。”
LUKE|23|43|耶稣对他说：“我实在告诉你，今日你要同我在乐园里了。”
LUKE|23|44|那时大约是正午，全地都黑暗了，直到下午三点钟，
LUKE|23|45|太阳变黑了，殿的幔子从当中裂为两半。
LUKE|23|46|耶稣大声喊着说：“父啊，我将我的灵交在你手里！”他说了这话，气就断了。
LUKE|23|47|百夫长看见所发生的事，就归荣耀给上帝，说：“这人真是个义人！”
LUKE|23|48|聚集观看这事的众人，见了所发生的事，都捶着胸回去了。
LUKE|23|49|所有与耶稣熟悉的人，和从 加利利 跟着他来的妇女们，都远远地站着，看这些事。
LUKE|23|50|有一个人名叫 约瑟 ，是个议员，为人善良正直，
LUKE|23|51|却没有附从别人的所谋所为。他是 犹太 的 亚利马太城 人，素常盼望着上帝的国。
LUKE|23|52|这人去见 彼拉多 ，请求要耶稣的身体。
LUKE|23|53|他把耶稣的身体取下来，用细麻布裹好，安放在凿岩而成的坟墓里；那坟墓从来没有葬过人。
LUKE|23|54|那日是预备日，安息日快到了。
LUKE|23|55|那些从 加利利 和耶稣同来的妇女跟在后面，看见了坟墓和他的身体怎样安放。
LUKE|23|56|她们就回去，预备了香料香膏。在安息日，她们遵照诫命安息了。
LUKE|24|1|七日的第一日，黎明的时候，那些妇女带着所预备的香料来到坟墓那里，
LUKE|24|2|发现石头已经从坟墓滚开了，
LUKE|24|3|她们就进去，只是不见主耶稣的身体。
LUKE|24|4|正在为这事困惑的时候，忽然有两个人站在旁边，衣服放光。
LUKE|24|5|妇女们非常害怕，就俯伏在地上。那两个人对她们说：“为什么在死人中找活人呢？
LUKE|24|6|他不在这里，已经复活了。要记得他还在 加利利 的时候怎样告诉你们的，
LUKE|24|7|他说：‘人子必须被交在罪人手里，钉在十字架上，第三天复活。’”
LUKE|24|8|她们就想起耶稣的话来。
LUKE|24|9|于是她们从坟墓那里回去，把这一切事告诉十一个使徒和其余的人。
LUKE|24|10|把这些事告诉使徒的有 抹大拉 的 马利亚 、 约亚拿 ，和 雅各 的母亲 马利亚 ，还有跟她们在一起的妇女。
LUKE|24|11|她们这些话，使徒以为是胡言，就不相信。
LUKE|24|12|彼得 起来，跑到坟墓前，俯身往里看，只见细麻布，就回去了，因所发生的事而心里惊讶。
LUKE|24|13|同一天，门徒中有两个人往一个村子去；这村子名叫 以马忤斯 ，离 耶路撒冷 约有二十五里 。
LUKE|24|14|他们彼此谈论所发生的这一切事。
LUKE|24|15|正交谈议论的时候，耶稣亲自走近他们，和他们同行，
LUKE|24|16|可是他们的眼睛模糊了，没认出他。
LUKE|24|17|耶稣对他们说：“你们一边走一边谈，彼此谈论的是什么事呢？”他们就站住，脸上带着愁容。
LUKE|24|18|两人中有一个名叫 革流巴 的回答：“你是在 耶路撒冷 的旅客中，惟一还不知道这几天在那里发生了什么事的人吗？”
LUKE|24|19|耶稣对他们说：“什么事呢？”他们对他说：“就是 拿撒勒 人耶稣的事。他是个先知，在上帝和众百姓面前，说话行事都大有能力。
LUKE|24|20|祭司长们和我们的官长竟把他解去，定了死罪，钉在十字架上。
LUKE|24|21|但我们素来所盼望要救赎 以色列 民的就是他。不但如此，这些事发生到现在已经三天了。
LUKE|24|22|还有，我们中间的几个妇女使我们惊奇：她们清早去了坟墓，
LUKE|24|23|不见他的身体，就回来告诉我们，说她们看见了天使显现，说他活了。
LUKE|24|24|又有我们的几个人往坟墓那里去，所发现的正如妇女们所说的，只是没有看见他。”
LUKE|24|25|耶稣对他们说：“无知的人哪，先知所说的一切话，你们的心信得太迟钝了。
LUKE|24|26|基督不是必须受这些苦难，然后进入他的荣耀吗？”
LUKE|24|27|于是，他从 摩西 和众先知起，凡经上所指着自己的话都给他们作了解释。
LUKE|24|28|他们走近所要去的村子，耶稣好像还要往前走，
LUKE|24|29|他们却强留他说：“时候晚了，天快黑了，请你同我们住下吧。”耶稣就进去，要同他们住下。
LUKE|24|30|坐下来和他们用餐的时候，耶稣拿起饼来，祝福了，擘开，递给他们。
LUKE|24|31|他们的眼睛开了，这才认出他来。耶稣却从他们眼前消失了。
LUKE|24|32|他们彼此说：“在路上他和我们说话，给我们讲解圣经的时候，我们的心在我们里面 岂不是火热的吗？”
LUKE|24|33|于是他们立刻起身，回 耶路撒冷 去，看见十一个使徒和与他们正在一起的人聚集在一处，
LUKE|24|34|说：“主果然复活了，已经显现给 西门 看了。”
LUKE|24|35|于是，两个人把路上所遇到，和耶稣擘饼的时候怎么被他们认出来的事，都述说了一遍。
LUKE|24|36|正说这些话的时候，耶稣亲自站在他们当中，说：“愿你们平安！”
LUKE|24|37|他们却惊慌害怕，以为所看见的是魂。
LUKE|24|38|耶稣对他们说：“你们为什么惊恐不安？为什么心里起疑惑呢？
LUKE|24|39|你们看我的手和我的脚，就知道实在是我了。摸摸我，看，因为魂无骨无肉，你们看，我是有的。”
LUKE|24|40|说了这话，他就把手和脚给他们看。
LUKE|24|41|他们还在又惊又喜、不敢相信的时候，耶稣对他们说：“你们这里有什么吃的没有？”
LUKE|24|42|他们给了他一片烤鱼，
LUKE|24|43|他接过来，在他们面前吃了。
LUKE|24|44|耶稣对他们说：“这就是我从前和你们同在时所告诉你们的话： 摩西 的律法、先知的书，和《 诗篇》 上所记一切指着我的话都必须应验。”
LUKE|24|45|于是耶稣开他们的心窍，使他们能明白圣经，
LUKE|24|46|又对他们说：“照经上所写的，基督必受害，第三天从死人中复活，
LUKE|24|47|并且人们要奉他的名传悔改、使罪得赦的道，从 耶路撒冷 起直传到万邦。
LUKE|24|48|你们就是这些事的见证。
LUKE|24|49|我要将我父所应许的降在你们身上，你们要在城里等候，直到你们领受从上面来的能力。”
LUKE|24|50|耶稣领他们出来，直到 伯大尼 附近，就举手给他们祝福。
LUKE|24|51|正祝福的时候，他离开他们，被带到天上去了。
LUKE|24|52|他们就拜他，带着极大的喜乐回 耶路撒冷 去，
LUKE|24|53|常在圣殿里称颂上帝。
JOHN|1|1|太初有道，道与上帝同在，道就是上帝。
JOHN|1|2|这道太初与上帝同在。
JOHN|1|3|万物都是藉着他造的，没有一样不是藉着他造的。凡被造的，
JOHN|1|4|在他里面有生命 ，这生命就是人的光。
JOHN|1|5|光照在黑暗里，黑暗却没有胜过光 。
JOHN|1|6|有一个人，是从上帝那里差来的，名叫 约翰 。
JOHN|1|7|这人来是为了作见证，是为那光作见证，要使众人藉着他而信。
JOHN|1|8|他不是那光，而是要为那光作见证。
JOHN|1|9|那光是真光，来到世上，照亮所有的人 。
JOHN|1|10|他在世界，世界是藉着他造的，世界却不认识他。
JOHN|1|11|他来到自己的地方，自己的人并不接纳他。
JOHN|1|12|凡接纳他的，就是信他名的人，他就赐他们权柄作上帝的儿女。
JOHN|1|13|这些人不是从血生的，不是从情欲生的，也不是从人的意愿生的，而是从上帝生的。
JOHN|1|14|道成了肉身，住在我们中间，充充满满地有恩典有真理，我们也见过他的荣光，正是父独一儿子 的荣光。
JOHN|1|15|约翰 为他作见证，喊着说：“这就是我曾说：‘那在我以后来的先于我，因为在我以前，他已经存在。’”
JOHN|1|16|从他的丰富里，我们都领受了恩典，而且恩上加恩。
JOHN|1|17|律法是藉着 摩西 颁布的；恩典和真理却是由耶稣基督来的。
JOHN|1|18|从来没有人见过上帝，只有在父怀里独一的儿子将他表明出来。
JOHN|1|19|这是 约翰 的见证： 犹太 人从 耶路撒冷 差祭司和 利未 人到 约翰 那里去问他：“你是谁？”
JOHN|1|20|他就承认，并不隐瞒，承认说：“我不是基督。”
JOHN|1|21|他们又问他：“那么，你是谁？是 以利亚 吗？”他说：“我不是。”“是那位先知吗？”他回答：“不是。”
JOHN|1|22|于是他们对他说：“你到底是谁，好让我们回覆差我们来的人。你说，你自己是谁？”
JOHN|1|23|他说： “我就是那在旷野呼喊的声音： 修直主的道。” 正如 以赛亚 先知所说的。
JOHN|1|24|那些人是法利赛人差来的。
JOHN|1|25|他们就问他：“你既不是基督，不是 以利亚 ，也不是那位先知，那么，你为什么施洗呢？”
JOHN|1|26|约翰 回答：“我是用水施洗，但有一位站在你们中间，是你们不认识的，
JOHN|1|27|就是那在我以后来的，我给他解鞋带也不配。”
JOHN|1|28|这些事发生在 约旦河 东边的 伯大尼 ， 约翰 施洗的地方。
JOHN|1|29|第二天， 约翰 看见耶稣来到他那里，就说：“看哪，上帝的羔羊，除去世人的罪的！
JOHN|1|30|这就是我曾说‘那在我以后来的先于我，因为在我以前，他已经存在’的那一位。
JOHN|1|31|我先前不认识他，如今我来用水施洗，为要使他显明给 以色列 人。”
JOHN|1|32|约翰 又作见证说：“我曾看见圣灵仿佛鸽子从天降下，停留在他的身上。
JOHN|1|33|我先前不认识他，可是那差我来用水施洗的对我说：‘你看见圣灵降下来，停留在谁的身上，谁就是用圣灵施洗的。’
JOHN|1|34|我看见了，所以作证：这一位是上帝的儿子。”
JOHN|1|35|又过了一天， 约翰 同两个门徒站在那里。
JOHN|1|36|他见耶稣走过，就说：“看哪，上帝的羔羊！”
JOHN|1|37|两个门徒听见他的话，就跟从了耶稣。
JOHN|1|38|耶稣转过身来，看见他们跟着，就对他们说：“你们要什么？”他们对他说：“拉比，你在哪里住？”（“拉比”翻出来就是老师。）
JOHN|1|39|耶稣说：“你们来看。”他们就去看他在哪里住。这一天他们就跟他同住；那时大约是下午四点钟。
JOHN|1|40|听了 约翰 的话而跟从耶稣的那两个人，其中一个是 西门．彼得 的弟弟 安得烈 。
JOHN|1|41|他先找到自己的哥哥 西门 ，对他说：“我们遇见弥赛亚了。”（“弥赛亚”翻出来就是基督。）
JOHN|1|42|于是 安得烈 领 西门 去见耶稣。耶稣看着他，说：“你是 约翰 的儿子 西门 ，你要称为 矶法 。”（“矶法”翻出来就是 彼得 。）
JOHN|1|43|又过了一天，耶稣想要往 加利利 去。他找到 腓力 ，就对他说：“来跟从我！”
JOHN|1|44|这 腓力 是 伯赛大 人，是 安得烈 和 彼得 的同乡。
JOHN|1|45|腓力 找到 拿但业 ，对他说：“ 摩西 在律法书上所写的，和众先知所记的那一位，我们遇见了，就是 约瑟 的儿子 拿撒勒 人耶稣。”
JOHN|1|46|拿但业 对他说：“ 拿撒勒 还能出什么好的吗？” 腓力 说：“你来看。”
JOHN|1|47|耶稣看见 拿但业 向他走来，就论到他说：“看哪，这真是个 以色列 人！他心里是没有诡诈的。”
JOHN|1|48|拿但业 对耶稣说：“你从哪里认识我的？”耶稣回答他说：“ 腓力 还没有呼唤你，你在无花果树底下，我就看见你了。”
JOHN|1|49|拿但业 回答他说：“拉比！你是上帝的儿子，你是 以色列 的王。”
JOHN|1|50|耶稣回答他说：“因为我说在无花果树底下看见你，你就信吗？你将看见比这些更大的事呢！”
JOHN|1|51|他又说：“我实实在在地告诉你们，你们将要看见天开了，上帝的使者在人子身上，上去下来。”
JOHN|2|1|第三日，在 加利利 的 迦拿 有一个婚宴，耶稣的母亲在那里。
JOHN|2|2|耶稣和他的门徒也被请去赴宴。
JOHN|2|3|酒用完了，耶稣的母亲对他说：“他们没有酒了。”
JOHN|2|4|耶稣说：“母亲 ，我与你何干呢？我的时候还没有到。”
JOHN|2|5|他母亲对用人说：“他告诉你们什么，你们就做吧。”
JOHN|2|6|照 犹太 人洁净礼的规矩，有六口石缸摆在那里，每口可以盛两三桶 水。
JOHN|2|7|耶稣对用人说：“把缸倒满水。”他们就倒满了，直到缸口。
JOHN|2|8|耶稣又说：“现在舀出来，送给宴会总管。”他们就送了去。
JOHN|2|9|宴会总管尝了那水变的酒，并不知道是哪里来的，只有舀水的用人知道。于是宴会总管叫新郎来，
JOHN|2|10|对他说：“人家都是先摆上好酒，等客人喝够了才摆上次的，你倒把好酒留到现在！”
JOHN|2|11|这是耶稣所行的第一个神迹，是在 加利利 的 迦拿 行的，显出了他的荣耀来，他的门徒就信他了。
JOHN|2|12|这事以后，耶稣与他的母亲、兄弟 和门徒 都下 迦百农 去，在那里住了不多几天。
JOHN|2|13|犹太 人的逾越节近了，耶稣上 耶路撒冷 去。
JOHN|2|14|他看见圣殿里有卖牛羊和鸽子的，还有兑换银钱的人坐着，
JOHN|2|15|耶稣就拿绳子做成鞭子，把所有的，包括牛羊都赶出圣殿，倒出兑换银钱之人的银钱，推翻他们的桌子，
JOHN|2|16|又对卖鸽子的说：“把这些东西拿走！不要把我父的殿当作买卖的地方。”
JOHN|2|17|他的门徒就想起经上记着：“我为你的殿心里焦急，如同火烧。”
JOHN|2|18|因此 犹太 领袖问他：“你能显什么神迹给我们看，表明你可以做这些事呢？”
JOHN|2|19|耶稣回答他们说：“你们拆毁这殿，我三日内要把它重建。”
JOHN|2|20|犹太 人问：“这殿造了四十六年，你三日内就能重建吗？”
JOHN|2|21|但耶稣所说的殿是指他的身体。
JOHN|2|22|所以他从死人中复活以后，门徒想起他曾说过这事，就信了圣经和耶稣所说的话。
JOHN|2|23|耶稣在 耶路撒冷 过逾越节的时候，有许多人看见他所行的神迹，就信了他的名。
JOHN|2|24|耶稣自己却不信任他们，因为他认识所有的人，
JOHN|2|25|也用不着谁来证明人是怎样的，因为他自己认识人的内心。
JOHN|3|1|有一个法利赛人，名叫 尼哥德慕 ，是 犹太 人的官。
JOHN|3|2|这人夜里来见耶稣，对他说：“拉比，我们知道你是由上帝那里来作老师的；因为你所行的神迹，若没有上帝同在，无人能行。”
JOHN|3|3|耶稣回答他说：“我实实在在地告诉你，人若不重生 ，就不能见上帝的国。”
JOHN|3|4|尼哥德慕 对他说：“人已经老了，如何能重生呢？岂能再进母腹生出来吗？”
JOHN|3|5|耶稣回答：“我实实在在地告诉你，人若不是从水和圣灵生的，就不能进上帝的国。
JOHN|3|6|从肉身生的就是肉身；从灵生的就是灵。
JOHN|3|7|我说‘你们必须重生’，你不要惊讶。
JOHN|3|8|风 随着意思吹，你听见风的声音，却不知道是从哪里来，往哪里去；凡从圣灵生的也是如此。”
JOHN|3|9|尼哥德慕 问他：“怎么能有这些事呢？”
JOHN|3|10|耶稣回答，对他说：“你是 以色列 人的老师，还不明白这些事吗？
JOHN|3|11|我实实在在地告诉你，我们所说的是我们知道的，我们所见证的是我们见过的，你们却不领受我们的见证。
JOHN|3|12|我对你们说地上的事，你们尚且不信，若对你们说天上的事，如何能信呢？
JOHN|3|13|除了从天降下 的人子，没有人升过天。
JOHN|3|14|摩西 在旷野怎样举蛇，人子也必须照样被举起来，
JOHN|3|15|要使一切信他的人都得永生。
JOHN|3|16|“上帝爱世人，甚至将他独一的儿子 赐给他们，叫一切信他的人不致灭亡，反得永生。
JOHN|3|17|因为上帝差他的儿子到世上来，不是要定世人的罪 ，而是要使世人因他得救。
JOHN|3|18|信他的人不被定罪；不信的人已经被定罪了，因为他不信上帝独一儿子的名。
JOHN|3|19|光来到世上，世人因自己的行为是恶的，不爱光，倒爱黑暗，这就定了他们的罪。
JOHN|3|20|凡作恶的人都恨恶光，不来接近光，恐怕他的行为被暴露。
JOHN|3|21|但实行真理的人就来接近光，为要显明他的行为是靠上帝而行的。”
JOHN|3|22|这些事以后，耶稣和门徒到了 犹太 地区，在那里他和他们同住，并且施洗。
JOHN|3|23|约翰 也在靠近 撒冷 的 哀嫩 施洗，因为那里水多，众人都去受洗。
JOHN|3|24|那时 约翰 还没有下在监里。
JOHN|3|25|约翰 的门徒和一个 犹太 人辩论洁净的礼仪，
JOHN|3|26|就来见 约翰 ，对他说：“拉比，从前同你在 约旦河 的东边，你所见证的那位，你看，他在施洗，众人都到他那里去了。”
JOHN|3|27|约翰 回答说：“若不是从天上赐的，人就不能得到什么。
JOHN|3|28|你们自己可以为我作见证，我曾说，我不是基督，只是奉差遣在他前面开路的。
JOHN|3|29|娶新娘的是新郎；新郎的朋友站在一旁听，一听见新郎的声音就欢喜快乐。因此，我这喜乐得以满足了。
JOHN|3|30|他必兴旺；我必衰微。”
JOHN|3|31|“从上头来的是在万有之上；出于地的是属于地，他所说的也是属于地。从天上来的是在万有之上。
JOHN|3|32|他把所见所闻的见证出来，只是没有人领受他的见证。
JOHN|3|33|那领受他见证的，就印证上帝是真实的。
JOHN|3|34|上帝所差来的说上帝的话，因为上帝所赐给他的圣灵是没有限量的。
JOHN|3|35|父爱子，已把万有交在他手里。
JOHN|3|36|信子的人有永生；不信子的人得不到永生，而且上帝的愤怒常在他身上。”
JOHN|4|1|耶稣 知道法利赛人听见他收门徒和施洗比 约翰 还多， （
JOHN|4|2|其实不是耶稣亲自施洗，而是他的门徒施洗，）
JOHN|4|3|他就离开 犹太 ，又回 加利利 去。
JOHN|4|4|他必须经过 撒玛利亚 ，
JOHN|4|5|于是到了 撒玛利亚 的一座城，名叫 叙加 ，靠近 雅各 给他儿子 约瑟 的那块地。
JOHN|4|6|雅各井 就在那里；耶稣因旅途疲乏，坐在井旁。那时约是正午。
JOHN|4|7|有一个 撒玛利亚 妇人来打水。耶稣对她说：“请给我水喝。”
JOHN|4|8|因为那时门徒进城买食物去了。
JOHN|4|9|撒玛利亚 妇人对他说：“你是 犹太 人，怎么向我一个 撒玛利亚 女人要水喝呢？”因为 犹太 人和 撒玛利亚 人没有来往。
JOHN|4|10|耶稣回答她说：“你若知道上帝的恩赐，和对你说‘请给我水喝’的是谁，你早就会求他，他也早就会给了你活水。”
JOHN|4|11|妇人对耶稣说：“先生，你没有打水的器具，井又深，哪里去取活水呢？
JOHN|4|12|我们的祖宗 雅各 把这井留给我们，他自己和儿女以及牲畜都喝这井里的水，难道你比他还大吗？”
JOHN|4|13|耶稣回答，对她说：“凡喝这水的，还要再渴；
JOHN|4|14|谁喝我所赐的水，就永远不渴。我所赐的水要在他里面成为泉源，直涌到永生。”
JOHN|4|15|妇人对他说：“先生，请把这水赐给我，使我不渴，也不用到这里来打水。”
JOHN|4|16|耶稣对她说：“你去，叫你的丈夫，再到这里来。”
JOHN|4|17|妇人回答，对耶稣说：“我没有丈夫。”耶稣说：“你说没有丈夫是对的。
JOHN|4|18|你已经有过五个丈夫，你现在有的并不是你的丈夫。你这话是真的。”
JOHN|4|19|妇人对他说：“先生，我看你是一位先知。
JOHN|4|20|我们的祖宗在这山上敬拜上帝，你们倒说，应当敬拜的地方是在 耶路撒冷 。”
JOHN|4|21|耶稣对她说：“妇人，你要信我。时候将到，你们敬拜父，既不在这山上，也不在 耶路撒冷 。
JOHN|4|22|你们所敬拜的，你们不知道；我们所敬拜的，我们知道，因为救恩是从 犹太 人出来的。
JOHN|4|23|时候将到，现在就是了，那真正敬拜父的，要用心灵和诚实敬拜他，因为父要这样的人敬拜他。
JOHN|4|24|上帝是灵，所以敬拜他的必须用心灵和诚实敬拜他。”
JOHN|4|25|妇人对他说：“我知道弥赛亚—就是那称为基督的—要来；他来了，会把一切的事都告诉我们。”
JOHN|4|26|耶稣对她说：“我就是，正在跟你说话呢！”
JOHN|4|27|正在这时，门徒回来了。他们对耶稣正在和一个妇人说话感到惊讶，可是没有人说：“你要什么？”或说：“你为什么和她说话？”
JOHN|4|28|那妇人留下水罐，往城里去，对众人说：
JOHN|4|29|“你们来看！有一个人把我素来所做的一切事都说了出来，难道这个人就是基督吗？”
JOHN|4|30|他们就出城，来到耶稣那里。
JOHN|4|31|就在这个时候，门徒求耶稣说：“拉比，请吃吧。”
JOHN|4|32|耶稣对他们说：“我有食物吃，是你们不知道的。”
JOHN|4|33|门徒就彼此说：“难道有人拿什么给他吃了吗？”
JOHN|4|34|耶稣对他们说：“我的食物就是要遵行差我来那位的旨意，完成他的工作。
JOHN|4|35|你们不是说‘到收割的时候还有四个月’吗？我告诉你们，举目向田观看，庄稼熟了，可以收割了。
JOHN|4|36|收割的人已经得工钱 ，为永生储存五谷，使撒种的和收割的一同快乐。
JOHN|4|37|‘那人撒种，这人收割’，这话可见是真的。
JOHN|4|38|我差你们去收你们所没有辛劳的；别人辛劳，你们享受他们辛劳的成果。”
JOHN|4|39|那城里有好些 撒玛利亚 人信了耶稣，因为那妇人作见证，说：“他把我素来所做的一切事都说了出来。”
JOHN|4|40|于是 撒玛利亚 人来见耶稣，求他在他们那里住下，他就在那里住了两天。
JOHN|4|41|因为耶稣的话，信的人就更多了。
JOHN|4|42|他们对那妇人说：“现在我们信，不再是因为你的话，而是我们亲自听见了，知道这人真是世界的救主。”
JOHN|4|43|过了那两天，耶稣离开那地方，往 加利利 去。
JOHN|4|44|因为耶稣自己作过见证说：“先知在自己的家乡是没有人尊敬的。”
JOHN|4|45|到了 加利利 ， 加利利 人都欢迎他，因为他们也上 耶路撒冷 去过节，曾经看过他在节期间所做的一切事。
JOHN|4|46|耶稣又到了 加利利 的 迦拿 ，就是他从前变水为酒的地方。有一个大臣，他的儿子在 迦百农 病了。
JOHN|4|47|他听见耶稣从 犹太 到了 加利利 ，就来见他，求他下去医治他的儿子，因为他儿子快要死了。
JOHN|4|48|耶稣对他说：“若不看见神迹奇事，你们总是不信。”
JOHN|4|49|那大臣对他说：“先生，求你趁着我的孩子还没有死就下去吧。”
JOHN|4|50|耶稣对他说：“回去吧，你的儿子会活！”那人信耶稣所说的话，就回去了。
JOHN|4|51|正下去的时候，他的仆人迎面而来，说他的儿子活了。
JOHN|4|52|他就问什么时候见好的。他们对他说：“昨天下午一点钟热就退了。”
JOHN|4|53|他就知道这正是耶稣对他说“你的儿子会活”的时候；他自己和全家就都信了。
JOHN|4|54|这是耶稣从 犹太 回到 加利利 后所行的第二个神迹。
JOHN|5|1|这些事以后，到了 犹太 人的一个节期，耶稣上 耶路撒冷 去。
JOHN|5|2|在 耶路撒冷 ，靠近 羊门 有一个池子， 希伯来 话叫 毕士大 ，旁边有五个柱廊；
JOHN|5|3|里面躺着许多病人，有失明的、瘸腿的、瘫痪的 。
JOHN|5|4|
JOHN|5|5|在那里有一个人，病了三十八年。
JOHN|5|6|耶稣看见他躺着，知道他病了很久，就问他：“你要痊愈吗？”
JOHN|5|7|病人回答他：“先生，水动的时候，没有人把我放在池子里；我正要去的时候，别人比我先下去了。”
JOHN|5|8|耶稣对他说：“起来，拿起你的褥子走吧！”
JOHN|5|9|那人立刻痊愈，就拿起自己的褥子走了。 那天是安息日，
JOHN|5|10|所以 犹太 人对那被治好了的人说：“今天是安息日，你拿褥子是不合法的。”
JOHN|5|11|他却回答他们：“那使我痊愈的人对我说：‘拿起你的褥子走吧！’”
JOHN|5|12|他们问他：“对你说‘拿起褥子走’的是什么人？”
JOHN|5|13|那治好了的人不知道那人是谁，因为那里人很多，耶稣已经躲开了。
JOHN|5|14|后来耶稣在圣殿里找到他，对他说：“你已经痊愈了，不要再犯罪，免得你的遭遇更坏。”
JOHN|5|15|那人就去告诉 犹太 人，使他痊愈的是耶稣。
JOHN|5|16|所以 犹太 人迫害耶稣，因为他在安息日做了这些事。
JOHN|5|17|耶稣就回答他们：“我父做事直到如今，我也做事。”
JOHN|5|18|为了这缘故， 犹太 人越发想要杀他，因为他不但犯了安息日，而且称上帝为他的父，把自己和上帝看为同等。
JOHN|5|19|于是耶稣回答，对他们说：“我实实在在地告诉你们，子凭着自己不能做什么，惟有看见父所做的，他才做；父所做的事，子也照样做。
JOHN|5|20|父爱子，将自己所做的一切事指示给他看，还要将比这更大的事给他看，使你们惊讶。
JOHN|5|21|父怎样叫死人复活，赐他们生命，子也照样随自己的意愿赐人生命。
JOHN|5|22|父不审判任何人，而是把审判的事全交给子，
JOHN|5|23|为要使人都尊敬子，如同尊敬父一样。不尊敬子的，就是不尊敬差子来的父。
JOHN|5|24|“我实实在在地告诉你们，那听我话又信差我来那位的，就有永生，不至于被定罪，而是已经出死入生了。
JOHN|5|25|我实实在在地告诉你们，时候将到，现在就是了，死人要听见上帝儿子的声音，听见的人就要活了。
JOHN|5|26|因为父怎样自己里面有生命，也照样赐给他儿子自己里面有生命，
JOHN|5|27|并且赐给他施行审判的权柄，因为他是人子。
JOHN|5|28|你们不要对这事感到惊讶，因为时候将到，凡在坟墓里的，都要听见他的声音，
JOHN|5|29|并且要出来：行善的，复活得生命；作恶的，复活被定罪。
JOHN|5|30|“我凭着自己不能做什么。我怎么听见就怎么审判，而我的审判是公平的，因为我不寻求自己的意愿，只寻求差我来那位的旨意。”
JOHN|5|31|“我若为自己作见证，我的见证就不真。
JOHN|5|32|另有一位为我作见证，我也知道他为我作的见证是真的。
JOHN|5|33|你们曾差人到 约翰 那里，他为真理作过见证。
JOHN|5|34|其实，我所受的见证不是从人来的；然而，我说这些话是为了使你们得救。
JOHN|5|35|约翰 是点亮的明灯，你们情愿因他的光欢欣一时。
JOHN|5|36|但我有比 约翰 更大的见证：父交给我去完成的工作，就是我正在做的，为我作证是父差遣了我。
JOHN|5|37|那差我来的父也为我作了见证。你们从来没有听见他的声音，也没有看见他的形像。
JOHN|5|38|你们并没有他的道存在心里，因为你们不信他所差来的那一位。
JOHN|5|39|你们查考圣经，因你们以为其中有永生；而这经正是为我作见证的。
JOHN|5|40|然而，你们不肯到我这里来得生命。
JOHN|5|41|“我不接受从人来的荣耀，
JOHN|5|42|但我知道，你们没有爱上帝的心。
JOHN|5|43|我奉我父的名来了，你们并不接纳我；若有别人奉自己的名来，你们倒会接纳他。
JOHN|5|44|你们互相受荣耀，却不寻求从独一上帝来的荣耀，怎能信我呢？
JOHN|5|45|不要以为我会在父面前告你们；有一位告你们的，就是你们所仰望的 摩西 。
JOHN|5|46|如果你们信 摩西 ，也会信我，因为他写过关于我的事。
JOHN|5|47|你们若不信他的书，怎能信我的话呢？”
JOHN|6|1|这些事以后，耶稣渡过 加利利海 ，就是 提比哩亚海 。
JOHN|6|2|有一大群人因为看见他在病人身上所行的神迹，就跟随他。
JOHN|6|3|耶稣上了山，和门徒一同坐在那里。
JOHN|6|4|那时 犹太 人的逾越节近了。
JOHN|6|5|耶稣举目看见一大群人来，就对 腓力 说：“我们到哪里去买饼给这些人吃呢？”
JOHN|6|6|他说这话是要考验 腓力 ，他自己原知道要怎样做。
JOHN|6|7|腓力 回答他：“就是两百个银币的饼也不够给他们每人吃一点点。”
JOHN|6|8|有一个门徒，就是 西门．彼得 的弟弟 安得烈 ，对耶稣说：
JOHN|6|9|“这里有一个孩子，带着五个大麦饼和两条鱼，但是分给这么多人还算什么呢？”
JOHN|6|10|耶稣说：“你们叫大家坐下。”那地方的草多，人们就坐下，男人的数目约有五千。
JOHN|6|11|耶稣拿起饼来，祝谢了，就分给坐着的人，也同样分了鱼，都照他们所要的来分。
JOHN|6|12|他们吃饱后，耶稣对门徒说：“把剩下的碎屑收拾起来，免得糟蹋了。”
JOHN|6|13|他们就把那五个大麦饼的碎屑，就是大家吃剩的，收拾起来，装满了十二个篮子。
JOHN|6|14|人们看见耶稣所行的神迹，就说：“这真是那要到世上来的先知！”
JOHN|6|15|耶稣知道他们要来强迫他作王，就独自又退到山上去了。
JOHN|6|16|到了晚上，他的门徒下到海边，
JOHN|6|17|上了船，要过海往 迦百农 去。天已经黑了，耶稣还没有来到他们那里。
JOHN|6|18|忽然狂风大作，海浪翻腾。
JOHN|6|19|门徒摇橹，约行了十里多 ，看见耶稣在海面上走，渐渐靠近了船，他们就害怕。
JOHN|6|20|耶稣对他们说：“是我，不要怕！”
JOHN|6|21|门徒就欣然接他上船，船立刻到了他们所要去的地方。
JOHN|6|22|第二天，留在海的对岸的众人发觉那里原来只有一条小船，而且耶稣没有同他的门徒上船，是门徒自己去的。
JOHN|6|23|另外有几条从 提比哩亚 来的小船，却停靠在主祝谢后给他们吃饼的地方附近。
JOHN|6|24|这时众人见耶稣和门徒都不在那里，就上了船，往 迦百农 去找耶稣。
JOHN|6|25|他们在海的对岸找到他后，对他说：“拉比，你几时到这里来的？”
JOHN|6|26|耶稣回答他们说：“我实实在在地告诉你们，你们找我，并不是因见了神迹，而是因吃饼吃饱了。
JOHN|6|27|不要为那会坏的食物操劳，而要为那存到永生的食物操劳。这食物是人子要赐给你们的，因为父上帝已印证了。”
JOHN|6|28|于是他们问他：“我们该做什么才算是做上帝的工作呢？”
JOHN|6|29|耶稣回答，对他们说：“信上帝所差来的，这就是上帝的工作。”
JOHN|6|30|于是他们对他说：“你行什么神迹，好让我们看见而信你呢？你到底要做什么呢？
JOHN|6|31|我们的祖宗在旷野吃过吗哪，如经上写着：‘他从天上赐下粮食来给他们吃。’”
JOHN|6|32|于是耶稣对他们说：“我实实在在地告诉你们，那从天上来的粮不是 摩西 赐给你们的，那从天上来的真粮是我父赐给你们的。
JOHN|6|33|因为上帝的粮就是那位从天上降下来，并且赐生命给世界的。”
JOHN|6|34|于是他们对他说：“主啊，请常常把这粮赐给我们！”
JOHN|6|35|耶稣对他们说：“我就是生命的粮。到我这里来的，绝不饥饿；信我的，永不干渴。
JOHN|6|36|可是，我告诉过你们，你们已经看见我 ，还是不信。
JOHN|6|37|凡父所赐给我的人，必到我这里来；到我这里来的，我总不丢弃他。
JOHN|6|38|因为我从天上降下来，不是要按自己的意愿行，而是要遵行差我来那位的旨意。
JOHN|6|39|差我来那位的旨意就是：他所赐给我的，要我一个也不失落，并且在末日使他复活。
JOHN|6|40|因为我父的旨意是要使每一个见了子而信的人得永生，并且在末日我要使他复活。”
JOHN|6|41|犹太 人因为耶稣说“我是从天上降下来的粮”，就私下议论他，
JOHN|6|42|说：“这不是 约瑟 的儿子耶稣吗？我们岂不认得他的父母吗？现在他怎么说‘我是从天上降下来的’呢？”
JOHN|6|43|耶稣回答，对他们说：“你们不要彼此私下议论。
JOHN|6|44|若不是差我来的父吸引人，就没有人能到我这里来；到我这里来的，在末日我要使他复活。
JOHN|6|45|在先知书上写着：‘他们都要蒙上帝教导。’凡听了父的教导而学习的，都到我这里来。
JOHN|6|46|这不是说有人看见过父，惟独从上帝来的，他才看见过父。
JOHN|6|47|我实实在在地告诉你们，信的人有永生。
JOHN|6|48|我就是生命的粮。
JOHN|6|49|你们的祖宗在旷野吃过吗哪，还是死了。
JOHN|6|50|这是从天上降下来的粮，使人吃了就不死。
JOHN|6|51|我就是从天上降下来生命的粮；人若吃这粮，必永远活着。我为世人的生命所赐下的粮就是我的肉。”
JOHN|6|52|因此， 犹太 人彼此争论说：“这个人怎能把他的肉给我们吃呢？”
JOHN|6|53|耶稣对他们说：“我实实在在地告诉你们，你们若不吃人子的肉，不喝人子的血，在你们里面就没有生命。
JOHN|6|54|吃我肉、喝我血的人就有永生，并且在末日我要使他复活。
JOHN|6|55|我的肉是真正可吃的；我的血是真正可喝的。
JOHN|6|56|吃我肉、喝我血的人常在我里面，我也常在他里面。
JOHN|6|57|永生的父怎样差我来，我又怎样因父活着，照样，吃我肉的人也要因我活着。
JOHN|6|58|这是从天上降下来的粮，不像你们的祖宗吃过吗哪还是死了；吃这粮的人将永远活着。”
JOHN|6|59|这些话是耶稣在 迦百农 会堂里教导人的时候说的。
JOHN|6|60|他的门徒中有好些人听见了，就说：“这话很难，谁听得进呢？”
JOHN|6|61|耶稣心里知道门徒为这话私下议论，就对他们说：“这话成了你们的绊脚石吗？
JOHN|6|62|如果你们看见人子升到他原来所在之处，会怎么样呢？
JOHN|6|63|圣灵赐人生命，肉体毫无用处。我对你们所说的话就是灵，就是生命。
JOHN|6|64|可是你们中间有些人不信。”耶稣起初就知道哪些人不信他，哪一个要出卖他。
JOHN|6|65|于是耶稣说：“所以，我对你们说过，若不是蒙我父的恩赐，没有人能到我这里来。”
JOHN|6|66|从此，他门徒中有很多退却了，不再和他同行。
JOHN|6|67|耶稣就对那十二使徒说：“你们也要离开吗？”
JOHN|6|68|西门．彼得 回答他：“主啊，你有永生之道，我们还跟从谁呢？
JOHN|6|69|我们已经信了，又知道你是上帝的圣者。”
JOHN|6|70|耶稣回答他们：“我不是拣选了你们十二个吗？但你们中间有一个是魔鬼。”
JOHN|6|71|耶稣这话是指着要出卖他的 加略 人 西门 的儿子 犹大 说的；他本是十二使徒里的一个。
JOHN|7|1|这些事以后，耶稣周游 加利利 ，不愿在 犹太 往来，因为 犹太 人想要杀他。
JOHN|7|2|这时 犹太 人的住棚节近了。
JOHN|7|3|耶稣的兄弟们对他说：“你离开这里上 犹太 去吧，好让你的门徒也看见你所做的事。
JOHN|7|4|因为人要扬名，没有在隐秘的地方行事的，如果你要做这些事，该把自己显明给世人看。”
JOHN|7|5|原来连他的兄弟们也不信他。
JOHN|7|6|于是耶稣对他们说：“我的时机还没有到，你们的时机却随时都有。
JOHN|7|7|世人不会恨你们，却是恨我，因为我指证他们的行为是恶的。
JOHN|7|8|你们上去过节吧！我现在不上去过这节 ，因为我的时机还没有成熟。”
JOHN|7|9|耶稣说了这些话，仍然留在 加利利 。
JOHN|7|10|但他的兄弟们上去过节以后，他也上去，不是公开去，却似乎 是秘密地去的。
JOHN|7|11|节期间， 犹太 人寻找耶稣，说：“他在哪里？”
JOHN|7|12|人群中有许多人对他议论纷纷，另有的说：“他是好人。”有的说：“不，他是迷惑群众的。”
JOHN|7|13|可是没有人公开谈论他，因为他们怕 犹太 人。
JOHN|7|14|节期已过了一半，耶稣上圣殿去教导人。
JOHN|7|15|犹太 人惊讶地说：“这个人没有学过，怎么那样熟悉经典呢？”
JOHN|7|16|于是耶稣回答他们，说：“我的教导不是我自己的，而是差我来那位的。
JOHN|7|17|人若立志要遵行上帝的旨意，就会知道这教导究竟是出于上帝，还是我凭着自己说的。
JOHN|7|18|凭着自己说的人是寻求自己的荣耀；但那寻求差他来那位的荣耀的人，他是真诚的，在他心里没有不义。
JOHN|7|19|摩西 不是传了律法给你们吗？你们却没有一个人守律法。为什么想要杀我呢？”
JOHN|7|20|众人回答：“你是被鬼附了！谁想要杀你呢？”
JOHN|7|21|耶稣回答，对他们说：“我做了一件事，你们都惊讶。
JOHN|7|22|摩西 传割礼给你们（其实割礼不是从 摩西 开始，而是从列祖开始的），你们就在安息日给人行割礼。
JOHN|7|23|人若在安息日受割礼，是为了不违背 摩西 的律法，我在安息日使一个人痊愈了，你们就向我发怒吗？
JOHN|7|24|不要凭外表断定是非，总要按公平断定是非。”
JOHN|7|25|于是 耶路撒冷 人中有的说：“这个人不是他们想要杀的吗？
JOHN|7|26|你看，他还公开讲道，他们也不对他说什么。难道官长真的认为这是基督吗？
JOHN|7|27|然而，我们知道这个人从哪里来；可是基督来的时候，没有人知道他从哪里来。”
JOHN|7|28|那时，耶稣在圣殿里教导人，喊着说：“你们认识我，也知道我从哪里来；我并不是凭着自己来的。但差我来的那位是真实的，你们不认识他。
JOHN|7|29|我却认识他，因为我从他那里来，是他差遣了我。”
JOHN|7|30|于是他们想要捉拿耶稣，只是没有人下手，因为他的时候还没有到。
JOHN|7|31|但人群中有好些人信他，他们说：“基督来的时候，他所行的神迹难道会比这人行的更多吗？”
JOHN|7|32|法利赛人听见群众对耶稣这样议论纷纷，祭司长和法利赛人就打发圣殿警卫去捉拿他。
JOHN|7|33|于是耶稣说：“我跟你们在一起的时候不会太久了，我要回到那差我来的那里去。
JOHN|7|34|你们要找我，却找不到；我所在的地方，你们不能去。”
JOHN|7|35|于是 犹太 人彼此问：“这人要往哪里去，使我们找不到他呢？难道他要往散居在 希腊 的 犹太 人那里去教导 希腊 人吗？
JOHN|7|36|他说‘你们要找我，却找不到；我所在的地方，你们不能去’这话是什么意思呢？”
JOHN|7|37|节期的最后一天，就是最隆重的一天，耶稣站着，喊着说：“人若渴了，到我这里来喝！
JOHN|7|38|信我的人，就如经上所说：‘从他腹中将流出活水的江河来。’”
JOHN|7|39|耶稣这话是指信他的人要受圣灵说的；那时还没有赐下圣灵，因为耶稣还没有得到荣耀。
JOHN|7|40|众人听见这些话，有的说：“这真是那先知。”
JOHN|7|41|另有的说：“这是基督。”但也有的说：“难道基督是出自 加利利 吗？
JOHN|7|42|经上不是说‘基督是 大卫 的后裔，出自 大卫 的本乡 伯利恒 ’吗？”
JOHN|7|43|于是众人因耶稣而分裂了。
JOHN|7|44|其中有人要捉拿他，只是没有人下手。
JOHN|7|45|警卫们回到祭司长和法利赛人那里。他们对警卫说：“你们为什么没有带他来呢？”
JOHN|7|46|警卫回答：“从来没有像他这样说话的！”
JOHN|7|47|于是法利赛人说：“你们也受了迷惑吗？
JOHN|7|48|难道官长或法利赛人中有信他的吗？
JOHN|7|49|但这些不明白律法的众人是被诅咒的！”
JOHN|7|50|其中有 尼哥德慕 ，就是从前去见过耶稣的，对他们说：
JOHN|7|51|“不先听本人的口供，查明他所做的事，难道我们的律法还定他的罪吗？”
JOHN|7|52|他们回答他说：“你也是出自 加利利 吗？你去查考就知道， 加利利 是不出先知的。” 〔
JOHN|7|53|于是各人都回家去了，
JOHN|8|1|耶稣却到 橄榄山 去。
JOHN|8|2|清早，他又回到圣殿里。众百姓都到他那里去，他就坐下，教导他们。
JOHN|8|3|文士和法利赛人带着一个犯奸淫时被捉的女人来，叫她站在当中，
JOHN|8|4|然后对耶稣说：“老师，这女人是正在犯奸淫的时候被捉到的。
JOHN|8|5|摩西 在律法书上命令我们把这样的女人用石头打死。那么，你怎么说呢？”
JOHN|8|6|他们说这话是要试探耶稣，要抓到控告他的把柄。耶稣却弯下腰，用指头在地上写字。
JOHN|8|7|他们还是不住地问他，耶稣就直起腰来，对他们说：“你们中间谁没有罪，谁就先拿石头打她！”
JOHN|8|8|于是他又弯着腰，用指头在地上写字。
JOHN|8|9|他们听见这话，从老的开始，一个一个都走开了，只剩下耶稣一人和那仍然站在中间的女人。
JOHN|8|10|耶稣就直起腰来，对她说：“妇人，那些人在哪里呢？没有任何人定你的罪吗？”
JOHN|8|11|她说：“主啊，没有。”耶稣说：“我也不定你的罪。去吧！从今以后不要再犯罪了。”〕
JOHN|8|12|耶稣又对众人说：“我就是世界的光。跟从我的，必不在黑暗里走，却要得着生命的光。”
JOHN|8|13|法利赛人对他说：“你是为自己作见证，你的见证不真。”
JOHN|8|14|耶稣回答他们，对他们说：“即使我为自己作见证，我的见证还是真的，因为我知道我从哪里来，到哪里去。你们却不知道我从哪里来，到哪里去。
JOHN|8|15|你们是以人的标准来判断人，我不判断任何人。
JOHN|8|16|即使我判断人，我的判断也是真确的，因为不是我独自在判断，而是差我来的父与我一同判断。
JOHN|8|17|你们的律法也记着说：‘两个人的见证才算为真’。
JOHN|8|18|我是为自己作见证，还有差我来的父也为我作见证。”
JOHN|8|19|于是他们问他：“你的父在哪里？”耶稣回答：“你们不认识我，也不认识我的父；若是认识我，也会认识我的父。”
JOHN|8|20|这些话是耶稣在圣殿的银库房里教导人的时候说的。当时没有人捉拿他，因为他的时候还没有到。
JOHN|8|21|于是耶稣又对他们说：“我去了，你们会找我，而你们会死在自己的罪中；我所去的地方，你们不能去。”
JOHN|8|22|犹太 人说：“他说‘我所去的地方，你们不能去’，难道他要自杀吗？”
JOHN|8|23|耶稣对他们说：“你们是从下面来的，我是从上面来的；你们是属这世界的，我不是属这世界的。
JOHN|8|24|所以我对你们说，你们会死在自己的罪中，你们若不信我就是那位，就会死在自己的罪中。”
JOHN|8|25|他们就问他：“你到底是谁？”耶稣对他们说：“我从起初就告诉你们了。
JOHN|8|26|我有许多事要讲论你们，判断你们；但差我来的那位是真实的，我从他那里所听见的，就告诉世人。”
JOHN|8|27|他们不明白耶稣是对他们讲父的事。
JOHN|8|28|所以耶稣说：“你们举起人子以后就会知道我就是那位了，并且知道我没有一件事是凭着自己做的。我说这些话是照着父所教导我的。
JOHN|8|29|差我来的那位与我同在；他没有撇下我独自一人，因为我一直行他所喜悦的事。”
JOHN|8|30|耶稣说这些话的时候，有许多人信了他。
JOHN|8|31|耶稣对信他的 犹太 人说：“你们若继续遵守我的道，就真是我的门徒了。
JOHN|8|32|你们将认识真理，真理会使你们自由。”
JOHN|8|33|他们回答他：“我们是 亚伯拉罕 的后裔，从来没有作过谁的奴隶，你怎么说‘会使你们自由’呢？”
JOHN|8|34|耶稣回答他们：“我实实在在地告诉你们，所有犯罪的人就是罪的奴隶。
JOHN|8|35|奴隶不能永远住在家里；儿子才永远住在家里。
JOHN|8|36|所以，上帝的儿子若使你们自由，你们就真正自由了。”
JOHN|8|37|“我知道，你们是 亚伯拉罕 的后裔，你们却想要杀我，因为你们心里容不下我的道。
JOHN|8|38|我所说的是在我父那里看见的；你们所做的是在你们的父那里听到的。”
JOHN|8|39|他们回答耶稣：“我们的父是 亚伯拉罕 。”耶稣对他们说：“你们若是 亚伯拉罕 的儿女，就会做 亚伯拉罕 所做的事。
JOHN|8|40|我把在上帝那里所听见的真理告诉了你们，现在你们却想要杀我； 亚伯拉罕 没有做过这样的事。
JOHN|8|41|你们是做你们父的工作。”他们就对他说：“我们不是从淫乱生的，我们只有一位父，就是上帝。”
JOHN|8|42|耶稣对他们说：“假如上帝是你们的父，你们会爱我，因为我本是出于上帝，也是从上帝而来，我不是凭着自己来，而是他差我来的。
JOHN|8|43|你们为什么不明白我的话呢？无非是你们听不进我的道。
JOHN|8|44|你们是出于你们的父魔鬼，你们宁愿随着你们父的欲念而行。他从起初就是杀人的，不守真理，因他心里没有真理。他说谎是出于自己的本性，因他本来是说谎的，也是说谎者之父。
JOHN|8|45|但是，因为我讲真理，你们就不信我。
JOHN|8|46|你们中间谁能指证我有罪呢？既然我讲真理，你们为什么不信我呢？
JOHN|8|47|出于上帝的，必听上帝的话；你们不听，因为你们不是出于上帝。”
JOHN|8|48|犹太 人回答他：“我们说你是 撒玛利亚 人，并且是被鬼附的，这话不是很对吗？”
JOHN|8|49|耶稣回答：“我没有被鬼附的；我尊敬我的父，你们却不尊敬我。
JOHN|8|50|我不寻求自己的荣耀，但有一位为我寻求荣耀，判断是非。
JOHN|8|51|我实实在在地告诉你们，人若遵守我的道，就永远不经历死亡。”
JOHN|8|52|于是 犹太 人对他说：“现在我们知道你是被鬼附了。 亚伯拉罕 死了，众先知也死了，你还说：‘人若遵守我的道，就永远不经历死亡。’
JOHN|8|53|难道你比我们的祖宗 亚伯拉罕 还大吗？他死了，众先知也死了，你把自己当作什么人呢？”
JOHN|8|54|耶稣回答：“我若荣耀自己，我的荣耀就算不了什么；荣耀我的是我的父，就是你们所说的你们的上帝。
JOHN|8|55|你们不认识他，我却认识他。我若说不认识他，我就是说谎的，像你们一样；但我认识他，也遵守他的道。
JOHN|8|56|你们的祖宗 亚伯拉罕 欢欢喜喜地仰望我的日子，他看见了，就快乐。”
JOHN|8|57|犹太 人就对他说：“你还没有五十岁，难道见过 亚伯拉罕 吗？”
JOHN|8|58|耶稣对他们说：“我实实在在地告诉你们，还没有 亚伯拉罕 我就存在了。”
JOHN|8|59|于是他们拿石头要打他，耶稣却躲开，走出了圣殿。
JOHN|9|1|耶稣往前走的时候，看见一个生来就失明的人。
JOHN|9|2|门徒问耶稣：“拉比，这人生来失明，是谁犯了罪？是这人还是他的父母呢？”
JOHN|9|3|耶稣回答：“既不是这人犯了罪，也不是他的父母，而是要在他身上显出上帝的作为来。
JOHN|9|4|趁着白日，我们 必须做差我 来的那位的工；黑夜来到，就没有人能做工了。
JOHN|9|5|我在世上的时候，是世上的光。”
JOHN|9|6|耶稣说了这些话，就吐唾沫在地上，用唾沫和了泥抹在盲人的眼睛上，
JOHN|9|7|对他说：“你到 西罗亚 池子里去洗。”（ 西罗亚 翻出来就是“奉差遣”。）于是他去，洗了，回来就看见了。
JOHN|9|8|他的邻舍和素常见他讨饭的人，就说：“这不是那从前坐着讨饭的人吗？”
JOHN|9|9|有的说：“是他”；又有的说：“不是，却是像他。”他自己说：“是我。”
JOHN|9|10|于是他们对他说：“你的眼睛是怎么开的呢？”
JOHN|9|11|那人回答：“有一个名叫耶稣的，他和了泥抹我的眼睛，对我说：‘你到 西罗亚 池子去洗。’我去一洗，就看见了。”
JOHN|9|12|他们对他说：“那个人在哪里？”他说：“我不知道。”
JOHN|9|13|他们把以前失明的那个人带到法利赛人那里。
JOHN|9|14|耶稣和泥开他眼睛的那一天是安息日。
JOHN|9|15|法利赛人又问他是怎么得看见的。他对他们说：“他把泥抹在我的眼睛上，我一洗，就看见了。”
JOHN|9|16|于是法利赛人中有的说：“这个人不是从上帝来的，因为他不守安息日。”另有的说：“一个罪人怎能行这样的神迹呢？”他们之间就产生了分裂。
JOHN|9|17|于是他们又对那盲人说：“他开了你的眼睛，你说他是怎样的人呢？”他说：“他是个先知。”
JOHN|9|18|犹太 人不信他以前是失明，后来能看见的，等到叫了他的父母来，
JOHN|9|19|问他们说：“这是你们的儿子吗？你们说他生来是失明的，现在怎么看见了呢？”
JOHN|9|20|他的父母就回答说：“他是我们的儿子，生来就失明，这是我们知道的。
JOHN|9|21|至于他现在怎么能看见，我们却不知道；是谁开了他的眼睛，我们也不知道。他已经是成人，你们问他吧，他自己会说。”
JOHN|9|22|他父母说这些话，是怕 犹太 人，因为 犹太 人已经商定，若有宣认耶稣是基督的，要把他赶出会堂。
JOHN|9|23|因此他父母说“他已经是成人，你们问他吧”。
JOHN|9|24|于是法利赛人第二次叫了那以前失明的人来，对他说：“你要将荣耀归给上帝，我们知道这人是个罪人。”
JOHN|9|25|那人就回答：“他是不是个罪人，我不知道；有一件事我知道，我本来是失明的，现在我看见了。”
JOHN|9|26|他们就问他：“他给你做了什么？是怎么开了你的眼睛？”
JOHN|9|27|他回答他们：“我已经告诉你们了，你们不听，为什么又要听呢？难道你们也要作他的门徒吗？”
JOHN|9|28|他们就骂他：“你是他的门徒，而我们是 摩西 的门徒。
JOHN|9|29|上帝对 摩西 说话是我们知道的，可是这个人，我们不知道他从哪里来。”
JOHN|9|30|那人回答，对他们说：“他开了我的眼睛，你们竟不知道他从哪里来，这真是奇怪！
JOHN|9|31|我们知道上帝不听罪人，惟有敬奉上帝、遵行他旨意的，上帝才听他。
JOHN|9|32|从创世以来，未曾听见有人开了生来就失明的人的眼睛。
JOHN|9|33|这人若不是从上帝来的，什么也不能做。”
JOHN|9|34|他们回答他说：“你完全是生在罪中的，还要来教训我们吗？”于是他们把他赶出去了。
JOHN|9|35|耶稣听说他们把他赶出去，就找到他，说：“你信人子 吗？”
JOHN|9|36|那人回答说：“主啊，人子是谁？告诉我，好让我信他。”
JOHN|9|37|耶稣对他说：“你已经看见他，现在和你说话的就是他。”
JOHN|9|38|他说：“主啊，我信！”他就拜耶稣。
JOHN|9|39|耶稣说：“我为审判到这世上来，使不能看见的看见，能看见的反而失明。”
JOHN|9|40|同他在那里的法利赛人听见这些话，就对他说：“难道我们也失明了吗？”
JOHN|9|41|耶稣对他们说：“你们若是失明的，就没有罪了；但现在你们说‘我们能看见’，你们的罪还在。”
JOHN|10|1|“我实实在在地告诉你们，那不从门进羊圈，倒从别处爬进去的，就是贼，就是强盗。
JOHN|10|2|那从门进去的才是羊的牧人。
JOHN|10|3|看门的给他开门，羊也听他的声音。他按著名叫自己的羊，把羊领出来。
JOHN|10|4|当他把自己的羊都放出来，就走在前面，羊也跟着他，因为它们认得他的声音。
JOHN|10|5|羊绝不跟陌生人，反而会逃走，因为不认得陌生人的声音。”
JOHN|10|6|耶稣把这比方告诉他们，但他们不明白他所说的是什么。
JOHN|10|7|所以，耶稣又对他们说：“我实实在在地告诉你们，我就是羊的门。
JOHN|10|8|凡在我以前 来的都是贼，是强盗；羊没有听从他们。
JOHN|10|9|我就是门，凡从我进来的，必得安全 ，并且可进出，找到草吃。
JOHN|10|10|盗贼来，无非要偷窃，杀害，毁坏；我来了，是要羊得生命，并且得的更丰盛。
JOHN|10|11|“我是好牧人，好牧人为羊舍命。
JOHN|10|12|雇工不是牧人，羊不是他自己的，他一看见狼来，就撇下羊群逃跑；狼抓住羊，把它们赶散。
JOHN|10|13|雇工逃走，因为他是雇工，对羊毫不关心。
JOHN|10|14|我是好牧人；我认识我的羊，我的羊也认识我，
JOHN|10|15|正如父认识我，我也认识父一样；并且我为羊舍命。
JOHN|10|16|我另外有羊，不属这圈里的，我必须领它们来，它们也要听我的声音，并且要合成一群，归一个牧人。
JOHN|10|17|为此，我父爱我，因为我把命舍去，好再取回来。
JOHN|10|18|没有人夺去我的命，是我自己舍的；我有权舍弃，也有权再取回。这是我从我父所受的命令。”
JOHN|10|19|犹太 人为这些话又起了分裂。
JOHN|10|20|其中有好些人说：“他是被鬼附了，而且疯了，为什么听他的呢？”
JOHN|10|21|另有的说：“这不是被鬼附的人所说的话。鬼岂能开盲人的眼睛呢？”
JOHN|10|22|那时正是冬天，在 耶路撒冷 有献殿节。
JOHN|10|23|耶稣在圣殿里的 所罗门 廊下行走。
JOHN|10|24|犹太 人围着他，对他说：“你让我们犹豫不定到几时呢？你若是基督，就明白地告诉我们。”
JOHN|10|25|耶稣回答他们：“我已经告诉你们，你们却不信。我奉我父的名所行的事可以为我作见证。
JOHN|10|26|但是你们不信，因为你们不是我的羊。
JOHN|10|27|我的羊听我的声音，我认识它们，它们也跟从我。
JOHN|10|28|并且，我赐给他们永生；他们永不灭亡，谁也不能从我手里把他们夺去。
JOHN|10|29|我父所赐给我的比万有都大 ，谁也不能从我父手里把他们夺去。
JOHN|10|30|我与父原为一。”
JOHN|10|31|犹太 人又拿起石头来要打他。
JOHN|10|32|耶稣回应他们：“我做了许多从父那里来的善事给你们看，你们是为哪一件拿石头打我呢？”
JOHN|10|33|犹太 人回答他：“我们不是为了善事拿石头打你，而是为了你说亵渎的话；因为你是个人，却把自己当作上帝。”
JOHN|10|34|耶稣回答他们：“你们的律法书上不是写着‘我曾说你们是诸神’吗？
JOHN|10|35|经上的话是不能废的；如果那些领受上帝的道的人，上帝尚且称他们为诸神，
JOHN|10|36|那么父所分别为圣又差到世上来的那位说‘我是上帝的儿子’，你们还对他说‘你说亵渎的话’吗？
JOHN|10|37|我若不做我父的工作，你们就不必信我；
JOHN|10|38|我若做了，你们即使不信我，也当信这些工作，好让你们知道并且明白父在我里面，我也在父里面。”
JOHN|10|39|于是，他们又要捉拿他，他却从他们手中逃脱了。
JOHN|10|40|耶稣又往 约旦河 的东边去，到了 约翰 起初施洗的地方，就住在那里。
JOHN|10|41|有许多人来到他那里，说：“ 约翰 没有行过一件神迹，但 约翰 所说有关这人的一切话都是真的。”
JOHN|10|42|在那里，许多人信了耶稣。
JOHN|11|1|有一个患病的人，名叫 拉撒路 ，住在 伯大尼 ，就是 马利亚 和她姐姐 马大 的村庄。
JOHN|11|2|这 马利亚 就是那用香膏抹主，又用头发擦他脚的；患病的 拉撒路 是她的弟弟。
JOHN|11|3|姊妹两个就打发人去见耶稣，说：“主啊，你所爱的人病了。”
JOHN|11|4|耶稣听见后却说：“这病不至于死，而是为了上帝的荣耀，为要使上帝的儿子藉此得荣耀。”
JOHN|11|5|耶稣素来爱 马大 和她妹妹，以及 拉撒路 。
JOHN|11|6|他听见 拉撒路 病了，仍在原地住了两天，
JOHN|11|7|然后对门徒说：“我们再到 犹太 去吧！”
JOHN|11|8|门徒对他说：“拉比， 犹太 人近来要拿石头打你，你还再到那里去吗？”
JOHN|11|9|耶稣回答：“白天不是有十二小时吗？人若在白天行走，就不致跌倒，因为他看见这世上的光。
JOHN|11|10|人若在黑夜行走，就会跌倒，因为他没有光。”
JOHN|11|11|耶稣说了这些话，随后对他们说：“我们的朋友 拉撒路 睡了，我去叫醒他。”
JOHN|11|12|门徒就说：“主啊，他若睡了，就会好的。”
JOHN|11|13|耶稣说这话是指 拉撒路 死了，他们却以为他是指通常的睡眠。
JOHN|11|14|于是耶稣就明白地告诉他们：“ 拉撒路 死了。
JOHN|11|15|为了你们的缘故，我不在那里反而欢喜，为要使你们信。现在我们到他那里去吧。”
JOHN|11|16|于是那称为 低土马 的 多马 对其他的门徒说：“我们也去和他同死吧！”
JOHN|11|17|耶稣到了，知道 拉撒路 在坟墓里已经四天了。
JOHN|11|18|伯大尼 离 耶路撒冷 不远，约有六里 路。
JOHN|11|19|有好些 犹太 人来看 马大 和 马利亚 ，要为她们弟弟的缘故安慰她们。
JOHN|11|20|马大 听见耶稣来了，就出去迎接他； 马利亚 却仍然坐在家里。
JOHN|11|21|马大 对耶稣说：“主啊，你若早在这里，我弟弟就不会死了。
JOHN|11|22|我也知道，即使现在，你无论向上帝求什么，上帝也必赐给你。”
JOHN|11|23|耶稣对她说：“你弟弟会复活的。”
JOHN|11|24|马大 对他说：“我知道在末日复活的时候，他会复活。”
JOHN|11|25|耶稣对她说：“复活...也在我 。信我的人虽然死了，也必复活；
JOHN|11|26|凡活着信我的人必永远不死。你信这话吗？”
JOHN|11|27|马大 对他说：“主啊，是的。我信你是基督，是上帝的儿子，就是那要临到世界的。”
JOHN|11|28|马大 说了这话就回去，叫她妹妹 马利亚 ，私下说：“老师来了，他在叫你。”
JOHN|11|29|马利亚 听见了，急忙起来，到耶稣那里去。
JOHN|11|30|那时，耶稣还没有进村子，仍在 马大 迎接他的地方。
JOHN|11|31|那些同 马利亚 在家里安慰她的 犹太 人，见她急忙起来，出去，就跟着她，以为她要往坟墓那里去哭。
JOHN|11|32|马利亚 到了耶稣那里，看见他，就俯伏在他脚前，对他说：“主啊，你若早在这里，我弟弟就不会死了。”
JOHN|11|33|耶稣看见她哭，并看见与她同来的 犹太 人也哭，就心里悲叹，又甚忧愁，
JOHN|11|34|就说：“你们把他安放在哪里？”他们对他说：“主啊，请你来看。”
JOHN|11|35|耶稣哭了。
JOHN|11|36|犹太 人就说：“你看，他多么爱他！”
JOHN|11|37|其中有人说：“他既然开了盲人的眼睛，难道不能叫这人不死吗？”
JOHN|11|38|耶稣又心里悲叹，来到坟墓前。那坟墓是个穴，有一块石头挡着。
JOHN|11|39|耶稣说：“把石头挪开！”那死者的姐姐 马大 对他说：“主啊，他现在必定臭了，因为他已经死了四天了。”
JOHN|11|40|耶稣对她说：“我不是对你说过，你若信就必看见上帝的荣耀吗？”
JOHN|11|41|于是他们把石头挪开。耶稣举目望天，说：“父啊，我感谢你，因为你已经听了我。
JOHN|11|42|我知道你常常听我，但我说这话是为了周围站着的众人，要使他们信是你差了我来的。”
JOHN|11|43|说了这些话，他大声呼叫说：“ 拉撒路 ，出来！”
JOHN|11|44|那死了的人就出来了，手脚都裹着布，脸上包着头巾。耶稣对他们说：“解开他，让他走！”
JOHN|11|45|于是来看 马利亚 的 犹太 人中，有很多人见了耶稣所做的事，就信了他。
JOHN|11|46|但其中也有人去见法利赛人，把耶稣所做的事告诉他们。
JOHN|11|47|祭司长和法利赛人召开议会，说：“这人行好些神迹，我们怎么办呢？
JOHN|11|48|若让他这样做，人人都要信他； 罗马 人也要来毁灭我们的圣殿 和我们的民族。”
JOHN|11|49|其中有一个人，名叫 该亚法 ，那年当大祭司，对他们说：“你们什么都不知道，
JOHN|11|50|也不想想，一个人替百姓死，免得整个民族灭亡，这对你们是有利的。”
JOHN|11|51|他这话不是出于自己的意思，而是因他那年当大祭司，所以预言耶稣将为这民族而死。
JOHN|11|52|他不但替这民族死，还要把上帝四散的儿女都聚集起来，合成一群。
JOHN|11|53|从那日起，他们就商议要杀耶稣。
JOHN|11|54|所以，耶稣不再公开在 犹太 人中走动，却离开那里，往靠近旷野的乡间去，到了一座城，名叫 以法莲 ，就在那里和门徒住下来。
JOHN|11|55|犹太 人的逾越节近了，有许多人从乡下上 耶路撒冷 去，要在过节前洁净自己。
JOHN|11|56|于是他们寻找耶稣，站在圣殿里彼此说：“你们认为怎样，他不会来过节吧？”
JOHN|11|57|那时，祭司长和法利赛人早已下令，若有人知道耶稣的下落，就要报告，他们好去捉拿他。
JOHN|12|1|逾越节前六天，耶稣来到 伯大尼 ，就是他使 拉撒路 从死人中复活的地方。
JOHN|12|2|有人在那里为耶稣预备宴席； 马大 伺候， 拉撒路 也在同耶稣坐席的人中间。
JOHN|12|3|马利亚 拿着一斤极贵的纯哪哒 香膏，抹耶稣的脚，又用自己头发去擦，屋里充满了膏的香气。
JOHN|12|4|有一个门徒，就是那将要出卖耶稣的 加略 人 犹大 ，说：
JOHN|12|5|“为什么不把这香膏卖三百个银币去周济穷人呢？”
JOHN|12|6|他说这话，并不是关心穷人，而是因为他是个贼，又管钱囊，常偷取钱囊中所存的。
JOHN|12|7|耶稣说：“由她吧！她这香膏本是为我的安葬之日留着的。
JOHN|12|8|因为常有穷人和你们在一起，但是你们不常有我。”
JOHN|12|9|有一大群 犹太 人知道耶稣在那里，就来了，不但是为耶稣的缘故，也是要看耶稣使他从死人中复活的 拉撒路 。
JOHN|12|10|于是众祭司长商议连 拉撒路 也要杀了，
JOHN|12|11|因为有许多 犹太 人为了 拉撒路 的缘故，开始背离他们，信了耶稣。
JOHN|12|12|第二天，有一大群上来过节的人听见耶稣要来 耶路撒冷 ，
JOHN|12|13|就拿着棕树枝出去迎接他，喊着： “和散那 ， 以色列 的王！ 奉主名来的是应当称颂的！”
JOHN|12|14|耶稣找到了一匹驴驹，就骑上，如经上所记：
JOHN|12|15|“ 锡安 的儿女 啊，不要惧怕！ 看哪，你的王来了； 他骑在驴驹上。”
JOHN|12|16|门徒当初不明白这些事，等到耶稣得了荣耀后才想起这些话是指他写的，并且人们果然对他做了这些事。
JOHN|12|17|当耶稣呼唤 拉撒路 ，使他从死人中复活出坟墓的时候，同耶稣在那里的众人就作见证。
JOHN|12|18|众人因听见耶稣行了这神迹，就去迎接他。
JOHN|12|19|法利赛人彼此说：“你们看，你们一事无成，世人都随着他去了。”
JOHN|12|20|那时，上来过节礼拜的人中，有几个 希腊 人。
JOHN|12|21|他们来见 加利利 的 伯赛大 人 腓力 ，请求他说：“先生，我们想见耶稣。”
JOHN|12|22|腓力 去告诉 安得烈 ，然后 安得烈 同 腓力 去告诉耶稣。
JOHN|12|23|耶稣回答他们说：“人子得荣耀的时候到了。
JOHN|12|24|我实实在在地告诉你们，一粒麦子不落在地里死了，仍旧是一粒；若是死了，就结出许多子粒来。
JOHN|12|25|爱惜自己性命的，就丧失性命；那恨恶自己在这世上的性命的，要保全性命到永生。
JOHN|12|26|若有人服事我，就当跟从我；我在哪里，服事我的人也要在哪里；若有人服事我，我父必尊重他。”
JOHN|12|27|“我现在心里忧愁，我说什么才好呢？说‘父啊，救我脱离这时候’吗？但我正是为这时候来的。
JOHN|12|28|父啊，愿你荣耀你的名！”于是有声音从天上来，说：“我已经荣耀了我的名，还要再荣耀。”
JOHN|12|29|站在旁边的众人听见，就说：“打雷了。”另有的说：“有天使对他说话。”
JOHN|12|30|耶稣回答说：“这声音不是为我，而是为你们来的。
JOHN|12|31|现在正是这世界受审判的时候；现在这世界的统治者要被赶出去。
JOHN|12|32|我从地上被举起来的时候，我要吸引万人来归我。”
JOHN|12|33|耶稣这话是指自己将要怎样死说的。
JOHN|12|34|众人就回答他：“我们听见律法书上说，基督是永存的；你怎么说，人子必须被举起来呢？这人子是谁呢？”
JOHN|12|35|耶稣对他们说：“光在你们中间为时不多了，应该趁着有光的时候行走，免得黑暗临到你们；那在黑暗里行走的，不知道往何处去。
JOHN|12|36|你们趁着有光，要信从这光，使你们成为光明之子。” 耶稣说了这些话，就离开他们隐藏了。
JOHN|12|37|他虽然在他们面前行了许多神迹，他们还是不信他。
JOHN|12|38|这是要应验 以赛亚 先知所说的话： “主啊，我们所传的有谁信呢？ 主的膀臂向谁显露呢？”
JOHN|12|39|他们所以不能信，因为 以赛亚 又说：
JOHN|12|40|“主使他们瞎了眼， 使他们硬了心， 免得他们眼睛看见， 他们心里明白，回转过来， 我会医治他们。”
JOHN|12|41|以赛亚 因看见了他的荣耀，就说了关于他的这话。
JOHN|12|42|虽然如此，官长中却有好些信他的，只因法利赛人的缘故不敢承认，恐怕被赶出会堂。
JOHN|12|43|这是因他们爱人给的尊荣过于爱上帝给的尊荣。
JOHN|12|44|耶稣喊着说：“信我的人不是信我，而是信差我来的那位。
JOHN|12|45|看见我的，就是看见差我来的那位。
JOHN|12|46|我就是来到世上的光，使凡信我的不住在黑暗里。
JOHN|12|47|若有人听见我的话而不遵守，我不审判他，因为我来不是要审判世人，而是要拯救世人。
JOHN|12|48|弃绝我、不领受我话的人自有审判他的；我所讲的道在末日要审判他。
JOHN|12|49|因为我没有凭着自己讲，而是差我来的父已经给我命令，叫我说什么，讲什么。
JOHN|12|50|我也知道他的命令就是永生。所以，我讲的正是照着父所告诉我的，我就这么讲了。”
JOHN|13|1|逾越节以前，耶稣知道自己离世归父的时候到了。他一向爱世间属自己的人，就爱他们到底。
JOHN|13|2|晚餐的时候，魔鬼已把出卖耶稣的意思放在 加略 人 西门 的儿子 犹大 心里。
JOHN|13|3|耶稣知道父已把万有交在他手里，且知道自己是从上帝出来的，又要回到上帝那里去，
JOHN|13|4|就离席站起来，脱了衣服，拿一条手巾束腰，
JOHN|13|5|随后把水倒在盆里，开始洗门徒的脚，并用束腰的手巾擦干。
JOHN|13|6|到了 西门．彼得 跟前， 彼得 对他说：“主啊，你洗我的脚吗？”
JOHN|13|7|耶稣回答他说：“我所做的，你现在不知道，但以后会明白。”
JOHN|13|8|彼得 对他说：“你绝对不可以洗我的脚！”耶稣回答他：“我若不洗你，你就与我无份了。”
JOHN|13|9|西门．彼得 对他说：“主啊，不仅是我的脚，连手和头也要洗！”
JOHN|13|10|耶稣对他说：“凡洗过澡的人不需要再洗，只要把脚一洗，全身就干净了。你们是干净的，然而不都是干净的。”
JOHN|13|11|耶稣已知道要出卖他的是谁，因此说“你们不都是干净的”。
JOHN|13|12|耶稣洗完了他们的脚，就穿上衣服，又坐下，对他们说：“我为你们所做的，你们明白吗？
JOHN|13|13|你们称呼我老师，称呼我主，你们说的不错，我本来就是。
JOHN|13|14|我是你们的主，你们的老师，尚且洗你们的脚，你们也应当彼此洗脚。
JOHN|13|15|我给你们作了榜样，为要你们照着我为你们所做的去做。
JOHN|13|16|我实实在在地告诉你们，仆人不大于主人；奉差的人也不大于差他的人。
JOHN|13|17|你们既知道这些事，若是去实行就有福了。
JOHN|13|18|我不是指着你们众人说的，我知道我所拣选的是谁；但是要应验经上的话：‘吃我饭的人 用脚踢我。’
JOHN|13|19|事情还没有发生，我现在先告诉你们，让你们到事情发生的时候好信我就是那位。
JOHN|13|20|我实实在在地告诉你们，接纳我所差遣的就是接纳我；接纳我的就是接纳差遣我的那位。”
JOHN|13|21|耶稣说了这些话，心里忧愁，于是明确地说：“我实实在在地告诉你们，你们中间有一个人要出卖我。”
JOHN|13|22|门徒彼此相看，猜不出他说的是谁。
JOHN|13|23|门徒中有一个人，是耶稣所爱的，侧身挨近耶稣的胸怀。
JOHN|13|24|西门．彼得 就对这个人示意，要问耶稣是指着谁说的。
JOHN|13|25|于是那人紧靠着耶稣的胸膛，问他：“主啊，是谁呢？”
JOHN|13|26|耶稣回答：“我蘸一点饼给谁，就是谁。”耶稣就蘸了一点饼，递给 加略 人 西门 的儿子 犹大 。
JOHN|13|27|他接 了那饼以后，撒但就进入他的心。于是耶稣对他说：“你要做的，快做吧！”
JOHN|13|28|同席的人没有一个知道耶稣为什么对他说这话。
JOHN|13|29|有人因 犹大 管钱囊，以为耶稣是对他说“你去买我们过节所需要的东西”，或是叫他拿些什么给穷人。
JOHN|13|30|犹大 受 了那点饼以后立刻出去。那时候是夜间了。
JOHN|13|31|犹大 出去后，耶稣说：“如今人子得了荣耀，上帝在人子身上也得了荣耀。
JOHN|13|32|如果上帝因人子得了荣耀 ，上帝也要因自己荣耀人子，并且要立刻荣耀他。
JOHN|13|33|孩子们！我与你们同在的时候不多了；你们会找我，但我所去的地方，你们不能去。这话我曾对 犹太 人说过，现在也照样对你们说。
JOHN|13|34|我赐给你们一条新命令，乃是叫你们彼此相爱；我怎样爱你们，你们也要怎样彼此相爱。
JOHN|13|35|你们若彼此相爱，众人因此就认出你们是我的门徒了。”
JOHN|13|36|西门．彼得 问耶稣：“主啊，你去哪里？”耶稣回答：“我所去的地方，你现在不能跟我去，以后却要跟我去。”
JOHN|13|37|彼得 对他说：“主啊，为什么我现在不能跟你去？我愿意为你舍命。”
JOHN|13|38|耶稣回答：“你愿意为我舍命吗？我实实在在地告诉你，鸡叫以前，你要三次不认我。”
JOHN|14|1|“你们心里不要忧愁；你们信上帝，也当信我。
JOHN|14|2|在我父的家里有许多住处；若是没有，我就早已告诉你们了。我去原是为你们预备地去方。
JOHN|14|3|我若去为你们预备了地方，就必再来接你们到我那里去，我在哪里，叫你们也在哪里。
JOHN|14|4|我往哪里去，你们知道那条路。”
JOHN|14|5|多马 对他说：“主啊，我们不知道你去哪里，怎么能知道那条路呢？”
JOHN|14|6|耶稣对他说：“我就是道路、真理、生命；若不藉着我，没有人能到父那里去。
JOHN|14|7|既然你们认识了我，也会认识我的父。从今以后，你们就认识他，并且已经看见他了。”
JOHN|14|8|腓力 对他说：“主啊，将父显给我们看，我们就知足了。”
JOHN|14|9|耶稣对他说：“ 腓力 ，我与你们在一起这么久了，你还不认识我吗？看见我的就是看见了父，你怎么还说‘将父显给我们看’呢？
JOHN|14|10|我在父里面，父在我里面，你不信吗？我对你们所说的话不是凭着自己说的，而是住在我里面的父在做他的工作。
JOHN|14|11|你们要信我，我在父里面，父在我里面；即使不信，也要因我所做的工作信我。
JOHN|14|12|我实实在在地告诉你们，我所做的工作，信我的人也要做，并且要做得比这些更大，因为我到父那里去。
JOHN|14|13|你们奉我的名无论求什么，我必成全，为了使父因儿子得荣耀。
JOHN|14|14|你们若奉我的名向我求什么，我必成全。”
JOHN|14|15|“你们若爱我，就会遵守我的命令。
JOHN|14|16|我要求父，父就赐给你们另外一位保惠师 ，使他永远与你们同在。
JOHN|14|17|他就是真理的灵，是世人不能接受的。因为他们既看不见他，也不认识他；你们却认识他，因他常与你们同在，也要在你们里面。
JOHN|14|18|我不会撇下你们为孤儿，我必到你们这里来。
JOHN|14|19|再过不久，世人不再看见我，你们却会看见我，因为我活着，你们也要活着。
JOHN|14|20|到那日，你们就会知道我在父里面，你们在我里面，我也在你们里面。
JOHN|14|21|有了我的命令而又遵守的人，就是爱我的；爱我的人，我父要爱他，我也要爱他，并且要亲自向他显现。”
JOHN|14|22|犹大 （不是 加略 人 犹大 ）问耶稣：“主啊，为什么亲自向我们显现，而不向世人显现呢？”
JOHN|14|23|耶稣回答他说：“凡爱我的人就会遵守我的道，我父也会爱他，并且我们要到他那里去，与他同住。
JOHN|14|24|不爱我的人就不遵守我的道。你们所听见的道不是我的，而是差我来之父的。
JOHN|14|25|“我还与你们在一起的时候，已对你们说了这些事。
JOHN|14|26|但保惠师，就是父因我的名所要差来的圣灵，他要把一切的事教导你们，并且要使你们想起我对你们所说的一切话。
JOHN|14|27|我留下平安给你们，我把我的平安赐给你们。我所赐给你们的，不像世人所赐的。你们心里不要忧愁，也不要胆怯。
JOHN|14|28|你们听见我对你们说过，我去了还要回到你们这里来。你们若爱我，就会因我到父那里去而喜乐，因为父比我大。
JOHN|14|29|现在事情还没有发生，我预先告诉你们，使你们在事情发生的时候会信。
JOHN|14|30|我不再和你们多说了，因为这世界的统治者将到，他在我身上一无所能。
JOHN|14|31|我这么做是照着父命令我的，为了让世人知道我爱父。起来，我们走吧！”
JOHN|15|1|“我就是真葡萄树，我父是栽培的人。
JOHN|15|2|凡属我不结果子的枝子，他就剪掉；凡结果子的，他就修剪干净，使枝子结果子更多。
JOHN|15|3|现在你们因我讲给你们的道已经洁净了。
JOHN|15|4|你们要常在我里面，我也常在你们里面。枝子若不常在葡萄树上，自己就不能结果子；你们若不常在我里面，也是这样。
JOHN|15|5|我就是葡萄树，你们是枝子。常在我里面的，我也常在他里面，这人就多结果子，因为离了我，你们就不能做什么。
JOHN|15|6|人若不常在我里面，就像枝子被丢在外面，枯干了，人捡起来，扔进火里烧了。
JOHN|15|7|你们若常在我里面，我的话也常在你们里面，凡你们想要的，祈求，就给你们成全。
JOHN|15|8|你们多结果子，我父就因此得荣耀，你们也就是 我的门徒了。
JOHN|15|9|我爱你们，正如父爱我一样；你们要常在我的爱里。
JOHN|15|10|你们若遵守我的命令，就会常在我的爱里，正如我遵守了我父的命令，常在他的爱里。
JOHN|15|11|“我已对你们说了这些事，是要让我的喜乐存在你们心里，并让你们的喜乐得以满足。
JOHN|15|12|你们要彼此相爱，像我爱你们一样，这是我的命令。
JOHN|15|13|人为朋友舍命，人的爱心没有比这个更大的了。
JOHN|15|14|你们若遵行我所命令的，就是我的朋友。
JOHN|15|15|以后我不再称你们为仆人，因为仆人不知道主人所做的事；但我称你们为朋友，因为我从我父所听见的一切都已经让你们知道了。
JOHN|15|16|不是你们拣选了我，而是我拣选了你们，并且派你们去结果子，让你们的果子得以长存，好使你们奉我的名，无论向父求什么，他会赐给你们。
JOHN|15|17|我这样命令你们，是要你们彼此相爱。”
JOHN|15|18|“世人若恨你们，你们要知道，他们在恨你们以前已经恨我了。
JOHN|15|19|你们若属世界，世界会爱属自己的；只因你们不属世界，而是我从世界中拣选了你们，所以世界就恨你们。
JOHN|15|20|你们要记得我对你们说过的话：‘仆人不大于主人。’他们若迫害了我，也会迫害你们，他们若遵守了我的话，也会遵守你们的话。
JOHN|15|21|但他们要因我的名向你们做这一切的事，因为他们不认识差我来的那位。
JOHN|15|22|我若没有来教导他们，他们就没有罪；但如今他们的罪无可推诿了。
JOHN|15|23|恨我的也恨我的父。
JOHN|15|24|我若没有在他们中间做过别人未曾做的事，他们就没有罪；但如今连我与我的父，他们也看见了，也恨恶了。
JOHN|15|25|这是要应验他们律法上所写的话：‘他们无故地恨我。’
JOHN|15|26|“但我要从父那里差保惠师来，就是从父出来的那真理的灵，他来的时候要为我作见证。
JOHN|15|27|你们也要作见证，因为你们从起初就与我同在。”
JOHN|16|1|“我对你们说了这些事，是要使你们不至于跌倒。
JOHN|16|2|人要把你们赶出会堂，而且时候将到，凡杀你们的还以为是在事奉上帝。
JOHN|16|3|他们这样做，是因为没有认识父，也没有认识我。
JOHN|16|4|我对你们说了这些事，是要在他们做这些事的时候，你们会想起我对你们说过的话。” “我起先没有对你们说这些事，因为我一直与你们同在。
JOHN|16|5|现在我要到差我来的父那里去，你们中间却没有人问我‘你去哪里？’
JOHN|16|6|只因我对你们说了这些事，你们就满心忧愁。
JOHN|16|7|然而，我把真情告诉你们，我去对你们是有益的。我若不去，保惠师就不会到你们这里来；我若去，就差他到你们这里来。
JOHN|16|8|他来的时候，要为罪、为义，为审判，指证世人；
JOHN|16|9|为罪，是因他们不信我；
JOHN|16|10|为义，是因我到父那里去，你们将不再见到我；
JOHN|16|11|为审判，是因这世界的统治者已受了审判。
JOHN|16|12|“我还有好些事要告诉你们，但你们现在担当不了 。
JOHN|16|13|但真理的灵来的时候，他要引导你们进入一切真理。因为他不是凭着自己说的，而是把他所听见的都说出来，并且要把将要来的事向你们传达。
JOHN|16|14|他要荣耀我，因为他要把从我领受的向你们传达。
JOHN|16|15|凡父所有的都是我的，所以我说，他要把从我领受的向你们传达。”
JOHN|16|16|“不久，你们将不再见到我；再过不久，你们还要见到我。”
JOHN|16|17|有几个门徒彼此说：“他对我们说‘不久，你们将不再见到我；再过不久，你们还要见到我’；又说‘因我到父那里去’。这是什么意思呢？”
JOHN|16|18|于是门徒说：“他说 ‘不久’到底是什么意思呢？我们不明白他说什么。”
JOHN|16|19|耶稣看出他们要问他，就对他们说：“我说‘不久，你们将不再见到我；再过不久，你们还要见到我’，你们为这话彼此询问吗？
JOHN|16|20|我实实在在地告诉你们，你们将要痛哭，哀号，世人反要欢喜。你们将要忧愁，然而你们的忧愁要变成喜乐。
JOHN|16|21|妇人生产的时候会忧愁，因为她的时候到了；但孩子一生出来，就不再记得那痛苦了，因为欢喜有一个人生在世上了。
JOHN|16|22|你们现在也是忧愁，但我要再见到你们，你们的心就会有喜乐了；这喜乐没有人能夺去。
JOHN|16|23|到那日，你们什么也不会问我了。我实实在在地告诉你们，你们奉我的名无论向父求什么，他会赐给你们 。
JOHN|16|24|直到现在，你们没有奉我的名求什么，如今你们求就必得着，使你们的喜乐得以满足。”
JOHN|16|25|“这些事，我是用比方对你们说的；时候将到，我不再用比方对你们说，而是要把父的事明白地告诉你们。
JOHN|16|26|到那日，你们要奉我的名祈求；我并不对你们说，我要为你们向父祈求。
JOHN|16|27|父自己爱你们，因为你们已经爱我，又信我是从上帝 而来的。
JOHN|16|28|我从父而来，到了世界 ，又离开世界，到父那里去。”
JOHN|16|29|门徒说：“你看，如今你是明说，不用比方了。
JOHN|16|30|现在我们晓得你凡事都知道，也不需要有人问你；从此我们信你是从上帝而来的。”
JOHN|16|31|耶稣回答他们：“现在你们信了吗？
JOHN|16|32|看哪，时候将到，其实已经到了，你们要分散，各归自己的地方，留下我独自一人；然而我不是独自一人，因为有父与我同在。
JOHN|16|33|我对你们说了这些事，是要使你们在我里面有平安。在世上你们有苦难，但你们要有勇气 ，我已经胜过世界。”
JOHN|17|1|耶稣说了这些话，就举目望天，说：“父啊，时候到了，愿你荣耀你的儿子，使儿子也荣耀你；
JOHN|17|2|因为你曾赐给他权柄掌管凡血肉之躯的，使他把永生赐给你所赐给他的人。
JOHN|17|3|认识你—独一的真神，并且认识你所差来的耶稣基督，这就是永生。
JOHN|17|4|我在地上已经荣耀你，你交给我做的工作，我已完成了。
JOHN|17|5|父啊，现在求你使我在你面前得荣耀，就是在未有世界以前，我同你享有的荣耀。
JOHN|17|6|“你从世上赐给我的人，我已把你的名显明给他们。他们本是你的，你把他们赐给我，他们也遵守了你的道。
JOHN|17|7|现在他们知道，你所赐给我的一切都是从你那里来的；
JOHN|17|8|因为你所赐给我的话，我已经赐给他们，他们也领受了，又确实知道，我是从你出来的，并且信你差了我来。
JOHN|17|9|我为他们祈求，不为世人祈求，却为你所赐给我的人祈求，因他们本是你的。
JOHN|17|10|凡是我的都是你的，你的也是我的，并且我因他们得了荣耀。
JOHN|17|11|我到你那里去；我不再留在世上，他们却在世上。圣父啊，求你因你的名，就是你所赐给我的名，保守他们，使他们像我们一样合而为一。
JOHN|17|12|我与他们同在的时候，我奉你的名，就是你所赐给我的名，保守了他们，我也护卫了他们；其中除了那灭亡之子，没有一个灭亡的，好使经上的话得以应验。
JOHN|17|13|现在我到你那里去，我在世上说这些话，是要他们心里充满了我的喜乐。
JOHN|17|14|我已把你的道赐给他们；世界恨他们，因为他们不属世界，正如我不属世界一样。
JOHN|17|15|我不求你把他们从世上接走，只求你保全他们，使他们脱离那恶者。
JOHN|17|16|他们不属世界，正如我不属世界一样。
JOHN|17|17|求你用真理使他们成圣；你的道就是真理。
JOHN|17|18|你怎样差我到世上，我也照样差他们到世上。
JOHN|17|19|我为他们的缘故使自己分别为圣，为要使他们也因真理成圣。
JOHN|17|20|“我不但为这些人祈求，也为那些藉着他们的话信我的人祈求，
JOHN|17|21|使他们都合而为一。正如父你在我里面，我在你里面，使他们也在我们里面，好让世人信是你差我来的。
JOHN|17|22|你所赐给我的荣耀，我已赐给他们，使他们合而为一，像我们合而为一。
JOHN|17|23|我在他们里面，你在我里面，使他们完完全全合而为一，让世人知道是你差我来的，也知道你爱他们，如同爱我一样。
JOHN|17|24|父啊，我在哪里，愿你所赐给我的人也同我在哪里，使他们看见你所赐给我的荣耀，因为创世以前，你已经爱我了。
JOHN|17|25|公义的父啊，世人未曾认识你，我却认识你，这些人也知道是你差我来的。
JOHN|17|26|我已让他们认识你的名，还要让他们认识，好让你爱我的爱在他们里面，我也在他们里面。”
JOHN|18|1|耶稣说了这些话，就同门徒出去，过了 汲沦溪 。在那里有一个园子，他和门徒进去了。
JOHN|18|2|出卖耶稣的 犹大 也知道那地方，因为耶稣和门徒屡次在那里聚集。
JOHN|18|3|犹大 领了一队兵，以及祭司长和法利赛人的圣殿警卫，拿着灯笼、火把和兵器来到园里。
JOHN|18|4|耶稣知道将要临到自己的一切事，就出来对他们说：“你们找谁？”
JOHN|18|5|他们回答他：“ 拿撒勒 人耶稣。”耶稣对他们说：“我就是。”出卖他的 犹大 也同他们站在一起。
JOHN|18|6|耶稣一对他们说“我就是”，他们就退后，倒在地上。
JOHN|18|7|他又问他们：“你们找谁？”他们说：“ 拿撒勒 人耶稣。”
JOHN|18|8|耶稣回答：“我已经告诉你们，我就是。你们若找的是我，就让这些人走吧。”
JOHN|18|9|这要应验耶稣说过的话：“你所赐给我的人，我一个也不失落。”
JOHN|18|10|西门．彼得 带着一把刀，就拔出来，把大祭司的仆人砍了一刀，削掉了他的右耳，那仆人名叫 马勒古 。
JOHN|18|11|于是耶稣对 彼得 说：“收刀入鞘吧！我父给我的杯，我岂可不喝呢？”
JOHN|18|12|那队兵、千夫长和 犹太 人的警卫拿住耶稣，把他捆绑了，
JOHN|18|13|先带到 亚那 面前，因为他是那年的大祭司 该亚法 的岳父。
JOHN|18|14|这 该亚法 就是从前向 犹太 人忠告说“一个人替百姓死是有利的”那个人。
JOHN|18|15|西门．彼得 跟着耶稣，另一个门徒也跟着；那门徒是大祭司所认识的，他就同耶稣进了大祭司的院子。
JOHN|18|16|彼得 却站在门外。大祭司所认识的那个门徒出来，对看门的使女说了一声，就领 彼得 进去。
JOHN|18|17|那看门的使女对 彼得 说：“你不也是这人的门徒吗？”他说：“我不是。”
JOHN|18|18|仆人和警卫因为天冷生了炭火，站在那里取暖； 彼得 也同他们站着取暖。
JOHN|18|19|于是，大祭司盘问耶稣有关他的门徒和他教导的事。
JOHN|18|20|耶稣回答他：“我一向都是公开地对世人讲话，我常在会堂和圣殿里，就是 犹太 人聚集的地方教导人，我私下并没有讲什么。
JOHN|18|21|你为什么问我呢？去问那些听过我讲话的人，我所说的，他们都知道。”
JOHN|18|22|耶稣说了这些话，旁边站着的一个警卫打了他一耳光，说：“你这样回答大祭司吗？”
JOHN|18|23|耶稣回答他：“假如我说的不对，你指证不对的地方；假如我说的对，你为什么打我呢？”
JOHN|18|24|于是 亚那 把耶稣绑着押解到大祭司 该亚法 那里。
JOHN|18|25|西门．彼得 正站着取暖，有人对他说：“你不也是他的门徒吗？” 彼得 不承认，说：“我不是。”
JOHN|18|26|大祭司的一个仆人，是被 彼得 削掉耳朵那人的亲属，说：“我不是看见你同他在园子里吗？”
JOHN|18|27|彼得 又不承认，立刻鸡就叫了。
JOHN|18|28|他们把耶稣从 该亚法 那里押解到总督府。那时是清早。他们自己却不进总督府，恐怕染了污秽，不能吃逾越节的宴席。
JOHN|18|29|于是 彼拉多 出来，到他们那里，说：“你们告这人是为什么事呢？”
JOHN|18|30|他们回答他说：“这人若不作恶，我们就不会把他交给你了。”
JOHN|18|31|彼拉多 对他们说：“你们自己带他去，按着你们的律法问他吧！” 犹太 人说：“我们没有杀人的权柄。”
JOHN|18|32|这是要应验耶稣所说，指自己将要怎样死的话。
JOHN|18|33|于是 彼拉多 又进了总督府，叫耶稣来，对他说：“你是 犹太 人的王吗？”
JOHN|18|34|耶稣回答：“这话是你说的，还是别人论到我时对你说的呢？”
JOHN|18|35|彼拉多 回答：“难道我是 犹太 人吗？你的同胞和祭司长把你交给我。你做了什么事呢？”
JOHN|18|36|耶稣回答：“我的国不属于这世界；我的国若属于这世界，我的部下就会为我战斗，使我不至于被交给 犹太 人。只是我的国不属于这世界。”
JOHN|18|37|于是 彼拉多 对他说：“那么，你是王了？”耶稣回答：“是你说我是王。我为此而生，也为此来到世界，为了给真理作见证。凡属真理的人都听我的话。”
JOHN|18|38|彼拉多 对他说：“真理是什么呢？” 说了这话， 彼拉多 又出来到 犹太 人那里，对他们说：“我查不出他有什么罪状。
JOHN|18|39|但你们有个规矩，在逾越节要我给你们释放一个人，你们要我给你们释放这 犹太 人的王吗？”
JOHN|18|40|他们又再喊着说：“不要这人！要 巴拉巴 ！”这 巴拉巴 是个强盗。
JOHN|19|1|于是， 彼拉多 命令把耶稣带去鞭打了。
JOHN|19|2|士兵用荆棘编了冠冕，戴在他头上，给他穿上紫袍，
JOHN|19|3|又走到他面前，说：“万岁， 犹太 人的王！”他们就打他耳光。
JOHN|19|4|彼拉多 又出来对众人说：“看，我带他出来见你们，让你们知道我查不出他有什么罪状。”
JOHN|19|5|耶稣出来，戴着荆棘冠冕，穿着紫袍。 彼拉多 对他们说：“看哪，这个人！”
JOHN|19|6|祭司长和圣殿警卫看见他，就喊着说：“钉十字架！钉十字架！” 彼拉多 对他们说：“你们自己把他带去钉十字架吧！我查不出他有什么罪状。”
JOHN|19|7|犹太 人回答他：“我们有律法，按照律法，他是该死的，因为他自以为是上帝的儿子。”
JOHN|19|8|彼拉多 听见这话，越发害怕，
JOHN|19|9|又进了总督府，对耶稣说：“你是哪里来的？”耶稣却不回答。
JOHN|19|10|于是 彼拉多 对他说：“你不对我说话吗？难道你不知道我有权柄释放你，也有权柄把你钉十字架吗？”
JOHN|19|11|耶稣回答他：“若不是从上头赐给你的，你就毫无权柄办我，所以，把我交给你的那人罪更重了。”
JOHN|19|12|从此， 彼拉多 想要释放耶稣，无奈 犹太 人喊着说：“你若释放这个人，你就不是凯撒的忠臣 。凡自立为王的就是背叛凯撒。”
JOHN|19|13|彼拉多 听见这些话，就带耶稣出来，到了一个地方，叫“铺华石处”， 希伯来 话叫 厄巴大 ，就在那里坐堂。
JOHN|19|14|那日是逾越节的预备日，约在正午。 彼拉多 对 犹太 人说：“看哪，你们的王！”
JOHN|19|15|他们就喊着：“除掉他！除掉他！把他钉十字架！” 彼拉多 对他们说：“要我把你们的王钉十字架吗？”祭司长回答：“除了凯撒，我们没有王。”
JOHN|19|16|于是 彼拉多 把耶稣交给他们去钉十字架。 他们就把耶稣带了去。
JOHN|19|17|耶稣背着自己的十字架出来，到了一个地方，名叫“髑髅地”， 希伯来 话叫 各各他 。
JOHN|19|18|他们就在那里把他钉在十字架上，还有两个人和他一同被钉，一边一个，耶稣在中间。
JOHN|19|19|彼拉多 又写了一个牌子，钉在十字架上，写的是：“ 犹太 人的王， 拿撒勒 人耶稣。”
JOHN|19|20|有许多 犹太 人念这牌子，因为耶稣被钉十字架的地方靠近城，而且牌子是用 希伯来 、 罗马 、 希腊 三种文字写的。
JOHN|19|21|犹太 人的祭司长就对 彼拉多 说：“不要写‘ 犹太 人的王’，要写‘那人说：我是 犹太 人的王’。”
JOHN|19|22|彼拉多 回答：“我写了就写了。”
JOHN|19|23|士兵把耶稣钉在十字架上以后，把他的衣服拿来分为四份，每人一份。他们又拿他的内衣，这件内衣没有缝，是上下一片织成的。
JOHN|19|24|他们就彼此说：“我们不要撕开，我们抽签，看是谁的。”这要应验经上的话说： “他们分了我的外衣， 为我的内衣抽签。” 士兵果然做了这些事。
JOHN|19|25|站在耶稣十字架旁边的，有他的母亲、姨母、 革罗罢 的妻子 马利亚 ，和 抹大拉 的 马利亚 。
JOHN|19|26|耶稣见母亲和他所爱的那门徒站在旁边，就对母亲说：“母亲 ，看，你的儿子！”
JOHN|19|27|又对那门徒说：“看，你的母亲！”从那刻起，那门徒就接她到自己家里去了。
JOHN|19|28|这事以后，耶稣知道各样的事已经成了，为使经上的话应验，就说：“我渴了。”
JOHN|19|29|有一个盛满了醋的罐子放在那里，他们就拿海绵蘸满了醋，绑在牛膝草上，送到他嘴边。
JOHN|19|30|耶稣尝了那醋，说：“成了！”就低下头，断了气 。
JOHN|19|31|因为这日是预备日，又因为那安息日是个大日子， 犹太 人就来求 彼拉多 叫人打断他们的腿，把他们搬走，免得尸首在安息日留在十字架上。
JOHN|19|32|于是士兵来，把第一个人的腿，和与耶稣同钉的另一个人的腿，都打断了。
JOHN|19|33|当他们来到耶稣那里，见他已经死了，就没有打断他的腿。
JOHN|19|34|然而有一个士兵拿枪扎他的肋旁，立刻有血和水流出来。
JOHN|19|35|看见这事的人作了见证—他的见证是真的，他知道自己所说的是真的—好让你们也信。
JOHN|19|36|这些事发生，为要应验经上的话：“他的骨头一根也不可折断。”
JOHN|19|37|另有经文也说：“他们要仰望自己所扎的人。”
JOHN|19|38|这些事以后， 亚利马太 的 约瑟 来求 彼拉多 ，要把耶稣的身体领去。他是耶稣的门徒，只因怕 犹太 人，就暗地里作门徒。 彼拉多 准许了，他就把耶稣的身体领走。
JOHN|19|39|尼哥德慕 也来了，就是先前夜里去见耶稣的那位，他带着约一百斤的没药和沉香。
JOHN|19|40|他们照 犹太 人丧葬的规矩，用细麻布加上香料，把耶稣的身体裹好了。
JOHN|19|41|在耶稣钉十字架的地方有一个园子，园子里有一座新墓穴，是从来没有葬过人的。
JOHN|19|42|因为那天是 犹太 人的预备日，而那坟墓又在附近，他们就把耶稣安放在那里。
JOHN|20|1|七日的第一日清早，天还黑的时候， 抹大拉 的 马利亚 来到坟墓，看见石头已从坟墓挪开了，
JOHN|20|2|就跑来见 西门．彼得 和耶稣所爱的那个门徒，对他们说：“有人从坟墓里把主移走了，我们不知道他们把他放在哪里。”
JOHN|20|3|彼得 和那门徒就出来，往坟墓去。
JOHN|20|4|两个人同跑，那门徒比 彼得 跑得快，先到了坟墓，
JOHN|20|5|低头往里看，看见细麻布还放在那里，只是没有进去。
JOHN|20|6|西门．彼得 随后也到了，进了坟墓，看见细麻布放在那里，
JOHN|20|7|又看见耶稣的裹头巾没有和细麻布放在一起，是另在一处卷着。
JOHN|20|8|然后先到坟墓的那门徒也进去，他看见就信了。
JOHN|20|9|他们还不明白圣经所说耶稣必须从死人中复活的意思。
JOHN|20|10|于是两个门徒回自己的住处去了。
JOHN|20|11|马利亚 却站在坟墓外面哭。她哭的时候，低头往坟墓里看，
JOHN|20|12|看见两个天使穿着白衣，在安放耶稣身体的地方坐着，一个在头，一个在脚。
JOHN|20|13|天使对她说：“妇人，你为什么哭？”她对他们说：“因为有人把我主移走了，我不知道他们把他放在哪里。”
JOHN|20|14|说了这些话，她转过身来，看见耶稣站在那里，却不知道他是耶稣。
JOHN|20|15|耶稣问她：“妇人，你为什么哭？你找谁？” 马利亚 以为他是看园子的，就对他说：“先生，若是你把他移了去，请告诉我，你把他放在哪里，我去把他移回来。”
JOHN|20|16|耶稣对她说：“ 马利亚 。” 马利亚 转过身来，用 希伯来 话对他说：“拉波尼！”（“拉波尼”就是老师的意思。）
JOHN|20|17|耶稣对她说：“不要拉住我，因为我还没有升上去见我的父。你到我弟兄那里去告诉他们，我要升上去见我的父，也是你们的父，见我的上帝，也是你们的上帝。”
JOHN|20|18|抹大拉 的 马利亚 就向门徒报信：“我已经看见了主。”她又把主对她说的话告诉他们。
JOHN|20|19|那日（就是七日的第一日）晚上，门徒因怕 犹太 人，所在的地方门都关了。耶稣来，站在当中，对他们说：“愿你们平安！”
JOHN|20|20|说了这话，他把手和肋旁给他们看。门徒一看见主就喜乐了。
JOHN|20|21|于是耶稣又对他们说：“愿你们平安！父怎样差遣了我，我也照样差遣你们。”
JOHN|20|22|说了这话，他向他们吹一口气，说：“领受圣灵吧！
JOHN|20|23|你们赦免谁的罪，谁的罪就得赦免；你们不赦免谁的罪，谁的罪就不得赦免。”
JOHN|20|24|那十二使徒中，有个叫 低土马 的 多马 ，耶稣来的时候，他没有和他们在一起。
JOHN|20|25|其他的门徒就对他说：“我们已经看见主了。” 多马 却对他们说：“除非我看见他手上的钉痕，用我的指头探入那钉痕，用我的手探入他的肋旁，我绝不信。”
JOHN|20|26|过了八日，门徒又在屋里， 多马 也和他们在一起。门都关了，耶稣来，站在当中，说：“愿你们平安！”
JOHN|20|27|然后他对 多马 说：“把你的指头伸到这里来，看看我的手；把你的手伸过来，探入我的肋旁。不要疑惑，总要信！”
JOHN|20|28|多马 回答，对他说：“我的主！我的上帝！”
JOHN|20|29|耶稣对他说：“你因为看见了我才信吗？那没有看见却信的有福了。”
JOHN|20|30|耶稣在他门徒面前另外行了许多神迹，没有记录在这书上。
JOHN|20|31|但记载这些事是要使你们信 耶稣是基督，是上帝的儿子，并且使你们信他，好因着他的名得生命。
JOHN|21|1|这些事以后，耶稣在 提比哩亚 海边又向门徒显现。他怎样显现记在下面。
JOHN|21|2|西门．彼得 、叫 低土马 的 多马 、 加利利 的 迦拿 人 拿但业 、 西庇太 的两个儿子，和另外两个门徒，都在一起。
JOHN|21|3|西门．彼得 对他们说：“我打鱼去。”他们对他说：“我们也和你一起去。”他们就出去，上了船；那一夜并没有打着什么。
JOHN|21|4|天刚亮的时候，耶稣站在岸上，门徒却不知道他是耶稣。
JOHN|21|5|耶稣就对他们说：“孩子们！你们有吃的没有？”他们回答他：“没有。”
JOHN|21|6|耶稣对他们说：“你们把网撒在船的右边，就会得到。”于是他们撒下网去，竟拉不上来了，因为鱼很多。
JOHN|21|7|耶稣所爱的那门徒对 彼得 说：“是主！”那时 西门．彼得 赤着身子，一听见是主，就束上外衣，跳进海里。
JOHN|21|8|其余的门徒因离岸不远，约有二百肘，就坐着小船把那网鱼拉过来。
JOHN|21|9|他们上了岸，看见那里有炭火，上面有鱼和饼。
JOHN|21|10|耶稣对他们说：“把刚才打的鱼拿几条来。”
JOHN|21|11|西门．彼得 就上船，把网拉到岸上，网里满了大鱼，共一百五十三条；虽然鱼这样多，网却没有破。
JOHN|21|12|耶稣对他们说：“你们来吃早饭。”门徒中没有一个敢问他：“你是谁？”因为他们知道他是主。
JOHN|21|13|耶稣走过来，拿饼给他们，也照样拿鱼给他们。
JOHN|21|14|耶稣从死人中复活后向门徒显现，这是第三次。
JOHN|21|15|他们吃完了早饭，耶稣对 西门．彼得 说：“ 约翰 的儿子 西门 ，你爱我比这些更深吗？” 彼得 对他说：“主啊，是的，你知道我爱你。”耶稣对他说：“你喂养我的小羊。”
JOHN|21|16|耶稣第二次又对他说：“ 约翰 的儿子 西门 ，你爱我吗？” 彼得 对他说：“主啊，是的，你知道我爱你。”耶稣说：“你牧养我的羊。”
JOHN|21|17|耶稣第三次对他说：“ 约翰 的儿子 西门 ，你爱我吗？” 彼得 因为耶稣第三次对他说“你爱我吗”，就忧愁，对耶稣说：“主啊，你无所不知，你知道我爱你。”耶稣说：“你喂养我的羊。
JOHN|21|18|我实实在在地告诉你，你年轻的时候，自己束上带子，随意往来；但年老的时候，你要伸出手来，别人要把你束上，带你到不愿意去的地方。”
JOHN|21|19|耶稣说这话，是指 彼得 会怎样死来荣耀上帝。说了这话，耶稣对他说：“你跟从我吧！”
JOHN|21|20|彼得 转过身来，看见耶稣所爱的那门徒跟着，就是在晚餐时靠着耶稣胸膛说“主啊，出卖你的是谁”的那门徒。
JOHN|21|21|彼得 看见他，就问耶稣：“主啊，这个人怎样呢？”
JOHN|21|22|耶稣对他说：“假如我要他等到我来的时候还在，跟你有什么关系呢？你跟从我吧！”
JOHN|21|23|于是这话在弟兄中间流传，说那门徒不死。其实，耶稣不是说他不死，而是对 彼得 说：“假如我要他等到我来的时候还在，跟你有什么关系呢？ ”
JOHN|21|24|这门徒就是为这些事作见证、并且记载这些事的，我们知道他的见证是真的。
JOHN|21|25|耶稣所行的事还有许多，若是一一都写出来，我想，就是全世界也容不下所要写的书。
ACTS|1|1|提阿非罗 啊，我在第一本书中已论到耶稣从开头所做和所教导的一切事，
ACTS|1|2|直到他藉着圣灵吩咐所拣选的使徒后，被接上升的日子为止。
ACTS|1|3|他受害以后，用许多确据向使徒显明自己是活着的，在四十天之中向他们显现，并讲说上帝国的事。
ACTS|1|4|耶稣和他们聚集的时候，嘱咐他们说：“不要离开 耶路撒冷 ，但要等候父的应许，就是你们听见我说过的。
ACTS|1|5|约翰 是用水施洗，但过了不多几天，你们要在圣灵里受洗。”
ACTS|1|6|他们聚集的时候，问耶稣：“主啊，你就要在这时候复兴 以色列 国吗？”
ACTS|1|7|耶稣对他们说：“父凭着自己的权柄所定的时候和日期，不是你们可以知道的。
ACTS|1|8|但圣灵降临在你们身上，你们就必得着能力，并要在 耶路撒冷 、 犹太 全地和 撒玛利亚 ，直到地极，作我的见证。”
ACTS|1|9|说了这些话，他们正看的时候，他被接上升，有一朵云彩从他们眼前把他接去。
ACTS|1|10|他升上去的时候，他们定睛望天，看哪，有两个人身穿白衣站在他们旁边，
ACTS|1|11|说：“ 加利利 人哪，你们为什么站着望天呢？这离开你们被接升天的耶稣，你们见他怎样升上天去，他也要怎样来临。”
ACTS|1|12|有一座山，名叫 橄榄山 ，离 耶路撒冷 不远，有安息日可行走的路程 。那时，门徒从那里回 耶路撒冷 去，
ACTS|1|13|他们一进城，就上了所住的楼房；在那里有 彼得 、 约翰 、 雅各 、 安得烈 、 腓力 、 多马 、 巴多罗买 、 马太 、 亚勒腓 的儿子 雅各 、激进党的 西门 ，和 雅各 的儿子 犹大 。
ACTS|1|14|这些人和几个妇人，包括耶稣的母亲 马利亚 ，和耶稣的兄弟，都同心合意地恒切祷告。
ACTS|1|15|那时，有许多人聚会，约有一百二十名， 彼得 在弟兄中间站起来，说：
ACTS|1|16|“诸位弟兄，圣经的话必须应验。圣经中，圣灵曾藉 大卫 的口预先说到那领人来拿耶稣的 犹大 ；
ACTS|1|17|他本来算是我们中的一个，并且得了这一份使徒的职任。
ACTS|1|18|这人用他不义的代价买了一块田，以后身子仆倒，肚腹崩裂，肠子都流出来。
ACTS|1|19|住在 耶路撒冷 的人都知道这事，所以按着他们当地的话把那块田叫 亚革大马 ，就是“血田”的意思。
ACTS|1|20|因为《诗篇》上写着： “愿他的住处变为废墟， 无人在内居住。” 又说： “愿别人得他的职分。”
ACTS|1|21|所以，主耶稣在我们中间出入的整段时间，就是从 约翰 施洗起，直到主离开我们被接上升的日子为止，必须从那常与我们一起的人中，立一位与我们同作耶稣复活的见证。”
ACTS|1|22|
ACTS|1|23|于是他们推举两个人，就是那叫 巴撒巴 ，又称为 犹士都 的 约瑟 ，和 马提亚 。
ACTS|1|24|众人祷告说：“主啊，你知道万人的心，求你从这两个人中指明你所拣选的是哪一位，
ACTS|1|25|去得这使徒的职任；这职位 犹大 已经丢弃，往自己的地方去了。”
ACTS|1|26|于是众人为他们摇签，摇出 马提亚 来；他就和十一个使徒同列。
ACTS|2|1|五旬节那日到了，他们全都聚集在一起。
ACTS|2|2|忽然，有响声从天上下来，好像一阵大风吹过，充满了他们所坐的整座屋子；
ACTS|2|3|又有舌头如火焰向他们显现，分开落在他们每个人身上。
ACTS|2|4|他们都被圣灵充满，就按着圣灵所赐的口才说起别国的话来。
ACTS|2|5|那时，有从天下各国来的虔诚的 犹太 人，住在 耶路撒冷 。
ACTS|2|6|这声音一响，许多人都来聚集，各人因为听见门徒用他们各自的乡谈说话，就甚纳闷，
ACTS|2|7|都诧异惊奇说：“看哪，这些说话的不都是 加利利 人吗？
ACTS|2|8|我们每个人怎么听见他们说我们生来所用的乡谈呢？
ACTS|2|9|我们 帕提亚 人、 玛代 人、 以拦 人，和住在 美索不达米亚 、 犹太 、 加帕多家 、 本都 、 亚细亚 、
ACTS|2|10|弗吕家 、 旁非利亚 、 埃及 的人，并靠近 古利奈 的 利比亚 一带地方的人，侨居的 罗马 人，
ACTS|2|11|包括 犹太 人和皈依 犹太 教的人， 克里特 人和 阿拉伯 人，都听见他们用我们的乡谈讲论上帝的大作为。”
ACTS|2|12|众人就都惊奇困惑，彼此说：“这是什么意思呢？”
ACTS|2|13|还有人讥诮，说：“他们是灌满了新酒吧！”
ACTS|2|14|彼得 和十一个使徒站起来，他就高声向众人说：“ 犹太 人和所有住在 耶路撒冷 的人哪，这件事你们要知道，要侧耳听我的话。
ACTS|2|15|这些人并不像你们所想的喝醉了，因为现在才早晨九点钟。
ACTS|2|16|这正是藉着先知 约珥 所说的：
ACTS|2|17|‘上帝说： 在末后的日子， 我要将我的灵浇灌凡血肉之躯的。 你们的儿女要说预言； 你们的少年要见异象； 你们的老人要做异梦。
ACTS|2|18|在那些日子，我要把我的灵浇灌， 甚至给我的仆人和婢女， 他们要说预言。
ACTS|2|19|在天上，我要显出奇事， 在地下，我要显出神迹， 有血，有火，有烟雾。
ACTS|2|20|太阳要变为黑暗， 月亮要变为血， 这都在主大而光荣的日子未到以前。
ACTS|2|21|那时，凡求告主名的都必得救。’
ACTS|2|22|“ 以色列 人哪，你们要听我这些话： 拿撒勒 人耶稣就是上帝以异能、奇事、神迹向你们证明出来的人，这些事是上帝藉着他在你们中间施行，正如你们自己知道的。
ACTS|2|23|他既按着上帝确定的旨意和预知被交与人，你们就藉着不法之人的手把他钉在十字架上，杀了。
ACTS|2|24|上帝却将死的痛苦解除，使他复活了，因为他原不能被死拘禁。
ACTS|2|25|大卫 指着他说： ‘我看见 主常在我眼前， 他在我右边，使我不至于动摇。
ACTS|2|26|所以我心里欢喜，我的舌头快乐， 而且我的肉身要安居在指望中。
ACTS|2|27|因你必不将我的灵魂撇在阴间， 也不让你的圣者见朽坏。
ACTS|2|28|你已将生命的道路指示我， 必使我在你面前充满快乐。’
ACTS|2|29|“诸位弟兄，先祖 大卫 的事，我可以坦然地对你们说：他死了，也埋葬了，而且他的坟墓直到今日还在我们这里。
ACTS|2|30|既然 大卫 是先知，他知道上帝曾向他起誓，要从他的后裔中立一位坐在他的宝座上。
ACTS|2|31|他预先看见了，就讲论基督的复活，说： ‘他不被撇在阴间； 他的肉身也不见朽坏。’
ACTS|2|32|这耶稣，上帝已经使他复活了，我们都是这事的见证人。
ACTS|2|33|他既被高举在上帝的右边，又从父受了所应许的圣灵，就把你们所看见所听见的，浇灌下来。
ACTS|2|34|大卫 并没有升到天上，但他自己说： ‘主对我主说： 你坐在我的右边，
ACTS|2|35|等我使你的仇敌作你的脚凳。’
ACTS|2|36|故此， 以色列 全家当确实知道，你们钉在十字架上的这位耶稣，上帝已经立他为主，为基督了。”
ACTS|2|37|众人听见这话，觉得扎心，就对 彼得 和其余的使徒说：“诸位弟兄，我们该怎样做呢？”
ACTS|2|38|彼得 对他们说：“你们各人要悔改，奉耶稣基督的名受洗，使你们的罪得赦免，就会领受所赐的圣灵。
ACTS|2|39|因为这应许是给你们和你们的儿女，并一切在远方的人，就是给所有主—我们的上帝所召来的人。”
ACTS|2|40|彼得 还用更多别的话作见证，劝勉他们说：“你们当救自己脱离这弯曲的世代。”
ACTS|2|41|于是领受他话的人，都受了洗；那一天，门徒约添了三千人。
ACTS|2|42|他们都专注于使徒的教导和彼此的团契，擘饼和祈祷。
ACTS|2|43|众人都心存敬畏；使徒们 又行了许多奇事神迹。
ACTS|2|44|信的人都聚在一处，凡物公用，
ACTS|2|45|又卖了田产和家业，照每一个人所需要的分给他们。
ACTS|2|46|他们天天同心合意恒切地在圣殿里敬拜，且在家中 擘饼，存着欢喜坦诚的心用饭，
ACTS|2|47|赞美上帝，得全体百姓的喜爱。主将得救的人天天加给他们。
ACTS|3|1|下午三点钟祷告的时候， 彼得 和 约翰 上圣殿去。
ACTS|3|2|一个从母腹里就是瘸腿的人正被人抬来，他们天天把他放在圣殿的一个叫 美门 的门口，求进圣殿的人施舍。
ACTS|3|3|他看见 彼得 、 约翰 将要进圣殿，就求他们施舍。
ACTS|3|4|彼得 和 约翰 定睛看他， 彼得 说：“看着我们！”
ACTS|3|5|那人就注目看他们，指望从他们得着什么。
ACTS|3|6|彼得 却说：“金银我都没有，但我把我有的给你：奉 拿撒勒 人耶稣基督的名起来 行走！”
ACTS|3|7|于是 彼得 拉着他的右手，扶他起来；他的脚和踝骨立刻健壮了，
ACTS|3|8|就跳起来，站着，又开始行走。他跟他们进了圣殿，边走边跳，赞美上帝。
ACTS|3|9|百姓都看见他又行走，又赞美上帝，
ACTS|3|10|认得他是那素常坐在圣殿的 美门 口求人施舍的，就因他所遇到的事满心惊讶诧异。
ACTS|3|11|那人正在称为 所罗门 的廊下，拉住 彼得 和 约翰 ，大家都觉得很惊讶，一齐跑到他们那里。
ACTS|3|12|彼得 看见，就对百姓说：“ 以色列 人哪，为什么因这事而惊讶呢？为什么定睛看我们，以为我们凭自己的能力和虔诚使这人行走呢？
ACTS|3|13|亚伯拉罕 的上帝、 以撒 的上帝、 雅各 的上帝，就是我们列祖的上帝，已经荣耀了他的仆人耶稣，这耶稣就是你们交付官府的那位， 彼拉多 决定要释放他时，你们却在 彼拉多 面前弃绝了他。
ACTS|3|14|你们弃绝了那圣洁公义者，反而要求释放一个凶手给你们。
ACTS|3|15|你们杀了那生命的创始者，上帝却叫他从死人中复活；我们都是这事的见证人。
ACTS|3|16|因信他的名，他的名使你们所看见所认识的这人健壮了；正是他所赐的信心使这人在你们众人面前完全好了。
ACTS|3|17|“如今，弟兄们，我知道你们做这事是出于无知，你们的官长也是如此。
ACTS|3|18|但上帝藉着众先知的口预先宣告过基督将要受害的事，就这样应验了。
ACTS|3|19|所以，你们当悔改归正，使你们的罪得以涂去，
ACTS|3|20|这样，那安舒的日子就必从主面前来到；主也必差遣所预定给你们的基督耶稣来临。
ACTS|3|21|他必须留在天上，直到万物复兴的时候，就是上帝自古藉着圣先知的口所说的。
ACTS|3|22|摩西 曾说：‘主—你们 的上帝要从你们弟兄中给你们兴起一位先知像我，凡他向你们所说的一切，你们都要听从。
ACTS|3|23|凡不听从那先知的，必将从民中灭绝。’
ACTS|3|24|从 撒母耳 以来和后继的众先知，凡说预言的，也都曾宣告这些日子。
ACTS|3|25|你们是先知的子孙，也是上帝与你们 祖宗所立之约的子孙，就是对 亚伯拉罕 说：‘地上万族都将因你的后裔得福。’
ACTS|3|26|上帝既兴起他的仆人，就先差他到你们这里来，赐福给你们，使各人回转，离开你们的邪恶。”
ACTS|4|1|彼得 和 约翰 正向百姓说话的时候，祭司们、守殿官和撒都该人来了，
ACTS|4|2|就很烦恼，因为使徒们教导百姓，传扬在耶稣的事上证明有死人复活，
ACTS|4|3|于是下手拿住他们；因为天已经晚了，就把他们押在拘留所到第二天。
ACTS|4|4|但听道的人有许多信了，男人的数目约有五千。
ACTS|4|5|第二天，官长、长老和文士在 耶路撒冷 聚集，
ACTS|4|6|又有 亚那 大祭司、 该亚法 、 约翰 、 亚历山大 ，和大祭司的亲族都在那里。
ACTS|4|7|他们叫使徒站在中间，问他们：“你们凭什么能力，奉谁的名做这事呢？”
ACTS|4|8|那时， 彼得 被圣灵充满，对他们说：“民间的官长和长老啊，
ACTS|4|9|倘若今日我们被查问是因为在残障的人身上所行的善事，就是这人怎么得了痊愈，
ACTS|4|10|那么，你们大家和 以色列 全民都当知道，站在你们面前的这人得痊愈，是因你们所钉在十字架、上帝使他从死人中复活的 拿撒勒 人耶稣基督的名。
ACTS|4|11|这位耶稣是： ‘你们匠人所丢弃的石头， 已成了房角的头块石头。’
ACTS|4|12|除他以外，别无拯救，因为在天下人间，没有赐下别的名，我们可以靠着得救。”
ACTS|4|13|他们见 彼得 、 约翰 的胆量，又看出他们原是没有学问的平民，就很惊讶，认出他们曾是跟耶稣一起的；
ACTS|4|14|又看见那治好了的人和他们一同站着，就无话可驳。
ACTS|4|15|于是他们吩咐他们两人从议会退出，就彼此商议，
ACTS|4|16|说：“我们当怎样办这两个人呢？因为他们诚然行了一件明显的神迹，凡住在 耶路撒冷 的人都知道，我们也不能否认。
ACTS|4|17|但为避免这事越发在民间传扬，我们必须威吓他们，叫他们不可再奉这名对任何人讲论。”
ACTS|4|18|于是他们叫了两人来，禁止他们，再不可奉耶稣的名讲论或教导人。
ACTS|4|19|彼得 和 约翰 回答他们说：“听从你们，不听从上帝，在上帝面前合理不合理，你们自己判断吧！
ACTS|4|20|我们所看见所听见的，我们不能不说。”
ACTS|4|21|官长为百姓的缘故，想不出任何法子惩罚他们，只好威吓一番就把他们释放了；这是因众人为了所行的奇事都归荣耀与上帝。
ACTS|4|22|原来经历这神迹医好的人有四十多岁了。
ACTS|4|23|二人既被释放，就到自己的人那里去，把祭司长和长老所说的话都告诉他们。
ACTS|4|24|他们听见了，就同心合意地高声向上帝说：“主宰啊！你是那创造天、地、海和其中万物的；
ACTS|4|25|你曾藉着圣灵托你仆人—我们祖宗 大卫 的口说： ‘外邦为什么扰动？ 万民为什么谋算虚妄的事？
ACTS|4|26|地上的君王都站稳， 臣宰也聚集一处， 要对抗主，对抗主的受膏者 ’。
ACTS|4|27|希律 和 本丢．彼拉多 ，同外邦人和 以色列 民，果然在这城里聚集，要攻打你所膏的圣仆耶稣，
ACTS|4|28|做了你手和你旨意所预定必成就的事。
ACTS|4|29|主啊，现在求你鉴察，他们的威吓，使你仆人放胆讲你的道，
ACTS|4|30|伸出你的手来，让医治、神迹、奇事藉着你圣仆耶稣的名行出来。”
ACTS|4|31|他们祷告完了，聚会的地方震动；他们都被圣灵充满，放胆传讲上帝的道。
ACTS|4|32|许多信徒都一心一意，没有一人说他的任何东西是自己的，都是大家公用。
ACTS|4|33|使徒以大能见证主耶稣 复活；众人也都蒙了大恩。
ACTS|4|34|他们当中没有一个缺乏的，因为凡有田产房屋的都卖了，把所卖的钱拿来，
ACTS|4|35|放在使徒脚前，照每人所需要的，分给每人。
ACTS|4|36|有一个 利未 人，名叫 约瑟 ，使徒称他为 巴拿巴 （ 巴拿巴 翻出来就是安慰之子），生在 塞浦路斯 。
ACTS|4|37|他有田地，也卖了，把钱拿来，放在使徒脚前。
ACTS|5|1|有一个人，名叫 亚拿尼亚 ，同他的妻子 撒非喇 ，卖了田产，
ACTS|5|2|把钱私自留下一部分，他的妻子也知道，其余的部分拿来放在使徒脚前。
ACTS|5|3|彼得 说：“ 亚拿尼亚 ！为什么撒但充满了你的心，使你欺骗圣灵，把卖田地的钱私自留下一部分呢？
ACTS|5|4|田地还没有卖，不是你自己的吗？既卖了，钱不是你作主吗？你怎么心里会想这样做呢？你不是欺骗人，是欺骗上帝！”
ACTS|5|5|亚拿尼亚 一听见这些话，就仆倒，断了气；所有听见的人都非常惧怕。
ACTS|5|6|有些年轻人起来，把他裹好，抬出去埋葬了。
ACTS|5|7|约过了三小时，他的妻子进来，还不知道所发生的事。
ACTS|5|8|彼得 对她说：“你告诉我，你们卖田地的钱就是这些吗？”她说：“就是这些。”
ACTS|5|9|彼得 对她说：“你们为什么同谋来试探主的灵呢？你看，埋葬你丈夫之人的脚已到门口，他们也要把你抬出去。”
ACTS|5|10|她立刻仆倒在 彼得 脚前，断了气。那些年轻人进来，见她已经死了，就把她抬出去，埋在她丈夫旁边。
ACTS|5|11|全教会和所有听见这些事的人都非常惧怕。
ACTS|5|12|主藉使徒的手在民间行了许多神迹奇事；他们都同心合意地聚集在 所罗门 的廊下。
ACTS|5|13|其余的人没有一个敢接近他们，百姓却尊重他们。
ACTS|5|14|信主的人越发增添，连男带女都很多，
ACTS|5|15|甚至有人将病人抬到街上，放在床上或褥子上，好让 彼得 走过来的时候，或者影子投在一些人身上。
ACTS|5|16|还有许多人带着病人和被污灵缠磨的，从 耶路撒冷 四围的城镇来，他们全都得了医治。
ACTS|5|17|于是，大祭司采取行动，他和他所有一起的人，就是撒都该派的人，满心忌恨，
ACTS|5|18|就下手拿住使徒，把他们押在公共拘留所内。
ACTS|5|19|但在夜间主的使者开了监门，领他们出来，说：
ACTS|5|20|“你们去，站在圣殿里，把这生命的一切话讲给百姓听。”
ACTS|5|21|使徒听了这话，天将亮的时候就进圣殿里去教导人。大祭司和他一起的人来了，叫齐议会的人和 以色列 人的众长老，然后派人到监牢里去把使徒提出来。
ACTS|5|22|但差役到了，不见他们在监里，就回来禀报，
ACTS|5|23|说：“我们看见监牢关得很紧，警卫也站在门外，但打开门来，里面一个人都不见。”
ACTS|5|24|守殿官和祭司长听了这些话，心里困惑，不知这事将来如何。
ACTS|5|25|有一个人来禀报说：“你们押在监里的人，现在站在圣殿里教导百姓。”
ACTS|5|26|于是守殿官和差役去带使徒来，并没有用暴力，因为怕百姓用石头打他们。
ACTS|5|27|他们把使徒带来了，就叫他们站在议会前。大祭司问他们，
ACTS|5|28|说：“我们不是严严地禁止你们，不可奉这名教导人吗？ 看，你们倒把你们的道理充满了 耶路撒冷 ，想要叫这人的血归到我们身上！”
ACTS|5|29|彼得 和众使徒回答：“我们必须顺从上帝，胜于顺从人。
ACTS|5|30|你们挂在木头上杀害的耶稣，我们祖宗的上帝已经使他复活了。
ACTS|5|31|上帝把他高举在自己的右边，使他作元帅，作救主，使 以色列 人得以悔改，并且罪得赦免。
ACTS|5|32|我们是这些事的见证人；上帝赐给顺从的人的圣灵也为这些事作见证。”
ACTS|5|33|议会的人听了极其恼怒，想要杀他们。
ACTS|5|34|但有一个法利赛人，名叫 迦玛列 ，是众百姓所敬重的律法教师，他在议会中站起来，吩咐人把使徒暂且带到外面去，
ACTS|5|35|然后对众人说：“ 以色列 人哪，对于这些人，你们应当小心怎样处理。
ACTS|5|36|从前 杜达 出现，自命不凡，附从他的人数约有四百；他被杀后，附从他的人全都散了，归于无有。
ACTS|5|37|此后，登记户籍的时候，又有 加利利 的 犹大 出现，引诱百姓跟从他，他也灭亡，附从他的人也都四散了。
ACTS|5|38|现在，我劝你们不要管这些人，任凭他们吧！他们所谋所为若是出于人，必要败坏；
ACTS|5|39|若是出于上帝，你们就不能败坏他们，恐怕你们倒是攻击上帝了。” 议会的人被他说服了，
ACTS|5|40|就叫使徒来，把他们打了，又吩咐他们不可奉耶稣的名讲道，然后把他们释放了。
ACTS|5|41|他们欢欢喜喜地离开议会，因他们算配为这名受辱。
ACTS|5|42|他们就每日在圣殿里，在家里 ，不住地教导人，传耶稣是基督的福音。
ACTS|6|1|那些日子，门徒增多，有说希腊话的 犹太 人向 希伯来 人发怨言，因为在日常的供给上忽略了他们的寡妇。
ACTS|6|2|十二使徒叫众门徒来，说：“我们撇下上帝的道去管理饭食，是不合宜的。
ACTS|6|3|所以弟兄们，当从你们中间选出七个有好名声、满有圣灵和智慧，我们派他们管理这事。
ACTS|6|4|至于我们，我们要专注于祈祷和传道的事奉。”
ACTS|6|5|这话使全会众都喜悦，就拣选了 司提反 —他是一个满有信心和圣灵的人；他们又拣选了 腓利 、 伯罗哥罗 、 尼迦挪 、 提门 、 巴米拿 ，并皈依 犹太 教的 安提阿 人 尼哥拉 ，
ACTS|6|6|叫他们站在使徒面前，使徒祷告后，就为他们按手。
ACTS|6|7|上帝的道兴旺起来；在 耶路撒冷 门徒数目增加得很多，也有许多祭司听从了这信仰。
ACTS|6|8|司提反 满有恩惠和能力，在民间行了大奇事和神迹。
ACTS|6|9|当时有从称为“自由人”会堂，并 古利奈 、 亚历山大 会堂来的人，还有些从 基利家 、 亚细亚 来的人，起来和 司提反 辩论。
ACTS|6|10|司提反 是以智慧和圣灵说话，众人抵挡不住，
ACTS|6|11|就收买人来说：“我们听见他说亵渎 摩西 和上帝的话。”
ACTS|6|12|他们又煽动百姓、长老和文士，就突然来捉拿他，把他带到议会去，
ACTS|6|13|设下假见证，说：“这个人不断地说话，侮辱神圣的地方和律法。
ACTS|6|14|我们曾听见他说，这 拿撒勒 人耶稣要毁坏这地方，也要改变 摩西 所交给我们的规矩。”
ACTS|6|15|在议会里坐着的人都定睛看他，见他的面貌好像天使的面貌。
ACTS|7|1|大祭司说：“果真有这些事吗？”
ACTS|7|2|司提反 说：“诸位父老弟兄请听！从前我们的祖宗 亚伯拉罕 在 美索不达米亚 ，还没有住在 哈兰 的时候，荣耀的上帝向他显现，
ACTS|7|3|对他说：‘你要离开本地和亲族，往我所要指示你的地去。’
ACTS|7|4|他就离开 迦勒底 人的地方，住在 哈兰 。他父亲死了以后，上帝使他从那里搬到你们现在所住的地方。
ACTS|7|5|在这里上帝并没有给他产业，连立足的地方都没有，但应许要将这地赐给他和他的后裔为业，虽然那时他还没有儿子。
ACTS|7|6|上帝这样说：‘他的后裔必寄居外邦，那里的人要使他们作奴隶，苦待他们四百年。’
ACTS|7|7|上帝又说：‘但我要惩罚使他们作奴隶的那国。以后他们要出来，在这地方事奉我。’
ACTS|7|8|上帝又赐他割礼的约。于是 亚伯拉罕 生了 以撒 ，在第八日给他行了割礼；后来 以撒 生 雅各 ， 雅各 生十二位先祖。
ACTS|7|9|“先祖嫉妒 约瑟 ，把他卖到 埃及 去，上帝却与他同在，
ACTS|7|10|救他脱离一切苦难，又使他在 埃及 王法老面前蒙恩，又有智慧。法老派他作 埃及 国的宰相兼管法老的全家。
ACTS|7|11|后来全 埃及 和 迦南 遭遇饥荒和大灾难，我们的祖宗绝了粮。
ACTS|7|12|雅各 听见在 埃及 有粮，就打发我们的祖宗初次往那里去。
ACTS|7|13|第二次 约瑟 与兄弟们相认，法老才认识他的家族。
ACTS|7|14|约瑟 就打发人，请父亲 雅各 和全族七十五个人都来。
ACTS|7|15|于是 雅各 下了 埃及 ，后来他和我们的祖宗都死在那里；
ACTS|7|16|他们又被迁到 示剑 ，葬于 亚伯拉罕 在 示剑 用银子从 哈抹 子孙 买来的坟墓里。
ACTS|7|17|“当上帝应许 亚伯拉罕 的日期将到的时候， 以色列 人在 埃及 人丁兴旺，
ACTS|7|18|直到另一位不认识 约瑟 的王兴起统治 埃及 。
ACTS|7|19|他用诡计待我们的宗族，苦待我们的祖宗，强迫他们丢弃婴孩，使婴孩不能存活。
ACTS|7|20|就在那时， 摩西 生了下来，上帝看为俊美，在父亲家里被抚养了三个月。
ACTS|7|21|他被丢弃的时候，法老的女儿拾了去，当自己的儿子抚养。
ACTS|7|22|摩西 学了 埃及 人一切的学问，说话办事都有才能。
ACTS|7|23|“他到了四十岁，心中起意去看望他的弟兄 以色列 人。
ACTS|7|24|他见他们中的一个人受冤屈，就庇护他，为那被压迫的人报仇，打死了那 埃及 人。
ACTS|7|25|他以为他的弟兄们必明白上帝是藉他的手搭救他们，他们却不明白。
ACTS|7|26|第二天，他遇见有人在打架，就想劝他们和好，说：‘二位，你们是弟兄，为什么彼此欺负呢？’
ACTS|7|27|那欺负邻舍的人把他推开，说：‘谁立你作我们的领袖和审判官呢？
ACTS|7|28|难道你要杀我像昨天杀那 埃及 人一样吗？’
ACTS|7|29|摩西 听见这话就逃走了，寄居于 米甸 地，在那里生了两个儿子。
ACTS|7|30|“过了四十年，在 西奈山 的旷野，有一位天使在荆棘的火焰中向 摩西 显现。
ACTS|7|31|摩西 见了那异象，觉得很惊讶，正往前观看的时候，有主的声音说：
ACTS|7|32|‘我是你列祖的上帝，就是 亚伯拉罕 、 以撒 、 雅各 的上帝。’ 摩西 战战兢兢，不敢观看。
ACTS|7|33|主对他说：‘把你脚上的鞋脱下来，因为你所站的地方是圣地。
ACTS|7|34|我的百姓在 埃及 所受的困苦，我确实看见了；他们悲叹的声音，我也听见了。我下来要救他们。现在，你来，我要差你往 埃及 去。’
ACTS|7|35|“这 摩西 就是有人曾弃绝他说‘谁立你作我们的领袖和审判官’的，上帝却藉那在荆棘中显现的天使的手差派他作领袖，作解救者。
ACTS|7|36|这人领 以色列 人出来，在 埃及 地，在 红海 ，在旷野的四十年间行了奇事神迹。
ACTS|7|37|这人是 摩西 ，就是那曾对 以色列 人说‘上帝要从你们弟兄中给你们兴起一位先知像我’的。
ACTS|7|38|这人是那曾在旷野的会众中和 西奈山 上，与那对他说话的天使同在，又与我们祖宗同在的，他领受了活泼的圣言传给我们。
ACTS|7|39|我们的祖宗不肯听从，反弃绝他，他们的心转向 埃及 ，
ACTS|7|40|对 亚伦 说：‘你为我们造神明，在我们前面引路，因为领我们出 埃及 地的这个 摩西 ，我们不知道他遭遇了什么事。’
ACTS|7|41|那时，他们造了一个牛犊，又拿祭物献给那像，为自己手所做的工作欢跃。
ACTS|7|42|但是上帝转脸不顾，任凭他们祭拜天上的日月星辰，正如先知书上所写的： ‘ 以色列 家啊，你们四十年间在旷野， 何曾将牺牲和祭物献给我？
ACTS|7|43|你们抬着 摩洛 的帐幕 和 理番 ──你们神明的星， 就是你们所造为要敬拜的像。 因此，我要把你们迁到 巴比伦 外去。’
ACTS|7|44|“我们的祖宗在旷野，有作证的会幕，是上帝吩咐 摩西 照着他所看见的样式做的。
ACTS|7|45|这帐幕，我们的祖宗同 约书亚 相继承受了，当上帝在他们面前赶走外邦人的时候，他们把这帐幕搬进承受为业之地，直存到 大卫 的日子。
ACTS|7|46|大卫 在上帝面前蒙恩，祈求为 雅各 的家 预备居所。
ACTS|7|47|但却是 所罗门 为上帝造成殿宇。
ACTS|7|48|其实，至高者并不住人手所造的，就如先知所言：
ACTS|7|49|‘主说：天是我的宝座， 地是我的脚凳。 你们要为我造怎样的殿宇？ 哪里是我安歇的地方呢？
ACTS|7|50|这一切不都是我手所造的吗？’
ACTS|7|51|“你们这硬着颈项，心与耳未受割礼的人哪，时常抗拒圣灵！你们的祖宗怎样，你们也怎样。
ACTS|7|52|先知中有哪一个不是受你们祖宗的迫害呢？他们把预先宣告那义者要来的人杀了。如今你们成了那义者的出卖者和凶手了。
ACTS|7|53|你们领受了天使所传布的律法，竟不遵守。”
ACTS|7|54|众人听见这些话，心中极其恼怒，向 司提反 咬牙切齿。
ACTS|7|55|但 司提反 满有圣灵，定睛望天，看见上帝的荣耀，又看见耶稣站在上帝的右边，
ACTS|7|56|就说：“我看见天开了，人子站在上帝的右边。”
ACTS|7|57|众人大声喊叫，捂着耳朵，齐心冲向他，
ACTS|7|58|把他推到城外，用石头打他。作见证的人把他们的衣裳放在一个名叫 扫罗 的青年脚前。
ACTS|7|59|他们正用石头打 司提反 的时候，他呼求说：“主耶稣啊，求你接纳我的灵魂！”
ACTS|7|60|然后他跪下来，大声喊着：“主啊，不要将这罪归于他们！”说了这话，就长眠了。
ACTS|8|1|扫罗 也赞同处死他。从那一天开始， 耶路撒冷 的教会遭受到大迫害，除了使徒以外，众门徒都分散在 犹太 和 撒玛利亚 各处。
ACTS|8|2|有些虔诚的人把 司提反 埋葬了，为他大大哀哭。
ACTS|8|3|扫罗 却残害教会，挨家挨户地进去，拉着男女关在监里。
ACTS|8|4|那些分散的人往各地去传福音的道。
ACTS|8|5|腓利 下 撒玛利亚城 去 ，向当地人宣讲基督。
ACTS|8|6|众人都聚精会神，同心合意地听 腓利 所说的话，一边听他的话，一边看他所行的神迹。
ACTS|8|7|因为有许多人被污灵附着，那些污灵大声呼叫，从他们身上出来；还有许多瘫痪的、瘸腿的都得了医治。
ACTS|8|8|那城里，有极大的喜乐。
ACTS|8|9|有一个人名叫 西门 ，向来在那城里行邪术，自命为大人物，使 撒玛利亚 的居民惊奇。
ACTS|8|10|所有的人，从小到大都听从他，说：“这个人就是上帝的能力，那称为大能者的。”
ACTS|8|11|他们听从他，因他很久以来用邪术使他们惊奇。
ACTS|8|12|当他们信了 腓利 所传上帝国的福音和耶稣基督的名，连男带女都受了洗。
ACTS|8|13|西门 自己也信了；既受了洗，就常与 腓利 在一处，看见他所行的神迹和大异能，就觉得很惊奇。
ACTS|8|14|在 耶路撒冷 的使徒听见 撒玛利亚 人领受了上帝的道，就打发 彼得 和 约翰 到他们那里去。
ACTS|8|15|两个人下去，就为他们祷告，要让他们领受圣灵，
ACTS|8|16|因为圣灵还没有降在他们任何一个人身上，他们只奉主耶稣的名受了洗。
ACTS|8|17|于是使徒按手在他们头上，他们就领受了圣灵。
ACTS|8|18|西门 看见使徒一按手，就有圣灵赐下，就拿钱给使徒，
ACTS|8|19|说：“请把这权柄也给我，使我手按着谁，谁就可以领受圣灵。”
ACTS|8|20|彼得 对他说：“你的银子和你一同灭亡吧！因为你想上帝的恩赐是可以用钱买的。
ACTS|8|21|你在这道上无份无关；因为你在上帝面前心怀不正。
ACTS|8|22|你要为你这样的恶而悔改，祈求主，或者你心里的意念可得赦免。
ACTS|8|23|我看出你正在苦胆之中，被不义捆绑着。”
ACTS|8|24|西门 回答说：“请你们为我求主，使你们所说的，没有一样临到我身上。”
ACTS|8|25|使徒既作了见证，并且宣讲了主的道，就回 耶路撒冷 去，一路在 撒玛利亚 好些村庄传扬福音。
ACTS|8|26|有主的一个使者对 腓利 说：“起来！向南走，往那从 耶路撒冷 下 迦萨 的路上去。”那路是旷野。
ACTS|8|27|腓利 就起身去了。不料，有一个 埃塞俄比亚 人，是个有大权的太监，在 埃塞俄比亚 女王 甘大基 的手下总管银库，他上 耶路撒冷 去礼拜。
ACTS|8|28|回程中，他坐在车上，正念着 以赛亚 先知的书，
ACTS|8|29|圣灵对 腓利 说：“你去！靠近那车走。”
ACTS|8|30|腓利 就跑到太监那里，听见他正在念 以赛亚 先知的书，就说：“你明白你所念的吗？”
ACTS|8|31|他说：“没有人指教我，怎能明白呢？”于是他请 腓利 上车，与他同坐。
ACTS|8|32|他所念的那段经文是这样： “他像羊被牵去宰杀， 又像羔羊在剪毛的人手下无声， 他也是这样不开口。
ACTS|8|33|他卑微的时候，得不到公义的审判， 谁能述说他的身世？ 因为他的生命从地上被夺去。”
ACTS|8|34|太监回答 腓利 说：“请问，先知说这话是指谁，是指自己，还是指别人呢？”
ACTS|8|35|腓利 就开口，从这段经文开始，对他传讲耶稣的福音。
ACTS|8|36|二人正沿路往前走，到了有水的地方，太监说：“看哪！这里有水，有什么能阻止我受洗呢？”
ACTS|8|37|
ACTS|8|38|于是他吩咐把车停下来， 腓利 和太监二人一同下到水里， 腓利 就给他施洗。
ACTS|8|39|他们从水里上来，主的灵把 腓利 提了去，太监再也看不见他了，就欢欢喜喜地上路。
ACTS|8|40|后来有人在 亚锁都 遇见 腓利 ；他走遍那地方，在各城宣扬福音，一直到 凯撒利亚 。
ACTS|9|1|扫罗 不断用威吓凶悍的口气向主的门徒说话。他去见大祭司，
ACTS|9|2|要求发信给 大马士革 的各会堂，若是找着信奉这道的人，无论男女，都准他捆绑带到 耶路撒冷 。
ACTS|9|3|扫罗 在途中，将到 大马士革 的时候，忽然有一道光从天上下来，四面照射着他，
ACTS|9|4|他就仆倒在地，听见有声音对他说：“ 扫罗 ！ 扫罗 ！你为什么迫害我？”
ACTS|9|5|他说：“主啊！你是谁？”主说：“我就是你所迫害的耶稣。
ACTS|9|6|起来！进城去，你应该做的事，必有人告诉你。”
ACTS|9|7|同行的人站在那里，说不出话来，因为他们听见声音，却看不见人。
ACTS|9|8|扫罗 从地上起来，睁开眼睛，竟不能看见什么。有人拉他的手，领他进了 大马士革 。
ACTS|9|9|他三天什么都看不见，也不吃也不喝。
ACTS|9|10|那时，在 大马士革 有一个门徒，名叫 亚拿尼亚 。主在异象中对他说：“ 亚拿尼亚 ！”他说：“主啊，我在这里。”
ACTS|9|11|主对他说：“起来！往那叫 直街 的路去，在 犹大 的家里，去找一个 大数 人，名叫 扫罗 ；他正在祷告，
ACTS|9|12|在异象中 看见了一个人，名叫 亚拿尼亚 ，进来为他按手，让他能再看得见。”
ACTS|9|13|亚拿尼亚 回答：“主啊，我听见许多人讲到这个人，说他怎样在 耶路撒冷 多多苦待你的圣徒，
ACTS|9|14|并且他在这里有从祭司长得来的权柄，要捆绑一切求告你名的人。”
ACTS|9|15|主对他说：“你只管去。他是我所拣选的器皿，要在外邦人、君王和 以色列 人面前宣扬我的名。
ACTS|9|16|我也要指示他，为我的名必须受许多的苦难。”
ACTS|9|17|亚拿尼亚 就去了，进入那家，把手按在 扫罗 身上，说：“ 扫罗 弟兄，在你来的路上向你显现的主，就是耶稣，打发我来，叫你能再看得见，又被圣灵充满。”
ACTS|9|18|扫罗 的眼睛上立刻好像有鳞一般的东西掉下来，他就能再看得见，于是他起来，受了洗，
ACTS|9|19|吃过饭体力就恢复了。 扫罗 和 大马士革 的门徒一起住了些日子，
ACTS|9|20|立刻在各会堂里传扬耶稣，说他是上帝的儿子。
ACTS|9|21|凡听见的人都很惊奇，说：“在 耶路撒冷 残害求告这名的不就是这个人吗？他不是到这里来要捆绑他们，带到祭司长那里去吗？”
ACTS|9|22|但 扫罗 越发有能力，驳倒住在 大马士革 的 犹太 人，证明耶稣是基督。
ACTS|9|23|过了好些日子， 犹太 人商议要杀 扫罗 ，
ACTS|9|24|但他们的计谋被 扫罗 知道了。他们昼夜在城门守候着要杀他。
ACTS|9|25|他的门徒就在夜间用筐子把他从城墙上缒了下去。
ACTS|9|26|扫罗 到了 耶路撒冷 ，想与门徒结交，大家却都怕他，不信他是门徒。
ACTS|9|27|只有 巴拿巴 接待他，领他去见使徒，把他在路上怎么看见主，主怎么向他说话，他在 大马士革 怎么奉耶稣的名放胆传道，都述说出来。
ACTS|9|28|于是 扫罗 在 耶路撒冷 同门徒出入来往，奉主的名放胆传道，
ACTS|9|29|并和说 希腊 话的 犹太 人讲论辩驳，他们却想法子要杀他。
ACTS|9|30|弟兄们知道了，就带他下 凯撒利亚 ，送他往 大数 去。
ACTS|9|31|那时， 犹太 、 加利利 、 撒玛利亚 各处的教会都得平安，建立起来，凡事敬畏主，蒙圣灵的安慰，人数逐渐增多。
ACTS|9|32|彼得 在众信徒中到处奔波的时候，也到了住在 吕大 的圣徒那里。
ACTS|9|33|他在那里遇见一个人，名叫 以尼雅 ，得了瘫痪，在褥子上躺了八年。
ACTS|9|34|彼得 对他说：“ 以尼雅 ，耶稣基督医好你了，起来！整理你的褥子吧。”他立刻就起来了。
ACTS|9|35|凡住 吕大 和 沙仑 的人都看见了他，就归向主。
ACTS|9|36|在 约帕 有一个女门徒，名叫 大比大 ，翻出来的意思是 多加 ；她广行善事，多施周济。
ACTS|9|37|当时，她患病死了，有人把她清洗后，停在楼上。
ACTS|9|38|吕大 原与 约帕 相近；门徒听见 彼得 在那里，就派两个人去见他，央求他说：“请快到我们那里去，不要耽延。”
ACTS|9|39|彼得 就起身和他们同去。他到了，就有人领他上楼。众寡妇都站在 彼得 旁边哭，拿 多加 与她们同在时所做的内衣外衣给他看。
ACTS|9|40|彼得 叫她们都出去，然后跪下祷告，转身对着尸体说：“ 大比大 ，起来！”她就睁开眼睛，看见 彼得 ，就坐了起来。
ACTS|9|41|彼得 伸手扶她起来，叫那些圣徒和寡妇都进来，把 多加 活活地交给他们。
ACTS|9|42|这事传遍了 约帕 ，就有许多人信了主。
ACTS|9|43|此后， 彼得 在 约帕 一个皮革匠 西门 的家里住了好些日子。
ACTS|10|1|在 凯撒利亚 有一个人名叫 哥尼流 ，是 意大利 营的百夫长。
ACTS|10|2|他是个虔诚人，他和全家都敬畏上帝。他多多周济百姓，常常向上帝祷告。
ACTS|10|3|有一天，约在下午三点钟，他在异象中清楚看见上帝的一个使者进来，到他那里，对他说：“ 哥尼流 。”
ACTS|10|4|哥尼流 定睛看他，惊惶地说：“主啊，什么事？”天使对他说：“你的祷告和你的周济已达到上帝面前，蒙记念了。
ACTS|10|5|现在你要派人往 约帕 去，请一位称为 彼得 的 西门 来。
ACTS|10|6|他住在一个皮革匠 西门 的家里，房子就在海边。”
ACTS|10|7|向他说话的天使离开后， 哥尼流 叫了两个仆人和常伺候他的一个虔诚的兵来，
ACTS|10|8|把一切的事都讲给他们听，然后就派他们往 约帕 去。
ACTS|10|9|第二天，他们走路将近那城，约在正午， 彼得 上房顶去祷告。
ACTS|10|10|他觉得饿了，想要吃。那家的人正预备饭的时候， 彼得 魂游象外，
ACTS|10|11|看见天开了，有一块好像大布的东西降下，四角 吊着缒在地上，
ACTS|10|12|里面有地上各样四脚的走兽、爬虫和天上的飞鸟。
ACTS|10|13|又有声音对他说：“ 彼得 ，起来！宰了吃。”
ACTS|10|14|彼得 却说：“主啊，绝对不可！凡污俗和不洁净的东西，我从来没有吃过。”
ACTS|10|15|第二次有声音再对他说：“上帝所洁净的，你不可当作污俗的。”
ACTS|10|16|这样一连三次，那东西随即收回天上去了。
ACTS|10|17|正当 彼得 心里困惑，不知所看见的异象是什么意思时， 哥尼流 所差来的人已经找到了 西门 的家，站在门外，
ACTS|10|18|喊着问有没有一位称为 彼得 的 西门 住在这里。
ACTS|10|19|彼得 还在思考那异象的时候，圣灵对他说：“有三个人来找你。
ACTS|10|20|起来，下去，跟他们同去，不要疑惑，因为是我差他们来的。”
ACTS|10|21|于是 彼得 下去见那些人，说：“我就是你们要找的人，你们是为了什么缘故在这里？”
ACTS|10|22|他们说：“百夫长 哥尼流 是个义人，敬畏上帝，为 犹太 全民族所称赞。他蒙一位圣天使指示，叫他请你到他家里去，要听你讲话。”
ACTS|10|23|彼得 就请他们进去住宿。 次日，他起身和他们同去，还有 约帕 的几个弟兄跟他一起去。
ACTS|10|24|又次日，他 进入 凯撒利亚 ， 哥尼流 已经请了他的亲朋好友在等候他们。
ACTS|10|25|彼得 一进去， 哥尼流 就迎接他，俯伏在他脚前拜他。
ACTS|10|26|但是 彼得 拉他起来，说：“你起来，我自己也不过是人。”
ACTS|10|27|彼得 和他一边说话一边进去，见有好些人聚集，
ACTS|10|28|就对他们说：“你们知道， 犹太 人和别国的人结交来往本是不合规矩的，但上帝已经指示我，无论什么人都不可看作污俗或不洁净的。
ACTS|10|29|所以，我一被邀请，没有推辞就来了。现在请问，你们为什么叫我来呢？”
ACTS|10|30|哥尼流 说：“四天前，这个时候，我在家中守着下午三点钟的祷告，忽然有一个人穿着明亮的衣裳站在我面前，
ACTS|10|31|说：‘ 哥尼流 ，你的祷告已蒙垂听，你的周济在上帝面前已蒙记念了。
ACTS|10|32|你要派人往 约帕 去，请那称为 彼得 的 西门 来，他住在海边一个皮革匠 西门 的家里。’
ACTS|10|33|所以我立刻派人去请你。你来了真好。现在我们都在上帝面前，要听主 吩咐你的一切话。”
ACTS|10|34|彼得 开口说：“我真的看出上帝是不偏待人的。
ACTS|10|35|不但如此，在各国中那敬畏他而行义的人都为他所悦纳。
ACTS|10|36|上帝藉着耶稣基督—他是万有的主—传和平的福音，把这道传给 以色列 人。
ACTS|10|37|这话在 约翰 传扬洗礼以后，从 加利利 起，传遍了 犹太 。上帝怎样以圣灵和能力膏了 拿撒勒 人耶稣，这都是你们知道的。他到处奔波，行善事，医好凡被魔鬼压制的人，因为上帝与他同在。
ACTS|10|38|
ACTS|10|39|他在 犹太 人之地和 耶路撒冷 所行的一切事，有我们作见证人。他们竟把他挂在木头上杀了。
ACTS|10|40|第三天，上帝使他复活，使他显现出来；
ACTS|10|41|不是显现给所有的人看，而是显现给上帝预先所拣选为他作见证的人看，就是我们这些在他从死人中复活以后和他同吃同喝的人。
ACTS|10|42|他吩咐我们传道给众人，证明他是上帝所立定，要作审判活人、死人的审判者。
ACTS|10|43|众先知也为这人作见证：凡信他的人，必藉着他的名得蒙赦罪。”
ACTS|10|44|彼得 还在说这些话的时候，圣灵降在一切听道的人身上。
ACTS|10|45|那些奉割礼的信徒和 彼得 同来，见圣灵的恩赐也浇在外邦人身上，就都惊奇；
ACTS|10|46|因听见他们说方言 ，称赞上帝为大。于是 彼得 回答：
ACTS|10|47|“这些人既受了圣灵，跟我们一样，谁能阻止用水给他们施洗呢？”
ACTS|10|48|他就吩咐奉耶稣基督的名给他们施洗。于是他们请 彼得 住了几天。
ACTS|11|1|使徒和在 犹太 的众弟兄听到外邦人也领受了上帝的道。
ACTS|11|2|等到 彼得 上了 耶路撒冷 ，那些奉割礼的信徒和他争辩，
ACTS|11|3|说：“你竟进入未受割礼之人当中，和他们一同吃饭！”
ACTS|11|4|彼得 就开始把这事逐一向他们解释，说：
ACTS|11|5|“我在 约帕城 里祷告的时候，魂游象外，看见异象，有一块好像大布的东西降下，四角吊着从天缒下，直来到我跟前。
ACTS|11|6|我定睛观看，见内中有地上四脚的牲畜、野兽、爬虫和天上的飞鸟。
ACTS|11|7|我还听见有声音对我说：‘ 彼得 ，起来！宰了吃。’
ACTS|11|8|我说：‘主啊，绝对不可！凡污俗或不洁净的东西从来没有进过我的口。’
ACTS|11|9|第二次，有声音从天上回答：‘上帝所洁净的，你不可当作污俗的。’
ACTS|11|10|这样一连三次，然后一切就都收回天上去了。
ACTS|11|11|正当那时，有三个从 凯撒利亚 差来见我的人，站在我们 所住的屋子门前。
ACTS|11|12|圣灵吩咐我和他们同去，不要疑惑，还有这六位弟兄也跟我一起去，我们进了那人的家。
ACTS|11|13|那人就告诉我们，他如何看见一位天使站在他家里，说：‘你派人往 约帕 去，请那称为 彼得 的 西门 来，
ACTS|11|14|他有话要告诉你，因这些话你和你的全家都可以得救。’
ACTS|11|15|我一开始讲话，圣灵就降在他们身上，正像当初降在我们身上一样。
ACTS|11|16|我就想起主的话如何说：‘ 约翰 用水施洗，但你们要在圣灵里受洗。’
ACTS|11|17|既然上帝给他们恩赐，像在我们信主耶稣基督的时候给了我们一样，我是谁，能拦阻上帝吗？”
ACTS|11|18|众人听见这些话，就不说话了，只归荣耀给上帝，说：“这样看来，上帝也赐恩给外邦人，使他们悔改得生命了。”
ACTS|11|19|那些因 司提反 的事遭患难而四处分散的门徒，直走到 腓尼基 、 塞浦路斯 和 安提阿 。他们不向别人讲道，只向 犹太 人讲。
ACTS|11|20|但内中有 塞浦路斯 和 古利奈 人，他们到了 安提阿 也向 希腊 人传讲主耶稣的福音 。
ACTS|11|21|主的手与他们同在，信而归主的人数很多。
ACTS|11|22|这风声传到 耶路撒冷 教会的人耳中，他们就打发 巴拿巴 到 安提阿 去。
ACTS|11|23|他到了那里，看见上帝所赐的恩就欢喜，劝勉众人要立定心志，恒久靠主。
ACTS|11|24|这 巴拿巴 原是个好人，满有圣灵和信心，于是有许多人归服了主。
ACTS|11|25|他又往 大数 去找 扫罗 ，
ACTS|11|26|找着了，就带他到 安提阿 去。他们足有一年和教会一同聚集，教导了许多人。门徒称为“基督徒”是从 安提阿 开始的。
ACTS|11|27|当那些日子，有几位先知从 耶路撒冷 下到 安提阿 。
ACTS|11|28|内中有一位，名叫 亚迦布 ，站起来，藉着圣灵指示普天下将有大饥荒；这事在 克劳第 年间果然实现了。
ACTS|11|29|于是门徒决定，照各人的力量捐钱，送去供给住在 犹太 的弟兄。
ACTS|11|30|他们就这样做了，托 巴拿巴 和 扫罗 的手送到众长老那里。
ACTS|12|1|约在那时候， 希律 王下手苦待教会中的一些人，
ACTS|12|2|用刀杀了 约翰 的哥哥 雅各 。
ACTS|12|3|他见 犹太 人喜欢这事，也去拿住 彼得 。那时候正是除酵节期间。
ACTS|12|4|希律 捉了 彼得 ，押在监里，交给四班士兵看守，每班四个人，企图要在逾越节后把他提出来，当着百姓办他。
ACTS|12|5|于是 彼得 被囚在监里，教会却为他切切祷告上帝。
ACTS|12|6|希律 将要提他出来的前一夜， 彼得 被两条铁链锁着，睡在两个士兵当中；门前还有警卫看守。
ACTS|12|7|忽然，有主的一个使者显现，牢房里有光照耀；天使拍 彼得 的肋旁，叫醒了他，说：“快起来！”铁链就从他手上脱落下来。
ACTS|12|8|天使对他说：“束上腰带，穿上鞋子。”他就照着做了。天使又对他说：“披上外衣，跟我来。”
ACTS|12|9|彼得 就出来跟着他走，不知道天使所做是真的，以为见了异象。
ACTS|12|10|他们经过了第一层和第二层监牢，就来到往城内的铁门，那门就自动给他们开了。他们出来，走过一条街，忽然天使离开他去了。
ACTS|12|11|彼得 清醒过来，说：“现在我真知道主差遣他的使者，救我脱离 希律 的手，和 犹太 人所期待的一切。”
ACTS|12|12|他明白了，就到那称为 马可 的 约翰 的母亲 马利亚 家去，在那里已有好些人聚集祷告。
ACTS|12|13|彼得 敲外门时，有一个使女，名叫 罗大 ，出来应门，
ACTS|12|14|认出是 彼得 的声音，欢喜得顾不了开门，就跑进去报信，说 彼得 站在门外。
ACTS|12|15|他们对她说：“你疯了！”使女坚持真有其事。他们说：“那是他的天使。”
ACTS|12|16|彼得 不停地敲门；他们开了门，一见是他，就很惊奇。
ACTS|12|17|彼得 做个手势，要他们不作声，就告诉他们主怎样领他出监；又说：“你们要把这些事告诉 雅各 和众弟兄。”然后，他离开往别处去了。
ACTS|12|18|到了天亮，士兵中起了不少骚动，不知道 彼得 到哪里去了。
ACTS|12|19|希律 找他，找不着，就审问警卫，下令带走他们处死。后来 希律 离开 犹太 ，下 凯撒利亚 去，住在那里。
ACTS|12|20|希律 向 推罗 和 西顿 的人发怒。他们那一带地方是从王的土地供应粮食的，因此就托了王的内侍大臣 伯拉斯都 的情，一心来求和。
ACTS|12|21|希律 在所定的日子，穿上朝服，坐在位上，对他们演讲。
ACTS|12|22|民众一直喊着：“这是神明的声音，不是人的声音。”
ACTS|12|23|希律 不归荣耀给上帝，所以主的使者立刻击打他，他被虫咬，就断了气。
ACTS|12|24|上帝的道日见兴旺，越发广传。
ACTS|12|25|巴拿巴 和 扫罗 完成了供给的事，就回到 耶路撒冷 ，带著称为 马可 的 约翰 同去。
ACTS|13|1|在 安提阿 的教会中，有几位先知和教师，就是 巴拿巴 和称为 尼结 的 西面 、 古利奈 人 路求 ，与 希律 分封王一起长大的 马念 ，和 扫罗 。
ACTS|13|2|他们在事奉主和禁食的时候，圣灵说：“要为我分派 巴拿巴 和 扫罗 去做我召他们做的工作。”
ACTS|13|3|于是他们禁食祷告后，给 巴拿巴 和 扫罗 按手，然后派遣他们走了。
ACTS|13|4|他们既蒙圣灵差遣，就下到 西流基 ，从那里坐船往 塞浦路斯 去，
ACTS|13|5|到了 撒拉米 ，就在 犹太 人各会堂里宣讲上帝的道，也有 约翰 作他们的帮手。
ACTS|13|6|他们走遍全岛，直到 帕弗 ，在那里遇见一个术士— 犹太 人的假先知，名叫 巴耶稣 。
ACTS|13|7|这人常和 士求．保罗 省长在一起。 士求．保罗 是个通达人，他请 巴拿巴 和 扫罗 来，要听上帝的道。
ACTS|13|8|只是术士 以吕马 (他的名字翻出来就是行法术的意思)敌对使徒，设法使省长远离这信仰。
ACTS|13|9|扫罗 ，又名 保罗 ，被圣灵充满，定睛看他，
ACTS|13|10|说：“你这充满各样诡诈奸恶，魔鬼的儿子，一切正义的仇敌，你还不停止扭曲主的正道吗？
ACTS|13|11|现在你看，主的手临到你身上，你会瞎眼，暂时看不见日光。”立刻迷濛和黑暗笼罩着他，他到处摸索，求人拉着手领他。
ACTS|13|12|省长看见所发生的事就信了，因对主的教导感到惊奇。
ACTS|13|13|保罗 和他的同伴从 帕弗 开船，来到 旁非利亚 的 别加 ， 约翰 却离开他们，回 耶路撒冷 去了。
ACTS|13|14|他们从 别加 往前行，来到 彼西底 的 安提阿 。在安息日，他们进了会堂就坐下。
ACTS|13|15|在读完了律法和先知的书，会堂主管们叫人过去，对他们说：“二位弟兄，你们若有什么劝勉众人的话，请说。”
ACTS|13|16|保罗 就站起来，做个手势，说：“诸位 以色列 人和一切敬畏上帝的人，请听。
ACTS|13|17|这 以色列 民的上帝拣选了我们的祖宗，当百姓寄居 埃及 的时候抬举他们，用大能的手领他们从那地出来。
ACTS|13|18|他在旷野容忍 他们，约有四十年。
ACTS|13|19|他消灭了 迦南 地七族的人后，把那地分给他们为业，
ACTS|13|20|约有四百五十年。此后 ，他给他们设立士师，直到 撒母耳 先知的时候。
ACTS|13|21|从那时起，他们要求立一个王，上帝就将 便雅悯 支派中 基士 的儿子 扫罗 给他们作王，共四十年。
ACTS|13|22|他废了 扫罗 之后，就兴起 大卫 作他们的王，又为他作见证说：‘我寻得 耶西 的儿子 大卫 ，他是合我心意的人，他要遵行我一切的旨意。’
ACTS|13|23|从这人的后裔中，上帝已经照着所应许的为 以色列 人兴起一位救主，就是耶稣。
ACTS|13|24|在他没有出来以前， 约翰 已向 以色列 全民宣讲悔改的洗礼。
ACTS|13|25|约翰 快走完他的人生路程时，说：‘你们以为我是谁？我不是 ；但是有一位在我以后来的，我就是解他脚上的鞋带也不配。’
ACTS|13|26|“诸位弟兄— 亚伯拉罕 的子孙和你们中间敬畏上帝的人哪，这救世的道是传给我们的。
ACTS|13|27|耶路撒冷 的居民和他们的官长，因为不认识这基督，也不明白每安息日所读的先知的书，把他定了死罪，正应验了先知的预言。
ACTS|13|28|虽然他们查不出他有该死的罪状，还是要求 彼拉多 把他杀了。
ACTS|13|29|他们既实现了经上指着他所记的一切话，就从木头上把他取下来，放在坟墓里。
ACTS|13|30|上帝却使他从死人中复活。
ACTS|13|31|有许多日子，他向那些从 加利利 同他上 耶路撒冷 的人显现，这些人如今在民间成为他的见证人。
ACTS|13|32|我们报好信息给你们，就是那应许祖宗的话，
ACTS|13|33|上帝已经向我们这些作他们儿女的 应验，使耶稣复活了。正如《诗篇》第二篇上记着： ‘你是我的儿子， 我今日生了你。’
ACTS|13|34|论到上帝使他从死人中复活，不再归于朽坏，他曾这样说： ‘我必将所应许 大卫 那圣洁、 可靠的恩典赐给你们。’
ACTS|13|35|所以他也在另一篇说： ‘你必不让你的圣者见朽坏。’
ACTS|13|36|大卫 在世的时候，遵行了上帝的旨意就长眠了 ，归到他祖宗那里，已见朽坏；
ACTS|13|37|惟独上帝使他复活的那一位，他并未见朽坏。
ACTS|13|38|所以弟兄们，你们当知道：赦罪的道是由这人传给你们的，
ACTS|13|39|你们靠 摩西 的律法在不得称义的一切事上，每一个信靠这位耶稣的都得称义了。
ACTS|13|40|所以，你们要小心，免得先知书上所说的临到你们：
ACTS|13|41|‘要观看，你们这些藐视的人， 要惊讶，要灭亡， 因为在你们的日子，我行一件事， 虽有人告诉你们，你们总是不信。’”
ACTS|13|42|他们走出会堂的时候，众人请他们在下一个安息日再讲这些话给他们听。
ACTS|13|43|散会以后，有许多 犹太 人和敬虔的皈依 犹太 教的人跟从了 保罗 和 巴拿巴 。二人对他们讲话，劝他们务要恒久倚靠上帝的恩典。
ACTS|13|44|到下一个安息日，全城的人几乎都聚集起来，要听主的道 。
ACTS|13|45|但 犹太 人看见这么多的人，就满心嫉妒，辩驳 保罗 所说的话，并且毁谤他。
ACTS|13|46|于是 保罗 和 巴拿巴 放胆说：“上帝的道本应先传给你们；只因你们弃绝这道，断定自己不配得永生，我们就转向外邦人。
ACTS|13|47|因为主曾这样吩咐我们： ‘我已经立你作万邦之光， 使你施行我的救恩，直到地极。’”
ACTS|13|48|外邦人听见这话很欢喜，赞美主的道，凡被指定得永生的人都信了。
ACTS|13|49|于是主的道传遍了那一带地方。
ACTS|13|50|但 犹太 人挑唆虔敬尊贵的妇女和城内有名望的人，迫害 保罗 和 巴拿巴 ，把他们赶出境外。
ACTS|13|51|二人对着众人跺掉脚上的尘土，然后往 以哥念 去了。
ACTS|13|52|门徒满心喜乐，又被圣灵充满。
ACTS|14|1|同样的事也发生在 以哥念 。 保罗 和 巴拿巴 进了 犹太 人的会堂，在那里讲道，所以有很多 犹太 人和 希腊 人都信了。
ACTS|14|2|但那不顺从的 犹太 人煽动外邦人，使他们心里仇恨弟兄。
ACTS|14|3|二人在那里住了好些日子，倚靠主放胆讲道，主藉他们的手施行神迹奇事，证明他恩惠的道。
ACTS|14|4|城里的众人却分裂了：有依附 犹太 人的，有依附使徒的。
ACTS|14|5|那时，外邦人、 犹太 人和他们的官长，一齐拥上来，要凌辱使徒，用石头打他们。
ACTS|14|6|使徒知道了，就逃到 吕高尼 的 路司得 和 特庇 两个城，以及周围地方去，
ACTS|14|7|在那里继续传福音。
ACTS|14|8|路司得城 里有一个两脚无力的人，他从母腹里就是瘸腿的，老是坐着，从来没有走过。
ACTS|14|9|他听 保罗 讲道； 保罗 定睛看他，见他有信心，可得痊愈，
ACTS|14|10|就大声说：“起来！两脚站直。”那人就跳起来，开始行走。
ACTS|14|11|众人看见 保罗 所做的事，就用 吕高尼 话大声说：“有神明藉着人形降临在我们中间了。”
ACTS|14|12|于是他们称 巴拿巴 为 宙斯 ，称 保罗 为 希耳米 ，因为他总是带头说话。
ACTS|14|13|城外有 宙斯 庙的祭司牵着牛，拿着花环，来到门前，要同众人一起献祭。
ACTS|14|14|巴拿巴 和 保罗 二位使徒听见，就撕开衣裳，跳进众人中间，喊着：
ACTS|14|15|“诸位，为什么做这些事呢？我们也是人，性情和你们一样。我们传福音给你们，是要你们离弃这些虚妄的事，归向那创造天、地、海和其中万物的永生的上帝。
ACTS|14|16|他在从前的世代，任凭万国各行其道；
ACTS|14|17|然而他未尝不为自己留下证据来，就如常行善事，从天降雨，赏赐丰年，使你们饮食饱足，满心喜乐。”
ACTS|14|18|二人说了这些话，总算拦住众人不献祭给他们。
ACTS|14|19|但有些 犹太 人，从 安提阿 和 以哥念 来，挑唆众人，并且用石头打 保罗 ，以为他死了，就把他拖到城外。
ACTS|14|20|当门徒围着他的时候，他站了起来，走进城去。第二天， 保罗 同 巴拿巴 往 特庇 去。
ACTS|14|21|保罗 和 巴拿巴 对那城里的人传了福音，使好些人成为门徒后，又回 路司得 、 以哥念 、 安提阿 去，
ACTS|14|22|坚固门徒的心，劝他们持守他们的信仰，说：“我们进入上帝的国，必须经历许多艰难。”
ACTS|14|23|二人在各教会中选立了长老，禁食祷告后，把他们交托给他们所信的主。
ACTS|14|24|二人经过 彼西底 来到 旁非利亚 ，
ACTS|14|25|在 别加 讲了道，就下 亚大利 去，
ACTS|14|26|从那里坐船回 安提阿 去。当初，众人就在这地方，把他们交托在上帝的恩典中，要完成现在所做的工。
ACTS|14|27|他们一到那里，就聚集了会众，述说上帝藉他们所行的一切事，并且上帝怎样为外邦人开了信道的门。
ACTS|14|28|二人在那里同门徒住了一段日子。
ACTS|15|1|有几个人从 犹太 下来，教导弟兄们说：“你们若不按照 摩西 的规矩受割礼，不能得救。”
ACTS|15|2|保罗 和 巴拿巴 跟他们发生了激烈的争执和辩论；大家就决定指派 保罗 、 巴拿巴 和本会的几个人，为所辩论的事上 耶路撒冷 去见使徒和长老。
ACTS|15|3|于是教会为他们送行。他们经过 腓尼基 、 撒玛利亚 ，沿途叙说外邦人归主的事，使众弟兄都非常欢喜。
ACTS|15|4|他们到了 耶路撒冷 ，教会、使徒和长老都接待他们，他们就述说上帝同他们所做的一切事。
ACTS|15|5|惟有几个法利赛派的信徒起来，说：“必须给外邦人行割礼，吩咐他们遵守 摩西 的律法。”
ACTS|15|6|使徒和长老聚集商议这事。
ACTS|15|7|辩论了许久后， 彼得 站起来，对他们说：“诸位弟兄，你们知道上帝早已在你们中间拣选了我，让外邦人从我口中得听福音之道，而且相信。
ACTS|15|8|知道人心的上帝也为他们作了见证，赐圣灵给他们，正如给我们一样；
ACTS|15|9|又藉着信洁净了他们的心，他们和我们之间并没有什么分别。
ACTS|15|10|现在你们为什么试探上帝，要把我们祖宗和我们所不能负的轭放在门徒的颈项上呢？
ACTS|15|11|相反地，我们相信，我们得救是因主耶稣的恩典，和他们一样。”
ACTS|15|12|众人都默默无声，听 巴拿巴 和 保罗 述说上帝藉着他们在外邦人中所行的神迹和奇事。
ACTS|15|13|他们讲完了， 雅各 回答说：“诸位弟兄，请听我说。
ACTS|15|14|刚才 西门 述说上帝当初怎样眷顾外邦人，从他们中间选取人民归于自己的名下；
ACTS|15|15|众先知的话也与这意思相符合。
ACTS|15|16|正如经上所写的： ‘此后，我要回来， 重新修造 大卫 倒塌了的帐幕， 从废墟中重新修造， 把它建立起来，
ACTS|15|17|使剩余的人， 就是凡称我名的外邦人， 都寻求主。 这话是自古以来显明这些事的主说的。’
ACTS|15|18|
ACTS|15|19|所以，我的意见是不可难为那归向上帝的外邦人；
ACTS|15|20|但是要写信吩咐他们禁戒偶像所玷污的东西、血和勒死的牲畜 ，禁戒淫乱。
ACTS|15|21|因为历代以来， 摩西 的书在各城都有人宣讲，每逢安息日，也在会堂里诵读。”
ACTS|15|22|那时，使徒、长老和全教会认为应从他们中间拣选人，差他们和 保罗 、 巴拿巴 一同到 安提阿 去，所拣选的就是称为 巴撒巴 的 犹大 和 西拉 。这二人在弟兄中是领袖。
ACTS|15|23|他们带去的信说：“使徒和作长老的弟兄们向 安提阿 、 叙利亚 、 基利家 外邦众弟兄问安。
ACTS|15|24|我们听说，有几个人从我们这里出去 ，用一些话骚扰你们，使你们的心困惑， 其实我们并没有吩咐他们。
ACTS|15|25|我们认为，既然我们同心定意，就拣选几个人，派他们同我们所亲爱的 巴拿巴 和 保罗 到你们那里去。
ACTS|15|26|这二人曾为我主耶稣基督的名不顾自己的性命。
ACTS|15|27|所以我们派 犹大 和 西拉 去，他们也会亲口述说这些事。
ACTS|15|28|因为圣灵和我们决定除了这几件重要的事，不将别的重担放在你们身上，
ACTS|15|29|就是禁戒偶像所玷污的东西、血和勒死的牲畜，禁戒淫乱。这几件你们若能自己禁戒就好了。祝你们安康！”
ACTS|15|30|他们既奉了差遣就下 安提阿 去，聚集会众，把书信交给他们。
ACTS|15|31|众人念了，因为信上鼓励的话而感到欣慰。
ACTS|15|32|犹大 和 西拉 自己也是先知，就用许多话劝勉弟兄，坚固他们。
ACTS|15|33|二人住了些日子，弟兄们打发他们平平安安地回到差遣他们的人那里去。
ACTS|15|34|
ACTS|15|35|但 保罗 和 巴拿巴 仍留在 安提阿 ，和许多别的人一同教导，并传扬主的道。
ACTS|15|36|过了些日子， 保罗 对 巴拿巴 说：“让我们回到从前宣扬主道的各城，看看弟兄们的情况如何。”
ACTS|15|37|巴拿巴 有意要带称为 马可 的 约翰 同去；
ACTS|15|38|但 保罗 认为不宜带他去，因为 马可 从前在 旁非利亚 离开他们，不和他们一起工作。
ACTS|15|39|于是二人起了争执，甚至彼此分手。 巴拿巴 带着 马可 ，坐船往 塞浦路斯 去；
ACTS|15|40|保罗 则拣选了 西拉 ，也出发了，蒙弟兄们把他交于主的恩典中。
ACTS|15|41|他就走遍了 叙利亚 、 基利家 ，坚固众教会。
ACTS|16|1|后来， 保罗 来到 特庇 ，又到 路司得 。在那里有一个门徒，名叫 提摩太 ，是信主的 犹太 妇人的儿子，他父亲却是 希腊 人。
ACTS|16|2|路司得 和 以哥念 的弟兄都称赞他。
ACTS|16|3|保罗 要带他同去，只因那些地方的 犹太 人都知道他父亲是 希腊 人，就给他行了割礼。
ACTS|16|4|他们经过各城，把 耶路撒冷 使徒和长老所决定的规条交给门徒遵守。
ACTS|16|5|于是众教会信心越发坚固，人数天天增加。
ACTS|16|6|因为圣灵禁止他们在 亚细亚 讲道，他们就经过 弗吕家 、 加拉太 一带地方。
ACTS|16|7|到了 每西亚 的边界，他们想要往 庇推尼 去，耶稣的灵却不许。
ACTS|16|8|他们就越过 每西亚 ，下 特罗亚 去。
ACTS|16|9|夜间，有异象向 保罗 显现。有一个 马其顿 人站着求他说：“请你过来，到 马其顿 来帮助我们！”
ACTS|16|10|保罗 既看见这异象，我们就立即设法往 马其顿 去，认为上帝呼召我们传福音给那里的人。
ACTS|16|11|我们从 特罗亚 开船，直行驶到 撒摩特喇 ，第二天到了 尼亚坡里 ；
ACTS|16|12|从那里来到 腓立比 ，就是 马其顿 这一带的一个重要城市 ，也是 罗马 的驻防城。我们在这城里住了几天。
ACTS|16|13|在安息日，我们出城门，到了河边，知道那里有一个祷告的地方 ，我们就坐下来对那些聚会的妇女讲道。
ACTS|16|14|有一个卖紫色布的妇人，名叫 吕底亚 ，是 推雅推喇城 的人，素来敬拜上帝。她在听着，主就开导她的心，使她留心听 保罗 所讲的话。
ACTS|16|15|她和她一家都领了洗，就求我们说：“你们若以为我是真心信主的 ，请到我家里来住。”于是她坚决请我们留下。
ACTS|16|16|后来，我们往那祷告的地方去时，有一个被占卜的灵附身的使女迎面走来，她使用法术使她的主人们发了大财。
ACTS|16|17|她跟随 保罗 和我们，喊着说：“这些人是至高上帝的仆人，对你们传讲救人的道路。”
ACTS|16|18|她一连好几天这样喊叫， 保罗 就心中厌烦，转身对那灵说：“我奉耶稣基督的名吩咐你从她身上出来！”那灵立刻出来了。
ACTS|16|19|使女的主人们见发财的指望没有了，就揪住 保罗 和 西拉 ，拉他们到市上去见官；
ACTS|16|20|又带他们到行政官长们面前，说：“这些骚扰我们城的，他们是 犹太 人，
ACTS|16|21|竟传布我们 罗马 人所不可接受、不可遵守的规矩。”
ACTS|16|22|群众就一齐起来攻击他们。官长们吩咐撕开他们的衣裳，用棍子打；
ACTS|16|23|打了许多棍，就把他们下在监里，嘱咐狱警严紧看守。
ACTS|16|24|狱警领了这样的命令，就把他们下在内监，两脚拴在木架上。
ACTS|16|25|约在半夜， 保罗 和 西拉 正在祷告，唱诗赞美上帝，众囚犯也侧耳听着的时候，
ACTS|16|26|忽然，地大震动，甚至监牢的地基都摇动了，监门立刻全开，众囚犯的锁链也都解开了。
ACTS|16|27|狱警一醒，看见监门全开，以为囚犯已经逃走，就拔刀要自杀。
ACTS|16|28|保罗 大声呼叫：“不要伤害自己！我们都在这里。”
ACTS|16|29|狱警叫人拿灯来，就冲进去，战战兢兢地俯伏在 保罗 和 西拉 面前。
ACTS|16|30|然后狱警领他们出来，说：“二位先生，我必须做什么才可以得救？”
ACTS|16|31|他们说：“当信主耶稣，你和你一家都必得救 。”
ACTS|16|32|他们就把主的道讲给他和他全家的人听。
ACTS|16|33|当夜，就在那时候，狱警把他们带去，洗他们的伤；他和他所有的家人立刻都受了洗。
ACTS|16|34|于是狱警领他们上自己的家里去，给他们摆上饭。他和全家的人，因为信了上帝，都满心喜乐。
ACTS|16|35|到了天亮，官长们打发差役来，说：“释放那两个人吧。”
ACTS|16|36|狱警就把这些话告诉 保罗 ：“官长们打发人来，要释放你们，现在可以出监，平平安安去吧。”
ACTS|16|37|保罗 却说：“我们是 罗马 人，并没有定罪，他们竟在公众面前打了我们，又把我们下在监里；现在要私下赶我们出去吗？这不行！叫他们自己来领我们出去吧！”
ACTS|16|38|差役把这些话回禀官长们；官长们听见他们是 罗马 人，就害怕了，
ACTS|16|39|于是来劝他们，领他们出来，请他们离开那城。
ACTS|16|40|二人出了监牢，往 吕底亚 家里去，见了弟兄们，劝慰他们一番，就离开了。
ACTS|17|1|保罗 和 西拉 经过 暗妃坡里 、 亚波罗尼亚 ，来到 帖撒罗尼迦 ，在那里有 犹太 人的会堂。
ACTS|17|2|保罗 照他素常的规矩进去，一连三个安息日，根据圣经与他们辩论，
ACTS|17|3|讲解和说明基督必须受害，从死人中复活；又说：“我所传给你们的这位耶稣就是基督。”
ACTS|17|4|他们中间有些人听了劝，就跟从 保罗 和 西拉 ，还有许多虔敬的 希腊 人，尊贵的妇女也不少。
ACTS|17|5|但不信的 犹太 人心里嫉妒，聚集了些市井流氓，搭伙成群，煽动全城的人闯进 耶孙 的家，要把 保罗 和 西拉 带到民众那里。
ACTS|17|6|那些人找不着他们，就把 耶孙 和几个弟兄拉到地方官那里，喊叫着：“这些搅乱天下的人也到这里来了，
ACTS|17|7|耶孙 竟收留他们。这些人都违背凯撒的命令，说另有一个王耶稣。”
ACTS|17|8|众人和地方官听见这些话，就惶恐了，
ACTS|17|9|于是收了 耶孙 和其余的人的保证金后，释放了他们。
ACTS|17|10|当夜，弟兄们立刻送 保罗 和 西拉 往 庇哩亚 去；二人到了，就进入 犹太 人的会堂。
ACTS|17|11|这地方的 犹太 人比 帖撒罗尼迦 的人开明，热心领受这道，天天查考圣经，要知道这道是否真实。
ACTS|17|12|所以，他们中间有许多信了，又有 希腊 的尊贵妇人，男人也不少。
ACTS|17|13|但 帖撒罗尼迦 的 犹太 人知道 保罗 又在 庇哩亚 传上帝的道，就往那里去，煽动挑拨群众。
ACTS|17|14|于是，弟兄们立刻送 保罗 到海边去， 西拉 和 提摩太 却仍留在 庇哩亚 。
ACTS|17|15|护送 保罗 的人带他到了 雅典 ，他们领了 保罗 的命令，叫 西拉 和 提摩太 赶快到他那里来，然后回去了。
ACTS|17|16|保罗 在 雅典 等候他们的时候，看见满城都是偶像，就心里非常难过。
ACTS|17|17|于是他在会堂里与 犹太 人和虔敬的人，以及每日在市场上所遇见的人辩论。
ACTS|17|18|还有 伊壁鸠鲁 和 斯多亚 两派的哲学家也与他争辩。有的说：“这胡言乱语的要说什么？”有的说：“他似乎是宣传外邦鬼神的。”这是因 保罗 传讲耶稣与复活的福音。
ACTS|17|19|他们就把他带到 亚略巴古 ，说：“你所讲的这新学说，我们也可以知道吗？
ACTS|17|20|因为你有些奇怪的事传到我们耳中，我们想知道这些事是什么意思。”
ACTS|17|21|原来所有的 雅典 人和居住在那里的外国人都无暇管别的事，只是谈谈或听听新闻。
ACTS|17|22|保罗 站在 亚略巴古 当中，说：“诸位 雅典 人！我看你们凡事很敬畏鬼神。
ACTS|17|23|我到处走走的时候，仔细观察你们所敬拜的，发现一座坛，上面写着‘献给未识之神明’。你们所不认识而敬拜的，我现在向你们宣告：
ACTS|17|24|他是创造宇宙和其中万物的上帝；他既是天地的主，就不住在人手所造的殿宇里，
ACTS|17|25|也不用人手去服侍，好像缺少什么似的；自己倒将生命、气息、万物赐给万人。
ACTS|17|26|他从一人 造出万族，居住在全地面上，并且预先定准他们的年限和所住的疆界，
ACTS|17|27|为要使他们寻求上帝，或者可以揣摩而找到他，其实他离我们各人不远。
ACTS|17|28|我们生活、行动、存在都在于他。就如你们的诗人也有人说：‘我们也是他所生的。’
ACTS|17|29|既然我们是上帝所生的，就不应该以为上帝的神性像人用手艺和心思所雕刻的金、银、石像一般。
ACTS|17|30|世人蒙昧无知的时候，上帝并不追究，如今却吩咐各处的人都要悔改。
ACTS|17|31|因为他已经定了日子，要藉着他所设立的人按公义审判天下，并且使他从死人中复活，给万人作可信的凭据。”
ACTS|17|32|众人听见死人复活的话，就有人讥诮他；又有人说：“我们会再听你讲这事。”
ACTS|17|33|于是 保罗 从他们当中出去了。
ACTS|17|34|但有几个人依附他，信了主，其中有 亚略巴古 的议员 丢尼修 ，和一个名叫 大马哩 的妇人，还有几个与他们一起的人。
ACTS|18|1|这些事以后， 保罗 离开 雅典 ，来到 哥林多 。
ACTS|18|2|他遇见一个生在 本都 的 犹太 人，名叫 亚居拉 。不久前，他带着妻子 百基拉 从 意大利 来，因为 克劳第 命令所有的 犹太 人都离开 罗马 。 保罗 去投靠他们。
ACTS|18|3|他们本是制造帐棚为业。 保罗 因与他们同业，就和他们同住，一同做工。
ACTS|18|4|每逢安息日， 保罗 在会堂里辩论，劝导 犹太 人和 希腊 人。
ACTS|18|5|西拉 和 提摩太 从 马其顿 来的时候， 保罗 正专心传道，向 犹太 人证明耶稣是基督。
ACTS|18|6|当他们抗拒他、毁谤他的时候，他就抖掉衣裳的灰尘，对他们说：“你们的罪归到你们自己的头上，与我无干。从今以后，我要往外邦人那里去。”
ACTS|18|7|于是他离开那里，到了一个人的家里，他名叫 提多．犹士都 ，是敬拜上帝的人，他的家靠近会堂。
ACTS|18|8|会堂的主管 基利司布 和全家都信了主，还有许多 哥林多 人听了就信，而且受了洗。
ACTS|18|9|夜间，主在异象中对 保罗 说：“不要怕，只管讲，不要沉默，
ACTS|18|10|有我与你同在，没有人会下手害你，因为在这城里有许多属我的人。”
ACTS|18|11|保罗 在那里住了一年六个月，将上帝的道教导他们。
ACTS|18|12|到 迦流 作 亚该亚 省长的时候， 犹太 人齐心起来攻击 保罗 ，拉他到法庭，
ACTS|18|13|说：“这个人教唆人不按着律法敬拜上帝。”
ACTS|18|14|保罗 刚要开口， 迦流 对 犹太 人说：“你们这些 犹太 人哪！如果是为冤枉或奸恶的事，我理当耐性听你们。
ACTS|18|15|既然你们所争论的是关乎用字、名目和你们的律法，你们自己去办吧！这样的事我不愿意审问。”
ACTS|18|16|于是，他把他们逐出法庭。
ACTS|18|17|众人就揪住会堂的主管 所提尼 ，在法庭前打他。这些事 迦流 都不管。
ACTS|18|18|保罗 又住了好些日子，就辞别了弟兄，坐船到 叙利亚 去。 百基拉 、 亚居拉 和他同去。他因为许过愿，就在 坚革哩 剃了头发。
ACTS|18|19|到了 以弗所 ， 保罗 就把他们留在那里，自己进了会堂，和 犹太 人辩论。
ACTS|18|20|众人请他多住些日子，他没有答应，
ACTS|18|21|就辞别他们，说：“上帝若许可，我还要回到你们这里来。”于是他上船离开 以弗所 。
ACTS|18|22|他在 凯撒利亚 下了船，上 耶路撒冷 去问候教会，随后下 安提阿 去。
ACTS|18|23|他在那里住了些日子，又离开了那里，逐一经过 加拉太 和 弗吕家 各地方，坚固众门徒。
ACTS|18|24|有一个生在 亚历山大 的 犹太 人，名叫 亚波罗 ，来到 以弗所 ，他很有口才，很会讲解圣经。
ACTS|18|25|这人已经在主的道路上受了训练，心里火热，精确地讲论和教导耶稣的事；可是他只知道 约翰 的洗礼。
ACTS|18|26|他开始在会堂里放胆讲道； 百基拉 、 亚居拉 听见，就接他来，将上帝的道路 给他更精确地讲解。
ACTS|18|27|他想要往 亚该亚 去，弟兄们就勉励他，并写信请门徒们接待他，他到了那里，多多帮助那些蒙恩信主的人，
ACTS|18|28|因为他在公众面前极力驳倒 犹太 人，引圣经证明耶稣是基督。
ACTS|19|1|亚波罗 在 哥林多 的时候， 保罗 经过了内陆地区，来到 以弗所 ，在那里他遇见几个门徒，
ACTS|19|2|问他们：“你们信的时候领受了圣灵没有？”他们说：“没有，我们连什么是圣灵都没有听过。”
ACTS|19|3|保罗 说：“这样，你们受的是什么洗呢？”他们说：“是受了 约翰 的洗。”
ACTS|19|4|保罗 说：“ 约翰 所施的是悔改的洗礼，他告诉百姓当信那在他以后要来的那位，就是耶稣。”
ACTS|19|5|他们听见这话以后，就奉主耶稣的名受洗。
ACTS|19|6|保罗 给他们按手，圣灵就降在他们身上，他们开始说方言 和说预言。
ACTS|19|7|他们约有十二个人。
ACTS|19|8|保罗 进会堂，一连三个月放胆讲道，辩论上帝国的事，劝导众人。
ACTS|19|9|后来，有些人心里刚硬不信，在众人面前毁谤这道； 保罗 就离开他们，也叫门徒与他们分开，就在 推喇奴 的讲堂天天辩论。
ACTS|19|10|这样有两年之久，使一切住在 亚细亚 的，无论是 犹太 人是 希腊 人，都听见主的道。
ACTS|19|11|上帝藉 保罗 的手行了些奇异的神迹，
ACTS|19|12|甚至有人从 保罗 身上拿走手巾或围裙放在病人身上，病就消除了，邪灵也出去了。
ACTS|19|13|那时，有几个巡回各处念咒赶鬼的 犹太 人，擅自利用主耶稣的名，向那些被邪灵所附的人说：“我奉 保罗 所传的耶稣命令你们出来！”
ACTS|19|14|做这事的是 犹太 祭司长 士基瓦 的七个儿子。
ACTS|19|15|但邪灵回答他们：“耶稣我知道， 保罗 我也认识，你们却是谁呢？”
ACTS|19|16|被邪灵所附的人就扑到他们身上，制伏他们，胜过他们，使他们赤着身子，受了伤，从那房子里逃出去了。
ACTS|19|17|凡住在 以弗所 的，无论是 犹太 人是 希腊 人，都知道这件事，也都惧怕；主耶稣的名从此就更被尊为大了。
ACTS|19|18|许多已经信的人来承认并公开自己所行的事。
ACTS|19|19|又有许多平素行邪术的人把他们的书都拿来，堆积在众人面前焚烧。他们计算书价，得知共值五万块银钱。
ACTS|19|20|这样，主的道大大兴旺，而且普遍传开了。
ACTS|19|21|这些事过后， 保罗 心里决定要经过 马其顿 、 亚该亚 ，就往 耶路撒冷 去。他说：“我到了那里以后，也必须到 罗马 去看看。”
ACTS|19|22|于是他差遣两个助手 提摩太 和 以拉都 往 马其顿 去，自己暂时留在 亚细亚 。
ACTS|19|23|那时，因这道路而起的骚动不小。
ACTS|19|24|有一个银匠，名叫 底米丢 ，是制造 亚底米 神银龛的，他使从事这手艺的人生意发达。
ACTS|19|25|他聚集他们和同行的工人，说：“诸位，你们知道我们是倚靠这生意发财的。
ACTS|19|26|你们看到，也听见这 保罗 不但在 以弗所 ，也几乎在 亚细亚 全地，引诱迷惑了许多人，说：‘人手所做的不是神明。’
ACTS|19|27|这样，不仅我们这行业陷入被藐视的危险，就是大女神 亚底米 的庙也要被人轻看，连 亚细亚 全地和普天下所敬拜的女神的威望也受损害了。”
ACTS|19|28|众人听见，就怒气冲冲，喊着说：“大哉， 以弗所 人的 亚底米 ！”
ACTS|19|29|于是满城都骚动起来。众人抓住与 保罗 同行的 马其顿 人 该犹 和 亚里达古 ，齐心冲进剧场。
ACTS|19|30|保罗 想要进到民众那里，门徒却不许他去。
ACTS|19|31|连 亚细亚 的几位官员，是 保罗 的朋友，也打发人来劝他不要冒险到剧场里去。
ACTS|19|32|聚集的人乱成一团，有的喊这个，有的喊那个，大半不知道为了什么聚集。
ACTS|19|33|犹太 人把 亚历山大 推出去，人群中有人怂恿他，他就做手势，要向民众申诉。
ACTS|19|34|但他们一认出他是 犹太 人，大家就异口同声喊着：“大哉， 以弗所 人的 亚底米 ！”约喊了两小时。
ACTS|19|35|城里的书记官安抚了群众后，说：“ 以弗所 人哪，谁不知道 以弗所 人的城是看守大 亚底米 的庙和从 宙斯 那里落下来的像的守护者呢？
ACTS|19|36|既然这些事是驳不倒的，你们就要安静下来，不可妄动。
ACTS|19|37|你们把这些人带来，他们并没有偷窃庙中之物，也没有亵渎我们的女神。
ACTS|19|38|如果 底米丢 和他同行的手艺人有控告的事，自有公堂，也有省长，他们可以彼此控告。
ACTS|19|39|你们若有别的事请求，可以在合法的集会里解决。
ACTS|19|40|今日的扰乱本是无缘无故的，有被控告的危险。这次的骚动，我们也说不出理由来。”
ACTS|19|41|他说完这些话，就叫众人散会。
ACTS|20|1|骚乱平定以后， 保罗 请门徒来，劝勉了他们，就辞别他们，往 马其顿 去。
ACTS|20|2|他走遍那一带地方，用许多话劝勉门徒，然后来到 希腊 ，
ACTS|20|3|在那里住了三个月。他快要坐船往 叙利亚 去的时候， 犹太 人设计害他，他就决定从 马其顿 回去。
ACTS|20|4|同他到 亚细亚 去的，有 庇哩亚 人 毕罗斯 的儿子 所巴特 ， 帖撒罗尼迦 人 亚里达古 和 西公都 ，还有 特庇 人 该犹 和 提摩太 ，又有 亚细亚 人 推基古 和 特罗非摩 。
ACTS|20|5|这些人先走，在 特罗亚 等候我们。
ACTS|20|6|过了除酵节的日子，我们从 腓立比 开船，五天以后到了 特罗亚 ，和他们相会，在那里住了七天。
ACTS|20|7|七日的第一日，我们聚会擘饼的时候， 保罗 因次日要起行，就为他们讲道，直讲到半夜。
ACTS|20|8|我们聚会的那座楼上有好些灯火。
ACTS|20|9|有一个少年，名叫 犹推古 ，坐在窗口上，沉沉入睡。 保罗 讲了多时，少年睡熟了，从三层楼上掉下去，扶起来时已经死了。
ACTS|20|10|保罗 下去，伏在他身上，抱着他，说：“你们不要慌乱，他还有气呢！”
ACTS|20|11|保罗 又上楼去，擘饼，吃了，再讲了许久，直到天亮才离开。
ACTS|20|12|他们把那活过来的孩子带走，大家得到很大的安慰。
ACTS|20|13|我们先上船，起航往 亚朔 去，想要在那里接 保罗 ；因为他是这样安排的，他自己本来打算要走陆路。
ACTS|20|14|他既在 亚朔 与我们相会，我们就接他上船，来到 米推利尼 。
ACTS|20|15|我们从那里开船，第二天到了 基阿 的对岸；再下一天，在 撒摩 靠岸，又过了一天，到了 米利都 。
ACTS|20|16|因为 保罗 早已决定要越过 以弗所 ，免得在 亚细亚 耽延，他急忙前行，假如可能的话，在五旬节前能赶到 耶路撒冷 。
ACTS|20|17|保罗 从 米利都 打发人往 以弗所 去，请教会的长老来。
ACTS|20|18|他们来了， 保罗 对他们说：“你们自己知道，自从我到 亚细亚 的第一天，我怎样跟你们相处，
ACTS|20|19|怎样凡事谦卑，以眼泪服侍主，又因 犹太 人的谋害经历试炼。
ACTS|20|20|你们也知道，凡对你们有益的，我没有一样隐瞒不说的，或在公众面前，或在每一个人的家里，我都教导你们，
ACTS|20|21|不论 犹太 人和 希腊 人，我都已证明他们当在上帝面前悔改，信靠我们的主耶稣。
ACTS|20|22|现在我被圣灵催迫 要往 耶路撒冷 去，虽然不知道在那里会遭遇什么事，
ACTS|20|23|但知道圣灵在各城里向我指证，说有捆锁与患难等着我。
ACTS|20|24|我却不以性命为念，只要走完我的路程，完成我从主耶稣所领受的职分，为上帝恩典的福音作见证。
ACTS|20|25|“我素常在你们中间到处传讲上帝的国；现在我知道，你们众人以后不会再见到我的面了。
ACTS|20|26|所以我今日向你们作证，你们中间无论何人死亡，罪不在我。
ACTS|20|27|因为上帝一切的旨意，我并没有退缩不传给你们的。
ACTS|20|28|圣灵立你们作全群的监督，你们就当为自己谨慎，也为全群谨慎，牧养上帝 的教会，就是他用自己血所买来的 。
ACTS|20|29|我知道，在我离开以后必有凶暴的豺狼进入你们中间，不顾惜羊群。
ACTS|20|30|就是你们中间也必有人起来，说悖谬的话，要引诱门徒跟从他们。
ACTS|20|31|所以你们要警醒，记念我三年之久，昼夜不断地流泪劝戒你们各人。
ACTS|20|32|现在我把你们交托给上帝和他恩惠的道；这道能建立你们，使你们和一切成圣的人同得基业。
ACTS|20|33|我未曾贪图一个人的金、银或衣服。
ACTS|20|34|你们自己知道，我靠两只手工作来供给我和同工的需用。
ACTS|20|35|我凡事给你们作榜样，叫你们知道应当这样劳苦，扶助软弱的人，又当记念主耶稣的话，说：‘施比受更为有福。’”
ACTS|20|36|保罗 说完了这些话，就和大家跪下来祷告。
ACTS|20|37|众人痛哭，抱着 保罗 的颈项跟他亲吻。
ACTS|20|38|叫他们最伤心的，就是他说“以后不会再见到我的面”那句话。于是他们送他上船去了。
ACTS|21|1|我们离别了众人，就开船直航到 哥士 ，第二天到了 罗底 ，又从那里到 帕大喇 。
ACTS|21|2|我们遇见一只船要往 腓尼基 去，就上船起航。
ACTS|21|3|我们望见 塞浦路斯 ，就从南边行过，往 叙利亚 去，在 推罗 上岸，因为船要在那里卸货。
ACTS|21|4|我们在那里找到了一些门徒，就住了七天。他们藉着圣灵的感动，告诉 保罗 不要上 耶路撒冷 去。
ACTS|21|5|几天之后，我们又出发前行。他们众人同妻子儿女都送我们到城外，我们都跪在滩上祷告，彼此辞别。
ACTS|21|6|我们上了船，他们就回家去了。
ACTS|21|7|我们从 推罗 行完航程，来到了 多利买 ，问候那里的弟兄，和他们同住了一天。
ACTS|21|8|第二天，我们离开那里，来到 凯撒利亚 ，就进了传福音的 腓利 家里，和他同住；他是那七个执事里的一个。
ACTS|21|9|他有四个女儿，都是未出嫁的，都会说预言。
ACTS|21|10|我们在那里多住了好几天，有一个先知，名叫 亚迦布 ，从 犹太 下来。
ACTS|21|11|他到了我们这里，就拿 保罗 的腰带，捆上自己的手脚，说：“圣灵这样说：‘ 犹太 人在 耶路撒冷 要如此捆绑这腰带的主人，把他交在外邦人手里。’”
ACTS|21|12|我们听见这些话，就跟当地的人苦劝 保罗 不要上 耶路撒冷 去。
ACTS|21|13|于是 保罗 回答：“你们为什么这样痛哭，使我心碎呢？我为主耶稣的名，不但被人捆绑，就是死在 耶路撒冷 也是愿意的。”
ACTS|21|14|既然 保罗 不听劝，我们就住了口，只说：“愿主的旨意成就。”
ACTS|21|15|过了这几天，我们收拾行李上 耶路撒冷 去。
ACTS|21|16|有 凯撒利亚 的几个门徒和我们同去，带我们到一个早期的门徒 塞浦路斯 人 拿孙 的家里，请我们与他同住。
ACTS|21|17|我们到了 耶路撒冷 ，弟兄们欢欢喜喜地接待我们。
ACTS|21|18|第二天， 保罗 同我们去见 雅各 ；所有的长老也都在场。
ACTS|21|19|保罗 向他们问安，然后将上帝用他在外邦人中所做的事奉，一一述说了。
ACTS|21|20|他们听见了，就归荣耀给上帝，对 保罗 说：“弟兄，你看 犹太 人中有数以万计的信徒，而他们都是热心于律法的人。
ACTS|21|21|他们曾听见人说，你教导所有在外邦的 犹太 人离弃 摩西 ，对他们说，不要给孩子行割礼，也不要遵守规矩。
ACTS|21|22|众人必听见你来了，这可怎么办呢？
ACTS|21|23|你就照着我们的话做吧！我们这里有四个人，都有愿在身。
ACTS|21|24|你带他们去，与他们一同行洁净的礼，替他们缴纳规费，让他们得以剃头。这样，众人就会知道，先前所听见关于你的事都是假的；而且也知道，你自己为人循规蹈矩，遵行律法。
ACTS|21|25|至于信主的外邦人， 我们已经根据我们的决议写信，叫他们要禁戒偶像所玷污的东西、血和勒死的牲畜，禁戒淫乱。”
ACTS|21|26|于是 保罗 带着那四个人，第二天与他们一同行了洁净礼，进了圣殿，报告洁净期满的日子，等候祭司为他们各人献上祭物。
ACTS|21|27|那七日将完，从 亚细亚 来的 犹太 人看见 保罗 在圣殿里，就煽动所有的群众，下手拿住他，
ACTS|21|28|喊着：“ 以色列 人哪，来帮忙！这就是在各处教导众人糟蹋我们百姓、律法和这地方的人。不但如此，他还带了 希腊 人进圣殿，污秽了这圣地。”
ACTS|21|29|这话是因他们曾看见 以弗所 人 特罗非摩 跟 保罗 一起在城里，以为 保罗 带他进了圣殿。
ACTS|21|30|于是全城都骚动，百姓一齐跑来，拿住 保罗 ，拉他出圣殿，殿门立刻都关了。
ACTS|21|31|他们正想要杀他，有人报信给营里的千夫长，说 耶路撒冷 全城都乱了。
ACTS|21|32|千夫长立刻带着士兵和几个百夫长，跑下去到他们那里。他们见了千夫长和士兵，就停下来不打 保罗 。
ACTS|21|33|于是千夫长上前拿住他，吩咐用两条铁链捆锁，又问他是什么人，做了什么事。
ACTS|21|34|群众中有的喊这个，有的喊那个；因为这样乱嚷，千夫长无法知道实情，就下令将 保罗 带进营楼去。
ACTS|21|35|保罗 一走上台阶，群众挤得凶猛，士兵只得将 保罗 抬起来。
ACTS|21|36|一群人跟在后面，喊着：“除掉他！”
ACTS|21|37|保罗 快要被带进营楼时，对千夫长说：“我可以对你说句话吗？”千夫长说：“你懂得 希腊 话吗？
ACTS|21|38|那你就不是从前作乱、带领四千凶徒往旷野去的那 埃及 人了。”
ACTS|21|39|保罗 说：“我本是 犹太 人，生在 基利家 的 大数 ，并不是无名小城的公民。求你准我对百姓说话。”
ACTS|21|40|千夫长准了。 保罗 就站在台阶上，向百姓做了个手势，要他们静下来， 保罗 就用 希伯来 话对他们说：
ACTS|22|1|“诸位父老弟兄，请听我现在对你们的申辩。”
ACTS|22|2|他们听 保罗 说的是 希伯来 话，就更加安静了。
ACTS|22|3|保罗 说：“我原是 犹太 人，生在 基利家 的 大数 ，但在这城里长大，在 迦玛列 门下按着我们祖宗严紧的律法受教，热心事奉上帝，就如你们大家今日一样。
ACTS|22|4|我也曾迫害信奉这道路的人，置他们于死地，无论男女都捆绑，关在监里。
ACTS|22|5|这是大祭司和议会的众长老都可以给我作证的。我又从他们那里领了致弟兄们的书信，往 大马士革 去，要把在那里的信徒绑起来，带到 耶路撒冷 受刑。”
ACTS|22|6|“当我走近 大马士革 的时候，约在中午，忽然有一道大光从天上下来，照射在我周围。
ACTS|22|7|我就仆倒在地，听见有声音对我说：‘ 扫罗 ！ 扫罗 ！你为什么迫害我？’
ACTS|22|8|我回答：‘主啊！你是谁？’他对我说：‘我就是你所迫害的 拿撒勒 人耶稣。’
ACTS|22|9|跟我一起的人看见了那光，却没有听见那位对我说话的声音。
ACTS|22|10|我说：‘主啊，我该做什么？’主说：‘起来，进 大马士革 去，在那里有人会把指派你做的一切事告诉你。’
ACTS|22|11|我因那光的闪耀不能看见，跟我一起的人就拉着我的手进了 大马士革 。
ACTS|22|12|“那里有一个人，名叫 亚拿尼亚 ，按着律法是虔诚人，为所有住在那里的 犹太 人所称赞。
ACTS|22|13|他来见我，站在旁边，对我说：‘ 扫罗 弟兄，你看见吧！’就在那时，我恢复视觉，看见了他。
ACTS|22|14|他又说：‘我们祖宗的上帝拣选了你，让你明白他的旨意，又看见那义者，听见他口中所出的声音。
ACTS|22|15|因为你要将所看见的、所听见的，对着万人作他的见证人。
ACTS|22|16|现在你为什么耽延呢？起来，受洗，求告他的名，洗去你的罪。’”
ACTS|22|17|“后来，我回到 耶路撒冷 ，在圣殿里祷告的时候，魂游象外，
ACTS|22|18|看见主对我说：‘你赶紧离开 耶路撒冷 ，越快越好，因为这里的人不接受你为我作的见证。’
ACTS|22|19|我就说：‘主啊，他们都知道，我从前在各会堂里把信你的人监禁，又鞭打他们。
ACTS|22|20|当你的见证人 司提反 被害流血的时候，我也站在一旁赞同；又为打死他的人看守衣裳。’
ACTS|22|21|主对我说：‘你去吧！我要差你到远方外邦人那里去。’”
ACTS|22|22|众人听他说到这句话，就高声说：“这样的人，从地上除掉他吧！他是该死的。”
ACTS|22|23|大家一边喧嚷一边摔衣裳，向空中撒灰尘。
ACTS|22|24|千夫长下令把 保罗 带进营楼，叫人用鞭子拷问他，要知道他们向他这样喧嚷是什么缘故。
ACTS|22|25|他们刚用皮条把他捆上的时候， 保罗 对站在旁边的百夫长说：“一个 罗马 人，又未被定罪，你们就鞭打他是合法的吗？”
ACTS|22|26|百夫长听见这话，就去见千夫长，报告说：“你要怎么办呢？这个人是 罗马 人。”
ACTS|22|27|千夫长就来问 保罗 ：“你告诉我，你是 罗马 人吗？” 保罗 说：“是。”
ACTS|22|28|千夫长回答：“我用了许多银子才得到 罗马 公民的身份。” 保罗 说：“我生来就是。”
ACTS|22|29|于是那些要拷问 保罗 的人立刻离开他走了。千夫长一知道他是 罗马 人，又因为曾捆绑了他，也害怕起来。
ACTS|22|30|第二天，千夫长为要知道 犹太 人控告 保罗 的实情，就解开他，下令祭司长们和全议会的人都聚集，然后将 保罗 带下来，叫他站在他们面前。
ACTS|23|1|保罗 定睛看着议会的人，说：“诸位弟兄，我在上帝面前，行事为人都是凭着清白的良心，直到今日。”
ACTS|23|2|亚拿尼亚 大祭司就吩咐旁边站着的人打他的嘴。
ACTS|23|3|这时， 保罗 对他说：“你这粉饰的墙，上帝要打你！你坐堂是要按律法审问我，你竟违背律法，命令人打我吗？”
ACTS|23|4|站在旁边的人说：“你竟敢辱骂上帝的大祭司吗？”
ACTS|23|5|保罗 说：“弟兄们，我不知道他是大祭司；因为经上记着：‘不可毁谤你百姓的官长。’”
ACTS|23|6|保罗 看出他们一部分是撒都该人，一部分是法利赛人，就在议会中喊着：“诸位弟兄，我是法利赛人，也是法利赛人的子孙。我现在受审问是为有关死人复活的盼望。”
ACTS|23|7|说了这话，法利赛人和撒都该人争论起来，会众分为两派。
ACTS|23|8|因为撒都该人一方面说没有复活，另一方面没有天使和鬼魂；法利赛人却承认两方面都有。
ACTS|23|9|于是大大地争吵起来；有几个法利赛派的文士站起来争辩说：“我们看不出这人有什么错处；说不定有鬼魂或者天使对他说过话呢！”
ACTS|23|10|那时争辩越来越大，千夫长恐怕 保罗 被他们扯碎了，就命令士兵下去，把他从众人当中抢出来，带进营楼去。
ACTS|23|11|当夜，主站在 保罗 旁边，说：“放心吧！你怎样在 耶路撒冷 为我作见证，也必怎样在 罗马 为我作见证。”
ACTS|23|12|到了天亮， 犹太 人同谋起誓，说“若不先杀 保罗 就不吃不喝”。
ACTS|23|13|参与这阴谋的有四十多人。
ACTS|23|14|他们来见祭司长和长老，说：“我们已经发了重誓，若不先杀 保罗 就什么也不吃。
ACTS|23|15|现在你们和议会要通知千夫长，叫他把 保罗 带到你们这里来，假装要详细调查他的事；我们已经预备好，在他来到这里以前就杀掉他。”
ACTS|23|16|保罗 的外甥听见他们设下埋伏，就来到营楼里告诉 保罗 。
ACTS|23|17|保罗 请一个百夫长来，说：“你领这青年去见千夫长，他有事告诉他。”
ACTS|23|18|于是百夫长把他领去见千夫长，说：“被囚的 保罗 请我到他那里，求我领这青年来见你；他有事告诉你。”
ACTS|23|19|千夫长就拉着他的手，走到一旁，私下问他：“你有什么事告诉我呢？”
ACTS|23|20|他说：“ 犹太 人已经约定，要求你明天把 保罗 带到议会去，假装要详细查问他的事。
ACTS|23|21|你切不要随从他们，因为他们有四十多人埋伏，已经起誓，若不先杀掉 保罗 就不吃不喝。现在都预备好了，只等你的允准。”
ACTS|23|22|于是千夫长打发那青年走，嘱咐他：“不要告诉人，你已将这些事报告我了。”
ACTS|23|23|于是，千夫长叫了两个百夫长来，说：“预备步兵二百、骑兵七十、长枪手二百，今夜九点往 凯撒利亚 去；
ACTS|23|24|也要预备牲口让 保罗 骑上，护送到 腓力斯 总督那里去。”
ACTS|23|25|千夫长又写了公文，大略说：
ACTS|23|26|“ 克劳第．吕西亚 向 腓力斯 总督大人请安。
ACTS|23|27|这个人被 犹太 人拿住，快被杀害时，我得知他是 罗马 人，就带士兵下去，把他救了出来。
ACTS|23|28|因为我要知道他们告他的罪状，就带他下到他们的议会去。
ACTS|23|29|我查知他被告发是因他们律法上的争论，并没有什么该死或该监禁的罪名。
ACTS|23|30|后来有人把要害他的计谋告诉我，我立刻把他解到你那里去，又命令告他的人在你面前告他。 ”
ACTS|23|31|于是士兵照所命令他们的，连夜把 保罗 带到 安提帕底 。
ACTS|23|32|第二天，由骑兵护送 保罗 ，他们就回营楼去。
ACTS|23|33|骑兵来到 凯撒利亚 ，把公文呈给总督，就叫 保罗 站在他面前。
ACTS|23|34|总督读了公文，问 保罗 是哪一省的人；一知道他是 基利家 人，
ACTS|23|35|就说：“等告你的人来到，我才详细听你。”于是他命令把 保罗 拘留在 希律 的衙门里。
ACTS|24|1|过了五天， 亚拿尼亚 大祭司、几个长老和一个叫 帖土罗 的律师下来，向总督控告 保罗 。
ACTS|24|2|保罗 一被传来， 帖土罗 就开始控告他，说：“ 腓力斯 大人，我们因你得以享受国泰民安，并且这一国的弊病，因着你的远见得以改革。
ACTS|24|3|我们随时随地都满心感激不尽。
ACTS|24|4|为了不敢耽搁你太久，我只求你宽容一下，听我们说几句话。
ACTS|24|5|我们看这个人如同瘟疫一般，是鼓动普天下所有的 犹太 人作乱的人，又是 拿撒勒 教派里的一个头目。
ACTS|24|6|他甚至连圣殿也要污秽，我们就把他捉拿了。
ACTS|24|7|
ACTS|24|8|你自己审问他，就可以知道我们所控告他的一切事了。”
ACTS|24|9|众 犹太 人也随着控告他，说：“这些事情确是这样。”
ACTS|24|10|总督示意叫 保罗 说话， 保罗 就回答：“我知道你在本国作法官多年，所以我乐意为自己申辩。
ACTS|24|11|你查问就可以知道，从我上 耶路撒冷 去礼拜到今日不过十二天。
ACTS|24|12|他们并没有看见我在圣殿里跟人辩论，或在会堂里、在城里煽动群众。
ACTS|24|13|也不能对你证实他们现在所控告我的事。
ACTS|24|14|但有一件事我向你承认，就是我正按着他们所称为异端的道事奉我祖宗的上帝，又信合乎律法和先知书上所记载的一切。
ACTS|24|15|我对上帝存着这些人自己也接受的盼望，就是义人和不义的人都要复活。
ACTS|24|16|因此，我勉励自己，对上帝对人，时常存着无亏的良心。
ACTS|24|17|过了几年，我带着周济本国的捐项和供物上去。
ACTS|24|18|正献的时候，他们看见我在圣殿里已经洁净了，并没有聚众，也没有吵嚷，
ACTS|24|19|惟有几个从 亚细亚 来的 犹太 人—他们若有控告我的事，应当到你面前来告我。
ACTS|24|20|不然，让这些人自己说，他们看出我站在议会前的时间，有什么不对的地方。
ACTS|24|21|纵然有，也不过是为了一句话，就是我站在他们中间喊说：‘我今日在你们面前受审，是为了死人复活。’”
ACTS|24|22|腓力斯 本是详细认识这道，就拖延他们，说：“且等 吕西亚 千夫长下来，我再审判你们的案。”
ACTS|24|23|于是他下令百夫长看守 保罗 ，要从宽待他，不可拦阻他的亲友来供给他。
ACTS|24|24|过了几天， 腓力斯 和他夫人 犹太 女子 土西拉 一同来到，就叫 保罗 来，听他讲论信基督耶稣的事。
ACTS|24|25|保罗 讲论公义、节制和将来的审判， 腓力斯 害怕起来，就回答：“你暂且去吧！等我有机会时再来叫你。”
ACTS|24|26|腓力斯 又指望 保罗 送他银钱，所以屡次叫他来，和他谈论。
ACTS|24|27|过了两年， 波求．非斯都 接了 腓力斯 的任； 腓力斯 要讨 犹太 人的喜欢，就把 保罗 留在监里。
ACTS|25|1|非斯都 到省里上任，过了三天，就从 凯撒利亚 上 耶路撒冷 去。
ACTS|25|2|祭司长和 犹太 人的领袖向他控告 保罗 ；又央求他，
ACTS|25|3|向他求情要对付 保罗 ，把他提到 耶路撒冷 来，他们要在路上埋伏杀害他。
ACTS|25|4|非斯都 就回答：“ 保罗 押在 凯撒利亚 ，我自己快要往那里去。”
ACTS|25|5|他又说：“所以，你们中间有权的人与我一同下去，那人若有什么不是，就让他们控告他。”
ACTS|25|6|非斯都 在他们那里住了不超过八天或十天，就下 凯撒利亚 去；第二天开庭，下令把 保罗 提上来。
ACTS|25|7|保罗 来了，那些从 耶路撒冷 下来的 犹太 人周围站着，提出许多严重而不能证实的事控告他。
ACTS|25|8|保罗 申辩说：“无论 犹太 人的律法，或是圣殿，或是凯撒，我都没有干犯。”
ACTS|25|9|但 非斯都 要讨 犹太 人的喜欢，就回答 保罗 说：“你愿意上 耶路撒冷 去，在那里为这些事受我的审判吗？”
ACTS|25|10|保罗 说：“我现在站在凯撒的审判台前，这就是我应当受审的地方。我并没有对 犹太 人做过什么不对的事，这也是你明明知道的。
ACTS|25|11|我若做了不对的事，犯了什么该死的罪，就是死我也不辞。他们所控告我的事若都不实，就没有人能把我交给他们。我要向凯撒上诉。”
ACTS|25|12|非斯都 和议会商量了，就回答：“既然你要向凯撒上诉，你就到凯撒那里去吧。”
ACTS|25|13|过了些日子， 亚基帕 王和 百妮基 来到 凯撒利亚 ，拜访 非斯都 。
ACTS|25|14|他们在那里住了好些日子， 非斯都 将 保罗 的案件向王陈述，说：“这里有一个人，是 腓力斯 留在监里的。
ACTS|25|15|我在 耶路撒冷 的时候，祭司长和 犹太 的长老把他的事禀报了，要求定他的罪。
ACTS|25|16|我回覆他们，无论什么人，被告还没有和原告当面对质，没有机会为所控告的事申辩，就先定他罪的，这不是 罗马 人的规矩。
ACTS|25|17|及至他们都来到这里，我没有耽误，第二天就开庭，下令把那人提上来。
ACTS|25|18|控告他的人站起来告他，所控告的并没有任何我所预料的那等恶 事。
ACTS|25|19|不过，有几样辩论是有关他们自己敬鬼神的事，以及一个名叫耶稣的人，他已经死了， 保罗 却说他是活着的。
ACTS|25|20|我对这些事不知该怎样处理，所以问他是否愿意上 耶路撒冷 去，在那里为这些事接受审判。
ACTS|25|21|但 保罗 要求我留下他，要听皇上判断，我就下令把他留下，等我解他到凯撒那里去。”
ACTS|25|22|亚基帕 对 非斯都 说：“我也愿意亲自听听这个人。” 非斯都 说：“明天你就可以听他。”
ACTS|25|23|第二天， 亚基帕 和 百妮基 大张旗鼓而来，与众千夫长和城里的显要进了大厅。 非斯都 一声令下，就有人将 保罗 带进来。
ACTS|25|24|非斯都 说：“ 亚基帕 王和在这里的诸位，你们看这个人，他就是所有在 耶路撒冷 和这里的 犹太 人曾向我恳求呼叫，说不可容他再活着的。
ACTS|25|25|但我查明他并没有犯什么该死的罪，并且他自己也已向皇帝上诉了，所以我决定把他解去。
ACTS|25|26|论到这个人，我没有确实的事可以奏明主上。因此，我带他到你们面前，尤其到你 亚基帕 王面前，为要在查问之后有所呈奏。
ACTS|25|27|因为据我看，解送囚犯而不指明他的罪状是不合理的。”
ACTS|26|1|亚基帕 对 保罗 说：“准你为自己申诉。”于是 保罗 伸手辩护说：
ACTS|26|2|“ 亚基帕 王啊， 犹太 人所控告我的一切事，今日得以在你面前辩护，实为万幸。
ACTS|26|3|更庆幸的是你熟悉 犹太 人的规矩和他们的争论；所以，求你耐心听我。
ACTS|26|4|“我自幼为人如何，从起初在本国的同胞中，以及在 耶路撒冷 ，所有的 犹太 人都知道。
ACTS|26|5|他们若肯作见证，就知道我从起初是按着我们教中最严紧的教门作了法利赛人。
ACTS|26|6|现在我站在这里受审，是为了对上帝向我们祖宗的应许存着盼望。
ACTS|26|7|这应许，我们十二个支派，昼夜切切地事奉上帝，都指望得着。王啊，我正是因这指望被 犹太 人控告。
ACTS|26|8|上帝使死人复活，你们为什么判断为不可信呢？
ACTS|26|9|“从前我自己认为必须竭力反对 拿撒勒 人耶稣的名，
ACTS|26|10|我在 耶路撒冷 也曾这样做过；我不但从祭司长得了权柄，把许多圣徒收在监里，而且他们被杀，我也表示 赞成。
ACTS|26|11|在各会堂，我屡次用刑强迫他们说亵渎的话，我非常厌恶他们，甚至追逼他们，直到外邦的城镇。”
ACTS|26|12|“那时，我带着祭司长的权柄和命令往 大马士革 去。
ACTS|26|13|王啊！我在路上，中午的时候，看见从天上有一道光，比太阳还亮，四面照射着我和跟我同行的人。
ACTS|26|14|我们都仆倒在地，我就听见有声音用 希伯来 话对我说：‘ 扫罗 ！ 扫罗 ！你为什么迫害我？你用脚踢刺棒是自找苦吃的！’
ACTS|26|15|我说：‘主啊，你是谁？’主说：‘我就是你所迫害的耶稣。
ACTS|26|16|起来，站着，我向你显现的目的是要派你作仆役，为你所看见我 的事，和我将要指示你的事作见证人。
ACTS|26|17|我也要救你脱离百姓和外邦人的手。我差你到他们那里去，
ACTS|26|18|要开他们的眼睛，使他们从黑暗中转向光明，从撒但权下归向上帝；使他们因信我而得蒙赦罪，和一切成圣的人同得基业。’”
ACTS|26|19|“因此， 亚基帕 王啊！我没有违背那从天上来的异象；
ACTS|26|20|我先在 大马士革 ，后在 耶路撒冷 和 犹太 全地，以及外邦，劝勉他们应当悔改归向上帝，行事与悔改的心相称。
ACTS|26|21|为这缘故， 犹太 人在圣殿里拿住我，想要杀我。
ACTS|26|22|然而，我蒙上帝的帮助，直到今日还站立得稳，向尊贵的和卑微的作见证。我所讲的，并不外乎众先知和 摩西 所说将来必成的事，
ACTS|26|23|就是基督必须受害，并且首先从死人中复活，把亮光传给 犹太 人和外邦人。”
ACTS|26|24|保罗 这样申诉时， 非斯都 大声说：“ 保罗 ，你疯了！你的学问太大，反使你疯了！”
ACTS|26|25|保罗 说：“ 非斯都 大人，我不是疯了，我说的乃是真实和清醒的话。
ACTS|26|26|王也知道这些事，所以对王大胆直言，我深信这些事没有一件能向王隐瞒的，因为都不是在背地里做的。
ACTS|26|27|亚基帕 王啊，你信先知吗？我知道你是信的。”
ACTS|26|28|亚基帕 对 保罗 说：“你想稍微劝一劝就能说服我作基督徒了吗？”
ACTS|26|29|保罗 说：“无论少劝还是多劝，我向上帝所求的，不但你一个人，就是今天所有听我说话的人都要像我一样，只是不要有这些锁链。”
ACTS|26|30|于是，王和总督以及 百妮基 跟同坐的人都站起来，
ACTS|26|31|退到里面，彼此谈论说：“这个人并没有犯什么该死该监禁的罪。”
ACTS|26|32|亚基帕 对 非斯都 说：“这人若没有向凯撒上诉，早就被释放了。”
ACTS|27|1|既然 非斯都 决定要我们坐船往 意大利 去，就将 保罗 和别的囚犯交给御营里的一个名叫 犹流 的百夫长。
ACTS|27|2|有一只 亚大米田 的船要开往 亚细亚 沿海一带地方去，我们上了那船，就起航了；有 马其顿 的 帖撒罗尼迦 人 亚里达古 和我们同去。
ACTS|27|3|第二天，我们到了 西顿 。 犹流 宽待 保罗 ，准他往朋友那里去，受他们的照应。
ACTS|27|4|我们又从那里开船，因为遇到逆风，就贴着 塞浦路斯 的背风岸航行，
ACTS|27|5|渡过了 基利家 、 旁非利亚 一带的海面，就到了 吕家 的 每拉 。
ACTS|27|6|在那里，百夫长找到一只 亚历山大 的船要往 意大利 去，就叫我们上了那船。
ACTS|27|7|一连多日，船行得很慢，我们好不容易才来到 革尼土 的对面；又因被风拦阻，我们就贴着 克里特岛 背风岸，从 撒摩尼 对面航行。
ACTS|27|8|我们沿岸前进，十分艰难，来到一个名叫 佳澳 的地方，离那里不远有 拉西亚城 。
ACTS|27|9|航行的日子久了，已经过了禁食的节期，行船又危险， 保罗 就建议，
ACTS|27|10|对众人说：“诸位，我看这次航行，不但货物和船要受损伤，大遭破坏，连我们的性命也难保。”
ACTS|27|11|但百夫长信从船长和船主，不信 保罗 所说的。
ACTS|27|12|且因在这港口不适宜过冬，船上大多数的人都主张开船离开这地方，或者能到 非尼基 去过冬。 非尼基 是 克里特 的一个港口，一面朝西南，一面朝西北。
ACTS|27|13|当南风微微吹起时，他们以为对目的地已有了把握，就起锚，贴近 克里特 开去。
ACTS|27|14|过了不久，有一股叫“友拉革罗”的东北巨风从岛上扑来，
ACTS|27|15|船被风抓住，无法顶风航行，我们只好任它漂流。
ACTS|27|16|我们贴着一个叫 高大 的小岛的背风岸急航，好不容易才保住了救生艇。
ACTS|27|17|既然把救生艇拉上来，他们就用缆索捆绑船底，又恐怕在 赛耳底 浅滩上搁浅，就落了篷，任船漂流。
ACTS|27|18|我们被风浪逼得很急，第二天众人就把货物抛在海里。
ACTS|27|19|第三天，他们又亲手把船上的器具抛弃了。
ACTS|27|20|许多天都没有看到太阳和星辰，又有狂风大浪催逼，我们获救的指望都放弃了。
ACTS|27|21|众人已有好几天没有吃东西， 保罗 就出来站在他们中间，说：“诸位，你们本该听我的话不离开 克里特 岛，就不致遭到这样的损失和破坏。
ACTS|27|22|现在我劝你们放心，除了损失这条船，你们中间没有一人会丧失性命。
ACTS|27|23|因为昨夜，我所属所事奉的上帝的使者站在我旁边，
ACTS|27|24|说：‘ 保罗 ，不要害怕，你必定站在凯撒面前；并且上帝已把安全赐给与你同船的人了。’
ACTS|27|25|所以，诸位可以放心，我信上帝怎样对我说，事情也要怎样成就；
ACTS|27|26|只是我们必须在一个岛上搁浅。”
ACTS|27|27|到了第十四天夜间，船在 亚得里亚海 漂来漂去。约在半夜，水手以为渐近旱地，
ACTS|27|28|就去探测深浅，探得有十二丈 ；稍往前行，又探深浅，探得有九丈。
ACTS|27|29|恐怕我们撞到礁石，他们就从船尾抛下四个锚，盼望天亮。
ACTS|27|30|水手想弃船逃走，把救生艇缒下海里，假装要从船头抛锚的样子。
ACTS|27|31|保罗 对百夫长和士兵说：“这些人若不留在船上，你们就不能获救。”
ACTS|27|32|于是士兵砍断救生艇的绳子，由它漂去。
ACTS|27|33|天快亮的时候， 保罗 劝众人都用餐，说：“你们一直捱饿等候，不吃什么，已经十四天了。
ACTS|27|34|所以我劝你们吃点东西，这是关乎你们获救的，因为你们各人连一根头发也不至于掉落。”
ACTS|27|35|保罗 说了这话，就拿起饼来，在众人面前祝谢了上帝，然后擘开来吃。
ACTS|27|36|于是他们都放心，就吃了。
ACTS|27|37|我们在船上的共有二百七十六个人。
ACTS|27|38|他们吃饱了，为要使船轻一点，就把船上的麦子抛到海里。
ACTS|27|39|天亮的时候，他们不认得那地方，只见一个有岸可登的海湾，就想法子看能不能把船靠岸。
ACTS|27|40|于是他们砍断缆索，把锚丢到海里，同时也松开舵绳，拉起头篷，顺风向着岸行去。
ACTS|27|41|但碰到两水夹流的地方，就搁了浅，船头胶住不动，船尾被浪的猛力冲坏了 。
ACTS|27|42|士兵的意思要把囚犯都杀了，免得有游水脱逃的。
ACTS|27|43|但百夫长要救 保罗 ，不准他们任意而行，就吩咐会游水的，跳下水去，先上岸；
ACTS|27|44|其余的人则用板子或船的碎片上岸。这样，众人都获救，上了岸。
ACTS|28|1|我们既已获救，才知道那岛名叫 马耳他 。
ACTS|28|2|当地人非常友善地接待我们；因为正在下雨，天气又冷，他们就生了火欢迎我们众人。
ACTS|28|3|那时， 保罗 拾起一捆柴，放在火中，有一条毒蛇，因为热的缘故钻了出来，缠住他的手。
ACTS|28|4|当地的人看见那毒蛇悬在他手上，就彼此说：“这人必是个凶手，虽然他从海里获救，天理仍不容他活着。”
ACTS|28|5|保罗 竟把那毒蛇甩在火里，并没有受伤。
ACTS|28|6|当地的人想他快要肿起来，或是忽然倒下死了，但等了好久，见他没有什么异样，就转念说他是个神明。
ACTS|28|7|离那地方不远有一些田产，是岛长 部百流 的。他接纳我们，尽情款待了我们三日。
ACTS|28|8|当时， 部百流 的父亲卧病不起，患了热病和痢疾。 保罗 进去见他，为他祷告按手，治好了他。
ACTS|28|9|从此，岛上其余的病人也都来，得了医治。
ACTS|28|10|他们又多方面尊敬我们，到了开船的时候，又把我们所需用的东西送到船上。
ACTS|28|11|过了三个月，我们上了 亚历山大 的船起航。这船以“ 宙斯 双子”为记，是在那海岛过冬的。
ACTS|28|12|我们到了 叙拉古 ，停泊了三日；
ACTS|28|13|又从那里起锚开船， 来到 利基翁 。过了一天，起了南风，第二天就来到 部丢利 。
ACTS|28|14|我们在那里遇见一些弟兄，他们请我们同住了七天。就这样，我们来到 罗马 。
ACTS|28|15|那里的弟兄们一听见我们的消息，就到 亚比乌 市和 三馆 来迎接我们。 保罗 见了他们，就感谢上帝，越发壮胆。
ACTS|28|16|我们进了 罗马城 ， 保罗 蒙准和那个看守他的兵另住在一处。
ACTS|28|17|过了三天， 保罗 请当地 犹太 人的领袖来。他们来了， 保罗 对他们说：“诸位弟兄，虽然我没有做什么事干犯本国的百姓和我们祖宗的规矩，却在 耶路撒冷 被囚禁，交在 罗马 人的手里。
ACTS|28|18|他们审问了我，有意要释放我，因为在我身上并没有该死的罪状。
ACTS|28|19|但 犹太 人反对，我不得已只好上诉于凯撒，并不是有什么事要控告我本国的百姓。
ACTS|28|20|为这缘故，我请你们来见我当面谈话，我原是为 以色列 人所指望的那位才被这铁链捆绑的。”
ACTS|28|21|他们对他说：“我们并没有接到从 犹太 寄来有关于你的信，也没有弟兄到这里来向我们报告，或说你有什么不好的地方。
ACTS|28|22|但我们愿意听听你的意见，因为我们知道这教门是到处遭人反对的。”
ACTS|28|23|他们和 保罗 约定了日子，就有许多人到他的住处来。 保罗 从早到晚向他们讲解这事，为上帝的国作证，并引 摩西 的律法和先知的书劝导他们信从耶稣。
ACTS|28|24|他所说的话，有的信，有的不信。
ACTS|28|25|他们间彼此不合，就分散了；未散以先， 保罗 说了一句话：“圣灵藉 以赛亚 先知向你们祖宗所说的话是对的。
ACTS|28|26|他说： ‘你去对这百姓说： 你们听了又听，却不明白； 看了又看，却看不清。
ACTS|28|27|因为这百姓的心麻木， 耳朵塞着， 眼睛闭着， 免得眼睛看见， 耳朵听见， 心里明白，回转过来， 我会医治他们。’
ACTS|28|28|所以，你们当知道，上帝这救恩已经传给外邦人；他们会听的。”
ACTS|28|29|
ACTS|28|30|保罗 在自己所租的房子里住了足足两年。凡来见他的人，他都接待，
ACTS|28|31|放胆传讲上帝的国，并教导主耶稣基督的事，没有人禁止。
ROM|1|1|基督耶稣的仆人 保罗 ，蒙召为使徒，奉派传上帝的福音。
ROM|1|2|这福音是上帝从前藉众先知，在圣经上所应许的。
ROM|1|3|论到他儿子－我主耶稣基督，按肉体说，是从 大卫 后裔生的；按神圣的灵说，因从死人中复活，用大能显明他是上帝的儿子。
ROM|1|4|
ROM|1|5|我们从他蒙恩受了使徒的职分，为他的名在万国中使人因信而顺服，
ROM|1|6|其中也有你们这蒙召属耶稣基督的人。
ROM|1|7|我写信给你们在 罗马 、为上帝所爱、蒙召作圣徒的众人。愿恩惠、平安 从我们的父上帝和主耶稣基督归给你们！
ROM|1|8|首先，我靠着耶稣基督，为你们众人感谢我的上帝，因你们的信德传遍了天下。
ROM|1|9|我在他儿子的福音上，用心灵所事奉的上帝可以见证，我怎样不住地提到你们，
ROM|1|10|在我的祷告中常常恳求，或许照上帝的旨意，最终我能毫无阻碍地往你们那里去。
ROM|1|11|因为我迫切地想见你们，要把一些属灵的恩赐分给你们，使你们得以坚固，
ROM|1|12|也可以说，我在你们中间，因你我彼此的信心而同得安慰。
ROM|1|13|弟兄们，我不愿意你们不知道，我屡次计划往你们那里去，要在你们中间得些果子，如同在其余的外邦人中一样，只是到如今仍有拦阻。
ROM|1|14|无论是 希腊 人、未开化的人、聪明人、愚拙人，我都欠他们的债，
ROM|1|15|所以愿意尽我的力量把福音也传给你们在 罗马 的人。
ROM|1|16|我不以福音为耻；这福音本是上帝的大能，要救一切相信的，先是 犹太 人，后是 希腊 人。
ROM|1|17|因为上帝的义正在这福音上显明出来；这义是本于信，以至于信。如经上所记：“义人必因信得生。”
ROM|1|18|原来，上帝的愤怒从天上显明在一切不虔不义的人身上，就是那些行不义压制真理的人。
ROM|1|19|上帝的事情，人所能知道的，原显明在人心里，因为上帝已经向他们显明。
ROM|1|20|自从造天地以来，上帝的永能和神性是明明可知的，虽然眼不能见，但藉着所造之物就可以了解看见，叫人无可推诿。
ROM|1|21|因为，他们虽然知道上帝，却不把他当作上帝荣耀他，也不感谢他。他们的思想变为虚妄，无知的心昏暗了。
ROM|1|22|他们自以为聪明，反成了愚昧，
ROM|1|23|将不能朽坏之上帝的荣耀变为偶像，仿照必朽坏的人、飞禽、走兽、爬虫的形像。
ROM|1|24|所以，上帝任凭他们随着心里的情欲行污秽的事，以致彼此羞辱自己的身体。
ROM|1|25|他们将上帝的真实变为虚谎，去敬拜事奉受造之物，不敬奉那造物的主—主是可称颂的，直到永远。阿们！
ROM|1|26|因此，上帝任凭他们放纵可羞耻的情欲。他们的女人把自然的关系变成违反自然的；
ROM|1|27|男人也是如此，放弃了和女人自然的关系，欲火攻心，男的和男的彼此贪恋，行可耻的事，就在自己身上受这逆性行为当得的报应。
ROM|1|28|他们既然故意不认识上帝，上帝就任凭他们存扭曲的心，做那些不该做的事，
ROM|1|29|装满了各样不义 、邪恶、贪婪、恶毒，满心是嫉妒、凶杀、纷争、诡诈、毒恨，又是毁谤的、
ROM|1|30|说人坏话的、怨恨上帝的 、侮辱人的、狂傲的、自夸的、制造是非的、忤逆父母的、
ROM|1|31|顽梗不化的、言而无信的、无情无义的、不怜悯人的。
ROM|1|32|他们虽知道上帝判定做这样事的人是该死的，然而他们不但自己去做，还赞同别人去做。
ROM|2|1|所以，你这评断人的人哪，无论你是谁，都无可推诿。你在什么事上评断人，就在什么事上定自己的罪。因你这评断人的，自己所做的却和别人一样。
ROM|2|2|我们知道这样做的人，上帝必公平地审判他。
ROM|2|3|你这个人哪，你评断做这样事的人，自己所做的却和别人一样，你以为能逃脱上帝的审判吗？
ROM|2|4|还是你藐视他丰富的恩慈、宽容、忍耐，不知道他的恩慈是领你悔改吗？
ROM|2|5|你竟放任你刚硬不悔改的心，为自己累积愤怒！在愤怒的日子，上帝公义的审判要显示出来。
ROM|2|6|他要照各人的行为报应各人。
ROM|2|7|凡恒心行善，寻求荣耀、尊贵和不能朽坏的，就有永生报偿他们；
ROM|2|8|但是那些自私自利、不顺从真理、反顺从不义的人，就有恼恨、愤怒报应他们。
ROM|2|9|他要把患难、困苦加给一切作恶的人，先是 犹太 人，后是 希腊 人；
ROM|2|10|却把荣耀、尊贵、平安加给一切行善的人，先是 犹太 人，后是 希腊 人。
ROM|2|11|因为上帝不偏待人。
ROM|2|12|凡在律法之外犯了罪的，将在律法之外灭亡；凡在律法之内犯了罪的，将按律法受审判。
ROM|2|13|原来在上帝面前，不是听律法的为义，而是行律法的称义。
ROM|2|14|没有律法的外邦人若顺着本性行律法上的事，他们虽然没有律法，自己就是自己的律法。
ROM|2|15|他们显明律法的功用刻在他们心里，他们的良心一同作证—他们的内心挣扎，有时自责，有时为自己辩护。
ROM|2|16|在那日，上帝要藉着基督耶稣 ，按照我所传的福音，审判人隐藏的事。
ROM|2|17|但是你，你既自称为 犹太 人，倚靠律法，以上帝夸口，
ROM|2|18|知道上帝的旨意，从律法受了教导而能分辨是非；
ROM|2|19|你既深信自己是给盲人领路的，是在黑暗中人的光，
ROM|2|20|是无知的人的师傅，是小孩子的老师，体现了律法中的知识和真理；
ROM|2|21|那么，你这教导别人的，还不教导自己吗？你这宣讲不可偷窃的，自己还偷窃吗？
ROM|2|22|你这说不可奸淫的，自己还奸淫吗？你这厌恶偶像的，自己还抢劫庙中之物吗？
ROM|2|23|你这以律法夸口的，自己倒违犯律法，羞辱上帝！
ROM|2|24|上帝的名在外邦人中因你们受了亵渎，正如经上所记的。
ROM|2|25|你若遵行律法，割礼固然于你有益；若违犯律法，你的割礼就算不得割礼。
ROM|2|26|所以，那未受割礼的，若遵守律法的要求，他虽然未受割礼，岂不算是受了割礼吗？
ROM|2|27|而且那本来未受割礼的，若能全守律法，岂不是要审判你这有仪文和割礼，竟违犯律法的人吗？
ROM|2|28|因为外表是 犹太 人的不是真 犹太 人；外表肉身的割礼也不是真割礼。
ROM|2|29|惟有内心作 犹太 人的才是真 犹太 人，真割礼也是心里的，在乎圣灵 ，不在乎仪文。这样的人所受的称赞不是从人来的，而是从上帝来的。
ROM|3|1|这样说来， 犹太 人有什么比别人强呢？割礼有什么益处呢？
ROM|3|2|很多，各方面都有。首先，上帝的圣言交托他们。
ROM|3|3|即使有不信的，这又何妨呢？难道他们的不信就废掉上帝的信实吗？
ROM|3|4|绝对不会！不如说，上帝是真实的，而人都是虚谎的。如经上所记： “以致你责备的时候显为公义； 你被指控的时候一定胜诉。”
ROM|3|5|我姑且照着人的看法来说，我们的不义若显出上帝的义来，我们要怎么说呢？上帝降怒是他不义吗？
ROM|3|6|绝对不是！若是这样，上帝怎能审判世界呢？
ROM|3|7|若上帝的真实因我的虚谎越发显出他的荣耀，为什么我还像罪人一样受审判呢？
ROM|3|8|为什么不说，我们可以作恶以成善呢？有人毁谤我们，说我们讲过这话；这等人被定罪是应该的。
ROM|3|9|那又怎么样呢？我们比他们强吗？绝不是！因我们已经指证： 犹太 人和 希腊 人都在罪恶之下。
ROM|3|10|就如经上所记： “没有义人，连一个也没有。
ROM|3|11|没有明白的， 没有寻求上帝的。
ROM|3|12|人人偏离正路，一同走向败坏。 没有行善的，连一个也没有 。
ROM|3|13|他们的喉咙是敞开的坟墓； 他们的舌头玩弄诡诈。 他们的嘴唇里有毒蛇的毒液，
ROM|3|14|满口是咒骂苦毒。
ROM|3|15|他们的脚为杀人流血飞跑；
ROM|3|16|他们的路留下毁坏和灾难。
ROM|3|17|和平的路，他们不认识；
ROM|3|18|他们眼中不怕上帝。”
ROM|3|19|我们知道律法所说的话都是对律法之下的人说的，好塞住各人的口，使普世的人都伏在上帝的审判之下。
ROM|3|20|所以，凡血肉之躯没有一个能因律法的行为而在上帝面前称义，因为律法本是要人认识罪。
ROM|3|21|但如今，上帝的义在律法之外已经显明出来，有律法和先知为证：
ROM|3|22|就是上帝的义，因信耶稣基督 加给一切信的人。这并没有分别，
ROM|3|23|因为世人都犯了罪，亏缺了上帝的荣耀，
ROM|3|24|如今却蒙上帝的恩典，藉着在基督耶稣里的救赎，就白白地得称为义。
ROM|3|25|上帝设立耶稣作赎罪祭，是凭耶稣的血，藉着信，要显明上帝的义；因为他用忍耐的心宽容人先前所犯的罪，好使今时显明他的义，让人知道他自己为义，也称信耶稣的人为义 。
ROM|3|26|
ROM|3|27|既是这样，哪里可夸口呢？没有可夸的。是藉什么法呢？功德吗？不是！是藉信主之法。
ROM|3|28|所以我们认定，人称义是因着信，不在于律法的行为。
ROM|3|29|难道上帝只是 犹太 人的吗？不也是外邦人的吗？是的，他也是外邦人的上帝。
ROM|3|30|既然上帝是一位，他就要本于信称那受割礼的为义，也要藉着信称那未受割礼的为义。
ROM|3|31|这样，我们藉着信废了律法吗？绝对不是！更是巩固律法。
ROM|4|1|这样，那按肉体作我们祖宗的 亚伯拉罕 ，我们要怎么说呢？
ROM|4|2|倘若 亚伯拉罕 是因行为称义，他就有可夸的，但是在上帝面前他一无可夸。
ROM|4|3|经上说什么呢？“ 亚伯拉罕 信了上帝，这就算他为义。”
ROM|4|4|做工的得工资不算是恩典，而是应得的；
ROM|4|5|但那不做工的，只信那位称不敬虔之人为义的，他的信就算为义。
ROM|4|6|正如 大卫 称那在行为之外蒙上帝算为义的人是有福的：
ROM|4|7|“过犯得赦免，罪恶蒙遮盖的人有福了！
ROM|4|8|主不算为有罪的，这样的人有福了！”
ROM|4|9|如此看来，这福只加给那受割礼的人吗？不也加给那未受割礼的人吗？我们说，因着信，就算 亚伯拉罕 为义。
ROM|4|10|那么，这是怎么算的呢？是在他受割礼的时候呢？还是在他未受割礼的时候呢？不是在受割礼的时候，而是在未受割礼的时候。
ROM|4|11|并且，他受了割礼的记号，作他未受割礼的时候因信称义的印证，为使他作一切未受割礼而信之人的父，使他们也算为义，
ROM|4|12|也使他作受割礼之人的父，就是那些不但受割礼，而且跟随我们的祖宗 亚伯拉罕 未受割礼而信的足迹的人。
ROM|4|13|因为上帝给 亚伯拉罕 和他后裔承受世界的应许不是藉着律法，而是藉着信而得的义。
ROM|4|14|若是属于律法的人才是后嗣，信就落空了，应许也就失效了。
ROM|4|15|因为律法是惹动愤怒的，哪里没有律法，哪里就没有过犯。
ROM|4|16|所以，人作后嗣是出于信，因此就属乎恩，以致应许保证归给所有的后裔，不但归给那属于律法的，也归给那效法 亚伯拉罕 之信的人。 亚伯拉罕 所信的是那叫死人复活、使无变为有的上帝，在这位上帝面前 亚伯拉罕 成为我们众人的父，如经上所记：“我已经立你作多国之父。”
ROM|4|17|
ROM|4|18|他在没有盼望的时候，仍存着盼望来相信，就得以作多国之父，正如先前所说：“你的后裔将要如此。”
ROM|4|19|他将近百岁的时候，虽然想到 自己的身体如同已死， 撒拉 也不可能生育，他的信心还是不软弱，
ROM|4|20|仍仰望上帝的应许，总没有因不信而起疑惑，反倒因信而刚强，将荣耀归给上帝，
ROM|4|21|且满心相信上帝所应许的必能成就。
ROM|4|22|所以这也 就算他为义。
ROM|4|23|“算他为义”这句话不是单为他写的，
ROM|4|24|也是为我们将来得算为义的人写的，就是为我们这些信上帝使我们的主耶稣从死人中复活的人写的。
ROM|4|25|耶稣被出卖，是为我们的过犯；他复活，是为使我们称义。
ROM|5|1|所以，我们既因信称义，就藉着我们的主耶稣基督得以与上帝和好。
ROM|5|2|我们又藉着他，因信 得以进入现在所站立的这恩典中，并且欢欢喜喜盼望上帝的荣耀。
ROM|5|3|不但如此，就是在患难中也是欢欢喜喜的，因为知道患难生忍耐，
ROM|5|4|忍耐生老练，老练生盼望，
ROM|5|5|盼望不至于落空，因为上帝的爱，已藉着所赐给我们的圣灵，浇灌在我们心里。
ROM|5|6|我们还软弱的时候，基督就在特定的时刻为不敬虔之人死。
ROM|5|7|为义人死，是少有的；为仁人死，或者有敢做的。
ROM|5|8|惟有基督在我们还作罪人的时候为我们死，上帝的爱就在此向我们显明了。
ROM|5|9|现在我们既靠着他的血称义，就更要藉着他得救，免受上帝的愤怒。
ROM|5|10|因为我们作仇敌的时候，尚且藉着上帝儿子的死得以与上帝和好，既已和好，就更要因他的生得救了。
ROM|5|11|不但如此，我们既藉着我们的主耶稣基督得以与上帝和好，也就藉着他以上帝为乐。
ROM|5|12|为此，正如罪是从一人进入世界，死又从罪而来，于是死就临到所有的人，因为人人都犯了罪。
ROM|5|13|没有律法之前，罪已经在世上，但没有律法，罪也不算罪。
ROM|5|14|然而，从 亚当 到 摩西 ，死就掌了权，连那些不与 亚当 犯一样罪过的，也在死的权下。 亚当 是那以后要来之人的预像。
ROM|5|15|但是过犯不如恩赐，若因一人的过犯，众人都死了，那么，上帝的恩典，与那因耶稣基督一人而来的恩典中的赏赐，岂不加倍地临到众人吗？
ROM|5|16|因一人犯罪而来的后果，也不如赏赐，原来审判是由一人而定罪，恩赐乃是由许多过犯而称义。
ROM|5|17|若因一人的过犯，死就因这一人掌权，那些受洪恩又蒙所赐之义的，岂不更要因耶稣基督一人在他们生命中掌权吗？
ROM|5|18|这样看来，因一次的过犯，所有的人都被定罪；照样，因一次的义行，所有的人也就被称义而得生命了。
ROM|5|19|因一人的悖逆，众人成为罪人；照样，因一人的顺从，众人也成为义了。
ROM|5|20|而且加添了律法，使得过犯增加，只是罪在哪里增加，恩典就在哪里越发丰盛了。
ROM|5|21|所以，正如罪藉着死掌权；照样，恩典也藉着义掌权，使人因我们的主耶稣基督得永生。
ROM|6|1|这样，我们要怎么说呢？我们可以仍在罪中使恩典增多吗？
ROM|6|2|绝对不可！我们向罪死了的人，岂可仍在罪中活着呢？
ROM|6|3|难道你们不知道，我们这受洗归入基督耶稣的人，就是受洗归入他的死吗？
ROM|6|4|所以，我们藉着洗礼归入死，和他一同埋葬，是要我们行事为人都有新生的样子，像基督藉着父的荣耀从死人中复活一样。
ROM|6|5|我们若与他合一，经历与他一样的死，也将经历与他一样的复活。
ROM|6|6|我们知道，我们的旧人和他同钉十字架，使罪身灭绝，叫我们不再作罪的奴隶，
ROM|6|7|因为已死的人是脱离了罪。
ROM|6|8|我们若与基督同死，我们信也必与他同活，
ROM|6|9|因为知道基督既从死人中复活，就不再死，死也不再作他的主了。
ROM|6|10|他死了，是对罪死，只这一次；他活，是对上帝活着。
ROM|6|11|这样，你们也要看自己对罪是死的，在基督耶稣里对上帝却是活的。
ROM|6|12|所以，不要让罪在你们必死的身上掌权，使你们顺从身体的私欲。
ROM|6|13|也不要把你们的肢体献给罪作不义的工具，倒要像从死人中活着的人，把自己献给上帝，并把你们的肢体献给上帝作义的工具。
ROM|6|14|罪必不能作你们的主，因你们不在律法之下，而是在恩典之下。
ROM|6|15|那又怎么样呢？我们在恩典之下，不在律法之下，就可以犯罪吗？绝对不可！
ROM|6|16|难道你们不知道，你们献自己作奴仆，顺从谁就作谁的奴仆吗？或作罪的奴隶，以至于死；或作顺服的奴仆，以至于成义。
ROM|6|17|感谢上帝！因为你们从前虽然作罪的奴隶，现在却从心里顺服了所传给你们教导的典范。
ROM|6|18|你们既从罪里得了释放，就作了义的奴仆。
ROM|6|19|我因你们肉体的软弱，就以人的观点来说。你们从前怎样把肢体献给不洁不法作奴隶，以至于不法；现在也要照样将肢体献给义作奴仆，以至于成圣。
ROM|6|20|因为你们作罪的奴隶时，不被义所约束。
ROM|6|21|那么，你们现在所看为羞耻的事，当时有什么果子呢？那些事的结局就是死。
ROM|6|22|但如今，你们既从罪里得了释放，作了上帝的奴仆，就结出果子，以至于成圣，那结局就是永生。
ROM|6|23|因为罪的工价乃是死；惟有上帝的恩赐，在我们的主基督耶稣里，乃是永生。
ROM|7|1|弟兄们，我对你们这些明白律法的人说，你们岂不知道律法约束人是在他活着的时候吗？
ROM|7|2|就如女人有了丈夫，丈夫还活着，她就被律法约束；丈夫若死了，她就从丈夫的律法中解脱了。
ROM|7|3|所以丈夫还活着，她若跟了别的男人，就叫淫妇；丈夫若死了，她就脱离了律法，虽然跟了别的男人，也不是淫妇。
ROM|7|4|我的弟兄们，这样说来，你们藉着基督的身体对律法也是死了，使你们归于另一位，就是归于那从死人中复活的，为要使我们结果子给上帝。
ROM|7|5|因为我们属肉体的时候，那因律法而生犯罪的欲望在我们肢体中发动，以致结出死亡的果子。
ROM|7|6|但如今，我们既然在捆绑我们的律法上死了，就从律法中解脱，使我们服侍主，要按着圣灵 的新样，不按着仪文的旧样。
ROM|7|7|这样，我们要怎么说呢？律法是罪吗？绝对不是！但是，若不是藉着律法，我就不知何为罪；若不是律法说“不可贪心”，我就不知何为贪心。
ROM|7|8|然而，罪趁着机会，藉着诫命，使各样的贪心在我里头发动，因为没有律法，罪是死的。
ROM|7|9|以前没有律法的时候，我是活的；但是诫命来到，罪活起来，
ROM|7|10|我就死了。那本该叫人活的诫命反而叫我死。
ROM|7|11|因为罪趁着机会，藉着诫命诱惑我，并且藉着诫命杀了我。
ROM|7|12|这样看来，律法是圣的，诫命也是圣的、义的、善的。
ROM|7|13|那么，那善的是叫我死吗？绝对不是！叫我死的是罪。罪藉着那善的叫我死，为要显出这真是罪，以致罪藉着诫命更显出是恶极了。
ROM|7|14|我们原知道律法是属灵的，我却是属肉体的，是已经卖给罪了。
ROM|7|15|因为我所做的，我自己不明白。我所愿意的，我并不做；我所恨恶的，我反而去做。
ROM|7|16|如果我所做的是我所不愿意的，我得承认律法是善的。
ROM|7|17|事实上，这不是我做的，而是住在我里面的罪做的。
ROM|7|18|我也知道，住在我里面的，就是我肉体之中，没有善。因为立志为善由得我，只是行出来由不得我。
ROM|7|19|我所愿意的善，我不去做；我所不愿意的恶，我反而去做。
ROM|7|20|如果我去做我不愿意做的，就不是我做的，而是住在我里面的罪做的。
ROM|7|21|我觉得有个律，就是我愿意行善的时候，就有恶缠着我。
ROM|7|22|因为，按着我里面的人，我喜欢上帝的律，
ROM|7|23|但我看出肢体中另有个律和我内心的律交战，把我掳去，使我附从那肢体中罪的律。
ROM|7|24|我真苦啊！谁能救我脱离这必死的身体呢？
ROM|7|25|感谢上帝，靠着我们的主耶稣基督就能！这样看来，一方面，我内心顺服上帝的律，另一方面，肉体却顺服罪的律了。
ROM|8|1|如今，那些在基督耶稣里的人就不被定罪了。
ROM|8|2|因为赐生命的圣灵的律，在基督耶稣里从罪和死的律中把你释放出来。
ROM|8|3|律法既因肉体软弱而无能为力，上帝就差遣自己的儿子成为罪身的样子，为了对付罪 ，在肉体中定了罪，
ROM|8|4|为要使律法要求的义，实现在我们这不随从肉体、只随从圣灵去行的人身上。
ROM|8|5|因为，随从肉体的人体贴肉体的事；随从圣灵的人体贴圣灵的事。
ROM|8|6|体贴肉体就是死；体贴圣灵就是生命和平安 。
ROM|8|7|因为体贴肉体就是与上帝为敌，对上帝的律法不顺服，事实上也无法顺服。
ROM|8|8|属肉体的人无法使上帝喜悦。
ROM|8|9|如果上帝的灵住在你们里面，你们就不属肉体，而是属圣灵了。人若没有基督的灵，就不是属基督的。
ROM|8|10|基督若在你们里面，身体就因罪而死，灵却因义而活。
ROM|8|11|然而，使耶稣从死人中复活的上帝的灵若住在你们里面，那使基督从死人中复活的，也必藉着住在你们里面的圣灵使你们必死的身体又活过来。
ROM|8|12|弟兄们，这样看来，我们不是欠肉体的债去顺从肉体而活。
ROM|8|13|你们若顺从肉体活着，必定会死；若靠着圣灵把身体的恶行处死，就必存活。
ROM|8|14|因为凡被上帝的灵引导的都是上帝的儿子。
ROM|8|15|你们所领受的不是奴仆的灵，仍旧害怕；所领受的是儿子名分的灵，因此我们呼叫：“阿爸，父！”
ROM|8|16|圣灵自己与我们的灵一同见证我们是上帝的儿女。
ROM|8|17|若是儿女，就是后嗣，是上帝的后嗣，和基督同作后嗣。如果我们和他一同受苦，是要我们和他一同得荣耀。
ROM|8|18|我认为，现在的苦楚，若比起将来要显示给我们的荣耀，是不足介意的。
ROM|8|19|受造之物切望等候上帝的众子显出来。
ROM|8|20|因为受造之物屈服在虚空之下，不是自己愿意，而是因那使它屈服的叫他如此。但受造之物仍然指望从败坏的辖制下得释放，得享上帝儿女荣耀的自由。
ROM|8|21|
ROM|8|22|我们知道，一切受造之物一同呻吟，一同忍受阵痛，直到如今。
ROM|8|23|不但如此，就是我们这有圣灵作初熟果子的，也是自己内心呻吟，等候得着儿子的名分，就是我们的身体得救赎。
ROM|8|24|我们得救是在于盼望；可是看得见的盼望就不是盼望。谁还去盼望他所看得见的呢？
ROM|8|25|但我们若盼望那看不见的，我们就耐心等候。
ROM|8|26|同样，我们的软弱有圣灵帮助。我们本不知道当怎样祷告，但是圣灵亲自用无可言喻的叹息替我们祈求。
ROM|8|27|那鉴察人心的知道圣灵所体贴的，因为圣灵照着上帝的旨意替圣徒祈求。
ROM|8|28|我们知道，万事 都互相效力，叫爱上帝的人得益处，就是按他旨意被召的人。
ROM|8|29|因为他所预知的人，他也预定他们效法他儿子的榜样，使他儿子在许多弟兄中作长子 。
ROM|8|30|他所预定的人，他又召他们来；所召来的人，他又称他们为义；所称为义的人，他又叫他们得荣耀。
ROM|8|31|既是这样，我们对这些事还要怎么说呢？上帝若帮助我们，谁能抵挡我们呢？
ROM|8|32|上帝既不顾惜自己的儿子，为我们众人舍了他，岂不也把万物和他一同白白地赐给我们吗？
ROM|8|33|谁能控告上帝所拣选的人呢？有上帝称他们为义了。
ROM|8|34|谁能定他们的罪呢？有基督耶稣 已经死了，而且复活了，现今在上帝的右边，也替我们祈求。
ROM|8|35|谁能使我们与基督的爱隔绝呢？难道是患难吗？是困苦吗？是迫害吗？是饥饿吗？是赤身露体吗？是危险吗？是刀剑吗？
ROM|8|36|如经上所记： “我们为你的缘故终日被杀； 人看我们如将宰的羊。”
ROM|8|37|然而，靠着爱我们的主，在这一切的事上，我们已经得胜有余了。
ROM|8|38|因为我深信，无论是死，是活，是天使，是掌权的，是有权能的 ，是现在的事，是将来的事，
ROM|8|39|是高处的，是深处的，是别的受造之物，都不能使我们与上帝的爱隔绝，这爱是在我们的主基督耶稣里的。
ROM|9|1|我在基督里说真话，不说谎话；我的良心被圣灵感动为我作证。
ROM|9|2|我非常忧愁，心里时常伤痛。
ROM|9|3|为我弟兄，我骨肉之亲，就是自己被诅咒，与基督分离，我也愿意。
ROM|9|4|他们是 以色列 人，那儿子的名分、荣耀、诸约、律法的颁布、敬拜的礼仪、应许都是给他们的。
ROM|9|5|列祖是他们的，基督按肉体说也是从他们出来的。愿在万有之上的上帝被称颂，直到永远 。阿们！
ROM|9|6|这不是说上帝的话落了空。因为从 以色列 生的不都是 以色列 人，
ROM|9|7|也不因为是 亚伯拉罕 的后裔就都是他的儿女；惟独“从 以撒 生的才要称为你的后裔。”
ROM|9|8|这就是说，肉身所生的儿女不是上帝的儿女，惟独那应许的儿女才算是后裔。
ROM|9|9|因为所应许的话是这样：“到明年这时候我要来， 撒拉 必会生一个儿子。”
ROM|9|10|不但如此， 利百加 也是这样。她从一个人，就是从我们的祖宗 以撒 怀了孕。
ROM|9|11|双胞胎还没有生下来，善恶还没有行出来，为要贯彻上帝拣选人的旨意，
ROM|9|12|不是凭着人的行为，而是凭着那呼召人的，上帝就对 利百加 说：“将来，大的要服侍小的。”
ROM|9|13|正如经上所记：“ 雅各 是我所爱的； 以扫 是我所恶的。”
ROM|9|14|这样，我们要怎么说呢？难道上帝有什么不义吗？绝对没有！
ROM|9|15|因他对 摩西 说： “我要怜悯谁就怜悯谁， 要恩待谁就恩待谁。”
ROM|9|16|由此看来，这不靠人的意愿，也不靠人的努力，只靠上帝的怜悯。
ROM|9|17|因为经上有话对法老说：“我将你兴起来，特要在你身上彰显我的权能，为要使我的名传遍全地。”
ROM|9|18|由此看来，上帝要怜悯谁就怜悯谁，要使谁刚硬就使谁刚硬。
ROM|9|19|这样，你会对我说：“那么，他为什么还指责人呢？有谁能抗拒他的旨意呢？”
ROM|9|20|你这个人哪，你是谁，竟敢向上帝顶嘴呢？受造之物岂会对造他的说：“你为什么把我造成这样呢？”
ROM|9|21|难道陶匠没有权从一团泥里拿一块做成贵重的器皿，又拿一块做成卑贱的器皿吗？
ROM|9|22|倘若上帝要显明他的愤怒，彰显他的权能，难道不可多多忍耐宽容那应受愤怒、预备遭毁灭的器皿吗？
ROM|9|23|这是为了要把他丰盛的荣耀彰显在那蒙怜悯、早预备得荣耀的器皿上。
ROM|9|24|这器皿也就是我们这些蒙上帝所召的，不但是从 犹太 人中，也是从外邦人中召来的。
ROM|9|25|正如上帝在《何西阿书》上说： “那本来不是我子民的， 我要称为‘我的子民’； 本来不是蒙爱的， 我要称为‘蒙爱的’。
ROM|9|26|从前在什么地方对他们说： 你们不是我的子民， 将来就在那里称他们为‘永生上帝的儿子’。”
ROM|9|27|关于 以色列 人， 以赛亚 喊着：“虽然 以色列 人多如海沙，得救的将是剩下的余数，
ROM|9|28|因为主要在地上施行他的话，彻底而又迅速。”
ROM|9|29|又如 以赛亚 先前说过： “若不是万军之主给我们存留余种， 我们早已变成 所多玛 ，像 蛾摩拉 一样了。”
ROM|9|30|这样，我们要怎么说呢？那不追求义的外邦人却获得了义，就是因信而获得的义。
ROM|9|31|但 以色列 人追求律法的义，反而达不到律法的义。
ROM|9|32|这是什么缘故呢？是因为他们不凭着信心，而是凭着行为，他们正跌在那绊脚石上。
ROM|9|33|就如经上所记： “我在 锡安 放一块绊脚的石头，使人跌倒的磐石； 信靠他的人必不蒙羞。”
ROM|10|1|弟兄们，我心里所渴望的和向上帝所求的，是要 以色列 人得救。
ROM|10|2|我为他们作证，他们对上帝有热心，但不是按着真知识。
ROM|10|3|因为不明白上帝的义，想要立自己的义，他们就不服上帝的义了。
ROM|10|4|律法的总结就是基督，使所有信他的人都得着义。
ROM|10|5|论到出于律法的义， 摩西 写着：“行这些事的人，就必因此得生。”
ROM|10|6|但出于信的义却如此说：“你不要心里说：谁要升到天上去呢？（就是说，把基督领下来。）
ROM|10|7|或说：谁要下到阴间去呢？（就是说，把基督从死人中领上来。）”
ROM|10|8|他到底怎么说呢？ “这话语就离你近， 就在你口中，在你心里，” （就是说，我们传扬所信的话语。）
ROM|10|9|你若口里宣认耶稣为主，心里信上帝叫他从死人中复活，就必得救。
ROM|10|10|因为，人心里信就可以称义，口里宣认就可以得救。
ROM|10|11|经上说：“凡信靠他的人必不蒙羞。”
ROM|10|12|犹太 人和 希腊 人并没有分别，因为人人都有同一位主，他也厚待求告他的每一个人。
ROM|10|13|因为“凡求告主名的就必得救”。
ROM|10|14|然而，人未曾信他，怎能求告他呢？未曾听见他，怎能信他呢？没有传道的，怎能听见呢？
ROM|10|15|若没有奉差遣，怎能传道呢？如经上所记：“报福音、传喜信的人，他们的脚踪何等佳美！”
ROM|10|16|但不是每一个人都听从福音，因为 以赛亚 说：“主啊，我们所传的有谁信呢？”
ROM|10|17|可见，信道是从听道来的，听道是从基督的话来的。
ROM|10|18|但我要问，人没有听见吗？当然听见了。 “他们的声音传遍全地； 他们的言语传到地极。”
ROM|10|19|我再问， 以色列 人不知道吗？先有 摩西 说： “我要以不成国的激起你们嫉妒； 我要以愚顽的国惹起你们发怒。”
ROM|10|20|又有 以赛亚 放胆说： “没有寻找我的，我要让他们寻见； 没有求问我的，我要向他们显现。”
ROM|10|21|关于 以色列 人，他说：“我整天向那悖逆顶嘴的百姓招手。”
ROM|11|1|那么，我要问，上帝弃绝了他的百姓吗？绝对没有！因为我也是 以色列 人， 亚伯拉罕 的后裔，属 便雅悯 支派的。
ROM|11|2|上帝并没有弃绝他预先所知道的百姓。你们岂不知道经上论到 以利亚 是怎么说的呢？他在上帝面前怎样控告 以色列 人说：
ROM|11|3|“主啊，他们杀了你的先知，拆了你的祭坛，只剩下我一个人，他们还要我的命。”
ROM|11|4|但上帝的指示是怎么对他说的呢？他说：“我为自己留下七千人，是未曾向 巴力 屈膝的。”
ROM|11|5|现在这时刻也是这样，照着出于恩典的拣选，还有所留的余数。
ROM|11|6|既是靠恩典，就不凭行为，不然，恩典就不再是恩典了。
ROM|11|7|那又怎么说呢？ 以色列 人所寻求的，他们没有得着。但是蒙拣选的人得着了，其余的人却成了顽梗不化的。
ROM|11|8|如经上所记： “上帝给他们昏沉的灵， 眼睛看不见， 耳朵听不到， 直到今日。”
ROM|11|9|大卫 也说： “愿他们的宴席变为罗网，变为陷阱， 变为绊脚石，作他们的报应。
ROM|11|10|愿他们的眼睛昏花，看不见； 愿你时常弯下他们的腰。”
ROM|11|11|那么，我再问，他们失足是要他们跌倒吗？绝对不是！因他们的过犯，救恩反而临到外邦人，要激起他们嫉妒的心。
ROM|11|12|如果他们的过犯成为世界的富足，他们的缺乏成为外邦人的富足，更何况他们全数得救呢？
ROM|11|13|我对你们外邦人说，正因为我是外邦人的使徒，我敬重我的职分，
ROM|11|14|希望可以激起我骨肉之亲的嫉妒，好救他们一些人。
ROM|11|15|如果他们被丢弃，世界因而得以与上帝和好；他们被收纳，岂不就是从死人中复生吗？
ROM|11|16|所献的新面若圣洁，整个面团都圣洁了；树根若圣洁，树枝也圣洁了。
ROM|11|17|若有几根枝子被折下来，你这野橄榄枝接上去，同享橄榄根的肥汁，
ROM|11|18|你就不可向旧枝子夸口；若是夸口，该知道不是你托着根，而是根托着你。
ROM|11|19|你会说，那些枝子被折下来是为了使我接上去。
ROM|11|20|不错。他们因为不信，所以被折下来；你因为信，所以立得住。你不可自高，反要战战兢兢。
ROM|11|21|上帝既然不顾惜原来的枝子，岂会顾惜你？
ROM|11|22|可见，上帝又恩慈又严厉：对那跌倒的人是严厉的；对你是恩慈的，只要你长久在他的恩慈里，不然，你也要被砍下来。
ROM|11|23|而且，他们若不是长久不信，仍要被接上，因为上帝能够重新把他们接上去。
ROM|11|24|你是从那天生的野橄榄上砍下来的，尚且违反自然地接在好橄榄上，何况这些原来的枝子岂不更要接在原树上吗？
ROM|11|25|弟兄们，我不愿意你们不知道这奥秘，恐怕你们自以为聪明。这奥秘就是有一部分 以色列 人是硬心的，等到外邦人的数目添满了，
ROM|11|26|以色列 全家都要得救。如经上所记： “必有一位救主从 锡安 出来， 要消除 雅各 家一切不虔不敬。”
ROM|11|27|“这就是我与他们所立的约， 那时我要除去他们的罪。”
ROM|11|28|就福音来说，他们为你们的缘故是仇敌；就拣选来说，他们因列祖的缘故是蒙爱的。
ROM|11|29|因为上帝的恩赐和选召是不会撤回的。
ROM|11|30|你们从前不顺服上帝，如今因他们的不顺服，你们倒蒙了怜悯。
ROM|11|31|同样，他们现在也是不顺服，叫他们因着施给你们的怜悯，现在 也就蒙怜悯。
ROM|11|32|因为上帝把众人都圈在不顺服中，为的是要怜悯众人。
ROM|11|33|深哉，上帝的丰富、智慧和知识！ 他的判断何其难测！ 他的踪迹何其难寻！
ROM|11|34|谁知道主的心？ 谁作过他的谋士？
ROM|11|35|谁先给了他， 使他后来偿还呢？
ROM|11|36|因为万有都是本于他， 倚靠他，归于他。 愿荣耀归给他，直到永远。阿们！
ROM|12|1|所以，弟兄们，我以上帝的慈悲劝你们，将身体献上当作活祭，是圣洁的，是上帝所喜悦的，你们如此事奉乃是理所当然的 。
ROM|12|2|不要效法这个世界，只要心意更新而变化，叫你们察验何为上帝的善良、纯全、可喜悦的旨意。
ROM|12|3|我凭着所赐我的恩对你们每一位说：不要把自己看得太高，要照着上帝所分给各人的信心来衡量，看得合乎中道。
ROM|12|4|正如我们一个身子上有好些肢体，肢体也不都有一样的用处。
ROM|12|5|这样，我们许多人在基督里是一个身体，互相联络作肢体。
ROM|12|6|按着所得的恩典，我们各有不同的恩赐：或说预言，要按着信心的程度说预言；
ROM|12|7|或服事的，要专一服事；或教导的，要专一教导；
ROM|12|8|或劝勉的，要专一劝勉；施舍的，要诚实；治理的，要殷勤；怜悯人的，要乐意。
ROM|12|9|爱，不可虚假；恶，要厌恶；善，要亲近。
ROM|12|10|爱弟兄，要相亲相爱；恭敬人，要彼此推让；
ROM|12|11|殷勤，不可懒惰。要灵里火热；常常服侍主。
ROM|12|12|在盼望中要喜乐；在患难中要忍耐；祷告要恒切。
ROM|12|13|圣徒有缺乏，要供给；异乡客，要殷勤款待。
ROM|12|14|要祝福迫害你们 的，要祝福，不可诅咒。
ROM|12|15|要与喜乐的人同乐；要与哀哭的人同哭。
ROM|12|16|要彼此同心，不要心高气傲，倒要俯就卑微的人。不要自以为聪明。
ROM|12|17|不要以恶报恶，众人以为美的事要留心去做。
ROM|12|18|若是可行，总要尽力与众人和睦。
ROM|12|19|各位亲爱的，不要自己伸冤，宁可给主的愤怒留地步，因为经上记着：“主说：‘伸冤在我，我必报应。’”
ROM|12|20|不但如此，“你的仇敌若饿了，就给他吃；若渴了，就给他喝。因为你这样做，就是把炭火堆在他的头上。”
ROM|12|21|不要被恶所胜，反要以善胜恶。
ROM|13|1|在上有权柄的，人人要顺服，因为没有权柄不是来自上帝的。掌权的都是上帝所立的。
ROM|13|2|所以，抗拒掌权的就是抗拒上帝所立的；抗拒的人必自招审判。
ROM|13|3|作官的原不是要使行善的惧怕，而是要使作恶的惧怕。你愿意不惧怕掌权的吗？只要行善，你就可得他的称赞；
ROM|13|4|因为他是上帝的用人，是与你有益的。你若作恶，就该惧怕，因为他不是徒然佩剑；他是上帝的用人，为上帝的愤怒，报应作恶的。
ROM|13|5|所以，你们必须顺服，不但是因上帝的愤怒，也是因着良心。
ROM|13|6|你们纳粮也为这个缘故，因他们是上帝的仆役，专管这事。
ROM|13|7|凡人所当得的，就给他。当得粮的，给他纳粮；当得税的，给他上税；当惧怕的，惧怕他；当恭敬的，恭敬他。
ROM|13|8|你们除了彼此相爱，对任何人都不可亏欠什么，因为那爱人的就成全了律法。
ROM|13|9|那不可奸淫，不可杀人，不可偷盗，不可贪婪，或别的诫命，都包括在“爱邻 如己”这一句话之内了。
ROM|13|10|爱是不对邻人作恶，所以爱就成全了律法。
ROM|13|11|还有，你们要知道，现在正是该从睡梦中醒来的时候了；因为我们得救，现在比初信的时候更近了。
ROM|13|12|黑夜已深，白昼将近。所以我们该除去暗昧的行为，带上光明的兵器。
ROM|13|13|行事为人要端正，好像在白昼行走。不可荒宴醉酒；不可好色淫荡；不可纷争嫉妒。
ROM|13|14|总要披戴主耶稣基督，不要只顾满足肉体，去放纵私欲。
ROM|14|1|信心软弱的，你们要接纳，不同的意见，不要争论。
ROM|14|2|有人信什么都可吃；但那软弱的，只吃蔬菜。
ROM|14|3|吃的人不可轻看不吃的人；不吃的人也不可评断吃的人，因为上帝已经接纳他了。
ROM|14|4|你是谁，竟评断别人的仆人呢？他或站立或跌倒，自有他的主人在，而且他也必会站立，因为主能使他站稳。
ROM|14|5|有人看这日比那日强；有人看日日都是一样。只是各人要在自己的心意上坚定。
ROM|14|6|守日子的人是为主守的。吃的人是为主吃的，因他感谢上帝；不吃的人是为主不吃的，他也感谢上帝。
ROM|14|7|我们没有一个人为自己而活，也没有一个人为自己而死。
ROM|14|8|我们若活，是为主而活；我们若死，是为主而死。所以，我们或死或活总是主的人。
ROM|14|9|为此，基督死了，又活了，为要作死人和活人的主。
ROM|14|10|可是你，你为什么评断弟兄呢？你又为什么轻看弟兄呢？因我们都要站在上帝的审判台前。
ROM|14|11|经上写着： “主说，我指着我的永生起誓： 万膝必向我跪拜； 万口必称颂上帝。”
ROM|14|12|这样看来，我们各人一定要把自己的事在上帝面前 交代。
ROM|14|13|所以，我们不可再彼此评断，宁可决意不给弟兄放置障碍或绊脚石。
ROM|14|14|我凭着主耶稣确知深信，凡物本来没有不洁净的，除非人以为不洁净的，在他就不洁净了。
ROM|14|15|你若因食物使弟兄忧愁，就不是按着爱心行事。基督已经为他死，你不可因你的食物使他败坏。
ROM|14|16|所以，不可让你们的善被人毁谤。
ROM|14|17|因为上帝的国不在乎饮食，而在乎公义、和平及圣灵中的喜乐 。
ROM|14|18|凡这样服侍基督的，就为上帝所喜悦，又为人所赞许。
ROM|14|19|所以，我们务要追求 和平与彼此造就的事。
ROM|14|20|不可因食物毁坏上帝的工作。一切都是洁净的，但有人因食物使人跌倒，这在他就是恶了。
ROM|14|21|无论是吃肉是喝酒，是什么别的事，使弟兄跌倒，一概不做，才是善的。
ROM|14|22|你有信心，就要在上帝面前持守。人能在自己以为可行的事上不自责就有福了。
ROM|14|23|若有人疑惑而吃的，就被定罪，因为他吃不是出于信心。凡不出于信心的都是罪。
ROM|15|1|我们坚强的人应该分担不坚强的人的软弱，不求自己的喜悦。
ROM|15|2|我们各人务必要让邻人喜悦，使他得益处，得造就。
ROM|15|3|因为基督也不求自己的喜悦，如经上所记：“辱骂你的人的辱骂都落在我身上。”
ROM|15|4|从前所写的圣经都是为教导我们写的，要使我们藉着忍耐和因圣经所生的安慰，得着盼望。
ROM|15|5|但愿赐忍耐和安慰的上帝使你们彼此同心，效法基督耶稣，
ROM|15|6|为使你们同心同声荣耀我们主耶稣基督的父上帝！
ROM|15|7|所以，你们要彼此接纳，如同基督接纳你们一样，归荣耀给上帝。
ROM|15|8|我说，基督是为上帝真理作了受割礼的人的执事，要证实所应许列祖的话，
ROM|15|9|并使外邦人，因他的怜悯，荣耀上帝。如经上所记： “因此，我要在外邦中称颂你， 歌颂你的名。”
ROM|15|10|又说： “外邦人哪，你们要与主的子民一同欢乐。”
ROM|15|11|又说： “列邦啊，你们要赞美主！ 万民哪，你们都要颂赞他！”
ROM|15|12|又有 以赛亚 说： “将来有 耶西 的根， 就是那兴起来要治理列邦的； 外邦人要仰望他。”
ROM|15|13|愿赐盼望的上帝，因你们的信把各样的喜乐、平安 充满你们的心，使你们藉着圣灵的能力大有盼望！
ROM|15|14|我的弟兄们，我本人也深信你们自己充满良善，有各种丰富的知识，也能彼此劝戒。
ROM|15|15|但我更大胆写信给你们，是要在一些事上提醒你们，我因上帝所赐我的恩，
ROM|15|16|使我为外邦人作基督耶稣的仆役，作上帝福音的祭司，使所献上的外邦人因着圣灵成为圣洁，可蒙悦纳。
ROM|15|17|所以，有关上帝面前的事奉，我在基督耶稣里是有可夸的。
ROM|15|18|除了基督藉我做的那些事，我什么都不敢提，只提他藉我的言语作为，用神迹奇事的能力，并上帝的灵 的能力，使外邦人顺服；甚至我从 耶路撒冷 ，直转到 以利哩古 ，到处传了基督的福音。
ROM|15|19|
ROM|15|20|这样，我立了志向，不在基督的名已经传扬过的地方传福音，免得建造在别人的根基上；
ROM|15|21|却如经上所记： “未曾传给他们的，他们必看见； 未曾听见过的事，他们要明白。”
ROM|15|22|因此我多次被拦阻，不能到你们那里去。
ROM|15|23|但如今，在这一带再没有可传的地方，而且这许多年来，我迫切想去你们那里，
ROM|15|24|盼望到 西班牙 去的时候经过，得见你们，先与你们彼此交往，心里稍得满足，然后蒙你们为我送行。
ROM|15|25|但如今我要到 耶路撒冷 去，供应圣徒的需要。
ROM|15|26|因为 马其顿 和 亚该亚 人乐意凑出一些捐款给 耶路撒冷 圣徒中的穷人。
ROM|15|27|这固然是他们乐意的，其实也算是所欠的债；因为外邦人既然分享了他们灵性上的好处，就当把肉体上的需用供给他们。
ROM|15|28|等我办完了这事，把这笔捐款 交付给他们，我就要路过你们那里，到 西班牙 去。
ROM|15|29|我也知道去你们那里的时候，我将带着基督丰盛的恩典去。
ROM|15|30|弟兄们，我藉着我们的主耶稣基督，又藉着圣灵的爱，劝你们与我一同竭力为我祈求上帝，
ROM|15|31|使我脱离在 犹太 不顺从的人，也让我在 耶路撒冷 的事奉可蒙圣徒悦纳，
ROM|15|32|并使我照着上帝的旨意欢欢喜喜地到你们那里，与你们同得安息。
ROM|15|33|愿赐平安的上帝与你们众人同在。阿们！
ROM|16|1|我对你们推荐我们的姊妹 非比 ，她是 坚革哩 教会中的执事。
ROM|16|2|请你们在主里用合乎圣徒的方式来接待她。她在任何事上需要你们帮助，你们就帮助她；因她素来帮助许多人，也帮助了我。
ROM|16|3|请向 百基拉 和 亚居拉 问安。他们在基督耶稣里作我的同工，
ROM|16|4|也为我的性命把自己的生死置之度外；不但我感谢他们，就是外邦的众教会也感谢他们。
ROM|16|5|又向在他们家中的教会问安。向我所亲爱的 以拜尼土 问安，他是 亚细亚 归于基督的初结果子。
ROM|16|6|又向 马利亚 问安，她为你们非常辛劳。
ROM|16|7|又向与我一同坐监的亲戚 安多尼古 和 犹尼亚 问安，他们在使徒中是有名望的，也是比我先在基督里的。
ROM|16|8|又向我在主里面所亲爱的 暗伯利 问安。
ROM|16|9|又向我们在基督里的同工 耳巴奴 和我所亲爱的 士大古 问安。
ROM|16|10|又向在基督里经过考验的 亚比利 问安。向 亚利多布 家里的人问安。
ROM|16|11|又向我亲戚 希罗天 问安。向 拿其数 家在主里的人问安。
ROM|16|12|又向为主辛劳的 土非拿 和 土富撒 问安。向所亲爱、为主非常辛劳的 彼息 问安。
ROM|16|13|又向在主里蒙拣选的 鲁孚 和他母亲问安，他的母亲就是我的母亲。
ROM|16|14|又向 亚逊其土 、 弗勒干 、 黑米 、 八罗巴 、 黑马 ，和跟他们在一起的弟兄们问安。
ROM|16|15|又向 非罗罗古 和 犹利亚 ， 尼利亚 和他姊妹， 阿林巴 和跟他们在一起的众圣徒问安。
ROM|16|16|你们要以圣洁的吻彼此问安。基督的众教会都向你们问安！
ROM|16|17|弟兄们，那些离间你们、使你们跌倒、违背所学之道的人，我劝你们要留意躲避他们。
ROM|16|18|因为这样的人不服侍我们的主基督，只服侍自己的肚腹，用花言巧语诱惑老实人的心。
ROM|16|19|你们的顺服已经传于众人，所以我为你们欢喜；但我愿你们在善上聪明，在恶上愚拙。
ROM|16|20|那赐平安 的上帝快要把撒但践踏在你们脚下。愿我们主耶稣基督的恩与你们同在！
ROM|16|21|我的同工 提摩太 ，和我的亲戚 路求 、 耶孙 、 所西巴德 ，向你们问安。
ROM|16|22|我这代笔写信的 德提 ，在主里向你们问安。
ROM|16|23|那接待我，也接待全教会的 该犹 ，向你们问安。城里的财务官 以拉都 和弟兄 括土 向你们问安。
ROM|16|24|
ROM|16|25|惟有上帝能照我所传的福音和所讲的耶稣基督，并照历代以来隐藏的奥秘的启示，坚固你们。
ROM|16|26|这奥秘如今显示出来，而且按着永生上帝的命令，藉众先知的书指示万民，使他们因信而顺服。
ROM|16|27|愿荣耀，藉着耶稣基督，归给独一全智的上帝，直到永远。阿们！
1COR|1|1|奉上帝旨意，蒙召作基督耶稣使徒的 保罗 ，同弟兄 所提尼 ，
1COR|1|2|写信给在 哥林多 上帝的教会—就是在基督耶稣里成圣、蒙召作圣徒的—以及所有在各处求告我主耶稣基督之名的人。基督是他们的主，也是我们的主。
1COR|1|3|愿恩惠、平安 从我们的父上帝并主耶稣基督归给你们！
1COR|1|4|我常为你们感谢我的上帝，因上帝在基督耶稣里所赐给你们的恩惠。
1COR|1|5|因为你们在他里面凡事富足，具有各种口才、各样知识，
1COR|1|6|正如我为基督作的见证在你们心里得以坚固，
1COR|1|7|以致你们在恩赐上一无欠缺，切切等候我们主耶稣基督的显现。
1COR|1|8|他也必坚固你们到底，使你们在我们主耶稣基督 的日子无可指责。
1COR|1|9|上帝是信实的，他呼召你们好与他儿子—我们的主耶稣基督—共享团契。
1COR|1|10|弟兄们，我藉我们主耶稣基督的名劝你们说话要一致。你们中间不可分裂，只要一心一意彼此团结。
1COR|1|11|我的弟兄们， 革来 氏家里的人曾对我提起你们，说你们中间有纷争。
1COR|1|12|我的意思是，你们各人说：“我是属 保罗 的”；“我是属 亚波罗 的”；“我是属 矶法 的”；“我是属基督的。”
1COR|1|13|基督是分裂的吗？ 保罗 为你们钉了十字架吗？你们是奉 保罗 的名受了洗吗？
1COR|1|14|我感谢上帝 ，除了 基利司布 和 该犹 以外，我没有给你们中的任何一个人施洗，
1COR|1|15|免得有人说你们是奉我的名受洗的。
1COR|1|16|我曾为 司提法那 家施过洗；此外我已记不清有没有给别人施过洗。
1COR|1|17|因为基督差遣我不是为施洗，而是为传福音；并不是用智慧的言论，免得基督的十字架落了空。
1COR|1|18|因为十字架的道理，在那灭亡的人是愚拙，在我们得救的人却是上帝的大能。
1COR|1|19|就如经上所记： “我要摧毁智慧人的智慧， 废弃聪明人的聪明。”
1COR|1|20|智慧人在哪里？文士在哪里？这世上的辩士在哪里？上帝岂不是已使这世上的智慧变成愚拙了吗？
1COR|1|21|既然世人凭自己的智慧不认识上帝，上帝就本着自己的智慧乐意藉着人所传愚拙的话拯救那些信的人。
1COR|1|22|犹太 人要的是神迹， 希腊 人求的是智慧，
1COR|1|23|我们却是传被钉十字架的基督，这对 犹太 人是绊脚石，对外邦人是愚拙；
1COR|1|24|但对那蒙召的，无论是 犹太 人、 希腊 人，基督总是上帝的大能，上帝的智慧。
1COR|1|25|因为，上帝的愚拙总比人智慧；上帝的软弱总比人强壮。
1COR|1|26|弟兄们哪，想一想你们的蒙召，按着人的观点，有智慧的不多，有能力的不多，有尊贵地位的也不多。
1COR|1|27|但是，上帝拣选了世上愚拙的，为了使有智慧的羞愧；又拣选了世上软弱的，为了使强壮的羞愧。
1COR|1|28|上帝也拣选了世上卑贱的，被人厌恶的，以及那一无所有的，为要废掉那样样都有的，
1COR|1|29|使凡血肉之躯的，在上帝面前，一个也不能自夸。
1COR|1|30|但你们得以在基督耶稣里是本乎上帝，他使基督成为我们的智慧，成为公义、圣洁、救赎。
1COR|1|31|如经上所记：“要夸耀的，该夸耀主。”
1COR|2|1|弟兄们，从前我到你们那里去，并没有用高言大智对你们宣讲上帝的奥秘。
1COR|2|2|因为我曾定了主意，在你们中间不知道别的，只知道耶稣基督并他钉十字架。
1COR|2|3|我在你们那里时，又软弱，又惧怕，又战战兢兢。
1COR|2|4|我说的话、讲的道不是用委婉智慧的言语 ，而是以圣灵的大能来证明，
1COR|2|5|为要使你们的信不靠着人的智慧，而是靠着上帝的大能。
1COR|2|6|然而，在成熟的人中，我们也讲智慧，但不是今世的智慧，也不是今世有权有位、将要灭亡的人的智慧。
1COR|2|7|我们讲的是从前隐藏的、上帝奥秘的智慧，就是上帝在万世以前预定使我们得荣耀的智慧；
1COR|2|8|这智慧，今世有权有位的人没有一个知道，若知道，他们就不会把荣耀的主钉在十字架上了。
1COR|2|9|如经上所记： “上帝为爱他的人所预备的 是眼睛未曾看见，耳朵未曾听见， 人心也未曾想到的。”
1COR|2|10|只有上帝藉着圣灵把这事向我们显明了；因为圣灵参透万事，就是上帝深奥的事也参透了。
1COR|2|11|除了在人里头的灵，谁知道人的事？照样，除了上帝的灵，也没有人知道上帝的事。
1COR|2|12|我们所领受的并不是世上的灵，而是从上帝来的灵，为使我们知道上帝把恩赐赏给我们的事。
1COR|2|13|我们也讲说这些事，不是用人的智慧所教的言语，而是用圣灵所教的言语，用属灵的话解释属灵的事 。
1COR|2|14|然而，属血气的人不接受上帝的灵的事，他反倒以这为愚拙，并且他不能了解，因为这些事惟有属灵的人才能领悟。
1COR|2|15|属灵的人能看透万事，却没有一人能看透他。
1COR|2|16|“谁曾知道主的心？ 谁会教导他？” 至于我们，我们有基督的心。
1COR|3|1|弟兄们，我从前对你们说话，还不能把你们当作属灵的，只能把你们当作属肉体的，你们在基督里仅是婴孩。
1COR|3|2|我用奶喂你们，没有用饭喂你们，因为那时你们不能吃。就是如今还是不能，
1COR|3|3|因为你们仍是属肉体的。你们中间有嫉妒、纷争，这岂不是属乎肉体，照着世人的样子生活吗？
1COR|3|4|有人说：“我是属 保罗 的”；有人说：“我是属 亚波罗 的”；这样你们岂不是和世人一样吗？
1COR|3|5|亚波罗 算什么？ 保罗 算什么？我们都是上帝的执事，藉着我们，你们信了；这不过是照着主给各人的恩赐去做罢了。
1COR|3|6|我栽种了， 亚波罗 浇灌了，惟有上帝使它生长。
1COR|3|7|可见，栽种的算不了什么，浇灌的也算不了什么；惟有上帝能使它生长。
1COR|3|8|栽种的和浇灌的都是一样，但将来各人要照自己的劳苦得到自己的报酬。
1COR|3|9|因为我们是上帝的同工，而你们是上帝的田地，上帝的房屋。
1COR|3|10|我照上帝所给我的恩典，好像一个聪明的工头，立好了根基，别人在上面建造；只是各人要谨慎怎样在上面建造。
1COR|3|11|因为，那已经立好的根基就是耶稣基督，此外没有人能立别的根基。
1COR|3|12|若有人用金银、宝石，草木、禾秸，在这根基上建造，
1COR|3|13|各人的工程必将显露，因为那日子要将它显明，有火把它暴露出来，这火要试炼各人的工程怎样。
1COR|3|14|人在那根基上所建造的工程若能保得住，他将要得赏赐。
1COR|3|15|人的工程若被烧了，他将损失，虽然他自己将得救，却要像从火里经过一样。
1COR|3|16|难道不知你们是上帝的殿，上帝的灵住在你们里面吗？
1COR|3|17|若有人毁坏上帝的殿，上帝一定要毁灭那人；因为上帝的殿是神圣的，这殿就是你们。
1COR|3|18|谁都不可自欺。你们中间若有人自以为在今世有智慧，倒不如变为愚拙，好成为有智慧的。
1COR|3|19|因为这世界的智慧在上帝看来是愚拙的。如经上记着： “主使有智慧的人中了自己的诡计；”
1COR|3|20|又说： “主知道智慧人的意念， 因为它们是虚妄的。”
1COR|3|21|所以，无论谁都不可夸耀人；因为万有都是你们的，
1COR|3|22|或 保罗 ，或 亚波罗 ，或 矶法 ，或世界，或生，或死，或现今的事，或将来的事，全是你们的，
1COR|3|23|而你们是属基督的，基督是属上帝的。
1COR|4|1|人应该把我们看为基督的执事，为上帝的奥秘的管家。
1COR|4|2|所求于管家的，是要他忠心。
1COR|4|3|我被你们评断，或被别人评断，我都以为是极小的事；连我自己也不评断自己。
1COR|4|4|虽然我不觉得自己有错，却也不能因此判为无罪；审断我的是主。
1COR|4|5|所以，时候未到，在主来以前什么都不要评断，他要照出暗中的隐情，揭发人的动机。那时，各人要从上帝那里得著称赞。
1COR|4|6|弟兄们，为你们的缘故，我拿这些事应用到我自己和 亚波罗 身上，让你们从我们学到“不可过于圣经所记”这话的意思，免得你们自高自大，看重这个，看轻那个。
1COR|4|7|使你与人不同的是谁呢？你所有的有哪一个不是领受的呢？若是领受的，为何自夸，仿佛不是领受的呢？
1COR|4|8|你们已经饱足了，已经富足了，用不着我们，自己就作王了。我愿意你们果真作王，让我们也可以与你们一同作王！
1COR|4|9|我想，上帝把我们作使徒的明显地列在末后，好像定死罪的囚犯，因为我们成了一台戏，给世界、天使和众人观看。
1COR|4|10|我们为基督的缘故成为愚拙的；你们在基督里倒是聪明的。我们软弱，你们倒强壮；你们有荣耀，我们倒被藐视。
1COR|4|11|直到如今，我们还是又饥又渴，又赤身露体，又挨打，又到处漂泊，
1COR|4|12|并且劳碌，亲手做工；被人咒骂，我们就祝福；被人迫害，我们就忍受；
1COR|4|13|被人毁谤，我们就劝导。直到如今，人还把我们看作世上的污秽，万物中的渣滓。
1COR|4|14|我写这些话，不是要使你们羞愧，而是要警戒你们，好像我所爱的儿女一样。
1COR|4|15|虽然你们在基督里有无数的导师，却没有许多父亲，因我是在基督耶稣里用福音生了你们。
1COR|4|16|所以，我求你们要效法我。
1COR|4|17|因此，我已差 提摩太 到你们那里去。他在主里面是我亲爱和忠心的儿子；他要提醒你们，我在基督耶稣 里怎样行事为人，在各处各教会中怎样教导人。
1COR|4|18|有些人以为我不到你们那里去而自高自大。
1COR|4|19|但是，主若准许，我会很快到你们那里去；我所要知道的，不是那些自高自大者的言语，而是他们的权能。
1COR|4|20|因为上帝的国不在乎言语，而在乎权能。
1COR|4|21|你们愿意怎么样呢？要我带着棍子到你们那里去呢，还是带着慈爱温柔的心呢？
1COR|5|1|我确实听说在你们中间有淫乱的事；这种淫乱连外邦人中也没有，就是有人和他的继母同居。
1COR|5|2|你们还自高自大！你们不是该觉得痛心，把做这事的人从你们中间赶出去吗？
1COR|5|3|我人虽然不在你们那里，心却在你们那里，好像亲自与你们同在。我奉我们主耶稣 的名，已经判断了做这事的人。你们聚会的时候，我的心和你们同在。你们藉着我们主耶稣的权能，
1COR|5|4|
1COR|5|5|要把这样的人交给撒但，使他的肉体败坏，好让他的灵魂在主的日子可以得救。
1COR|5|6|你们这样自夸是不好的。你们不知道一点面酵能使全团发起来吗？
1COR|5|7|既然你们是无酵的面，要把旧酵除净，好使你们成为新团；因为我们逾越节的羔羊—基督已经被杀献为祭牲了。
1COR|5|8|所以，我们来守这节，不可用旧酵，就是不可用恶毒、邪恶的酵，只用纯洁真实的无酵饼。
1COR|5|9|我先前写信告诉过你们，不可与淫乱的人交往。
1COR|5|10|此话不是泛指这世上所有行淫乱的，或贪婪的，勒索的，或拜偶像的；若是这样，你们非离开这世界不可。
1COR|5|11|但现在，我写信告诉你们，若有称为弟兄的人却仍犯淫乱，或贪婪，或拜偶像，或辱骂，或醉酒，或勒索，这样的人不可跟他交往，就是跟他吃饭都不可以。
1COR|5|12|因为审判教外的人与我何干？教内的人岂不是你们要审判吗？
1COR|5|13|至于外人有上帝审判他们。如经上说：“要从你们中间把那邪恶的人赶出去。”
1COR|6|1|你们中间有彼此争吵的事，怎敢告到不义的人面前，而不告到圣徒面前呢？
1COR|6|2|你们岂不知圣徒要审判世界吗？若世界要受你们的审判，难道你们不配审判这最小的事吗？
1COR|6|3|你们岂不知我们要审判天使吗？何况今生的事呢！
1COR|6|4|既是这样，你们若有今生当审判的事，会让教会所轻看的人来审判吗？
1COR|6|5|我说这话是要使你们惭愧。难道你们中间没有一个有智慧的人能审断弟兄中的事吗？
1COR|6|6|你们竟然有弟兄去告弟兄，而且告到不信主的人面前。
1COR|6|7|你们彼此告状，这已经是你们的大错了。为什么不情愿受冤屈呢？为什么不情愿吃亏呢？
1COR|6|8|你们反倒去冤枉人，亏负人，况且所冤枉所亏负的就是弟兄。
1COR|6|9|你们岂不知不义的人不能承受上帝的国吗？不要自欺！无论是淫乱的、拜偶像的、奸淫的、作娼妓 的，亲男色的、
1COR|6|10|偷窃的、贪婪的、醉酒的、辱骂的、勒索的，都不能承受上帝的国。
1COR|6|11|从前你们中间也有人是这样；但现在你们奉主耶稣基督 的名，并藉着我们上帝的灵，已经洗净，已经成圣，已经称义了。
1COR|6|12|“凡事我都可行”，但不是凡事都有益处。“凡事我都可行”，但无论哪一件，我都不受它的辖制。
1COR|6|13|“食物是为肚腹，肚腹是为食物”；但上帝要使这两样都毁坏。身体不是为淫乱，而是为主；主也是为身体。
1COR|6|14|上帝已经使主复活，也要用他自己的能力使我们复活。
1COR|6|15|你们岂不知道你们的身体是基督的肢体吗？我可以把基督的肢体作为娼妓的肢体吗？绝对不可！
1COR|6|16|你们岂不知道与娼妓苟合的，就是与她成为一体吗？因为主说：“二人要成为一体。”
1COR|6|17|但与主联合的，就是与主成为一灵。
1COR|6|18|你们要远避淫行。人所犯的，无论什么罪，都在身体以外；惟有行淫的，是得罪自己的身体。
1COR|6|19|你们岂不知道你们的身体是圣灵的殿吗？这圣灵是从上帝而来，住在你们里面的。而且你们不是属自己的人，
1COR|6|20|因为你们是重价买来的。所以，要在你们的身体上荣耀上帝。
1COR|7|1|关于你们信上所提的事，男人不亲近女人倒好。
1COR|7|2|但为了避免淫乱的事，男人当各有自己的妻子，女人也当各有自己的丈夫。
1COR|7|3|丈夫对妻子要尽本分；妻子对丈夫也要如此。
1COR|7|4|妻子对自己的身体没有主张的权柄，权柄在丈夫；丈夫对自己的身体也没有主张的权柄，权柄在妻子。
1COR|7|5|夫妻不可忽略对方的需求，除非为了要专心祷告，在两相情愿下暂时分房；以后仍要同房，免得撒但趁着你们情不自禁而引诱你们。
1COR|7|6|我说这话是出于容忍，不是命令。
1COR|7|7|我愿众人像我一样；但是各人都有来自上帝的恩赐，一个是这样，一个是那样。
1COR|7|8|我对没有嫁娶的和寡妇说，他们若能维持独身像我一样就好。
1COR|7|9|但他们若不能自制，就应该嫁娶，与其欲火攻心，倒不如结婚为妙。
1COR|7|10|至于那已经嫁娶的，我吩咐他们—其实不是我，而是主吩咐的：妻子不可离开丈夫，
1COR|7|11|若是离开了，不可再嫁，不然要跟丈夫复和；丈夫也不可离弃妻子。
1COR|7|12|我对其余的人说—是我，不是主说—倘若某弟兄有不信的妻子，妻子也情愿和他一起生活，他就不可离弃妻子。
1COR|7|13|妻子有不信的丈夫，丈夫也情愿和她一起生活，她就不可离弃丈夫。
1COR|7|14|因为不信的丈夫会因着妻子成了圣洁；不信的妻子也会因着丈夫 成了圣洁。不然，你们的儿女就不洁净了，但现在他们是圣洁的。
1COR|7|15|倘若那不信的人要离开，就由他离开吧！无论是弟兄是姊妹，遇着这样的事都不必拘束。上帝召你们原是要你们和睦。
1COR|7|16|你这作妻子的怎么知道不能救你的丈夫呢？你这作丈夫的怎么知道不能救你的妻子呢？
1COR|7|17|无论如何，要照主所分给各人的恩赐和上帝所召各人的情况生活。我在各教会里都是这样规定的。
1COR|7|18|有人受割礼后才蒙召，他就不必除去割礼的记号。有人未受割礼前蒙召，他就不必受割礼。
1COR|7|19|受割礼算不了什么，不受割礼也算不了什么，只要谨守上帝的诫命就是了。
1COR|7|20|各人蒙召的时候是什么身份，要守住这身份。
1COR|7|21|你是作奴隶时蒙召的吗？不要介意；若能获得自由，就争取自由更好。
1COR|7|22|因为，蒙主呼召的奴仆是主所释放的人；蒙主呼召的自由之人是基督的奴仆。
1COR|7|23|你们是重价买来的；不要作人的奴仆。
1COR|7|24|弟兄们，你们各人蒙召的时候是什么身份，要在上帝面前守住这身份。
1COR|7|25|关于未婚女子，我没有主的命令，但我既蒙主怜悯、作为一个可信靠的人，把自己的意见告诉你们。
1COR|7|26|因现今的艰难，据我看来，人不如安于现状。
1COR|7|27|你已经有了妻子，就不要求摆脱；你还没有妻子，就不要想娶妻。
1COR|7|28|你若娶妻，并不是犯罪；未婚女子若出嫁，也不是犯罪。然而，这等人会遭受肉身上的苦难，我宁愿你们免受这苦难。
1COR|7|29|弟兄们，我是说：时候不多了。从此以后，那有妻子的，要像没有一样；
1COR|7|30|哀哭的，不像在哀哭；快乐的，不像在快乐；购买的，像一无所得；
1COR|7|31|享受这世界的，不像在享受这世界；因为这世界的局面将要过去了。
1COR|7|32|我愿你们一无挂虑。没有结婚的是为主的事挂虑，想怎样令主喜悦；
1COR|7|33|结了婚的是为世上的事挂虑，想怎样让妻子喜悦，
1COR|7|34|于是，他就分心了。没有结婚的和未婚的女子是为主的事挂虑，为要身体和心灵都圣洁；已经出嫁的是为世上的事挂虑，想怎样让丈夫喜悦。
1COR|7|35|我说这话是为你们的益处，不是要限制你们，而是要你们做合宜的事，得以不分心地对主忠诚。
1COR|7|36|若有人认为自己待他的女儿 不合宜，女儿也过了适婚年龄 ，他可以随意处理，不算有罪，让两人结婚就是了。
1COR|7|37|倘若有人心里坚定，没有不得已的事，并且由得自己作主，心里又决定了不让女儿结婚 ，这样做也好。
1COR|7|38|这样看来，让自己的女儿结婚 固然是好，不让她结婚更好。
1COR|7|39|丈夫活着的时候，妻子是受约束的；丈夫若长眠了，妻子就自由了，可以随意再嫁，只是要嫁给主里面的人。
1COR|7|40|然而，按我的意见，她若能守节就更有福气。我想我自己也有上帝的灵的感动。
1COR|8|1|关于祭过偶像的食物，我们晓得“我们都有知识”，但知识使人自高自大，惟有爱心能造就人。
1COR|8|2|若有人自以为知道什么，他其实仍不知道他所应当知道的。
1COR|8|3|若有人爱上帝，他就是上帝所认识的人了。
1COR|8|4|关于吃祭过偶像的食物，我们知道“偶像在世上算不得什么”；也知道“上帝只有一位，没有别的”。
1COR|8|5|虽然在天上或地上有许多所谓的神明，就如他们中间有许多的神明，许多的主，
1COR|8|6|但是我们只有一位上帝，就是父，万物都出于他，我们也归于他；并只有一位主，就是耶稣基督，万物都是藉着他而有，我们也是藉着他而有。
1COR|8|7|可是，不是人人都有这知识。有人到现在因拜惯了偶像，仍以为所吃的是祭过偶像的食物；既然他们的良心软弱，也就污秽了。
1COR|8|8|其实，食物不能使我们更接近上帝，因为我们不吃也无损，吃也无益。
1COR|8|9|可是，你们要谨慎，免得你们这自由竟成了软弱人的绊脚石。
1COR|8|10|若有人见你这有知识的在偶像的庙里坐席，而这人的良心是软弱的，他岂不放胆去吃那祭过偶像的食物吗？
1COR|8|11|因此，基督为他死的那软弱弟兄，也就因你的知识沉沦了。
1COR|8|12|你们这样得罪弟兄，伤了他们软弱的良心，就是得罪基督。
1COR|8|13|所以，食物若使我的弟兄跌倒，我就永远不吃肉，免得使我的弟兄跌倒了。
1COR|9|1|我不是自由的吗？我不是使徒吗？我不是见过我们的主耶稣吗？你们不是我在主里面工作的成果吗？
1COR|9|2|假若对别人来说，我不是使徒，对你们来说，我总是使徒；因为你们在主里正是我作使徒的印证。
1COR|9|3|对那些质问我的人，这就是我的答辩。
1COR|9|4|难道我们没有权利靠着传福音吃喝吗？
1COR|9|5|难道我们没有权利带着信主的妻子一起出入，如同其余的使徒，和主的兄弟们，和 矶法 一样吗？
1COR|9|6|只有我和 巴拿巴 没有权利不做工吗？
1COR|9|7|有谁当兵而自备粮饷呢？有谁栽葡萄园而不吃园里的果子呢？有谁牧养牛羊而不喝牛羊的奶呢？
1COR|9|8|我说这些话岂是照一般人的看法？律法不也是这样说吗？
1COR|9|9|就如 摩西 的律法记着：“牛在踹谷的时候，不可笼住它的嘴。”难道上帝所挂念的是牛吗？
1COR|9|10|他不全是为我们说的吗？的确是为我们说的！因为耕种的要存着指望去耕种；收割的也要存着分享谷物的指望去收割。
1COR|9|11|我们既然把属灵的种子撒在你们中间，若从你们收取养生之物，这还算大事吗？
1COR|9|12|假如别人在你们身上享有这权利，何况我们呢？ 然而，我们并没有用过这权利，倒是凡事忍受，免得基督的福音受到阻碍。
1COR|9|13|你们岂不知在圣殿供职的人吃圣殿中的食物吗？在祭坛伺候的人分享坛上的供物吗？
1COR|9|14|主也是这样命令，要传福音的人靠着福音养生。
1COR|9|15|但这权利我全然没有用过。我写这些话，并非要你们这样待我，因为我宁可死也不让人使我所夸的落了空。
1COR|9|16|我传福音原没有可夸耀的，因为我是不得已的，若不传福音，我就有祸了。
1COR|9|17|我若甘心做这事，就有赏赐；若不甘心，责任却已经托付给我了。
1COR|9|18|这样，我的赏赐是什么呢？就是我传福音的时候，使人不花钱得福音，免得我用尽了传福音的权利。
1COR|9|19|我虽然是自由的，不受人管辖，但我甘心作了众人的仆人，为赢得更多的人。
1COR|9|20|对 犹太 人，我就作 犹太 人，为要赢得 犹太 人；对律法以下的人，我虽不在律法以下，还是作律法以下的人，为要赢得律法以下的人。
1COR|9|21|对没有律法的人，我就作没有律法的人，为要赢得没有律法的人；其实我在上帝面前，不是没有律法，而是在基督的律法之下。
1COR|9|22|对软弱的人，我就作软弱的人，为要赢得软弱的人。对什么样的人，我就作什么样的人。无论如何我总要救一些人。
1COR|9|23|凡我所做的，都是为福音的缘故，为要与人共享这福音的好处。
1COR|9|24|你们不知道在运动场上赛跑的，大家都跑，但得奖赏的只有一人？你们也要这样跑，好使你们得着奖赏。
1COR|9|25|凡参加竞赛的，在各方面都要有节制，他们不过是要得会朽坏的冠冕；我们却是要得不会朽坏的冠冕。
1COR|9|26|所以，我奔跑，不像无目标的；我斗拳，不像打空气的。
1COR|9|27|我克制己身，使它完全顺服，免得我传福音给别人，自己反而被淘汰了。
1COR|10|1|弟兄们，我不愿意你们不知道，我们的祖宗从前都在云下，都从海中经过，
1COR|10|2|都在云里、海里受洗 归了 摩西 ，
1COR|10|3|并且都吃了一样的灵粮，
1COR|10|4|也都喝了一样的灵水，所喝的是出于跟随着他们的灵磐石；那磐石就是基督。
1COR|10|5|但他们中间多半是上帝不喜欢的人，所以倒毙在旷野里了。
1COR|10|6|这些事都是我们的鉴戒，使我们不要贪恋恶事，像他们贪恋过的一样。
1COR|10|7|也不要拜偶像，像他们中有些人曾经拜过。如经上所记：“百姓坐下吃喝，起来玩乐。”
1COR|10|8|我们也不可犯奸淫，像他们中有些人曾经犯过，一天就倒毙了二万三千人。
1COR|10|9|也不可试探主 ，像他们中有些人曾试探主就被蛇咬死。
1COR|10|10|你们也不可发怨言，像他们中有些人曾经发过，就被毁灭者所灭。
1COR|10|11|这些事发生在他们身上，要作为鉴戒，而且写下来正是要警戒我们这末世的人。
1COR|10|12|所以，自以为站得稳的人必须谨慎，免得跌倒。
1COR|10|13|你们所受的考验无非是人所承受得了的。上帝是信实的，他不会让你们遭受无法承受的考验，在受考验的时候，总会给你们开一条出路，让你们能忍受得了。
1COR|10|14|所以，我亲爱的，你们要远避拜偶像的事。
1COR|10|15|我好像对精明人说的；你们要辨别我的话。
1COR|10|16|我们所祝谢的杯，岂不是同领基督的血吗？我们所擘开的饼，岂不是同领基督的身体吗？
1COR|10|17|因为饼只是一个，我们虽然人多，仍是一体，我们同享一个饼。
1COR|10|18|你们看那按肉体是 以色列 人的，那些吃祭物的人岂不是与祭坛有份吗？
1COR|10|19|那么，我怎么说呢？是说祭偶像之物算得了什么吗？或说偶像算得了什么吗？
1COR|10|20|不，我是说，他们 所献的祭是祭鬼，不是祭上帝；我不愿意你们与鬼来往。
1COR|10|21|你们不能喝主的杯，又喝鬼的杯；不能吃主的筵席，又吃鬼的筵席。
1COR|10|22|我们要惹主的嫉恨吗？我们比他更强吗？
1COR|10|23|“凡事都可行”，但不都有益处。“凡事都可行”，但不都造就人。
1COR|10|24|无论什么人，不要求自己的益处，而要求别人的益处。
1COR|10|25|凡市场上所卖的，你们只管吃，不要为良心的缘故问什么，
1COR|10|26|“因为地和其中所充满的都属于主”。
1COR|10|27|倘若有一个不信的人请你们吃饭，而你们也愿意去，凡摆在你们面前的，只管吃，不要为良心的缘故问什么。
1COR|10|28|若有人对你们说：“这是献过祭的物”，那么为了那告诉你们的人，并为了良心的缘故就不吃。
1COR|10|29|我说的良心不是你自己的，而是他的。我的自由为什么被别人的良心评断呢？
1COR|10|30|我若谢恩而吃，为什么因我谢恩的物被人毁谤呢？
1COR|10|31|所以，你们或吃或喝，无论做什么，都要为荣耀上帝而做。
1COR|10|32|你们不要使 犹太 人、 希腊 人，或上帝教会中的人跌倒；
1COR|10|33|但要像我一样，凡事都使众人喜欢，不求自己的益处，只求众人的益处，使他们得救。
1COR|11|1|你们该效法我，像我效法基督一样。
1COR|11|2|我称赞你们，因为你们凡事记得我，又坚守我所传授给你们的。
1COR|11|3|但是我要你们知道：基督是男人的头；男人是女人的头 ；上帝是基督的头。
1COR|11|4|凡男人祷告或讲道 ，若蒙着头，就是羞辱自己的头。
1COR|11|5|凡女人祷告或讲道，若不蒙着头，就是羞辱自己的头，因为这就如同剃了头发一样。
1COR|11|6|女人若不蒙着头，就该剪了头发；女人若以剪发剃发为羞愧，就该蒙着头。
1COR|11|7|男人本不该蒙着头，因为他是上帝的形像和荣耀；但女人是男人的荣耀。
1COR|11|8|起初，男人不是由女人而出，女人却是由男人而出。
1COR|11|9|而且男人不是为女人造的，女人却是为男人造的。
1COR|11|10|因此，女人为天使的缘故应当在头上有服权柄的记号。
1COR|11|11|然而，照主的安排，女人不可没有男人，男人也不可没有女人。
1COR|11|12|因为女人原是由男人而出，男人是藉着女人而生；但万有都是出于上帝。
1COR|11|13|你们自己要判断，女人祷告上帝，不蒙着头合宜吗？
1COR|11|14|你们的本性不也教导你们，男人若留长头发是他的羞辱吗？
1COR|11|15|但女人留长头发是她的荣耀，因为这头发是给她盖头的 。
1COR|11|16|若有人想要辩驳，我们却没有这样的规矩，上帝的众教会也没有。
1COR|11|17|我现在吩咐你们这话不是在称赞你们，因为你们聚会是有损无益的。
1COR|11|18|首先，我听说你们教会聚会的时候有分裂的事，我也有些相信这话。
1COR|11|19|在你们中间必然有分门结党的事，好使那些经得起考验的人显明出来。
1COR|11|20|你们聚会的时候，不是在吃主的晚餐，
1COR|11|21|因为吃的时候，各人先吃自己的饭，甚至有人饥饿，有人酒醉。
1COR|11|22|难道你们没有家可以吃喝吗？还是你们藐视上帝的教会，使那没有的羞愧呢？我该对你们说什么呢？我要称赞你们吗？在这事上我绝不称赞你们！
1COR|11|23|我当日传给你们的是从主所领受的。主耶稣被出卖的那一夜，拿起饼来，
1COR|11|24|祝谢了，就擘开，说：“这是我的身体，为你们舍 的；你们要如此行，为的是记念我。”
1COR|11|25|饭后，他也照样拿起杯来，说：“这杯是用我的血所立的新约；你们每逢喝的时候，要如此行，来记念我。”
1COR|11|26|你们每逢吃这饼，喝这杯，是宣告主的死，直到他来。
1COR|11|27|所以，任何不按规矩吃了主的饼，喝了主的杯，就是干犯主的身体和主的血了。
1COR|11|28|人应该省察自己，然后吃这饼，喝这杯。
1COR|11|29|因为人吃喝，若不分辨是主的身体，他的吃喝就是定自己的罪了。
1COR|11|30|因此，在你们中间有好些软弱的与患病的，长眠了的也不少。
1COR|11|31|我们若是先省察自己，就不至于受审判。
1COR|11|32|我们受审判的时候，就是被主管教，这样就免得和世人一同被定罪。
1COR|11|33|所以，我的弟兄们，你们聚会吃晚餐的时候，要彼此等待。
1COR|11|34|若有人饿了，要在家里先吃，免得你们聚会，反被定罪。其余的事等我来的时候再安排。
1COR|12|1|弟兄们，关于属灵的恩赐 ，我不愿意你们不明白。
1COR|12|2|你们知道，你们作外邦人的时候，随事被引诱，受了迷惑去拜不会出声的偶像。
1COR|12|3|所以，我要你们知道，被上帝的灵感动的，没有人会说“耶稣该受诅咒”；若不是被圣灵感动的，也没有人能说“耶稣是主”。
1COR|12|4|恩赐有许多种，却是同一位圣灵所赐。
1COR|12|5|事奉有许多种，却是事奉同一位主。
1COR|12|6|工作有许多种，却是同一位上帝在万人中运行万事。
1COR|12|7|圣灵彰显在各人身上，是要使人得益处。
1COR|12|8|有人藉着圣灵领受智慧的言语；有人也靠着同一位圣灵领受知识的言语；
1COR|12|9|又有人由同一位圣灵领受信心；还有人由同一位圣灵领受医病的恩赐；
1COR|12|10|又有人能行异能，又有人能作先知，又有人能辨别诸灵，又有人能说方言 ，又有人能翻方言。
1COR|12|11|这一切都是由惟一的、同一位圣灵所运行，随着自己的旨意分给各人的。
1COR|12|12|就如身体是一个，却有许多肢体，身体的肢体虽多，仍是一个身体；基督也是这样。
1COR|12|13|我们无论是 犹太 人是 希腊 人，是为奴的是自主的，都从一位圣灵受洗成了一个身体，并且共享这位圣灵。
1COR|12|14|身体原不只是一个肢体，而是许多肢体。
1COR|12|15|假如脚说：“我不是手，所以不属于身体”，它不能因此就不属于身体。
1COR|12|16|假如耳朵说：“我不是眼睛，所以不属于身体”，它也不能因此就不属于身体。
1COR|12|17|假如全身是眼睛，听觉在哪里呢？假如全身是耳朵，嗅觉在哪里呢？
1COR|12|18|但现在上帝随自己的意思把肢体一一安置在身体上了。
1COR|12|19|假如全都是一个肢体，身体在哪里呢？
1COR|12|20|但现在肢体虽多，身体还是一个。
1COR|12|21|眼睛不能对手说：“我用不着你。”头也不能对脚说：“我用不着你。”
1COR|12|22|不但如此，身上的肢体，人以为软弱的，更是不可缺少的；
1COR|12|23|身上的肢体，我们认为不体面的，越发给它加上体面；我们不雅观的，越发装饰得雅观。
1COR|12|24|我们雅观的肢体自然用不着装饰；但上帝配搭这身子，把加倍的体面给那有缺欠的肢体，
1COR|12|25|免得身体不协调，总要肢体彼此照顾。
1COR|12|26|假如一个肢体受苦，所有的肢体就一同受苦；假如一个肢体得光荣，所有的肢体就一同快乐。
1COR|12|27|你们是基督的身体，并且各自都是肢体。
1COR|12|28|上帝在教会所设立的：第一是使徒；第二是先知；第三是教师；其次是行异能的；再次是医病的恩赐，帮助人的，治理事的，说方言的。
1COR|12|29|难道个个都是使徒吗？难道个个都是先知吗？难道个个都是教师吗？难道个个都是行异能的吗？
1COR|12|30|难道个个都是有医病的恩赐吗？难道个个都是说方言的吗？难道个个都是翻方言的吗？
1COR|12|31|你们要追求那更大的恩赐。 我现今把最妙的道指示你们。
1COR|13|1|我若能说人间的方言，甚至天使的语言，却没有爱，我就成为鸣的锣、响的钹一般。
1COR|13|2|我若有先知讲道的能力，也明白各样的奥秘，各样的知识，而且有齐备的信心，使我能够移山，却没有爱，我就算不了什么。
1COR|13|3|我若将所有的财产救济穷人，又牺牲自己的身体让人夸赞 ，却没有爱，仍然对我无益。
1COR|13|4|爱是恒久忍耐；又有恩慈；爱是不嫉妒；爱是不自夸，不张狂，
1COR|13|5|不做害羞的事，不求自己的益处，不轻易发怒，不计算人的恶，
1COR|13|6|不喜欢不义，只喜欢真理；
1COR|13|7|凡事包容，凡事相信，凡事盼望，凡事忍耐。
1COR|13|8|爱是永不止息。先知讲道之能终必归于无有；说方言 之能终必停止；知识也终必归于无有。
1COR|13|9|我们现在所知道的有限，先知所讲的也有限，
1COR|13|10|等那完全的来到，这有限的必消逝。
1COR|13|11|我作孩子的时候，说话像孩子，心思像孩子，意念像孩子；既长大成人，就把孩子的事丢弃了。
1COR|13|12|我们现在是对着镜子观看，模糊不清 ；到那时，就要面对面了。我如今所认识的有限，到那时就全认识，如同主认识我一样。
1COR|13|13|如今常存的有信，有望，有爱这三样，其中最大的是爱。
1COR|14|1|你们要追求爱，也要切慕属灵的恩赐，尤其是作先知讲道 。
1COR|14|2|那说方言 的，不是对人说，而是对上帝说，因为没有人听得懂；他是藉着圣灵说各样的奥秘。
1COR|14|3|但作先知讲道的，是对人说，要造就、安慰、劝勉人。
1COR|14|4|说方言的，是造就自己；作先知讲道的，是造就教会。
1COR|14|5|我希望你们都说方言，更希望你们作先知讲道；因为说方言的，若不解释出来，使教会得造就，那作先知讲道的就比他强了。
1COR|14|6|弟兄们，我到你们那里去，若只说方言，不用启示，或知识，或预言，或教导，给你们讲解，我对你们有什么益处呢？
1COR|14|7|就连那有声而没有生命的东西，如箫，如琴，发出来的音若没有分别，怎能知道所吹所弹的是什么呢？
1COR|14|8|号角吹出来的音若不清楚，谁会预备打仗呢？
1COR|14|9|你们也是如此；若用舌头说听不懂的信息，怎能知道所说的是什么呢？你们就是向空气说话了。
1COR|14|10|世上有许多种语言，却没有一样是无意思的。
1COR|14|11|我若不明白那语言的意思，说话的人必以我为未开化的人，我也以他为未开化的人。
1COR|14|12|你们也是如此，既然你们切慕属灵的恩赐，就当追求多得造就教会的恩赐。
1COR|14|13|所以，那说方言的，就当祈求有翻方言的恩赐。
1COR|14|14|我若用方言祷告，是我的灵在祷告；但我的理智没有效果。
1COR|14|15|我应该怎么做呢？我要用灵祷告，也要用理智祷告；我要用灵歌唱，也要用理智歌唱。
1COR|14|16|不然，你用灵祝谢，那在座不通方言的人，既然不明白你的话，怎能在你感谢的时候说“阿们”呢？
1COR|14|17|你的感谢固然是好，不过不能造就别人。
1COR|14|18|我感谢上帝，我说方言比你们众人还多；
1COR|14|19|但在教会中，我宁可用理智说五句教导人的话，强过说万句方言。
1COR|14|20|弟兄们，在心志上不要作小孩子。但是，在恶事上要作婴孩，而在心志上总要作大人。
1COR|14|21|律法上记着：“主说： 我要用外邦人的舌头 和外邦人的嘴唇 向这百姓说话； 虽然如此，他们还是不听从我。”
1COR|14|22|这样看来，说方言不是为信的人作标记，而是为不信的人；作先知讲道不是为不信的人作标记，而是为信的人。
1COR|14|23|所以，全教会聚在一处的时候，若都说方言，偶然有不通方言的或是不信的人进来，岂不会说你们疯了吗？
1COR|14|24|若个个都作先知讲道，偶然有不信的或是不懂方言的人进来，就被众人劝戒，被众人审问，
1COR|14|25|他心里的隐情被显露出来，就必将脸伏地，敬拜上帝，宣告说：“上帝真的是在你们中间了。”
1COR|14|26|弟兄们，那么，你们该怎么做呢？你们聚会的时候，各人或有诗歌，或有教导，或有启示，或有方言，或有翻出来，凡事都应当造就人。
1COR|14|27|若有说方言的，只可有两个人，至多三个人，且要轮流着说，也要有一个人翻出来。
1COR|14|28|若没有人翻，就当在会中闭口，只对自己和上帝说就是了。
1COR|14|29|至于作先知讲道的，只可有两个人或是三个人，其余的人当慎思明辨。
1COR|14|30|假如旁边坐着的得了启示，那先说话的就当闭口不言。
1COR|14|31|因为你们都可以一个一个地作先知讲道，使众人都可以学习，使众人都得劝勉。
1COR|14|32|先知的灵是顺服先知的，
1COR|14|33|因为上帝不是叫人混乱，而是叫人和谐的上帝。 在圣徒的众教会中，
1COR|14|34|妇女应该闭口不言；因为，不准她们说话，总要顺服，正如律法所说的。
1COR|14|35|她们若要学什么，应该在家里问自己的丈夫，因为妇女在会中说话是可耻的。
1COR|14|36|难道上帝的话是从你们出来的吗？难道是单临到你们的吗？
1COR|14|37|若有人自以为是先知，或是属灵的，就应该知道，我所写给你们的是主的命令。
1COR|14|38|若有不理会的，你们也不必理会他。
1COR|14|39|所以，我的弟兄们，你们要切慕作先知讲道的恩赐，不要禁止说方言。
1COR|14|40|凡事都要规规矩矩地按着次序行。
1COR|15|1|弟兄们，我要你们认清我先前传给你们的福音；这福音你们领受了，又靠着它站立得住，
1COR|15|2|你们若能够持守我传给你们的信息，就必因这福音得救，否则你们是徒然相信。
1COR|15|3|我当日所领受又传给你们的，最重要的就是：照圣经所说，基督为我们的罪死了，
1COR|15|4|而且埋葬了；又照圣经所说，第三天复活了，
1COR|15|5|还显给 矶法 看，又显给十二使徒看，
1COR|15|6|后来一次显给五百多弟兄看，其中一大半到现在还在，却也有已经睡了的。
1COR|15|7|以后他显给 雅各 看，再显给众使徒看，
1COR|15|8|最后也显给我看；我如同未到产期而生的人一般。
1COR|15|9|我原是使徒中最小的，不配称为使徒，因为我曾迫害过上帝的教会。
1COR|15|10|然而，由于上帝的恩典，我才成了今日的我，并且他所赐给我的恩典不是徒然的。我比众使徒格外劳苦；其实不是我，而是上帝的恩典与我同在。
1COR|15|11|无论是我或是其他使徒，我们都如此传，你们也都如此信了。
1COR|15|12|既然我们传基督是从死人中复活了，怎么在你们中间有人说没有死人复活的事呢？
1COR|15|13|若没有死人复活的事，基督就没有复活了。
1COR|15|14|基督若没有复活，我们所传的就是枉然，你们所信的也是枉然。
1COR|15|15|这样，我们甚至被当作是为上帝妄作见证的，因为我们见证上帝是使基督复活了。如果死人真的没有复活，上帝就没有使基督复活了。
1COR|15|16|因为死人若不复活，基督也就没有复活了。
1COR|15|17|基督若没有复活，你们的信就是徒然，你们仍活在罪里。
1COR|15|18|就是在基督里睡了的人也灭亡了。
1COR|15|19|我们若靠基督只在今生有指望，就比所有的人更可怜了。
1COR|15|20|其实，基督已经从死人中复活，成为睡了之人初熟的果子。
1COR|15|21|既然死是因一人而来，死人复活也因一人而来。
1COR|15|22|在 亚当 里众人都死了；同样，在基督里众人也都要复活。
1COR|15|23|但各人是按着自己的次序复活：初熟的果子是基督；然后在他来的时候，是那些属于基督的。
1COR|15|24|再后，终结到了，那时基督既将一切执政的、掌权的、有权能的都毁灭了，就把国交给父上帝。
1COR|15|25|因为基督必须掌权，等上帝把一切仇敌都放在他的脚下。
1COR|15|26|他要毁灭的最后仇敌就是死亡。
1COR|15|27|因为经上说：“上帝使万物都服在他的脚下。”既然说万物都服了他，那使万物屈服的，很明显地是不在其内了。
1COR|15|28|既然万物服了他，那时，子也要自己顺服那叫万物服他的，好使上帝在万物之中，在万物之上。
1COR|15|29|不然，那些为死人受洗的，能做什么呢？如果死人不会复活，为什么替他们受洗呢？
1COR|15|30|我们为什么要时刻冒险呢？
1COR|15|31|弟兄们 ，我在我们的主基督耶稣里，指着你们—我所夸的极力地说，我天天冒死。
1COR|15|32|从人的观点看来，我当日在 以弗所 同野兽搏斗，对我有什么益处呢？如果死人没有复活， “让我们吃吃喝喝吧！ 因为明天要死了。”
1COR|15|33|不要被欺骗了； “滥交朋友败坏品德。”
1COR|15|34|你们要醒悟为善，不再犯罪；因为有人不认识上帝。我说这话是要使你们羞愧。
1COR|15|35|但是有人会问：“死人怎样复活呢？他们带着什么身体来呢？”
1COR|15|36|无知的人哪，你所种的若不死就不能生。
1COR|15|37|并且你所种的不是那将来要有的形体，无论是麦子或别样谷物，都不过是子粒。
1COR|15|38|但上帝随自己的意思给它一个形体，并叫各样子粒各有自己的形体。
1COR|15|39|不是所有的肉体都是同样的：人是一个样子，兽又是一个样子，鸟又是一个样子，鱼又是一个样子。
1COR|15|40|有天上的形体，也有地上的形体；但天上形体的荣光是一个样子，地上形体的荣光又是一个样子。
1COR|15|41|日有日的光辉，月有月的光辉，星有星的光辉；这星和那星的光辉也有区别。
1COR|15|42|死人复活也是这样。所种的是会朽坏的，复活的是不朽坏的；
1COR|15|43|所种的是羞辱的，复活的是荣耀的；所种的是软弱的，复活的是强壮的；
1COR|15|44|所种的是血肉的身体，复活的是灵性的身体。既有血肉的身体，也就有灵性的身体。
1COR|15|45|经上也是这样记着说：“首先的人 亚当 成了有生命的人”；末后的 亚当 成了赐生命的灵。
1COR|15|46|但是，不是属灵的在先，而是属血肉的在先，然后才是属灵的。
1COR|15|47|第一个人是出于地，是属于尘土；第二个人是出于天。
1COR|15|48|那属尘土的怎样，凡属尘土的也都怎样；属天的怎样，凡属天的也都怎样。
1COR|15|49|就如我们既有属尘土的形像，将来也必有属天的形像。
1COR|15|50|弟兄们，我要告诉你们的是：血肉之躯不能承受上帝的国，必朽坏的也不能承受不朽坏的。
1COR|15|51|我如今把一件奥秘的事告诉你们：我们不是都要睡觉，而是都要改变，
1COR|15|52|就在一刹那，眨眼之间，号筒末次吹响的时候。因号筒要吹响，死人要复活成为不朽坏的，我们也要改变。
1COR|15|53|这会朽坏的必须变成 不朽坏的；这会死的总要变成不会死的。
1COR|15|54|当这会朽坏的变成不朽坏的，这会死的变成不会死的，那时经上所记“死亡已被胜利吞灭了”的话就应验了。
1COR|15|55|“死亡啊！你得胜的权势在哪里？ 死亡啊！你的毒刺在哪里？”
1COR|15|56|死亡的毒刺就是罪，罪的权势就是律法。
1COR|15|57|感谢上帝，他使我们藉着我们的主耶稣基督得胜。
1COR|15|58|所以，我亲爱的弟兄们，你们务要坚固，不可动摇，常常竭力多做主工，因为你们知道，你们在主里的劳苦不是徒然的。
1COR|16|1|关于为圣徒捐款的事，我从前怎样吩咐 加拉太 的众教会，你们也该怎样做。
1COR|16|2|每逢七日的第一日，每人要照自己的收入抽出若干，保留起来，免得我来的时候现凑。
1COR|16|3|等到我来了，你们写信举荐谁，我就差遣他们，把你们的款项送到 耶路撒冷 去。
1COR|16|4|如果我也该去，他们可以和我同去。
1COR|16|5|我想穿越 马其顿 ；我经过了 马其顿 后，就到你们那里去，
1COR|16|6|可能会和你们同住一些时候，甚至和你们一起过冬。这样无论我往哪里去，你们可以给我送行。
1COR|16|7|我现在不愿意在路过的时候见你们；主若允许，我就指望和你们同住一些时候。
1COR|16|8|不过我要仍旧住在 以弗所 ，直到五旬节，
1COR|16|9|因为有又宽大又有效的门为我开了，虽然反对的人也多。
1COR|16|10|若是 提摩太 来到，你们要留心照顾他，使他在你们那里无所惧怕，因为他做主的工作像我一样。
1COR|16|11|所以，无论谁都不可藐视他。只要送他平安前行，让他到我这里来，因为我等着他和弟兄们同来。
1COR|16|12|至于 亚波罗 弟兄，我再三劝他同弟兄们到你们那里去；但现在他绝不愿意去，等有机会他就会去。
1COR|16|13|你们要警醒，在信仰上要站稳，要勇敢，要刚强。
1COR|16|14|你们所做的一切都要凭爱心而做。
1COR|16|15|弟兄们，你们知道 司提法那 一家，是 亚该亚 初结的果子；他们专以服事圣徒为念。
1COR|16|16|我劝你们顺服这样的人，和一切与他同工同劳的人。
1COR|16|17|司提法那 、 福徒拿都 和 亚该古 到这里来，我很高兴，因为他们补上了你们不在我身边的遗憾。
1COR|16|18|他们使我和你们心里都快慰；这样的人，你们务要敬重。
1COR|16|19|亚细亚 的众教会向你们问安。 亚居拉 、 百基拉 ，和在他们家里的教会，在主里热切地向你们问安。
1COR|16|20|众弟兄都向你们问安。要用圣洁的吻彼此问安。
1COR|16|21|我— 保罗 亲笔问安。
1COR|16|22|若有人不爱主，这人该受诅咒。主啊，愿你来！
1COR|16|23|愿主耶稣基督的恩常与你们众人同在。
1COR|16|24|我在基督耶稣里的爱与你们同在！
2COR|1|1|奉上帝旨意作基督耶稣使徒的 保罗 和弟兄 提摩太 ，写信给在 哥林多 上帝的教会和全 亚该亚 的众圣徒。
2COR|1|2|愿恩惠、平安 从我们的父上帝和主耶稣基督归给你们！
2COR|1|3|愿颂赞归于上帝—我们主耶稣基督的父；他是发慈悲的父，赐各样安慰的上帝。
2COR|1|4|我们在一切患难中，他安慰我们，使我们能用上帝所赐的安慰去安慰那些遭各样患难的人。
2COR|1|5|正如我们跟基督同受许多苦楚，我们也靠基督得许多安慰。
2COR|1|6|如果我们受患难，那是为使你们得安慰，得拯救；如果我们得安慰，那也是为使你们得安慰，这安慰能使你们忍受我们所受同样的苦楚。
2COR|1|7|我们为你们所存的盼望是确定的，因为知道你们分担了我们的痛苦，也要分享我们的安慰。
2COR|1|8|弟兄们，我们不要你们不知道，我们从前在 亚细亚 遭遇苦难，因受到无法忍受的压力，甚至连活命的指望都没有了。
2COR|1|9|自己心里也断定是必死无疑，这是要使我们不依靠自己，只依靠使死人复活的上帝。
2COR|1|10|他曾救我们脱离那极大的死亡，他要继续救我们，而且我们指望他将来还要救我们。
2COR|1|11|你们也要一同用祈祷来帮助我们，好使许多人为我们感恩，因着他们许多的祷告，我们获得了恩赐。
2COR|1|12|我们所夸的是：我们在世为人，特别是跟你们的关系，是凭着上帝所赐的坦率和真诚，不是靠人的聪明，而是靠上帝的恩惠；这是我们的良心可以作证的。
2COR|1|13|我们现在写给你们的话，无非是你们所能诵读、所能明白的，我也盼望你们真能彻底明白。
2COR|1|14|你们已经有几分认识我们，在我们主耶稣 的日子，你们会以我们为荣，正像我们也以你们为荣。
2COR|1|15|既然我这样深信，早就有意先到你们那里去，让你们得加倍的益处。
2COR|1|16|我要路过你们那里往 马其顿 去，再从 马其顿 回到你们那里，让你们给我送行往 犹太 去。
2COR|1|17|我有此意，难道是反覆不定吗？难道我的意愿是从私欲起的，以致我忽是忽非吗？
2COR|1|18|我指着信实的上帝说，我们向你们所传的道并非又是又非的。
2COR|1|19|因为，我、 西拉 和 提摩太 在你们中间传上帝的儿子耶稣基督，从没有“又是又非”的；在他只有一个“是”。
2COR|1|20|上帝的应许，不论有多少，在基督都是“是”的。所以，我们藉着他说“阿们”，使上帝因我们得荣耀。
2COR|1|21|那在基督里坚固我们和你们，并且膏抹我们的，就是上帝。
2COR|1|22|他在我们身上盖了印，并赐圣灵在我们心里作凭据。
2COR|1|23|我指着我的性命求告上帝作证，我没有再往 哥林多 去是为了要宽容你们。
2COR|1|24|我们并不是要控制你们的信心，而是要作你们的同工，让你们得快乐，因为你们在信仰上已经站得稳了。
2COR|2|1|我自己定了主意，下次不再带着悲伤到你们那里去。
2COR|2|2|我若使你们悲伤，除了因我而使他悲伤的那人以外，谁能使我喜乐呢？
2COR|2|3|我曾把这事写给你们，免得我到的时候，那该令我喜乐的人反倒令我悲伤。我也深信，你们众人都以我的喜乐为自己的喜乐。
2COR|2|4|我先前忧心忡忡、眼泪汪汪地给你们写了信，并非要使你们悲伤，而是要你们知道我格外疼爱你们。
2COR|2|5|如果有人使人悲伤，他不但使我悲伤，也是使你们众人有些悲伤。我说有些，恐怕说得太重了。
2COR|2|6|这样的人受了大多数人的责备也就够了，
2COR|2|7|倒不如赦免他，安慰他，免得他过分悲伤，甚至受不了啦！
2COR|2|8|所以，我劝你们，要向他肯定你们的爱心。
2COR|2|9|为此，我先前也写信给你们，正是要考验你们，看你们是否在一切事上都顺从我。
2COR|2|10|你们赦免谁，我也赦免谁。我若有所赦免，是在基督面前为你们的缘故赦免的，
2COR|2|11|免得撒但趁着机会胜过我们，因我们并非不知道他的诡计。
2COR|2|12|我从前为基督的福音到了 特罗亚 ，主给我开了门。
2COR|2|13|那时，因为没有遇见我的弟兄 提多 ，我心里不安，就辞别那里的人，往 马其顿 去了。
2COR|2|14|感谢上帝！他常率领我们在基督里得胜，并藉着我们在各处显扬那因认识基督而有的香气。
2COR|2|15|因为无论在得救的人或在灭亡的人当中，我们都是基督馨香之气，是献给上帝的。
2COR|2|16|对灭亡的人，这是死而又死的气味；对得救的人，这是生而又生的气味。这些事谁能当得起呢？
2COR|2|17|我们不像许多人，把上帝的道当商品贩卖，而是由于真诚，而是受命于上帝，在上帝面前凭着基督讲道。
2COR|3|1|难道我们又开始推荐自己吗？难道我们像某些人那样要用人的推荐信介绍给你们，或用你们的推荐信给人吗？
2COR|3|2|你们就是我们的推荐信，写在我们心里，被众人所知道、所诵读的，
2COR|3|3|而你们显明自己是基督的书信，藉着我们写成的。不是用墨写的，而是用永生上帝的灵写的；不是写在石版上，而是写在心版上的。
2COR|3|4|我们藉着基督才对上帝有这样的信心。
2COR|3|5|并不是我们凭自己配做什么事，我们之所以配做是出于上帝；
2COR|3|6|他使我们能配作新约的执事，不是文字上的约，而是圣灵的约；因为文字使人死，圣灵能使人活。
2COR|3|7|那用字刻在石头上属死的事奉尚且有荣光，以致 以色列 人因 摩西 脸上那逐渐褪色的荣光不能定睛看他的脸，
2COR|3|8|那属圣灵的事奉不是更有荣光吗？
2COR|3|9|若是那使人定罪的事奉有荣光，那使人称义的事奉的荣光就越发大了。
2COR|3|10|那从前有荣光的，因这更大的荣光，就算不得有荣光了；
2COR|3|11|若是那逐渐褪色的有荣光，这长存的就更有荣光了。
2COR|3|12|既然我们有这样的盼望，就大有胆量，
2COR|3|13|不像 摩西 将面纱蒙在脸上，使 以色列 人不能定睛看到那逐渐褪色的荣光的结局。
2COR|3|14|但他们的心地刚硬，直到今日诵读旧约的时候，这同样的面纱还没有揭去；因为这面纱在基督里才被废去。
2COR|3|15|然而直到今日，每逢诵读 摩西 书的时候，面纱还在他们心上。
2COR|3|16|但他们的心何时归向主，面纱就何时除去。
2COR|3|17|主就是那灵；主的灵在哪里，哪里就有自由。
2COR|3|18|既然我们众人以揭去面纱的脸得以看见 主的荣光，好像从镜子里返照，就变成了与主有同样的形像，荣上加荣，如同从主的灵 变成的。
2COR|4|1|所以，既然我们蒙怜悯受了这事奉的责任，就不丧胆，
2COR|4|2|反而把那些暗昧可耻的事弃绝了，不行诡诈，不曲解上帝的道，只将真理显扬出来，好在上帝面前把自己推荐给各人的良心。
2COR|4|3|即使我们的福音被遮蔽，那只是对灭亡的人遮蔽。
2COR|4|4|这些不信的人被这世界的神明弄瞎了心眼，使他们看不见基督荣耀的福音。基督本是上帝的像。
2COR|4|5|我们不是传自己，而是传耶稣基督为主，并且自己因耶稣作你们的仆人。
2COR|4|6|那吩咐光从黑暗里照出来的上帝已经照在我们心里，使我们知道上帝荣耀的光显在耶稣基督的脸上。
2COR|4|7|我们有这宝贝放在瓦器里，为要显明这莫大的能力是出于上帝，不是出于我们。
2COR|4|8|我们处处受困，却不被捆住；内心困扰，却没有绝望；
2COR|4|9|遭受迫害，却不被撇弃；击倒在地，却不致灭亡。
2COR|4|10|我们身上常带着耶稣的死，使耶稣的生也在我们身上显明。
2COR|4|11|因为我们这活着的人常为耶稣被置于死地，使耶稣的生命在我们这必死的人身上显明出来。
2COR|4|12|这样看来，死是在我们身上运作，生却在你们身上运作。
2COR|4|13|但我们既然有从同一位灵而来的信心，正如经上记着：“我信，故我说话”，我们也信，所以也说话；
2COR|4|14|因为知道，那使主耶稣复活的也必使我们与耶稣一同复活，并且使我们与你们一起站在他面前。
2COR|4|15|凡事都是为了你们，好使恩惠既藉着更多的人而加增，感恩也格外显多，好归荣耀给上帝。
2COR|4|16|所以，我们不丧胆。虽然我们外在的人日渐朽坏，内在的人却日日更新。
2COR|4|17|我们这短暂而轻微的苦楚要为我们成就极重、无比、永远的荣耀。
2COR|4|18|因为我们不是顾念看得见的，而是顾念看不见的；原来看得见的是暂时的，看不见的才是永远的。
2COR|5|1|因为我们知道，我们这地上的帐篷若拆毁了，我们将有上帝所造的居所，不是人手所造的，而是在天上永存的。
2COR|5|2|我们在这帐篷里叹息，渴望得到那从天上来的居所，好像穿上衣服；
2COR|5|3|倘若脱下也 不至于赤身了。
2COR|5|4|其实，我们在这帐篷里的人劳苦叹息，并不是愿意脱下地上的帐篷，而是愿意穿上天上的居所，好使这必死的被生命吞灭了。
2COR|5|5|那为我们安排这事的是上帝，他赐给我们圣灵作凭据 。
2COR|5|6|所以，我们总是勇敢的，并且知道，只要我们住在这身体内就是离开了主。
2COR|5|7|因为我们行事为人是凭着信心，不是凭着眼见。
2COR|5|8|我们勇敢，更情愿离开身体，与主同住。
2COR|5|9|所以，无论是住在身内或住在身外，我们都立了志向要得主的喜悦。
2COR|5|10|因为我们众人必须站在基督审判台前受审，为使各人按着本身所行的，或善或恶受报。
2COR|5|11|既然我们知道主是可畏的，就劝导人；但是上帝是认识我们的，我盼望你们的良心也认识我们。
2COR|5|12|我们不是向你们再推荐自己，而是要让你们有夸耀我们的机会，使你们好面对那凭外貌、不凭内心夸耀的人。
2COR|5|13|如果我们癫狂，是为上帝；如果我们清醒，是为你们。
2COR|5|14|原来基督的爱激励我们；因我们这样断定，一人既替众人死了，众人就都死了。
2COR|5|15|并且他替众人死，是叫那些活着的人不再为自己活，乃为替他们死而复活的主活。
2COR|5|16|所以，从今以后，我们不再按照人的看法来认识人，纵使我们曾经按照人的看法认识基督，如今却不再这样认识他了。
2COR|5|17|所以，若有人在基督里，他就是新造的人：旧事已过，都变成新的了。
2COR|5|18|一切都是出于上帝；他藉着基督使我们与他和好，又将劝人与他和好的使命赐给我们。
2COR|5|19|这就是：上帝在基督里使世人与自己和好，不将他们的过犯归到他们身上，并且将这和好的信息托付了我们。
2COR|5|20|所以，我们作基督的特使，就好像上帝藉我们劝你们一般。我们替基督求你们，与上帝和好吧！
2COR|5|21|上帝使那无罪 的，替我们成为罪，好使我们在他里面成为上帝的义。
2COR|6|1|我们与上帝同工的也劝你们，不可白受他的恩典；
2COR|6|2|因为他说： “在悦纳的时候，我应允了你； 在拯救的日子，我帮助了你。” 看哪，现在正是悦纳的时候！看哪，现在正是拯救的日子！
2COR|6|3|我们不在任何事上妨碍任何人，免得这使命被人毁谤；
2COR|6|4|反倒在各样的事上表明自己是上帝的用人：就如在持久的忍耐、患难、困苦、灾难、
2COR|6|5|鞭打、监禁、动乱、劳碌、失眠、饥饿、
2COR|6|6|廉洁、知识、坚忍、恩慈、圣灵的感化、无伪的爱心、
2COR|6|7|真实的言语、上帝的大能、藉着仁义的兵器在左在右、
2COR|6|8|荣誉或羞辱、恶名或美名。我们似乎是诱惑人的，却是诚实的；
2COR|6|9|似乎不为人所知，却是人所共知；似乎是死了，却是活着；似乎受惩罚，却没有被处死；
2COR|6|10|似乎忧愁，却常有喜乐；似乎贫穷，却使许多人富足；似乎一无所有，却样样都有。
2COR|6|11|哥林多 人哪，我们对你们，口是诚实的，心是宽宏的。
2COR|6|12|你们的狭窄不是由于我们，而是由于你们自己的心肠狭窄。
2COR|6|13|你们也要照样用宽宏的心报答我；我这话正像对自己的孩子说的。
2COR|6|14|你们不要和不信的人同负一轭。义和不义有什么相关？光明和黑暗有什么相连？
2COR|6|15|基督和 彼列 有什么相和？信主的和不信主的有什么相干？
2COR|6|16|上帝的殿和偶像有什么相同？因为我们是永生上帝的殿，就如上帝曾说： “我要在他们中间居住来往； 我要作他们的上帝， 他们要作我的子民。”
2COR|6|17|所以主说： “你们务要从他们中间出来， 跟他们分别； 不要沾不洁净的东西， 我就收纳你们。
2COR|6|18|我要作你们的父， 你们要作我的儿女。 这是全能的主说的。”
2COR|7|1|所以，亲爱的，既然我们有这样的应许，就当洁净自己，除去身体和灵魂一切的污秽，藉着敬畏上帝，得以成圣。
2COR|7|2|宽宏大量地接纳我们吧！我们未曾亏负谁，未曾败坏谁，未曾占谁的便宜。
2COR|7|3|我说这话，不是要定你们的罪，我已经说过，你们常在我们心里，我们情愿与你们同生共死。
2COR|7|4|我对你们很是放心，多多夸耀你们；我满有安慰，在我们一切患难中格外喜乐。
2COR|7|5|我们从前到了 马其顿 的时候，身体没有丝毫安宁，反而到处遭患难，外有纷争，内有惧怕。
2COR|7|6|但那安慰灰心之人的上帝藉着 提多 来安慰了我们；
2COR|7|7|不但藉着他来，也藉着他从你们所得的安慰安慰了我们，因为他把你们的思念，你们的哀恸，你们对我的热忱，都告诉了我，使我更加欢喜。
2COR|7|8|即使我先前那封信使你们忧愁，后来我曾懊悔，如今却不懊悔；因为我知道，那封信使你们忧愁，不过是暂时的。
2COR|7|9|如今我欢喜，不是因你们曾忧愁，而是因忧愁导致你们的悔改。你们依着上帝的意思忧愁，凡事就不至于因我们受亏损了。
2COR|7|10|因为依着上帝的意思而忧愁，就生出没有懊悔的悔改来，以致得救；但世俗的忧愁叫人死。
2COR|7|11|你看，你们依着上帝的意思而忧愁，这在你们当中产生了何等的殷勤、甚至辩白、甚至愤慨、甚至恐惧、甚至渴望、甚至热忱、甚至责罚。在这一切事上，你们都表明自己是无可指责的。
2COR|7|12|所以，虽然我从前写信给你们，却不是为那亏负人的，也不是为那受人亏负的，而是要在上帝面前把你们顾念我们的热忱表现出来。
2COR|7|13|因此，我们得了安慰。 在我们所得的安慰之外，又因你们众人使 提多 心里畅快喜乐，我们就更加欢喜了。
2COR|7|14|我若对 提多 夸奖过你们什么，也不觉得惭愧，因为我对 提多 夸奖你们的话是真的，正如我对你们所说的话也向来都是真的。
2COR|7|15|提多 一想起你们众人的顺服，怎样恐惧战兢地接待他，他爱你们的心就越发热切了。
2COR|7|16|我如今欢喜，因为我在一切事上对你们有信心。
2COR|8|1|弟兄们，我们要把上帝赐给 马其顿 众教会的恩惠告诉你们：
2COR|8|2|他们在患难中受大考验的时候，仍然满有喜乐，在极度贫穷中还格外显出他们乐捐的慷慨。
2COR|8|3|我可以证明，他们是按着能力，而且超过了能力来捐助，主动
2COR|8|4|再三恳求我们，准他们在这供给圣徒的善事上有份；
2COR|8|5|并且他们所做的，不但照我们所期望的，更照上帝的旨意先把自己献给主，又给了我们。
2COR|8|6|因此，我们劝 提多 ，既然在你们中间开始这慈善的事，就当把它办成。
2COR|8|7|既然你们在信心、口才、知识、万分的热忱，以及我们对你们 的爱心上，都胜人一等，那么，当在这慈善的事上也要胜人一等。
2COR|8|8|我说这话，并不是命令你们，而是藉着别人的热忱来考验你们爱心的真诚。
2COR|8|9|你们知道我们主耶稣基督的恩典：他本是富足，却为你们成了贫穷，好使你们因他的贫穷而成为富足。
2COR|8|10|我在这事上把我的意见告诉你们，是对你们有益，因为你们开始办这事，而且起此心意已经有一年了。
2COR|8|11|如今就当办成这事，既然有愿做的心，也当照你们所有的去办成。
2COR|8|12|因为人只要有愿做的心，必照他所有的蒙悦纳，并不是照他所没有的。
2COR|8|13|我不是要别人轻松，你们受累，而是要均匀：
2COR|8|14|就是要你们现在的富余补他们的不足，使他们的富余将来也可以补你们的不足，这就均匀了。
2COR|8|15|如经上所记： 多收的没有余， 少收的也没有缺。
2COR|8|16|感谢上帝，把我对你们的热忱同样放在 提多 心里。
2COR|8|17|他固然听了我的劝告，但自己更加热心，自愿往你们那里去。
2COR|8|18|我们还差遣一位弟兄和他同去，这人在传福音的事上得了众教会的称赞；
2COR|8|19|不但这样，他也被众教会选派跟我们同行，把所交托我们的这捐款送到了，为的是荣耀主，也表明我们的好意。
2COR|8|20|我们这样做，免得有人因我们收的捐款多而挑剔我们。
2COR|8|21|我们留心做好事，不但在主面前，就是在人面前也是这样。
2COR|8|22|我们又差遣一位弟兄同去。这人的热忱，我们在许多事上屡次考验过，现在他因为深深信任你们，就更加热心了。
2COR|8|23|至于 提多 ，他是我的伙伴，为服事你们作我的同工。至于那两位弟兄，他们是众教会的使者，是基督的荣耀。
2COR|8|24|所以，你们务要在众教会面前向他们显明你们的爱心和我所夸奖你们的凭据。
2COR|9|1|关于供给圣徒的事，我本来不必写信给你们；
2COR|9|2|因为我知道你们的好意，常对 马其顿 人夸奖你们，说 亚该亚 人预备好已经有一年了。你们的热心感动了许多人。
2COR|9|3|但我差遣那几位弟兄去，要使你们照我的话预备妥当，免得我们在这事上夸奖你们的话落了空。
2COR|9|4|万一有 马其顿 人与我同去，见你们没有预备好，就使我们所确信的反成了羞愧；你们的羞愧更不用说了。
2COR|9|5|因此，我想必须鼓励那几位弟兄先到你们那里去，把从前所应许的捐款预备妥当，好显出你们所捐的是出于乐意，不是出于勉强。
2COR|9|6|还有一点：“少种的少收；多种的多收。”
2COR|9|7|各人要随心所愿，不要为难，不要勉强，因为上帝爱乐捐的人。
2COR|9|8|上帝能将各样的恩惠多多加给你们，使你们凡事常常充足，能多做各样善事。
2COR|9|9|如经上所记： “他施舍，周济贫穷； 他的义行存到永远。”
2COR|9|10|那赐种子给撒种的，赐粮食给人吃的，必多多加给你们种地的种子，又增添你们仁义的果子。
2COR|9|11|你们必凡事富足，能多多施舍，使人藉着我们而生感谢上帝的心。
2COR|9|12|因为办这供给的事，不但补圣徒的缺乏，而且使许多人对上帝充满更多的感谢。
2COR|9|13|他们从这供给的事上得了凭据，知道你们宣认基督，顺服他的福音，慷慨捐助给他们和众人，把荣耀归给上帝。
2COR|9|14|他们也因上帝极大的恩赐显在你们身上而切切想念你们，为你们祈祷。
2COR|9|15|感谢上帝，因他有说不尽的恩赐！
2COR|10|1|我－ 保罗 与你们见面的时候是温和的，不在你们那里的时候向你们是勇敢的，如今亲自藉着基督的温柔和慈祥劝你们。
2COR|10|2|有人认为我们是凭着血气行事，我认为必须敢于对付这等人；我但求在那里的时候，不必这样勇敢。
2COR|10|3|我们虽然在血气中行事，却不凭着血气争战。
2COR|10|4|因为我们争战的兵器本不是属血气的，而是凭着上帝的能力，能够攻破坚固的营垒。我们攻破各样的计谋，
2COR|10|5|和各样拦阻人认识上帝的高垒，又夺回人心来顺服基督。
2COR|10|6|我已经预备好了，等你们完全顺服的时候来惩罚所有不顺服的人。
2COR|10|7|你们只看事情的外表。倘若有人自信是属基督的，他要再想想，他属基督，我们也属基督。
2COR|10|8|主赐给我们权柄，是要造就你们，并不是要拆毁你们；我就是为这权柄稍微夸口也不觉得惭愧。
2COR|10|9|我说这话，免得你们以为我写信是要恐吓你们。
2COR|10|10|因为有人说：“他信上的语气既严厉又强硬，他本人却软弱无能，言语粗俗。”
2COR|10|11|这等人当明白，我们不在那里时信上怎么说，见面时也必怎么做。
2COR|10|12|因为我们不敢将自己和某些自我推荐的人并列相比；他们用自己度量自己，用自己比较自己，是不明智的。
2COR|10|13|我们不愿意过分夸口，但是我们只在上帝划定的界限内夸口。这界限甚至扩展到你们那里。
2COR|10|14|我们扩展到你们那里时并没有越过了自己的界限，其实我们是首先到你们那里传基督福音的。
2COR|10|15|我们不靠别人所劳碌的过分夸口；我们只希望你们信心增长的时候，所划定给我们的范围也能够因着你们更加扩展，
2COR|10|16|使福音得以传到你们以外的地方，而不在别人的范围之内，以别人所成就的事夸口。
2COR|10|17|但“要夸耀的，该夸耀主”。
2COR|10|18|因为蒙悦纳的，不是自我称许的，而是主所称许的。
2COR|11|1|但愿你们容忍我小小的愚蠢；请你们务必容忍我。
2COR|11|2|我以上帝嫉妒的爱来爱你们，因为我曾把你们许配给一个丈夫，要把你们如同贞洁的童女献给基督。
2COR|11|3|我只怕你们的心偏邪了，失去那向基督所献诚恳贞洁 的心，就像蛇用诡诈诱惑了 夏娃 一样。
2COR|11|4|假如有人来，传另一个耶稣，不是我们所传过的；或者你们另受一个灵，不是你们所受过的圣灵；或者接纳另一个福音，不是你们所接纳过的；你们居然容忍了！
2COR|11|5|但我想，我一点也不在那些超级使徒以下。
2COR|11|6|虽然我不擅长说话，我的知识却不如此。这点我们已经在每一方面各样事上向你们表明了。
2COR|11|7|我贬低自己，为了使你们高升，因为我白白地传上帝的福音给你们，难道这算是我犯了错吗？
2COR|11|8|我剥夺了别的教会，向他们取了报酬来效劳你们。
2COR|11|9|我在你们那里有缺乏的时候，并没有连累你们一个人，因为我所缺乏的，那些从 马其顿 来的弟兄都补足了。我向来凡事谨慎，将来也必谨慎，总不要连累你们。
2COR|11|10|既有基督的真诚在我里面，在 亚该亚 一带地方就没有人能阻止我这样自夸。
2COR|11|11|为什么呢？是因我不爱你们吗？上帝知道，我爱你们！
2COR|11|12|我现在所做的，将来还要做，为要断绝那些寻机会之人的机会，不让他们在所夸耀的事上被人认为与我们一样。
2COR|11|13|那样的人是假使徒，行事诡诈，装作基督的使徒。
2COR|11|14|这也不足为奇，因为连撒但也装作光明的天使。
2COR|11|15|所以，他的差役若装作公义的差役也没有什么大不了。他们的结局必然跟他们的行为相符。
2COR|11|16|我再说，谁都不可把我看作愚蠢的；即使你们把我当作愚蠢人，那么，也让我稍微夸夸口吧。
2COR|11|17|我说的话不是奉主的权柄说的，而是像愚蠢人具有自信地放胆夸口。
2COR|11|18|既然有好些人凭着血气在夸口，我也要夸口了。
2COR|11|19|你们是聪明人，竟能甘心容忍愚蠢人！
2COR|11|20|假若有人奴役你们，或侵吞你们，或压榨你们，或侮辱你们，或打你们的脸，你们居然都能容忍。
2COR|11|21|说来惭愧，在这方面好像我们是太软弱了。 然而，我说句蠢话，人在什么事上敢夸口，我也敢夸口。
2COR|11|22|他们是 希伯来 人吗？我也是。他们是 以色列 人吗？我也是。他们是 亚伯拉罕 的后裔吗？我也是。
2COR|11|23|他们是基督的用人吗？我说句狂话，我更是。我比他们忍受更多劳苦，坐过更多次监牢，受过无数次的鞭打，常常冒死。
2COR|11|24|我被 犹太 人鞭打五次，每次四十减去一下；
2COR|11|25|被棍打了三次，被石头打了一次，遭海难三次，一昼一夜在深海里挣扎。
2COR|11|26|我又屡次行远路，遭江河的危险，盗贼的危险，同族人的危险，外族人的危险，城里的危险，旷野的危险，海中的危险，假弟兄的危险。
2COR|11|27|我劳碌困苦，常常失眠，又饥又渴，忍饥耐寒，赤身露体。
2COR|11|28|除了这些外表的事以外，我还有为众教会操心的事天天压在我身上。
2COR|11|29|有谁软弱，我不软弱呢？有谁跌倒，我不焦急呢？
2COR|11|30|我若必须夸口，就夸我软弱的事好了。
2COR|11|31|那永远可称颂之主耶稣的父上帝知道我不说谎。
2COR|11|32|在 大马士革 的 亚哩达 王手下的提督把守 大马士革城 ，要捉拿我，
2COR|11|33|我被人用筐子从城墙上的窗口缒下，逃脱了他的手。
2COR|12|1|虽然自夸无益，我还是不得不夸。我现在要提到主的异象和启示。
2COR|12|2|我认识一个在基督里的人，他在十四年前被提到第三层天上去；或在身内，我不知道，或在身外，我也不知道，只有上帝知道。
2COR|12|3|我认识的这样的一个人—或在身内，或在身外，我都不知道，只有上帝知道—
2COR|12|4|他被提到乐园里，听见隐秘的言语，是人不可说的。
2COR|12|5|为这人，我要夸口；但是为我自己，除了我的软弱以外，我并不夸口。
2COR|12|6|就是我愿意夸口也不算狂，因为我会说实话；只是我绝口不谈，恐怕有人把我看得太高了，过于他在我身上所看见所听见的；
2COR|12|7|又恐怕我因所得的启示太高深，就过于高抬自己，所以 有一根刺加在我身上，就是撒但的差役来折磨我，免得我过于高抬自己。
2COR|12|8|为了这事，我曾三次求主使这根刺离开我。
2COR|12|9|他对我说：“我的恩典是够你用的，因为我的能力是在人的软弱上显得完全。”所以，我更喜欢夸耀自己的软弱，好使基督的能力覆庇我。
2COR|12|10|为基督的缘故，我以软弱、凌辱、艰难、迫害、困苦为可喜乐的事；因为我什么时候软弱，什么时候就刚强了。
2COR|12|11|我成了愚蠢人，是被你们逼出来的，因为我本该被你们赞许才是。虽然我算不了什么，却没有一件事在那些超级使徒以下。
2COR|12|12|我在你们中间，用百般的忍耐，藉着神迹、奇事、异能显出使徒的凭据来。
2COR|12|13|除了我不曾连累你们这一件事，你们还有什么事不及别的教会呢？这不公平之处，请你们饶恕我吧。
2COR|12|14|如今，我准备第三次到你们那里去。我仍不会连累你们，因为我所求的是你们，不是你们的财物。儿女不该为父母积财，父母该为儿女积财。
2COR|12|15|我也甘心乐意为你们的灵魂费财费力。难道我越爱你们，就越少得你们的爱吗？
2COR|12|16|罢了，我自己并没有连累你们，你们却有人说，我施诡诈，用心计牢笼你们。
2COR|12|17|我所差遣到你们那里去的人，我何曾藉着他们中的任何人占过你们的便宜呢？
2COR|12|18|我劝 提多 到你们那里去，又差遣那位弟兄与他同去， 提多 占过你们的便宜吗？我们的行事为人不是同一心灵 吗？不是同一步伐吗？
2COR|12|19|你们一直认为我们是在你们面前为自己辩护吗？其实，我们本是在基督里当着上帝面前说话。亲爱的，一切的事都是为了造就你们。
2COR|12|20|我怕我再来的时候，见你们不合我所期望的，而你们见我也不合你们所期望的。我怕有纷争、嫉妒、愤怒、自私、毁谤、谗言、狂傲、动乱的事。
2COR|12|21|我怕我再来的时候，我的上帝使我在你们面前蒙羞，并且又因许多人从前犯罪，行污秽、淫乱、放荡的事，不肯悔改而悲伤。
2COR|13|1|这是我第三次要到你们那里去。“任何指控都要凭两个或三个证人的口述才能成立”。
2COR|13|2|对那些犯了罪的人和其余所有的人，正如我第二次见你们的时候曾说过，现在不在你们那里再次说：“我若再来，必不宽容。”
2COR|13|3|因为你们想求证基督是否藉着我说话。基督对你们并不是软弱的，而是在你们里面大有能力的。
2COR|13|4|他因软弱被钉在十字架上，却因上帝的大能仍然活着。我们在他里面也成为软弱的，但对你们，我们将因上帝的大能而与他一同活着。
2COR|13|5|你们总要省察自己是否在信仰中生活；你们要考验自己。除非你们经不起考验，你们自己岂不应该知道有耶稣基督在你们里面吗？
2COR|13|6|我希望你们知道，我们并不是经不起考验的人。
2COR|13|7|我们祈求上帝使你们不做任何恶事；这不是要显明我们是经得起考验的，而是要你们行事端正，即使我们似乎经不起考验也没有关系。
2COR|13|8|我们不能做任何对抗真理的事，只能维护真理。
2COR|13|9|当我们软弱而你们刚强时，我们也欢喜。我们所祈求的是：你们能成为完全人。
2COR|13|10|所以，我不在你们那里的时候，把这些话写给你们，好使我见你们的时候不用照主所给我的权柄严厉地待你们；这权柄原是为造就人，而不是为摧毁人。
2COR|13|11|末了，弟兄们，愿你们喜乐。要追求完全；要接受鼓励；要同心合意；要彼此和睦。如此，慈爱和平的上帝必与你们同在。
2COR|13|12|你们要用圣洁的吻彼此问安。众圣徒都向你们问安。
2COR|13|13|愿主耶稣基督的恩惠、上帝的慈爱、圣灵的感动常与你们众人同在！
GAL|1|1|我使徒 保罗 和所有跟我一起的弟兄，写信给 加拉太 的众教会。我作使徒不是由于人，也不是藉着人，而是藉着耶稣基督与使他从死人中复活的父上帝。
GAL|1|2|
GAL|1|3|愿恩惠、平安 从我们的父上帝和主耶稣基督归给你们！
GAL|1|4|基督照我们父上帝的旨意，为我们的罪舍己，要救我们脱离现今这罪恶的世代。
GAL|1|5|愿荣耀归给上帝，直到永永远远。阿们！
GAL|1|6|我很惊讶你们这么快就离开那位藉着基督之 恩呼召你们的上帝，而去随从别的福音；
GAL|1|7|其实并没有另一个福音，不过有些人骚扰你们，要把基督的福音更改了。
GAL|1|8|但无论是我们或是天上来的使者，若传福音给你们 ，与我们所传给你们的不同，他该受诅咒！
GAL|1|9|我们已经说了，现在我再说，若有人传福音给你们，与你们以往所领受的不同，他该受诅咒！
GAL|1|10|我现在是要得人的心，还是要得上帝的心呢？难道我在讨人的喜欢吗？我若仍旧想讨人的喜欢，我就不是基督的仆人了。
GAL|1|11|弟兄们，我要你们知道，我所传的福音不是按照人的意思；
GAL|1|12|因为我不是从人领受的，也不是人教导我的，而是藉着耶稣基督的启示而来。
GAL|1|13|你们听说过从前我在 犹太 教中的行径，我怎样竭力压迫残害上帝的教会。
GAL|1|14|在 犹太 教中，我比本国许多同辈的人更激进，为我祖宗的传统更热心。
GAL|1|15|然而，那位把我从母腹里分别出来、又施恩呼召我的上帝 ，既然乐意
GAL|1|16|把他儿子启示在我心里，让我在外邦人中传扬他，我就没有跟有血有肉的人商量，
GAL|1|17|也没有上 耶路撒冷 去见那些比我先作使徒的，惟独到 阿拉伯 去，后来又回到 大马士革 。
GAL|1|18|过了三年，我才上 耶路撒冷 去见 矶法 ，和他同住了十五天。
GAL|1|19|至于别的使徒，除了主的兄弟 雅各 ，我都没有见过。
GAL|1|20|我现在写给你们的是在上帝面前说的，不说谎话。
GAL|1|21|以后我到了 叙利亚 和 基利家 一带；
GAL|1|22|那时，在基督里的 犹太 各教会都没有见过我的面。
GAL|1|23|不过他们听说“那从前压迫我们的，现在竟传扬他原先所残害的信仰”。
GAL|1|24|他们就为我的缘故归荣耀给上帝。
GAL|2|1|过了十四年，我再上 耶路撒冷 去， 巴拿巴 同行，也带了 提多 一起去。
GAL|2|2|我是奉了启示上去的；我把在外邦人中所传的福音对弟兄们说明，我是私下对那些有名望的人说的，免得我现在或是从前都徒然奔跑了。
GAL|2|3|但跟我同去的 提多 ，虽是 希腊 人，也没有勉强他受割礼；
GAL|2|4|因为有偷着混进来的假弟兄，暗中窥探我们在基督耶稣里拥有的自由，要使我们作奴隶，
GAL|2|5|可是，为要使福音的真理仍存在你们中间，我们一点也没有让步顺服他们。
GAL|2|6|至于那些有名望的，不论他们是何等人，都与我无关；上帝不以外貌取人。那些有名望的，并没有加增我什么。
GAL|2|7|相反地，他们看见了主托付我传福音给未受割礼的人，正如主托付 彼得 传福音给受割礼的人；
GAL|2|8|那感动 彼得 、叫他为受割礼的人作使徒的，也感动我，叫我为外邦人作使徒。
GAL|2|9|那些被认为是教会柱石的 雅各 、 矶法 、 约翰 知道上帝所赐给我的恩典，就跟我和 巴拿巴 握右手以示合作，同意我们往外邦人那里去，他们往受割礼的人那里去。
GAL|2|10|他们只要求我们记念穷人，这也是我一向热心在做的。
GAL|2|11|后来， 矶法 到了 安提阿 ，因为他有可责之处，我就当面反对他。
GAL|2|12|从 雅各 那里来的人未到以前，他和外邦人一同吃饭，及至他们来到，他因怕奉割礼的人就退出，跟外邦人疏远了。
GAL|2|13|其余的 犹太 人也都随着他装假，甚至连 巴拿巴 也随伙装假。
GAL|2|14|但我一看见他们做得不对，与福音的真理不合，就在众人面前对 矶法 说：“你既是 犹太 人，却按照外邦人的样子，不按照 犹太 人的样子生活，怎么能勉强外邦人按照 犹太 人的样子生活呢？”
GAL|2|15|我们生来就是 犹太 人，不是外邦罪人；
GAL|2|16|可是我们知道，人称义不是因律法的行为，而是因信耶稣基督 ，我们也信了基督耶稣，为要使我们因信基督称义，不因律法的行为称义，因为，凡血肉之躯没有一个能因律法的行为称义。
GAL|2|17|我们若求在基督里称义，自己却还被视为罪人，那么，基督是罪的用人吗？绝对不是！
GAL|2|18|如果我重新建造我所拆毁的，这就证明自己是违犯律法的人。
GAL|2|19|我因律法而向律法死了，使我可以向上帝活着。我已经与基督同钉十字架，
GAL|2|20|现在活着的不再是我，乃是基督在我里面活着；并且我如今在肉身活着，是因信上帝的儿子而活；他是爱我，为我舍己。
GAL|2|21|我不废掉上帝的恩；如果义是藉着律法而获得，那么基督就白白死了。
GAL|3|1|无知的 加拉太 人哪，耶稣基督钉十字架，已经活现在你们眼前，谁又迷惑了你们呢？
GAL|3|2|这是我惟一要问你们的：你们领受了圣灵，是因律法的行为或是因听信福音呢？
GAL|3|3|你们既然以圣灵开始，如今竟要以肉身终结吗？你们是这样的无知吗？
GAL|3|4|你们受这么多的苦都是徒然的吗？如果真是徒然的，
GAL|3|5|那么，上帝赐给你们圣灵，又在你们中间行异能，是因律法的行为或是因听信福音呢？
GAL|3|6|正如 亚伯拉罕 “信了上帝，这就算他为义”。
GAL|3|7|所以，你们知道：有信心的人才是 亚伯拉罕 的子孙。
GAL|3|8|圣经既然预先看见上帝要使外邦人因信称义，预先传福音给 亚伯拉罕 ，说：“万国都必因你得福。”
GAL|3|9|可见，那有信心的人和有信心的 亚伯拉罕 一同得福。
GAL|3|10|凡出于律法的行为都是受诅咒的，因为经上记着：“凡不持守律法书上所记的一切而去行的，都是受诅咒的。”
GAL|3|11|没有一个人靠着律法在上帝面前称义，这是明显的，因为经上说：“义人必因信得生。”
GAL|3|12|律法并不出于信，而是说：“行这些事的就必因此得生。”
GAL|3|13|既然基督为我们成了诅咒，就把我们从律法的诅咒中赎出来。因为经上记着：“凡挂在木头上的都是受诅咒的。”
GAL|3|14|这是要使 亚伯拉罕 的福，因着基督耶稣临到外邦人，使我们能因信得着所应许的圣灵。
GAL|3|15|弟兄们，我照着人的观点说，人的遗嘱一经确定，没有人能废弃或加增。
GAL|3|16|那些应许原是向 亚伯拉罕 和他后裔说的，并不是说“和众后裔”，指许多人，而是说“和你那个后裔”，指一个人，就是基督。
GAL|3|17|我是这么说，上帝预先所立的约不能被四百三十年以后的律法废掉，使应许失效。
GAL|3|18|因为承受产业若是出于律法，就不再是出于应许；但上帝是凭着应许把产业赐给 亚伯拉罕 。
GAL|3|19|这样说来，为什么要有律法呢？律法是为过犯的缘故而加上去的，等候那蒙应许的子孙来到才结束，是藉着天使经中保之手而设立的。
GAL|3|20|但中保本不是为单方设立的；上帝却是一位。
GAL|3|21|这样，律法是与上帝的 应许对立吗？绝对不是！如果律法的颁布能使人得生命，义就诚然出于律法了。
GAL|3|22|但圣经把万物都圈在罪里，为要使因信耶稣基督 而来的应许归给信的人。
GAL|3|23|但这“信”还未来以前，我们被看守在律法之下，像被圈住，直到那将来的“信”显明出来。
GAL|3|24|这样，律法是我们的启蒙教师，直到基督来了 ，好使我们因信称义。
GAL|3|25|但这“信”既然来到，我们从此就不在启蒙教师的手下了。
GAL|3|26|其实，你们藉着信，在基督耶稣里都成为上帝的儿女。
GAL|3|27|你们凡受洗归入基督的都披戴基督了：
GAL|3|28|不再分 犹太 人或 希腊 人，不再分为奴的自主的，不再分男的女的，因为你们在基督耶稣里都成为一了。
GAL|3|29|既然你们属于基督，你们就是 亚伯拉罕 的子孙，是照着应许承受产业的了。
GAL|4|1|我说，虽然那承受产业的是整个产业的主人，但在未成年的时候却与奴隶毫无分别，
GAL|4|2|仍是在监护人和管家的手下，直等他父亲预定的时候来到。
GAL|4|3|我们也是一样，在未成年的时候，被世上粗浅的学说 所奴役，也是如此。
GAL|4|4|等到时候成熟，上帝就差遣他的儿子，为女子所生，且生在律法之下，
GAL|4|5|为要把律法之下的人赎出来，使我们获得儿子的名分。
GAL|4|6|因为你们是儿子，上帝就差他儿子的灵进入我们 的心，呼叫：“阿爸，父！”
GAL|4|7|可见，你不再是奴隶，而是儿子了，既然是儿子，就靠着上帝也成为后嗣了。
GAL|4|8|但从前不认识上帝的时候，你们是给那些本来不是上帝的神明作奴隶；
GAL|4|9|现在你们既然认识上帝，更可说是被上帝所认识的，怎么还要转回那懦弱无用的粗浅学说 ，情愿再给它们作奴隶呢？
GAL|4|10|你们竟又谨守日子、月份、节期、年份，
GAL|4|11|我为你们担心，惟恐我在你们身上是枉费工夫了。
GAL|4|12|弟兄们，我劝你们，要像我一样，因为我也像你们一样。你们一点没有亏负我。
GAL|4|13|你们知道，我因为身体有疾病才有第一次传福音给你们的机会。
GAL|4|14|虽然你们为我身体的缘故受试炼，却没有轻看我，也没有厌弃我，反倒接待我如同上帝的使者，如同基督耶稣。
GAL|4|15|你们当日的好意哪里去了呢？那时若办得到，你们就是把自己的眼睛挖出来给我，也都情愿。这是我可以给你们作证的。
GAL|4|16|如今我把真理告诉你们，倒成了你们的仇敌吗？
GAL|4|17|那些热心待你们的人，不怀好意，是要隔绝你们，好使你们热心待他们。
GAL|4|18|在善事上，时刻热心待别人原是好的，却不只是我与你们同在的时候才这样。
GAL|4|19|我的孩子们哪，我为你们再受生产之苦，直等到基督成形在你们心里 。
GAL|4|20|我期望现今就在你们那里，可以改变我的口气，因为我为你们心里难过。
GAL|4|21|你们这愿意在律法之下的人，请告诉我，你们没有听见律法吗？
GAL|4|22|因为律法上记着， 亚伯拉罕 有两个儿子，一个是使女生的，一个是自由的妇人生的。
GAL|4|23|那使女所生的是按着肉体生的；那自由的妇人所生的是凭着应许生的。
GAL|4|24|这是比方：那两个妇人就是两个约；一个妇人是出于 西奈山 ，生子为奴，就是 夏甲 。
GAL|4|25|这 夏甲 是指着 阿拉伯 的 西奈山 ，与现在的 耶路撒冷 同类，因为 耶路撒冷 和她的儿女都是为奴的。
GAL|4|26|但另一妇人就是在上的 耶路撒冷 ，是自由的，她是我们的母亲。
GAL|4|27|因为经上记着： 不怀孕、不生养的，你要欢乐； 未曾经过产难的，你要高声欢呼； 因为没有丈夫的，比有丈夫的有更多的儿女。
GAL|4|28|弟兄们，你们是凭着应许作儿女的，如同 以撒 一样。
GAL|4|29|当时，那按着肉体生的迫害了那按着圣灵生的，现在也是这样。
GAL|4|30|然而经上是怎么说的呢？是说：“把使女和她儿子赶出去！因为使女的儿子绝不能与自由妇人的儿子一同承受产业。”
GAL|4|31|弟兄们，这样看来，我们不是使女的儿女，而是自由妇人的儿女了。
GAL|5|1|基督释放了我们，为使我们得自由。所以要站稳了，不要再被奴隶的轭挟制。
GAL|5|2|我— 保罗 告诉你们，你们若受割礼，基督就对你们无益了。
GAL|5|3|我再指着凡受割礼的人确实地说，他有义务遵行全部的律法。
GAL|5|4|你们这要靠律法称义的是与基督隔绝，从恩典中坠落了。
GAL|5|5|至于我们，我们是靠着圣灵，凭着信心，等候所盼望的义。
GAL|5|6|因为在基督耶稣里，受割礼不受割礼都没有功效，惟独使人发出仁爱的信心才有功效。
GAL|5|7|你们向来跑得好，谁拦阻了你们，使你们不顺从真理呢？
GAL|5|8|这样的劝导不是出于那召你们的。
GAL|5|9|一点面酵能使全团都发起来。
GAL|5|10|我在主里深信你们必不怀别样的心；但骚扰你们的，无论是谁，必须承受惩罚。
GAL|5|11|弟兄们，我若仍旧传割礼，为什么还受迫害呢？若是这样，十字架绊倒人的地方就没有了。
GAL|5|12|恨不得那骚扰你们的人把自己阉割了。
GAL|5|13|弟兄们，你们蒙召是要得自由；只是不可把这自由当作放纵情欲的机会，总要用爱心互相服侍。
GAL|5|14|因为全部律法都包括在“爱邻 如己”这一句话之内了。
GAL|5|15|你们要谨慎，你们若相咬相吞，恐怕要彼此消灭了。
GAL|5|16|我说，你们要顺着圣灵而行，绝不可满足肉体的情欲。
GAL|5|17|因为肉体的情欲和圣灵相争，圣灵和肉体相争，这两个彼此敌对，使你们不能做所愿意做的。
GAL|5|18|但你们若被圣灵引导，就不在律法之下。
GAL|5|19|情欲的事都是显而易见的；就如淫乱、污秽、放荡、
GAL|5|20|拜偶像、行邪术、仇恨、纷争、忌恨、愤怒、自私、分派、结党、
GAL|5|21|嫉妒 、醉酒、荒宴等类。我从前告诉过你们，现在又告诉你们，做这样事的人必不能承受上帝的国。
GAL|5|22|圣灵的果子就是仁爱、喜乐、和平、忍耐、恩慈、良善、信实、
GAL|5|23|温柔、节制。这样的事没有律法禁止。
GAL|5|24|凡属基督耶稣 的人，是已经把肉体与肉体的邪情私欲同钉在十字架上了。
GAL|5|25|我们若靠着圣灵而活，也要靠着圣灵行事。
GAL|5|26|不要贪图虚名，彼此惹气，互相嫉妒。
GAL|6|1|弟兄们，若有人偶然被过犯所胜，你们属灵的人就要用温柔的心把他挽回过来；自己也要留意，免得也被引诱。
GAL|6|2|你们各人的重担要互相担当，这样就会成全 基督的律法。
GAL|6|3|人若没有什么了不起，还自以为了不起的，就是自欺。
GAL|6|4|各人要省察自己的行为；这样，他所夸口的只在自己，而不在别人。
GAL|6|5|因为人人必须担当自己的担子。
GAL|6|6|在真道上受教的，要把一切美好的东西与施教的人分享。
GAL|6|7|不要自欺；上帝是轻慢不得的，因为人种的是什么，收的也是什么。
GAL|6|8|顺着肉体撒种的，必从肉体收败坏；顺着圣灵撒种的，必从圣灵收永生。
GAL|6|9|我们行善不可丧志，因为若不灰心，到了适当的时候就有收成。
GAL|6|10|所以，一有机会就要向众人行善，向信徒一家的人更要这样。
GAL|6|11|你们看我亲手写给你们的字是何等的大！
GAL|6|12|那些想要炫耀外表的人才勉强你们受割礼，无非是怕自己为基督的十字架受迫害。
GAL|6|13|他们那些受割礼的，连自己也不守律法；他们要你们受割礼，不过是要拿你们的肉体夸口。
GAL|6|14|但我绝不以别的夸口，只夸我们主耶稣基督的十字架；因这十字架 ，就我而论，世界已经钉在十字架上；就世界而论，我已经钉在十字架上。
GAL|6|15|受割礼或不受割礼都无关紧要，要紧的就是作新造的人。
GAL|6|16|凡照这准则行的人，愿平安 怜悯，加给他们，和上帝的 以色列 民。
GAL|6|17|从今以后，不要有人再搅扰我，因为我身上带着耶稣的印记。
GAL|6|18|弟兄们，愿我们主耶稣基督的恩与你们的灵同在。阿们！
EPH|1|1|奉上帝旨意作基督耶稣使徒的 保罗 ，写信给在 以弗所 的 众圣徒，就是在基督耶稣里忠心的人。
EPH|1|2|愿恩惠、平安 从我们的父上帝和主耶稣基督归给你们！
EPH|1|3|愿颂赞归给我们主耶稣基督的父上帝。他在基督里曾把天上各样属灵的福气赐给我们。
EPH|1|4|因为他从创世以前，在基督里拣选了我们，使我们在他面前成为圣洁，没有瑕疵，满有爱心。
EPH|1|5|他按着自己旨意所喜悦的 ，预定我们藉着耶稣基督得儿子的名分，
EPH|1|6|使他荣耀的恩典得到称赞；这恩典是他在爱子里白白赐给我们的。
EPH|1|7|我们藉着这爱子的血得蒙救赎，过犯得以赦免，这是照他丰富的恩典，
EPH|1|8|充充足足地赏给我们的。他以诸般的智慧聪明，
EPH|1|9|照自己在基督里所立定的美意，使我们知道他旨意的奥秘，
EPH|1|10|要照着所安排的，在时机成熟的时候，使天上、地上、一切所有的，都在基督里面同归于一。
EPH|1|11|我们也在他里面得了基业；这原是那位随己意行万事的上帝照着自己的旨意所预定的，
EPH|1|12|为要使我们，这些首先把希望寄托在基督里的人，颂赞他的荣耀。
EPH|1|13|在基督里你们听见真理的道，就是那使你们得救的福音，你们也信了他，就受了所应许的圣灵为印记。
EPH|1|14|这圣灵是我们得基业的凭据，直等到上帝的子民得救赎，使他的荣耀得到称赞。
EPH|1|15|因此，我既然听见你们对主耶稣有信心，对众圣徒有爱心，
EPH|1|16|就不住地为你们感谢上帝，祷告的时候常常提到你们，
EPH|1|17|求我们主耶稣基督的上帝，荣耀的父，把那赐人智慧和启示的灵赐给你们，使你们真正认识他，
EPH|1|18|照亮你们心中的眼睛，使你们知道他呼召你们来得的指望是什么，他在圣徒中所得荣耀的基业是何等丰盛，
EPH|1|19|并知道他向我们这些信的人所显的能力是何等浩大，这是照他的大能大力运行的。
EPH|1|20|这大能曾运行在基督身上，使他从死人中复活，又使他在天上坐在自己的右边，
EPH|1|21|远超越一切执政的、掌权的、有权能的、统治的和一切有名号的；不但是今世的，连来世的也都超越了。
EPH|1|22|上帝使万有服在他的脚下，又使他为了教会作万有之首；
EPH|1|23|教会是他的身体，是那充满万有者所充满的。
EPH|2|1|从前，你们因着自己的过犯罪恶而死了。
EPH|2|2|那时，你们在过犯罪恶中生活，随从今世的风俗，顺服空中掌权者的领袖，就是现今在悖逆的人心中运行的邪灵。
EPH|2|3|我们从前也都生活在他们当中，放纵肉体的私欲，随着肉体和心中的意念去做，和别人一样，生来就是该受惩罚的人。
EPH|2|4|然而，上帝有丰富的怜悯，因着他爱我们的大爱，
EPH|2|5|竟在我们因过犯而死了的时候，使我们与基督一同活过来—可见你们得救是本乎恩—
EPH|2|6|他又使我们在基督耶稣里与他一同复活，一同坐在天上，
EPH|2|7|为要把他极丰富的恩典，就是他在基督耶稣里向我们所施的恩慈，显明给后来的世代。
EPH|2|8|你们得救是本乎恩，也因着信；这并不是出于自己，而是上帝所赐的；
EPH|2|9|也不是出于行为，免得有人自夸。
EPH|2|10|我们是他所造之物，在基督耶稣里创造的，为要使我们行善，就是上帝早已预备好要我们做的。
EPH|2|11|所以，你们要记得：从前你们按肉体是外邦人，是“没受割礼的”；这名字是那些凭人手在肉身上“受割礼的人”所取的。
EPH|2|12|要记得那时候，你们与基督无关，与 以色列 选民团体隔绝，在所应许的约上是局外人，而且在世上没有指望，没有上帝。
EPH|2|13|从前你们是远离上帝的人，如今却在基督耶稣里，靠着他的血，已经得以亲近了。
EPH|2|14|因为他自己是我们的和平 ，使双方合而为一，拆毁了中间隔绝的墙，而且以自己的身体终止了冤仇，
EPH|2|15|废掉那记在律法上的规条，为要使两方藉着自己造成一个新人，促成了和平；
EPH|2|16|既在十字架上消灭了冤仇，就藉这十字架使双方归为一体，与上帝和好，
EPH|2|17|并且来传和平的福音给你们远处的人，也传和平给那些近处的人，
EPH|2|18|因为我们双方藉着他，在同一位圣灵里得以进到父面前。
EPH|2|19|这样，你们不再是外人或客旅，是与圣徒同国，是上帝家里的人了，
EPH|2|20|被建造在使徒和先知的根基上，而基督耶稣自己为房角石，
EPH|2|21|靠着他整座房子连接得紧凑，渐渐成为在主里的圣殿。
EPH|2|22|你们也靠他同被建造，成为上帝藉着圣灵居住的所在。
EPH|3|1|因此，我— 保罗 为你们外邦人作了基督耶稣 囚徒的，替你们祈祷 。
EPH|3|2|想你们必曾听见上帝赐恩给我，把关切你们的职分托付我，
EPH|3|3|用启示让我知道福音的奥秘，正如我以前略略写过的。
EPH|3|4|你们读了，就会知道我深深了解基督的奥秘；
EPH|3|5|这奥秘在以前的世代没有让人知道，像如今藉着圣灵向他的圣使徒和先知启示一样，
EPH|3|6|就是外邦人在基督耶稣里，藉着福音，得以同为后嗣，同为一体，同为蒙应许的人。
EPH|3|7|我作了这福音的仆役，是照着上帝的恩赐，是照他运行的大能赐给我的。
EPH|3|8|虽然我比众圣徒中最小的还小，他还赐我这恩典，让我把基督那测不透的丰富传给外邦人，
EPH|3|9|又使众人都明白 什么是历代以来隐藏在创造万物之上帝里的奥秘，
EPH|3|10|为要在现今藉着教会使天上执政的、掌权的知道上帝百般的智慧。
EPH|3|11|这是照着上帝在我们主基督耶稣里所完成的永恒的计划。
EPH|3|12|我们因信耶稣 ，就在他里面放胆无惧，满有自信地进到上帝面前。
EPH|3|13|所以我求你们，不要因我为你们所受的患难丧胆；这原是你们的光荣。
EPH|3|14|因此，我在父面前屈膝—
EPH|3|15|天上地上的各家都是从他得名的－
EPH|3|16|为要他按着他丰盛的荣耀，藉着他的灵，使你们内心的力量刚强起来；
EPH|3|17|又要他使基督因着你们的信住在你们心里，使你们既在爱中生根立基，
EPH|3|18|能够和众圣徒一同明白基督的爱是何等的长、阔、高、深，并知道这爱是超过人的知识所能测度的，为要使你们充满上帝一切的丰盛。
EPH|3|19|
EPH|3|20|上帝能照着运行在我们心里的大能充充足足地成就一切，超过我们所求所想的。
EPH|3|21|愿他在教会中，并在基督耶稣里，得着荣耀，直到世世代代，永永远远。阿们！
EPH|4|1|我为主作囚徒的劝你们，既然蒙召，行事为人就要与你们所蒙的呼召相称。
EPH|4|2|凡事要谦虚、温柔、忍耐，用爱心互相宽容，
EPH|4|3|以和平彼此联系，竭力保持圣灵所赐的合一。
EPH|4|4|身体只有一个，圣灵只有一位，正如你们蒙召，是为同有一个指望而蒙召，
EPH|4|5|一主，一信，一洗，
EPH|4|6|一上帝－就是万人之父，超越万有之上，贯通万有，在万有之中。
EPH|4|7|我们每个人蒙恩都是照基督所量给每个人的恩赐。
EPH|4|8|所以有话说： “他升上高天的时候，掳掠了俘虏， 将各样的恩赐赏给人。”
EPH|4|9|既说“他升上”，岂不是指他曾降到地底下吗？
EPH|4|10|那降下的，就是高升远超越诸天之上的，为要充满万有。
EPH|4|11|他所赐的有使徒，有先知，有传福音的，有牧者和教师，
EPH|4|12|为要装备圣徒，做事奉的工作，建立基督的身体，
EPH|4|13|直等到我们众人在信仰上同归于一，认识上帝的儿子，得以长大成人，达到基督完全长成的身量。
EPH|4|14|这样，我们不再作小孩子，中了人的诡计和欺骗的法术，被一切邪说之风摇动，飘来飘去。
EPH|4|15|我们反而要用爱心说诚实话，各方面向着基督长进，连于元首基督，
EPH|4|16|靠着他全身都连接得紧凑，百节各按各职，照着各体的功用彼此相助，使身体渐渐增长，在爱中建立自己。
EPH|4|17|所以我这样说，且在主里郑重地说，你们行事为人，不要再像外邦人存虚妄的心而活。
EPH|4|18|他们心地昏昧，因自己无知，心里刚硬而与上帝所赐的生命隔绝了。
EPH|4|19|既然他们已经麻木，就放纵情欲，贪婪地行种种污秽的事。
EPH|4|20|但你们从基督学的不是这样。
EPH|4|21|如果你们听过他的道，领了他的教，因为真理就在耶稣里，
EPH|4|22|你们要脱去从前的行为，脱去旧我；这旧我是因私欲的迷惑而渐渐败坏的。
EPH|4|23|你们要把自己的心志更新，
EPH|4|24|并且穿上新我；这新我是照着上帝的形像造的，有从真理来的公义和圣洁。
EPH|4|25|所以，你们要弃绝谎言，每个人要与邻舍说诚实话，因为我们是互为肢体。
EPH|4|26|即使生气也不要犯罪；不可含怒到日落，
EPH|4|27|不可给魔鬼留地步。
EPH|4|28|偷窃的，不要再偷；总要勤劳，亲手 做正当的事，这样才可以把自己有的，分给有缺乏的人。
EPH|4|29|一句坏话也不可出口，只要随着需要说造就人的好话，让听见的人得益处。
EPH|4|30|不要使上帝的圣灵担忧，你们原是受了他的印记，等候得救赎的日子来到。
EPH|4|31|一切苦毒、愤怒、恼恨、嚷闹、毁谤，和一切的恶毒都要从你们中间除掉。
EPH|4|32|要仁慈相待，存怜悯的心，彼此饶恕，正如上帝在基督里饶恕了你们一样。
EPH|5|1|所以，作为蒙慈爱的儿女，你们该效法上帝。
EPH|5|2|要凭爱心行事，正如基督爱我们，为我们舍了自己，当作馨香的供物和祭物献给上帝。
EPH|5|3|至于淫乱和一切污秽，或是贪婪，在你们中间连提都不可，这才合乎圣徒的体统。
EPH|5|4|淫词、妄语和粗俗的俏皮话都不合宜；总要说感谢的话。
EPH|5|5|要确实知道，无论是淫乱的，是污秽的，是贪心的（贪心的就是拜偶像的），在基督和上帝的国里都得不到基业。
EPH|5|6|不要被人虚浮的话欺骗了，因这些事，上帝的愤怒必临到那些悖逆的人。
EPH|5|7|所以，不要与他们同伙。
EPH|5|8|从前你们是暗昧的，但如今在主里面是光明的，行事为人要像光明的子女—
EPH|5|9|光明所结的果子就是一切的良善、公义、诚实。
EPH|5|10|总要察验什么是主所喜悦的事。
EPH|5|11|那暗昧无益的事，不可参与，倒要把这种事揭发出来。
EPH|5|12|因为，他们暗中所做的，就是连提起来都是可耻的。
EPH|5|13|凡被光所照明的都显露出来，
EPH|5|14|因为使一切显露出来的就是光。所以有话说： “你这睡着的人醒过来吧！ 要从死人中复活， 基督要光照你了。”
EPH|5|15|你们要谨慎行事，不要像无知的人，要像智慧的人。
EPH|5|16|要把握时机 ，因为现今的世代邪恶。
EPH|5|17|不要作糊涂人，要明白主的旨意如何。
EPH|5|18|不要醉酒，酒能使人放荡；要被圣灵充满。
EPH|5|19|要用诗篇、赞美诗、灵歌彼此对说，口唱心和地赞美主。
EPH|5|20|凡事要奉我们主耶稣基督的名常常感谢父上帝。
EPH|5|21|要存敬畏基督的心彼此顺服。
EPH|5|22|作妻子的，你们要顺服自己的丈夫，如同顺服主。
EPH|5|23|因为丈夫是妻子的头，如同基督是教会的头；他又是这身体的救主。
EPH|5|24|教会怎样顺服基督，妻子也要怎样凡事顺服丈夫。
EPH|5|25|作丈夫的，你们要爱自己的妻子，正如基督爱教会，为教会舍己，
EPH|5|26|以水藉着道把教会洗净，使她成为圣洁，
EPH|5|27|好献给自己，作荣耀的教会，毫无玷污、皱纹等类的缺陷，而是圣洁没有瑕疵的。
EPH|5|28|丈夫也应当照样爱妻子，如同爱自己的身体；爱妻子就是爱自己了。
EPH|5|29|从来没有人恨恶自己的身体，总是保养爱惜，正像基督待教会一样，
EPH|5|30|因我们是他身体的肢体。
EPH|5|31|“为这个缘故，人要离开父母，与妻子结合，二人成为一体。”
EPH|5|32|这是极大的奥秘，而我是指基督和教会说的。
EPH|5|33|然而，你们每个人都要爱妻子，如同爱自己一样；妻子也要敬重她的丈夫。
EPH|6|1|作儿女的，你们要在主里 听从父母，这是理所当然的。
EPH|6|2|当孝敬父母，使你得福，在世长寿。这是第一条带应许的诫命。
EPH|6|3|
EPH|6|4|作父亲的，你们不要激怒儿女，但要照着主的教导和劝戒养育他们。
EPH|6|5|作仆人的，你们要惧怕战兢，用诚实的心听从你们肉身的主人，好像听从基督一般；
EPH|6|6|不要只在人的眼前这样做，像仅是讨人的喜欢，而是作基督的仆人，从心里遵行上帝的旨意，
EPH|6|7|甘心服侍，好像服侍主，不像服侍人，
EPH|6|8|因为知道每个人所做的善事，不论是为奴的或是自主的，都必按所做的从主得到赏赐。
EPH|6|9|作主人的，你们待仆人也是一样，不要威吓他们，因为知道他们和你们在天上同有一位主，他并不偏待人。
EPH|6|10|最后，你们要靠着主，依赖他的大能大力作刚强的人。
EPH|6|11|要穿戴上帝所赐的全副军装，好抵挡魔鬼的诡计。
EPH|6|12|因为我们的争战并不是对抗有血有肉的人，而是对抗那些执政的、掌权的、管辖这幽暗世界的，以及天空灵界的恶魔。
EPH|6|13|所以，要拿起上帝所赐的全副军装，好在邪恶的日子能抵挡仇敌，并且完成了一切后还能站立得住。
EPH|6|14|所以，要站稳了，用真理当作带子束腰，用公义当作护心镜遮胸，
EPH|6|15|又用和平的福音当作预备走路的鞋穿在脚上。
EPH|6|16|此外，要拿信德当作盾牌，用来扑灭那恶者一切烧着的箭。
EPH|6|17|要戴上救恩的头盔，拿着圣灵的宝剑—就是上帝的道。
EPH|6|18|要靠着圣灵，随时多方祷告祈求，并要为此警醒不倦，为众圣徒祈求。
EPH|6|19|也要为我祈求，让我有口才，能放胆开口讲明福音的奥秘，
EPH|6|20|我为这福音的奥秘作了带铁链的使者，让我能照着当尽的本分放胆宣讲。
EPH|6|21|今有亲爱、忠心服事主的弟兄 推基古 ，为了你们也明白我的事情和我的景况，他会让你们知道一切的事。
EPH|6|22|我特意打发他到你们那里去，好让你们知道我们的情况，又让他安慰你们的心。
EPH|6|23|愿平安 、慈爱、信心从父上帝和主耶稣基督归给弟兄们。
EPH|6|24|愿所有恒心爱我们主耶稣基督的人都蒙恩惠。
PHIL|1|1|基督耶稣的仆人 保罗 和 提摩太 写信给住 腓立比 、在基督耶稣里的众圣徒，以及诸位监督和执事。
PHIL|1|2|愿恩惠、平安 从我们的父上帝和主耶稣基督归给你们！
PHIL|1|3|我每逢想念你们，就感谢我的上帝，
PHIL|1|4|每逢为你们众人祈求的时候，总是欢欢喜喜地祈求，
PHIL|1|5|因为从第一天直到如今，你们都同心合意兴旺福音。
PHIL|1|6|我深信，那在你们心里动了美好工作的，到了耶稣基督的日子必完成这工作。
PHIL|1|7|我为你们众人有这样的想法原是应当的，因为你们常在我心里；无论我是在捆锁中，在辩明并证实福音的时候，你们都与我一同蒙恩。
PHIL|1|8|我以基督耶稣的心肠切切想念你们众人，这是上帝可以为我作证的。
PHIL|1|9|我所祷告的就是：要你们的爱心，在知识和各样见识上，不断增长，
PHIL|1|10|使你们能分辨是非，在基督的日子作真诚无可指责的人，
PHIL|1|11|更靠着耶稣基督结满仁义的果子，归荣耀称赞给上帝。
PHIL|1|12|弟兄们，我要你们知道，我所遭遇的事反而使福音更兴旺，
PHIL|1|13|以致御营全军和其余的人都知道我是为基督的缘故受捆锁的；
PHIL|1|14|而且那在主里的弟兄，多半都因我受的捆锁而笃信不疑，越发放胆无所惧怕地传道。
PHIL|1|15|有些人传基督是出于嫉妒纷争；有些人是出于好意。
PHIL|1|16|后者是出于爱心，知道我奉差遣是为福音辩护的。
PHIL|1|17|前者传基督是出于自私，动机不纯，企图要加增我捆锁的苦楚。
PHIL|1|18|这又何妨呢？或是假意或是真心，无论如何，只要基督被传开了，为此我就欢喜。 我还要欢喜，
PHIL|1|19|因为我知道，这事藉着你们的祈祷和耶稣基督的灵的帮助，终必使我得到释放。
PHIL|1|20|这就是我所切慕、所盼望的：没有一事能使我羞愧；反倒凡事坦然无惧，无论是生是死，总要让基督在我身上照常显大。
PHIL|1|21|因为我活着就是基督，死了就有益处。
PHIL|1|22|但是，我在肉身活着，若能有工作的成果，我就不知道该挑选什么。
PHIL|1|23|我处在两难之间：我情愿离世与基督同在，因为这是好得无比的；
PHIL|1|24|然而，我为你们肉身活着更加要紧。
PHIL|1|25|既然我这样深信，就知道仍要留在世间，且与你们众人一起存留，使你们在所信的道上又长进又喜乐，
PHIL|1|26|为了我再到你们那里时，你们在基督耶稣里的夸耀越发加增。
PHIL|1|27|最重要的是：你们行事为人要与基督的福音相称，这样，无论我来见你们，或不在你们那里，都可以听到你们的景况，知道你们同有一个心志，站立得稳，为福音的信仰齐心努力，
PHIL|1|28|丝毫不怕敌人的威胁；以此证明他们会沉沦，你们会得救，这是出于上帝。
PHIL|1|29|因为你们蒙恩，不但得以信服基督，而且要为他受苦。
PHIL|1|30|你们的争战，就与你们曾在我身上见过、现在所听到的是一样的。
PHIL|2|1|所以，在基督里若有任何劝勉，若有任何爱心的安慰，若有任何圣灵的团契，若有任何慈悲怜悯，
PHIL|2|2|你们就要意志相同，爱心相同，有一致的心思，一致的想法，使我的喜乐得以满足。
PHIL|2|3|凡事不可自私自利，不可贪图虚荣；只要心存谦卑，各人看别人比自己强。
PHIL|2|4|各人不要单顾自己的事，也要顾别人的事。
PHIL|2|5|你们当以基督耶稣的心为心：
PHIL|2|6|他本有上帝的形像， 却不坚持自己与上帝同等 ；
PHIL|2|7|反倒虚己， 取了奴仆的形像， 成为人的样式； 既有人的样子，
PHIL|2|8|就谦卑自己， 存心顺服，以至于死， 且死在十字架上。
PHIL|2|9|所以上帝把他升为至高， 又赐给他超乎万名之上的名，
PHIL|2|10|使一切在天上的、地上的和地底下的， 因耶稣的名， 众膝都要跪下，
PHIL|2|11|众口都要宣认： 耶稣基督是主， 归荣耀给父上帝。
PHIL|2|12|我亲爱的，这样看来，你们向来是顺服的，不但我在你们那里，就是我现在不在你们那里的时候更是顺服的，就当恐惧战兢完成你们自己得救的事；
PHIL|2|13|因为是上帝在你们心里运行，使你们又立志又实行，为要成就他的美意。
PHIL|2|14|你们无论做什么事，都不要发怨言起争论，
PHIL|2|15|好使你们无可指责，诚实无伪，在这弯曲悖谬的世代作上帝无瑕疵的儿女。你们在这世代中要像明光照耀，
PHIL|2|16|将生命的道显明出来，使我在基督的日子得以夸耀我没有白跑，也没有徒劳。
PHIL|2|17|我以你们的信心为供献的祭物，我若被浇献在其上也是喜乐，并且与你们众人一同喜乐。
PHIL|2|18|你们也要照样喜乐，并且与我一同喜乐。
PHIL|2|19|我靠主耶稣希望很快能差 提摩太 去见你们，好让我知道你们的事而心里得着安慰。
PHIL|2|20|因为我没有别人与我同心，真正关怀你们的事。
PHIL|2|21|其他的人都求自己的事，并不求耶稣基督的事。
PHIL|2|22|但你们知道 提摩太 是经得起考验的，他与我为了福音一同服侍，待我像儿子待父亲一样。
PHIL|2|23|所以，我一看出我的事怎样了结，我希望立刻差他去，
PHIL|2|24|但我靠着主自信我不久也会去。
PHIL|2|25|然而，我想必须差 以巴弗提 到你们那里去。他是我的弟兄、同工和战友，是你们差遣来供应我需要的。
PHIL|2|26|他很想念 你们众人，并且极其难过，因为你们听见他病了。
PHIL|2|27|他真的生病了，几乎要死。然而上帝怜悯他，不但怜悯他，也怜悯我，免得我忧上加忧。
PHIL|2|28|所以，我更要尽快送他回去，好让你们再见到他而喜乐，我也可以减少忧愁。
PHIL|2|29|故此，你们要在主里欢欢喜喜地接待他，而且要尊重这样的人，
PHIL|2|30|因他为做基督的工作不顾性命，几乎至死，为要补足你们供应我不够的地方。
PHIL|3|1|末了，我的弟兄们，你们要靠主喜乐。我把这些话再写给你们，对我并不困难，对你们却是妥当的。
PHIL|3|2|应当防备犬类，防备作恶的，防备妄自行割的。
PHIL|3|3|因为真受割礼的，就是我们这藉着上帝的灵敬拜、以基督耶稣为夸耀、不依靠肉体的。
PHIL|3|4|其实，我也可以靠肉体；若是别人以为他可以依靠肉体，我更可以。
PHIL|3|5|我出生后第八天受割礼；我是 以色列 族、 便雅悯 支派的人，是 希伯来 人所生的 希伯来 人。就律法说，我是法利赛人；
PHIL|3|6|就热心说，我是迫害教会的；就律法上的义说，我是无可指责的。
PHIL|3|7|只是我先前以为对我是有益的，我现在因基督的缘故而当作是有损的。
PHIL|3|8|不但如此，我已把万事当作是有损的，因我以认识我主基督耶稣为至宝。我为他已经丢弃万事，看作粪土，为要赢得基督，
PHIL|3|9|并且得以在他里面，不是有自己因律法而得的义，而是有信基督的义 ，就是基于信，从上帝而来的义，
PHIL|3|10|使我认识基督，知道他复活的大能，并且知道和他一同受苦，效法他的死，
PHIL|3|11|或许我也得以从死人中复活。
PHIL|3|12|这不是说我已经得着了，已经完全了；而是竭力追求，或许可以得着基督耶稣 所要我得着的 。
PHIL|3|13|弟兄们，我不是以为自己已经得着了；我只有一件事，就是忘记背后，努力面前的，
PHIL|3|14|向着标竿直跑，要得上帝在基督耶稣里从上面召我来得的奖赏。
PHIL|3|15|所以，我们中间凡是成熟的人，总要存这样的心；若在什么事上存别样的心，上帝也会把这些事指示你们。
PHIL|3|16|然而，我们达到什么地步，就当照这个地步行。
PHIL|3|17|弟兄们，你们要一同效法我，也当留意看那些效法我们榜样的人。
PHIL|3|18|因为，我屡次告诉你们，现在又流泪告诉你们：许多人行事是基督十字架的仇敌。
PHIL|3|19|他们的结局就是灭亡。他们的神明是自己的肚腹；他们以自己的羞辱为光荣，专以地上的事为念。
PHIL|3|20|我们却是天上的国民，并且等候救主，就是主耶稣基督从天上降临。
PHIL|3|21|他要按着那能使万有归服自己的大能，把我们这卑贱的身体改变形状，和他自己荣耀的身体相似。
PHIL|4|1|我所亲爱、所想念的弟兄们，你们就是我的喜乐，我的冠冕。我亲爱的，你们应当靠主站立得稳。
PHIL|4|2|我劝 友阿蝶 和 循都基 要在主里同心。
PHIL|4|3|我也求你这真实同负一轭的，要帮助这两个女人，因为她们在福音上曾与我、 革利免 和我其余的同工一同劳苦，他们的名字都在生命册上。
PHIL|4|4|你们要靠主常常喜乐。我再说，你们要喜乐。
PHIL|4|5|要让众人知道你们谦让的心。主已经近了。
PHIL|4|6|应当一无挂虑，只要凡事藉着祷告、祈求和感谢，将你们所要的告诉上帝。
PHIL|4|7|上帝所赐那超越人所能了解的平安 ，必在基督耶稣里，保守你们的心怀意念。
PHIL|4|8|末了，弟兄们，凡是真实的、凡是可敬的、凡是公义的、凡是清洁的、凡是可爱的、凡是有美名的，若有什么德行，若有什么称赞，你们都要留意。
PHIL|4|9|你们从我所学习的，所领受的，所听见的，所看见的事，你们都要继续去做，赐平安的上帝就必与你们同在。
PHIL|4|10|我靠主大大喜乐，因为你们关怀我的心如今又表现了出来；其实你们一直都关怀我，只是没有机会罢了。
PHIL|4|11|我并不是因缺乏而说这话，因为我已经学会无论在什么景况都可以知足。
PHIL|4|12|我知道怎样处卑贱，也知道怎样处丰富；或饱足或饥饿，或有余或缺乏，任何事情，任何景况，我都得了秘诀。
PHIL|4|13|我靠着那加给我力量的，凡事都能做。
PHIL|4|14|然而，你们能和我分担忧患是一件好事。
PHIL|4|15|腓立比 人哪，你们也知道我开始传福音、离开 马其顿 的时候，在收支的事上，除了你们以外，并没有别的教会和我分担。
PHIL|4|16|就是我在 帖撒罗尼迦 ，你们也一再差人来供给我的需用。
PHIL|4|17|我并不求什么馈赠，只求你们的果子不断增多，归在你们的账上。
PHIL|4|18|但我已经如数收到，并且有余；我已经充足，因我从 以巴弗提 受了你们的馈赠，当作极美的香气，为上帝所接纳、所喜悦的祭物。
PHIL|4|19|我的上帝必照他荣耀的丰富，在基督耶稣里，使你们一切所需用的都充足。
PHIL|4|20|愿荣耀归给我们的父上帝，直到永永远远。阿们！
PHIL|4|21|请问候在基督耶稣里的各位圣徒。跟我一起的众弟兄都问候你们。
PHIL|4|22|众圣徒都问候你们，特别在凯撒家里的人问候你们。
PHIL|4|23|愿主耶稣基督的恩与你们的灵同在！
COL|1|1|奉上帝旨意，作基督耶稣使徒的 保罗 ，和我们的弟兄 提摩太 ，
COL|1|2|写信给 歌罗西 的圣徒，在基督里忠心的弟兄。愿恩惠、平安 从我们的父上帝归给你们！
COL|1|3|我们为你们祷告的时候，常常感谢我们主耶稣基督的父上帝 ，
COL|1|4|因为听见你们对基督耶稣的信心，并对众圣徒有的爱心。
COL|1|5|这都是因着那给你们存在天上的盼望，它就是你们从前所听见真理的道，就是福音；
COL|1|6|这福音传到你们那里，也传到普天下，并且继续增长，不断结果，正如自从你们听见福音，真正知道上帝恩惠的日子起，在你们中间也是这样。
COL|1|7|这福音是你们从我们所亲爱、一同作仆人的 以巴弗 学到的。他为我们 作了基督的忠心仆役，
COL|1|8|也把圣灵赐给你们的爱告诉我们。
COL|1|9|因此，我们自从听见的日子就不住地为你们祷告和祈求，愿你们满有一切属灵的智慧和悟性，真正知道上帝的旨意，
COL|1|10|好使你们行事为人对得起主，凡事蒙他喜悦，在一切善事上结果子，对上帝的认识更有长进。
COL|1|11|愿你们从他荣耀的权能中，得以在一切事上力上加力，好使你们凡事欢欢喜喜地忍耐宽容，
COL|1|12|又感谢父，使你们配与众圣徒在光明中分享基业。
COL|1|13|他救了我们脱离黑暗的权势，迁移到他爱子的国度里。
COL|1|14|藉着他的爱子，我们得蒙救赎，罪得赦免。
COL|1|15|爱子是那看不见的上帝之像， 是首生的 ，在一切被造的以先。
COL|1|16|因为万有都是在他里面 造的， 无论是天上的、地上的， 能看见的、不能看见的， 或是有权位的、统治的， 或是执政的、掌权的， 一概都是藉着他为着他造的。
COL|1|17|他在万有之先； 万有也靠他而存在。
COL|1|18|他是身体（教会）的头； 他是元始， 是从死人中复活的首生者， 好让他在万有中居首位。
COL|1|19|因为上帝喜欢使一切的丰盛在他里面居住，
COL|1|20|藉着他 ，上帝使万有与自己和好， 无论是地上的、天上的， 都藉着他在十字架上所流的血促成了和平。
COL|1|21|从前你们与上帝隔绝，心思上与他为敌，行为邪恶；
COL|1|22|但如今，他藉着他儿子肉身的死，已经使你们与他自己和好了 ，把你们献在他的面前，成为圣洁，没有瑕疵，无可指责。
COL|1|23|只要你们持守信仰，根基稳固，坚定不移，不致动摇，离开了你们从前所听见的福音的盼望；这福音也是传给天下一切被造之物的，我— 保罗 作了这福音的仆役。
COL|1|24|现在我为你们受苦，倒很快乐；并且为基督的身体，就是为教会，我要在自己的肉身上补满基督未尽的苦难。
COL|1|25|我照上帝为你们所赐我的职分作了教会的仆役，要把上帝的道传得完满；
COL|1|26|这道就是历世历代所隐藏的奥秘，但如今向他的圣徒显明了。
COL|1|27|上帝要让他们知道，这奥秘在外邦人中有何等丰盛的荣耀；就是基督在你们心里 成了得荣耀的盼望。
COL|1|28|我们传扬他，是用诸般的智慧，劝戒各人，教导各人，要把各人在基督里完完全全地献上 。
COL|1|29|我也为此劳苦，照着他在我里面运用的大能尽心竭力。
COL|2|1|我要你们知道，我为你们和 老底嘉 人，和所有没有与我见过面的人，是何等地勤奋；
COL|2|2|为要使他们的心得安慰，因爱心互相联络，以致有从确实了解所产生的丰盛，好深知上帝的奥秘，就是基督；
COL|2|3|在他里面蕴藏着一切智慧和知识。
COL|2|4|我说这话，免得有人用花言巧语迷惑你们。
COL|2|5|虽然我身体不在你们那里，心却与你们同在，很高兴见你们循规蹈矩，对基督的信心也坚固。
COL|2|6|既然你们接受了主基督耶稣，就要靠着他而生活，
COL|2|7|照着你们所领受的教导，在他里面生根建造，信心坚固，充满着感谢的心。
COL|2|8|你们要谨慎，免得有人用他的哲学和虚空的废话，不照着基督，而是照人间的传统和世上粗浅的学说 ，把你们掳去。
COL|2|9|因为上帝本性一切的丰盛都有形有体地居住在基督里面；
COL|2|10|你们在他里面也已经成为丰盛。他是所有执政掌权者的元首。
COL|2|11|你们也在他里面受了不是人手所行的割礼，而是使你们脱去肉体情欲的基督的割礼。
COL|2|12|你们既受洗与他一同埋葬，也就在此礼上，因信那使他从死人中复活的上帝的作为跟他一同复活。
COL|2|13|你们从前在过犯和未受割礼的肉体中死了，上帝却赦免了你们一切的过犯，使你们与基督一同活过来，
COL|2|14|涂去了在律例上所写、敌对我们、束缚我们的字据，把它撤去，钉在十字架上。
COL|2|15|基督既将一切执政者、掌权者的权势解除了，就在凯旋的行列中，将他们公开示众，仗着十字架夸胜。
COL|2|16|所以，不要让任何人在饮食上，或节期、初一、安息日等事上评断你们。
COL|2|17|这些原是未来的事的影子，真体却是属基督的。
COL|2|18|不要让人藉着故作谦虚和敬拜天使夺去你们的奖赏。这等人拘泥在所见过的幻象 ，随着自己的欲望无故地自高自大，
COL|2|19|不紧随元首；其实，由于他全身藉着关节筋络才得到滋养，互相联络，靠上帝所赐的成长而成长。
COL|2|20|既然你们与基督同死而脱离了世上粗淺的学说，为什么仍像生活在世俗中一样，去服从那“不可拿、不可尝、不可摸”等类的规条呢？
COL|2|21|
COL|2|22|这些都是根据人的命令和教导，论到这一切都是一经使用就都败坏了。
COL|2|23|这些规条使人徒有智慧之名，用私意崇拜，自表谦卑，苦待己身，其实在克制肉体的情欲上毫无功效。
COL|3|1|所以，既然你们已经与基督一同复活，就当求上面的事；那里有基督，坐在上帝的右边。
COL|3|2|你们要思考上面的事，不要思考地上的事。
COL|3|3|因为你们已经死了，你们的生命与基督一同藏在上帝里面。
COL|3|4|基督是你们的生命，他显现的时候，你们也要与他一同在荣耀里显现。
COL|3|5|所以，要治死你们在地上的肢体；就如淫乱、污秽、邪情、恶欲和贪婪—贪婪就是拜偶像。
COL|3|6|因这些事，上帝的愤怒必临到那些悖逆的人 。
COL|3|7|当你们在这些事中活着的时候，你们的行为也曾是这样的。
COL|3|8|但现在你们要弃绝这一切的事，就是恼恨、愤怒、恶毒、毁谤和口中污秽的言语。
COL|3|9|不要彼此说谎，因为你们已经脱去旧人和旧人的行为，
COL|3|10|穿上了新人，这新人照着造他的主的形像在知识上不断地更新。
COL|3|11|在这事上并不分 希腊 人和 犹太 人，受割礼的和未受割礼的，未开化的人、 西古提 人、为奴的、自主的；惟独基督是一切，又在一切之内。
COL|3|12|所以，你们既是上帝的选民，圣洁、蒙爱的人，要穿上怜悯、恩慈、谦虚、温柔和忍耐。
COL|3|13|倘若这人与那人有嫌隙，总要彼此容忍，彼此饶恕；主 怎样饶恕了你们，你们也要怎样饶恕人。
COL|3|14|除此以外，还要穿上爱心，因为爱是贯通全德的。
COL|3|15|你们要让基督所赐的和平在你们心里作主，也为此蒙召，归为一体。你们还要存感谢的心。
COL|3|16|当用各样的智慧，把基督的道丰丰富富的存在心里，用诗篇、赞美诗、灵歌，彼此教导，互相劝戒，以感恩的心歌颂上帝。
COL|3|17|你们无论做什么，或说话或行事，都要奉主耶稣的名，藉着他感谢父上帝。
COL|3|18|你们作妻子的，要顺服自己的丈夫，这在主里面是合宜的。
COL|3|19|你们作丈夫的，要爱你们的妻子，不可虐待她们。
COL|3|20|你们作儿女的，要凡事听从父母，因为这是主所喜悦的。
COL|3|21|你们作父亲的，不要惹儿女生气，恐怕他们会灰心。
COL|3|22|你们作仆人的，要凡事听从你们肉身的主人，不要只在眼前服事，像是讨人喜欢的，总要心存诚实，因为你们敬畏主。
COL|3|23|你们无论做什么，都要从心里做，像是为主做的，不是为人做的；
COL|3|24|因为你们知道，从主那里必得着基业作为赏赐。你们要服侍的是主基督。
COL|3|25|行不义的人必受不义的报应；主并不偏待人。
COL|4|1|你们作主人的，待仆人要公正，因为知道，你们也有一位主在天上。
COL|4|2|你们要恒切祷告，在祷告中警醒感恩。
COL|4|3|同时，也要为我们祷告，求上帝给我们开传道的门，能宣讲基督的奥秘，
COL|4|4|使我能按着所该说的话将这奥秘显明出来，我为此而被捆锁。
COL|4|5|你们要把握时机，用智慧与外人来往。
COL|4|6|你们的言谈要时常带着温和，好像用盐调味，让你们知道该怎样应对每一个人。
COL|4|7|推基古 是我亲爱的弟兄，忠心的仆役，和我一同作主的仆人；他要把我一切的事都告诉你们。
COL|4|8|我特意打发他到你们那里去，好让你们知道我们的情况，又让他安慰你们的心。
COL|4|9|我又打发一位亲爱忠心的弟兄 阿尼西谋 同去；他也是你们那里的人。他们会把这里一切的事都告诉你们。
COL|4|10|与我一同坐牢的 亚里达古 问候你们。 巴拿巴 的表弟 马可 也问候你们。关于他，你们已经得到指示；他若到你们那里，你们要接待他。
COL|4|11|称为 犹士都 的 耶数 也问候你们。奉割礼的人中，只有这三个人是为上帝的国与我作同工的，也是使我心里得安慰的。
COL|4|12|有一位你们那里的人，作基督耶稣 仆人的 以巴弗 问候你们。他祷告的时候常为你们竭力祈求，愿你们能站稳而成熟，充分确信上帝一切的旨意。
COL|4|13|他为你们、 老底嘉 和 希拉坡里 的弟兄多多劳苦，这是我可以为他作见证的。
COL|4|14|亲爱的医生 路加 和 底马 问候你们。
COL|4|15|请问候 老底嘉 的弟兄以及 宁法 ，和她家里 的教会。
COL|4|16|你们宣读了这书信，也要交给 老底嘉 的教会宣读；你们也要宣读从 老底嘉 转来的书信。
COL|4|17|你们要对 亚基布 说：“务要完成你从主所领受的职分。”
COL|4|18|我— 保罗 亲笔问候你们。要记念我在捆锁中。愿恩惠与你们同在！
1THESS|1|1|保罗 、 西拉 、 提摩太 写信给 帖撒罗尼迦 在父上帝和主耶稣基督里的教会。愿恩惠、平安 归给你们！
1THESS|1|2|我们为你们众人常常感谢上帝，祷告的时候提到你们，
1THESS|1|3|在我们的父上帝面前，不住地记念你们因信心所做的工作，因爱心所受的劳苦，因盼望我们主耶稣基督所存的坚忍。
1THESS|1|4|上帝所爱的弟兄啊，我知道你们是蒙拣选的；
1THESS|1|5|因为我们的福音传到你们那里，不仅在言语，也在能力，也在圣灵和充足的确信。你们知道，我们在你们那里，为你们的缘故是怎样为人。
1THESS|1|6|你们成为效法我们，更效法主的人，因圣灵所激发的喜乐，在大患难中领受了真道，
1THESS|1|7|从此你们作了 马其顿 和 亚该亚 所有信主的人的榜样。
1THESS|1|8|因为主的道已经从你们那里传播出去，你们向上帝的信心不只在 马其顿 和 亚该亚 ，就是在各处也都传开了，所以不用我们说什么话。
1THESS|1|9|因为他们自己已经传讲我们是怎样进到你们那里，你们是怎样离弃偶像，归向上帝来服侍那又真又活的上帝，
1THESS|1|10|等候他儿子从天降临，就是上帝使他从死人中复活的那位救我们脱离将来愤怒的耶稣。
1THESS|2|1|弟兄们，你们自己知道我们来到你们那里并不是徒然的。
1THESS|2|2|我们从前在 腓立比 蒙难受辱，这是你们知道的，可是我们还是靠着上帝给我们的勇气，在强烈反对中把上帝的福音传给你们。
1THESS|2|3|我们的劝勉不是出于错误，也不是出于污秽，也不是用诡诈。
1THESS|2|4|但上帝既然认定我们经得起考验，把福音托付我们，我们就照着传讲，不是要讨人喜欢，而是要讨那考验我们的心的上帝喜欢。
1THESS|2|5|因为我们从来没有用过谄媚的话，这是你们知道的，也没有藏着贪心，这是上帝可以作证的。
1THESS|2|6|我们作为基督的使徒，虽然可以受人尊重，却没有向你们或向别人求荣耀，反而在你们当中心存温柔，如同母亲哺乳自己的孩子。
1THESS|2|7|
1THESS|2|8|既然我们这样爱你们，不但乐意将上帝的福音给你们，连自己的性命也乐意给你们，因为你们是我们所疼爱的。
1THESS|2|9|弟兄们，你们记念我们的辛苦劳碌，昼夜做工，传上帝的福音给你们，免得你们任何人受累。
1THESS|2|10|我们对你们信主的人是何等圣洁、正直、无可指责，这有你们作证，也有上帝作证。
1THESS|2|11|正如你们知道，我们待你们好像父亲待自己的儿女一样。
1THESS|2|12|我们劝勉你们，安慰你们，嘱咐你们，使你们行事对得起那召你们进他自己的国、得他荣耀的上帝。
1THESS|2|13|为此，我们也不断地感谢上帝，因为你们听见我们所传上帝的道的时候，你们领受了，不以为这是人的道，而以为这确实是上帝的道，而且在你们信主的人当中运行着。
1THESS|2|14|弟兄们，你们与 犹太 地区上帝的各教会，就是在基督耶稣里的各教会，有同样的遭遇，因为你们也受了同胞的迫害，像他们受了 犹太 人的迫害一样。
1THESS|2|15|这些 犹太 人不但杀了主耶稣和先知们，又把我们赶出去。他们令上帝不悦，且与众人为敌，
1THESS|2|16|阻挠我们传道给外邦人，使他们得救，以致常常恶贯满盈，但上帝的愤怒终于临到他们身上。
1THESS|2|17|弟兄们，我们被迫暂时与你们分离，身体离开，心却没有；我们极力想法子，渴望见你们的面。
1THESS|2|18|所以我们很想到你们那里去。我－ 保罗 有一两次要去，只是撒但阻挡了我们。
1THESS|2|19|当我们的主耶稣再来，我们站在他面前的时候，我们的盼望、喜乐和所夸的冠冕是什么呢？不正是你们吗？
1THESS|2|20|你们就是我们的荣耀和喜乐！
1THESS|3|1|既然我们不能再忍，就决定独自留在 雅典 ，
1THESS|3|2|于是差派我们在基督福音上作上帝同工的弟兄 提摩太 前去，在你们所信的道上坚固你们，劝勉你们，
1THESS|3|3|免得有人被这些患难动摇。因为你们自己知道，我们受患难原是命定的。
1THESS|3|4|我们在你们那里的时候，曾预先告诉你们，我们必受患难；你们知道，这果然发生了。
1THESS|3|5|为此，既然我不能再忍，就差派人去，要知道你们的信心如何，恐怕那诱惑人的果真诱惑了你们，以致我们的劳苦归于徒然。
1THESS|3|6|但是， 提摩太 刚从你们那里回来，将你们信心和爱心的好消息报给我们，又说你们常常记念我们，切切想见我们，如同我们想见你们一样。
1THESS|3|7|所以，弟兄们，我们在一切困苦患难中，因着你们的信心得到鼓励。
1THESS|3|8|如今你们若靠主站立得稳，我们就得生了。
1THESS|3|9|我们在上帝面前，因着你们满有喜乐。为这一切喜乐，我们能用怎样的感谢为你们报答上帝呢？
1THESS|3|10|我们昼夜切切祈求要见你们的面，来补足你们信心的不足。
1THESS|3|11|愿我们的父上帝自己和我们的主耶稣，为我们开路到你们那里去。
1THESS|3|12|又愿主使你们彼此相爱的心，和爱众人的心，都能增长，充足，如同我们爱你们一样，
1THESS|3|13|好坚固你们的心，使你们在我们的主耶稣同他众圣徒来临的时候，在我们父上帝面前，成为圣洁，无可指责。阿们！
1THESS|4|1|末了，弟兄们，我们靠着主耶稣求你们，劝你们，既然你们领受了我们的教导，知道该怎样行事为人，讨上帝的喜悦，其实你们也正这样行，我劝你们要更加努力。
1THESS|4|2|你们原知道，我们凭主耶稣传给你们什么命令。
1THESS|4|3|上帝的旨意就是要你们成为圣洁，远避淫行；
1THESS|4|4|要你们各人知道怎样用圣洁、尊贵控制自己的身体 ，
1THESS|4|5|不放纵私欲的邪情，像不认识上帝的外邦人。
1THESS|4|6|不准有人在这事上越轨，占他弟兄的便宜；因为这一类的事，主必报应，正如我预先对你们说过，又切切警告过你们的。
1THESS|4|7|上帝召我们本不是要我们沾染污秽，而是要我们圣洁。
1THESS|4|8|所以，那弃绝这教导的不是弃绝人，而是弃绝那把自己的圣灵赐给你们的上帝。
1THESS|4|9|有关弟兄间的手足之情，不用人写信给你们，因为你们自己蒙了上帝的教导要彼此相爱。
1THESS|4|10|你们向全 马其顿 的众弟兄固然是这样行，但我劝弟兄们要更加努力。
1THESS|4|11|要立志过安静的生活，管自己的事，亲手 做工，正如我们从前吩咐你们的，
1THESS|4|12|好使你们的行为能得外人的尊敬，同时也不依赖任何人。
1THESS|4|13|弟兄们，至于已睡了的人，我们不愿意你们不知道，恐怕你们忧伤，像那些没有指望的人一样。
1THESS|4|14|既然我们信耶稣死了，复活了，那些已经在耶稣里睡了的人，上帝也必将他们与耶稣一同带来。
1THESS|4|15|我们照主的话告诉你们一件事：我们这活着还存留到主来临的人，绝不会在那已经睡了的人之先。
1THESS|4|16|因为，召集令一发，天使长的呼声一叫，上帝的号角一吹，主必亲自从天降临；那在基督里死了的人必先复活，
1THESS|4|17|然后我们这些活着还存留的人必和他们一同被提到云里，在空中与主相会。这样，我们就要和主永远同在。
1THESS|4|18|所以，你们当用这些话彼此劝勉。
1THESS|5|1|弟兄们，关于那时候和日期，不用人写信给你们，
1THESS|5|2|因为你们自己明明知道，主的日子来到会像贼在夜间突然来到一样。
1THESS|5|3|人正说平安稳定的时候，灾祸忽然临到他们，如同阵痛临到怀胎的妇人一样，他们绝逃脱不了。
1THESS|5|4|弟兄们，你们并不在黑暗里，那日子不会像贼一样临到你们。
1THESS|5|5|你们都是光明之子，都是白昼之子；我们不属黑夜，也不属幽暗。
1THESS|5|6|所以，我们不要沉睡，像别人一样，总要警醒谨慎。
1THESS|5|7|因为睡了的人是在夜间睡，醉了的人是在夜间醉。
1THESS|5|8|但既然我们属于白昼，就应当谨慎，把信和爱当作护心镜遮胸，把得救的盼望当作头盔戴上。
1THESS|5|9|因为上帝不是预定我们受惩罚，而是预定我们藉着我们的主耶稣基督得救。
1THESS|5|10|他替我们死，让我们无论醒着、睡着，都与他同活。
1THESS|5|11|所以，你们该彼此劝勉，互相造就，正如你们素常做的。
1THESS|5|12|弟兄们，我们劝你们要敬重那些在你们中间劳苦的，就是在主里面督导你们、劝戒你们的人。
1THESS|5|13|又因他们所做的工作，要以爱心格外尊重他们。你们也要彼此和睦。
1THESS|5|14|弟兄们，我们劝你们，要警戒不守规矩的人，勉励灰心的人，扶助软弱的人，对众人要有耐心。
1THESS|5|15|你们要谨慎，无论是谁都不要以恶报恶，彼此间和对众人都要追求做好事。
1THESS|5|16|要常常喜乐，
1THESS|5|17|不住地祷告，
1THESS|5|18|凡事谢恩，因为这是上帝在基督耶稣里向你们所定的旨意。
1THESS|5|19|不要熄灭圣灵；
1THESS|5|20|不要藐视先知的讲论。
1THESS|5|21|但凡事要察验：美善的事要持守，
1THESS|5|22|各样恶事要禁戒。
1THESS|5|23|愿赐平安 的上帝亲自使你们完全成圣！愿你们的灵、魂、体得蒙保守，在我们的主耶稣基督来临的时候，完全无可指责。
1THESS|5|24|那召你们的本是信实的，他必成就这事。
1THESS|5|25|弟兄们，请也为 我们祷告。
1THESS|5|26|用圣洁的吻向众弟兄问安。
1THESS|5|27|我指着主嘱咐你们，要把这信宣读给众弟兄听。
1THESS|5|28|愿我们的主耶稣基督的恩惠与你们同在！
2THESS|1|1|保罗 、 西拉 和 提摩太 写信给 帖撒罗尼迦 、在我们的父上帝与主耶稣基督里的教会。
2THESS|1|2|愿恩惠、平安 从我们的 父上帝和主耶稣基督归给你们！
2THESS|1|3|弟兄们，我们该常常为你们感谢上帝，这本是合宜的；因为你们的信心格外增长，你们众人彼此相爱的心也都增加。
2THESS|1|4|所以，我们在上帝的各教会里为你们夸耀，因为你们在所受的一切压迫患难中仍牢守着耐心和信心。
2THESS|1|5|这正是上帝公义判断的明证，使你们配得上他的国，你们就是为这国受苦。
2THESS|1|6|既然上帝是公义的，他必以患难报复那加患难给你们的人，
2THESS|1|7|也必使你们这受患难的人与我们同得平安。那时，主耶稣同他有权能的天使从天上在火焰中显现，要报应那些不认识上帝和不听从我们的主耶稣福音的人。
2THESS|1|8|
2THESS|1|9|他们要受惩罚，永远沉沦，与主的面和他权能的荣光隔绝。
2THESS|1|10|这正是主再来，要在他圣徒的身上得荣耀，就是要使一切信的人感到惊讶的那日子，因为你们信了我们对你们作的见证。
2THESS|1|11|为此，我们常为你们祷告，愿我们的上帝看你们与他的呼召相配，又用大能成就你们一切良善的美意和因信心所做的工作，
2THESS|1|12|使我们主耶稣的名，照着我们的上帝和主耶稣基督的恩，在你们身上得荣耀，你们也在他身上得荣耀。
2THESS|2|1|弟兄们，关于我们主耶稣基督的来临和我们到他那里聚集，我劝你们：
2THESS|2|2|无论藉着灵，藉着言语，藉着冒我的名写的书信，说主的日子已经到了，不要轻易动心，也不要惊慌。
2THESS|2|3|不要让任何人用什么法子欺骗你们，因为那日子以前必有叛教的事，并有那不法的人，那沉沦之子出现。
2THESS|2|4|那抵挡者高抬自己超过一切称为神明的，和一切受人敬拜的，甚至坐在上帝的殿里，自称为上帝。
2THESS|2|5|我还在你们那里的时候曾把这些事告诉你们，你们不记得吗？
2THESS|2|6|现在你们也知道那拦阻他的是什么，为要使他到了时机才出现。
2THESS|2|7|因为那不法的隐秘已经运作，只是现在有一个阻挡的，要等到那阻挡的被除去才会发作，
2THESS|2|8|那时这不法的人必出现，主耶稣 要用口中的气灭绝他，以自己来临的光辉摧毁他。
2THESS|2|9|这不法的人来，是靠撒但的运作，行各样的异能、神迹和一切虚假的奇事，
2THESS|2|10|并且在那沉沦的人身上行各样不义的诡诈，因为他们不领受爱真理的心，好让他们得救。
2THESS|2|11|故此，上帝就给他们一个引发错误的心，叫他们信从虚谎，
2THESS|2|12|使一切不信真理、倒喜爱不义的人都被定罪。
2THESS|2|13|主所爱的弟兄们哪，我们本该常为你们感谢上帝，因为他拣选你们为初熟的果子 ，使你们因信真道，又蒙圣灵感化成圣，得到拯救。
2THESS|2|14|为此，上帝藉着我们所传的福音呼召你们，好得着我们主耶稣基督的荣光。
2THESS|2|15|所以，弟兄们，你们要站立得稳，凡所领受的教导，无论是我们口传的，是信上写的，都要坚守。
2THESS|2|16|愿我们主耶稣基督自己，和那爱我们、开恩将永远的安慰及美好的盼望赐给我们的父上帝，
2THESS|2|17|安慰你们的心，并且在一切善行善言上坚固你们！
2THESS|3|1|末了，弟兄们，请你们为我们祷告，好让主的道快快传开，得着荣耀，正如在你们中间一样，
2THESS|3|2|也让我们能脱离无理和邪恶人的手，因为不是人人都有信仰。
2THESS|3|3|但主是信实的，他要坚固你们，保护你们脱离那邪恶者。
2THESS|3|4|我们靠主对你们有信心，你们现在遵行，以后也必遵行我们所吩咐的。
2THESS|3|5|愿主引导你们的心去爱上帝，并学基督的忍耐！
2THESS|3|6|弟兄们，我们奉主耶稣基督的名吩咐你们，凡有弟兄懒散，不遵守我们所传授的教导，要远离他。
2THESS|3|7|你们自己知道该怎样效法我们。因为我们在你们当中从未懒散过，
2THESS|3|8|也从未白吃人的饭，倒是辛苦劳碌，昼夜做工，免得使你们中间有人受累。
2THESS|3|9|这并不是因我们没有权柄，而是要给你们作榜样，好让你们效法我们。
2THESS|3|10|我们在你们那里的时候曾吩咐你们，说若有人不肯做工，就不可吃饭。
2THESS|3|11|因为我们听说，在你们中间有人懒散，什么工都不做，反倒专管闲事。
2THESS|3|12|我们靠主耶稣基督吩咐并劝戒这样的人，要安分做工，自食其力。
2THESS|3|13|弟兄们，你们行善不可丧志。
2THESS|3|14|若有人不听从我们这信上的话，要把他记下，不和他交往，使他自觉羞愧；
2THESS|3|15|但不要把他当仇人，要劝他如劝弟兄。
2THESS|3|16|愿赐平安 的主随时随事亲自赐给你们平安！愿主与你们众人同在！
2THESS|3|17|我— 保罗 亲笔向你们问安。凡我的信都以此为记，我的笔迹就是这样。
2THESS|3|18|愿我们主耶稣基督的恩惠与你们众人同在！
1TIM|1|1|奉我们的救主上帝，和我们的盼望基督耶稣的命令，作基督耶稣使徒的 保罗 ，
1TIM|1|2|写信给那因信主作我真儿子的 提摩太 。愿恩惠、怜悯、平安 从父上帝和我们主基督耶稣归给你！
1TIM|1|3|我往 马其顿 去的时候，曾劝你留在 以弗所 ，好嘱咐某些人不可传别的教义，
1TIM|1|4|也不要听从无稽的传说和冗长的家谱；这样的事只会引起争论，无助于上帝的计划，这计划是凭着信才能了解的。
1TIM|1|5|但命令的目的就是爱；这爱是出于清洁的心、无愧的良心和无伪的信心。
1TIM|1|6|有人偏离了这些而转向空谈，
1TIM|1|7|想要作律法教师，却不明白自己所讲的是什么，也不知道所主张的是什么。
1TIM|1|8|我们知道，只要人善用律法，律法是好的；
1TIM|1|9|因为知道律法不是为义人订立的，而是为不法和叛逆的，不虔诚和犯罪的，不圣洁和恋世俗的，弑父母和杀人的，
1TIM|1|10|犯淫乱和亲男色的，拐卖人口和说谎话的，并起假誓的，或是为任何违背健全教义的事订立的。
1TIM|1|11|这是按照可称颂、荣耀之上帝交托我的福音说的。
1TIM|1|12|我感谢那赐给我力量的我们的主基督耶稣，因为他认为我可信任，派我服事他。
1TIM|1|13|我从前是亵渎、迫害、侮慢上帝的人；然而我还蒙了怜悯，因为我是在不信、不明白的时候做的。
1TIM|1|14|而且我们的主的恩典格外丰盛，使我在基督耶稣里有信心和爱心。
1TIM|1|15|这话可信，值得完全接受：“基督耶稣到世上来是要拯救罪人”，而在罪人中我是个罪魁。
1TIM|1|16|然而，我蒙了怜悯，好让基督耶稣在我这罪魁身上显明他完全的忍耐，给后来信他得永生的人作榜样。
1TIM|1|17|愿尊贵、荣耀归给永世的君王，那不朽坏、看不见、独一的上帝，直到永永远远。阿们！
1TIM|1|18|我儿 提摩太 啊，我照从前指着你的预言把这命令交托你，使你能藉着这些预言打那美好的仗，
1TIM|1|19|常存信心和无愧的良心。有些人丢弃良心，在信仰上触了礁；
1TIM|1|20|其中有 许米乃 和 亚历山大 ，我已经把他们交给撒但，让他们学会不再亵渎。
1TIM|2|1|所以，我劝你，首先要为人人祈求、祷告、代求、感谢；
1TIM|2|2|为君王和一切在位的，也要如此，使我们能够敬虔端正地过平稳宁静的生活。
1TIM|2|3|这是好的，在我们的救主上帝面前可蒙悦纳。
1TIM|2|4|他愿意人人得救，并得以认识真理。
1TIM|2|5|因为只有一位上帝， 在上帝和人之间也只有一位中保， 是成为人的基督耶稣。
1TIM|2|6|他献上自己作人人的赎价； 在适当的时候这事已经证实了。
1TIM|2|7|我为此奉派作传道，作使徒，在信仰和真理上作外邦人的教师。我说的是真话，不是说谎。
1TIM|2|8|我希望男人举起圣洁的手随处祷告，不发怒，不争论。
1TIM|2|9|我也希望女人以端正、克制和合乎体统的服装打扮自己，不以编发、金饰、珍珠和名贵衣裳来打扮。
1TIM|2|10|要有善行，这才与自称为敬畏上帝的女人相称。
1TIM|2|11|女人要事事顺服地安静学习。
1TIM|2|12|我不许女人教导，也不许她管辖男人，只要安静。
1TIM|2|13|因为 亚当 先被造，然后才是 夏娃 ；
1TIM|2|14|亚当 并没有受骗，而是女人受骗，陷在过犯里。
1TIM|2|15|然而，女人若持守信心、爱心，又圣洁克制，就必藉着生产而得救。
1TIM|3|1|“若有人想望监督的职分，他是在羡慕一件好事”，这话是可信的。
1TIM|3|2|监督必须无可指责，只作一个妇人的丈夫，有节制、克己、端正，乐意接待外人，善于教导，
1TIM|3|3|不酗酒，不打人；要温和，不好斗，不贪财。
1TIM|3|4|要好好管理自己的家，使儿女顺服，凡事庄重。
1TIM|3|5|人若不知道管理自己的家，怎能照管上帝的教会呢？
1TIM|3|6|刚信主的，不可作监督，恐怕他自高自大，落在魔鬼所受的惩罚里。
1TIM|3|7|监督也必须在教外有好名声，免得被人毁谤，落在魔鬼的罗网里。
1TIM|3|8|同样，执事也必须庄重，不一口两舌，不好酒，不贪不义之财；
1TIM|3|9|要存清白的良心固守信仰的奥秘。
1TIM|3|10|这些人也要先受考验，若没有可责之处，才让他们作执事。
1TIM|3|11|同样，女执事 也必须庄重，不说闲话，有节制，凡事忠心。
1TIM|3|12|执事只作一个妇人的丈夫，要好好管儿女和自己的家。
1TIM|3|13|因为善于作执事的，为自己得到美好的地位，并且无惧地坚信在基督耶稣里的信仰。
1TIM|3|14|我希望尽快到你那里去，所以先把这些事写给你；
1TIM|3|15|倘若我延误了，你也可以知道在上帝的家中该怎样做。这家就是永生上帝的教会，真理的柱石和根基。
1TIM|3|16|敬虔的奥秘是公认为伟大的： 上帝在肉身显现， 被圣灵称义， 被天使看见， 被传于外邦， 被世人信服， 被接在荣耀里。
1TIM|4|1|圣灵明说，在末后的时期必有人离弃信仰，去听信那诱惑人的邪灵和鬼魔的教训。
1TIM|4|2|这是出于撒谎者的假冒；这些人的良心如同被热铁烙了一般。
1TIM|4|3|他们禁止嫁娶，又禁戒食物—就是上帝所造、让那信而明白真理的人存感谢的心领受的。
1TIM|4|4|上帝所造之物样样都是好的，若存感谢的心领受，没有一样是不可吃的，
1TIM|4|5|都因上帝的话和人的祈祷而成为圣洁了。
1TIM|4|6|你若把这些事提醒弟兄们，就是基督耶稣的好执事，在信仰的话语和你向来所服从的正确教义上得到了栽培。
1TIM|4|7|要弃绝那世俗的言语和老妇的无稽传说。要在敬虔上操练自己：
1TIM|4|8|因操练身体有些益处；但敬虔在各方面都有益，它有现今和未来的生命的应许。
1TIM|4|9|这话可信，值得完全接受。
1TIM|4|10|我们劳苦，努力 正是为此，因为我们的指望在乎永生的上帝。他是人人的救主，更是信徒的救主。
1TIM|4|11|你要嘱咐和教导这些事。
1TIM|4|12|不可叫人小看你年轻，总要在言语、行为、爱心、信心、清洁上，都作信徒的榜样。
1TIM|4|13|要以宣读圣经，劝勉，教导为念，直等到我来。
1TIM|4|14|不要忽略你所得的恩赐，就是从前藉着预言、在众长老按手的时候赐给你的。
1TIM|4|15|这些事你要殷勤去做，并要在这些事上专心，让众人看出你的长进来。
1TIM|4|16|要谨慎自己和自己的教导，要在这些事上恒心，因为这样做，既能救自己，又能救听你的人。
1TIM|5|1|不可严责老年人，要劝他如同父亲。要待年轻人如同弟兄，
1TIM|5|2|年老妇女如同母亲。要清清洁洁地待年轻妇女如同姊妹。
1TIM|5|3|要尊敬真正守寡的妇人。
1TIM|5|4|寡妇若有儿女，或有孙儿女，要让儿孙先在自己家中学习行孝，报答亲恩，因为这在上帝面前是可蒙悦纳的。
1TIM|5|5|独居无靠的真寡妇只仰赖上帝，昼夜不住地祈求祷告。
1TIM|5|6|但好宴乐的寡妇活着也算是死了。
1TIM|5|7|这些事，你要嘱咐她们，让她们无可指责。
1TIM|5|8|若有人不照顾亲属，尤其是自己家里的人，就是背弃信仰，还不如不信的人。
1TIM|5|9|寡妇登记，年龄必须在六十岁以上，只作一个丈夫的妻子，
1TIM|5|10|又有行善的名声，就如养育儿女，收留外人，洗圣徒的脚，救济遭难的人，竭力行各样善事。
1TIM|5|11|至于年轻的寡妇，你要拒绝登记，因为她们情欲冲动、背弃基督的时候，就想嫁人，
1TIM|5|12|她们因废弃了当初所许的愿而被定罪。
1TIM|5|13|同时，她们又学了懒惰，习惯于挨家闲逛；不但懒惰，而且说长道短，好管闲事，说些不该说的话。
1TIM|5|14|所以，我希望年轻的寡妇嫁人，生养儿女，治理家务，不让敌人有辱骂的把柄，
1TIM|5|15|因为已经有一些人转去随从撒但了。
1TIM|5|16|信主的妇女若有亲戚是寡妇，要救济她们，不可拖累教会，好使教会能救济真正无助的寡妇。
1TIM|5|17|善于督导教会的长老，尤其是勤劳讲道教导人的，应该得到加倍的敬奉。
1TIM|5|18|因为经上说：“牛在踹谷的时候，不可笼住它的嘴”；又说：“工人得工资是应当的。”
1TIM|5|19|有控告长老的案件，非有两三个证人就不要受理。
1TIM|5|20|继续犯罪的人，要在众人面前责备他，使其余的人也有所惧怕。
1TIM|5|21|我在上帝、基督耶稣和蒙拣选的天使面前嘱咐你要遵守这些话，不可存成见，做事也不可偏心。
1TIM|5|22|不可急于给人行按手礼；也不可在别人的罪上有份，要保守自己纯洁。
1TIM|5|23|为了你的胃，又常患病，不要只喝水，要稍微喝点酒。
1TIM|5|24|有些人的罪是明显的，已先受审判了；有些人的罪是随后跟着来。
1TIM|5|25|同样，善行也有明显的，就是那不明显的也不能隐藏。
1TIM|6|1|凡负轭作奴隶的，要认为自己的主人配受各样的尊敬，免得上帝的名和教导被人亵渎。
1TIM|6|2|奴隶若有信主的主人，不可因他是主内弟兄就轻看他们，更要越发服侍他们，因为得到服侍的益处的正是信徒，是蒙爱的人。 你要教导人和劝勉这些事。
1TIM|6|3|若有人传别的教义，不符合我们主耶稣基督纯正的话语与合乎敬虔的教导，
1TIM|6|4|他是自高自大，一无所知，专好争辩，擅于舌战，因而生出嫉妒、纷争、毁谤、恶意猜疑，
1TIM|6|5|和心术不正与丧失真理的人不停地争吵，以敬虔为得利的门路。
1TIM|6|6|其实，敬虔加上知足就是大利。
1TIM|6|7|因为我们没有带什么到世上来， 也不能带什么去；
1TIM|6|8|只要有衣有食， 我们就该知足。
1TIM|6|9|但那些想要发财的人就陷在诱惑、罗网和许多无知有害的欲望中，使人沉沦，以致败坏和灭亡。
1TIM|6|10|贪财是万恶之根。有人因贪恋钱财而背离信仰，用许多愁苦把自己刺透了。
1TIM|6|11|但你这属上帝的人哪，要逃避这些事；要追求公义、敬虔、信心、爱心、忍耐、温柔。
1TIM|6|12|你要为信仰打那美好的仗；要持定永生，你为此被召，也已经在许多见证人面前作了那美好的见证。
1TIM|6|13|我在那赐生命给万物的上帝面前，并在向 本丢．彼拉多 作过那美好见证的基督耶稣面前嘱咐你 ：
1TIM|6|14|要守这命令，毫不玷污，无可指责，直到我们的主耶稣基督显现。
1TIM|6|15|到了适当的时候都要显明出来： 他是那可称颂、独一的权能者， 万王之王， 万主之主，
1TIM|6|16|就是那独一不死、 住在人不能靠近的光里， 是人未曾看见，也是不能看见的。 愿尊贵和永远的权能都归给他。阿们！
1TIM|6|17|至于那些今世富足的人，你要嘱咐他们不要自高，也不要倚赖靠不住的钱财；要倚靠那厚赐万物给我们享受的上帝。
1TIM|6|18|又要嘱咐他们行善，在好事上富足，甘心施舍，乐意分享，
1TIM|6|19|为自己积存财富，而为将来打美好的根基，好使他们能把握那真正的生命。
1TIM|6|20|提摩太 啊，要持守所给你的托付。要躲避世俗的空谈和那假冒知识的矛盾言论。
1TIM|6|21|有人自称有这知识而偏离了信仰。 愿恩惠与你们同在！
2TIM|1|1|奉上帝旨意，按照基督耶稣里所应许的生命，作基督耶稣使徒的 保罗 ，
2TIM|1|2|写信给我亲爱的儿子 提摩太 。愿恩惠、怜悯、平安 从父上帝和我们的主基督耶稣归给你！
2TIM|1|3|我感谢上帝，就是我接续祖先用纯洁的良心所事奉的上帝，在祈祷中昼夜不停地想念你。
2TIM|1|4|我一想起你的眼泪，就急切想见你，好让我满心快乐。
2TIM|1|5|我记得你无伪的信心，这信心先存在你外祖母 罗以 和你母亲 友妮基 的心里，我深信也存在你的心里。
2TIM|1|6|为这缘故，我提醒你要把上帝藉着我按手所给你的恩赐再如火挑旺起来。
2TIM|1|7|因为上帝赐给我们的不是胆怯的心，而是刚强、仁爱、自制的心。
2TIM|1|8|所以，不要以给我们的主作见证为耻，也不要以我这为主被囚的为耻；总要靠着上帝的大能，与我为福音同受苦难。
2TIM|1|9|上帝救了我们， 以圣召召我们， 不是按我们的行为， 而是按他的旨意和恩典； 这恩典是万古之先 在基督耶稣里赐给我们的，
2TIM|1|10|但如今 藉着我们的救主基督耶稣的显现已经表明出来； 他把死废去， 藉着福音，将不朽的生命彰显出来。
2TIM|1|11|我为这福音奉派作传道，作使徒，作教师。
2TIM|1|12|为这缘故，我也受这些苦难。然而，我不以为耻，因为我知道我所信的是谁，也深信他能保全他所交托我的 ，直到那日。
2TIM|1|13|你从我听到那健全的言论，要用在基督耶稣里的信心和爱心常常守着，作为规范。
2TIM|1|14|你要靠着那住在我们里面的圣灵，牢牢守住所交托给你那美好的事。
2TIM|1|15|你知道，所有在 亚细亚 的人都离弃了我，其中有 腓吉路 和 黑摩其尼 。
2TIM|1|16|愿主怜悯 阿尼色弗 一家的人，因为他屡次令我欣慰。他不以我的铁链为耻，
2TIM|1|17|反而一到 罗马 就急切寻找我，并且找到了。
2TIM|1|18|愿主使他在那日能蒙主的怜悯。他在 以弗所 怎样多服事我，你是清楚知道的。
2TIM|2|1|我儿啊，你要在基督耶稣的恩典上刚强起来。
2TIM|2|2|你在许多见证人面前听见我所教导的，也要交托给那忠心而又能教导别人的人。
2TIM|2|3|你要和我同受苦难，作基督耶稣的精兵。
2TIM|2|4|凡当兵的，不让世务缠身，好使那招他当兵的人喜悦。
2TIM|2|5|运动员在比赛的时候，不按规则就不能得冠冕。
2TIM|2|6|勤劳的农夫理当先得粮食。
2TIM|2|7|我所说的话，你要考虑，因为主必在凡事上给你聪明。
2TIM|2|8|要记得耶稣基督，他是 大卫 的后裔，从死人中复活；这就是我所传的福音。
2TIM|2|9|我为这福音受苦难，甚至像犯人一样被捆绑，然而上帝的话没有被捆绑。
2TIM|2|10|所以，我为了选民事事忍耐，为使他们也能得到那在基督耶稣里的救恩和永远的荣耀。
2TIM|2|11|这话是可信的： 我们若与基督同死，也必与他同活；
2TIM|2|12|我们若忍耐到底，也必和他一同作王。 我们若不认他，他也必不认我们；
2TIM|2|13|我们纵然失信，他仍是可信的， 因为他不能否认自己。
2TIM|2|14|你要向众人提醒这些事，在上帝 面前嘱咐他们不可在言词上争辩；这是没有益处的，只能伤害听的人。
2TIM|2|15|你当竭力在上帝面前作一个经得起考验、无愧的工人，按着正意讲解真理的话。
2TIM|2|16|要远避世俗的空谈，因为这等空谈会使人进到更不敬虔的地步。
2TIM|2|17|他们的话如同毒疮越烂越大；其中有 许米乃 和 腓理徒 ，
2TIM|2|18|他们偏离了真理，说复活的事已过去，败坏了好些人的信心。
2TIM|2|19|然而，上帝坚固的根基屹立不移；上面有这印记说：“主认得他自己的人”，又说：“凡称呼主名的人总要离开不义。”
2TIM|2|20|大户人家不但有金器银器，也有木器瓦器；有作为贵重之用的，有作为卑贱之用的。
2TIM|2|21|人若自洁，脱离卑贱的事，必成为贵重的器皿，成为圣洁，合乎主用，预备行各样的善事。
2TIM|2|22|你要逃避年轻人的私欲，同那以纯洁的心求告主的人追求公义、信实、仁爱、和平。
2TIM|2|23|但要弃绝那愚拙无知的辩论，因为你知道这等事只会引起争辩。
2TIM|2|24|主的仆人不可争辩，只要温和待人，善于教导，恒心忍耐，
2TIM|2|25|用温柔劝导反对的人。也许上帝会给他们悔改的心能明白真理，
2TIM|2|26|让他们这些已被魔鬼掳去顺从他诡计的人能醒悟过来，脱离他的罗网。
2TIM|3|1|你该知道，末世必有艰难的日子来到。
2TIM|3|2|那时人会专爱自己，贪爱钱财，自夸，狂傲，毁谤，违背父母，忘恩负义，心不圣洁，
2TIM|3|3|没有亲情，抗拒和解，好说谗言，不能节制，性情凶暴，不爱良善，
2TIM|3|4|卖主卖友，任意妄为，自高自大，爱好宴乐，不爱上帝，
2TIM|3|5|有敬虔的外貌，却背弃了敬虔的实质，这等人你要避开。
2TIM|3|6|他们当中有人潜入别人家里，操纵无知的妇女；这些妇女被罪恶压制，被各样的私欲引诱，
2TIM|3|7|虽然常常学习，终久无法达到明白真理的地步。
2TIM|3|8|从前 雅尼 和 佯庇 怎样反对 摩西 ，这等人也怎样抵挡真理；他们的心地败坏，信仰经不起考验。
2TIM|3|9|然而，他们没有进步，因为他们的愚昧必在众人面前显露出来，像那两人一样。
2TIM|3|10|但你已经追随了我的教导、行为、志向、信心、宽容、爱心、忍耐，
2TIM|3|11|以及我在 安提阿 、 以哥念 、 路司得 所遭遇的迫害和苦难。我忍受了何等的迫害！但从这一切苦难中，主都把我救了出来。
2TIM|3|12|其实，凡立志在基督耶稣里敬虔度日的，也都将受迫害。
2TIM|3|13|只是作恶的和骗人的将变本加厉，迷惑人也被人迷惑。
2TIM|3|14|至于你，你要持守所学习的和所确信的，因为你知道是跟谁学的，
2TIM|3|15|并且知道你从小明白圣经，这圣经能使你因在基督耶稣里的信 有得救的智慧。
2TIM|3|16|圣经都是上帝所默示的 ，于教训、督责、使人归正、教导人学义都是有益的，
2TIM|3|17|叫属上帝的人得以完全，预备行各样的善事。
2TIM|4|1|我在上帝面前，并在将来审判活人死人的基督耶稣面前，凭着他的显现和他的国度郑重地劝戒你：
2TIM|4|2|务要传道；无论得时不得时总要专心，并以百般的忍耐和各样的教导责备人，警戒人，劝勉人。
2TIM|4|3|因为时候将到，那时人会厌烦健全的教导，耳朵发痒，就随心所欲地增添好些教师，
2TIM|4|4|并且掩耳不听真理，偏向无稽的传说。
2TIM|4|5|至于你，凡事要谨慎，忍受苦难，做传福音的工作，尽你的职分。
2TIM|4|6|至于我，我已经被浇献，离世的时候到了。
2TIM|4|7|那美好的仗我已经打过了，当跑的路我已经跑尽了，该信的道我已经守住了。
2TIM|4|8|从此以后，有公义的冠冕为我存留，就是按着公义审判的主到了那日要赐给我的；不但赐给我，也赐给凡爱慕他显现的人。
2TIM|4|9|你要赶紧到我这里来。
2TIM|4|10|因为 底马 贪爱现今的世界，已经离弃我，往 帖撒罗尼迦 去了； 革勒士 往 加拉太 去； 提多 往 挞马太 去；
2TIM|4|11|只有 路加 在我这里。你来的时候把 马可 带来，因为他在服事 上于我有益。
2TIM|4|12|我已经打发 推基古 往 以弗所 去。
2TIM|4|13|我在 特罗亚 留给 加布 的那件外衣，你来的时候要带来，那些书也带来，特别是那几卷羊皮的书。
2TIM|4|14|铜匠 亚历山大 多方害我；主必照他所行的报应他。
2TIM|4|15|你也要防备他，因为他极力抗拒我们的话。
2TIM|4|16|我初次上诉时，没有人前来帮助，竟都离弃了我，但愿这罪不归在他们身上。
2TIM|4|17|惟有主站在我身边，加给我力量，使我能把福音完整地传开，让所有的外邦人都听见；我也从狮子口里被救出来。
2TIM|4|18|主必救我脱离一切的凶恶，也必救我进他的天国。愿荣耀归给他，直到永永远远。阿们！
2TIM|4|19|请向 百基拉 、 亚居拉 和 阿尼色弗 一家的人问安。
2TIM|4|20|以拉都 在 哥林多 住下了。 特罗非摩 病了，我把他留在 米利都 。
2TIM|4|21|你要赶紧在冬天以前到我这里来。 友布罗 、 布田 、 利奴 、 革老底亚 和众弟兄都向你问安。
2TIM|4|22|愿主与你的灵同在！愿恩惠与你们同在！
TITUS|1|1|上帝的仆人、耶稣基督的使徒 保罗 ，为了使上帝的选民信从与认识合乎敬虔的真理—
TITUS|1|2|这真理是在盼望那无谎言的上帝在万古之先所应许的永生，
TITUS|1|3|到了适当的时机，藉着传扬福音，把他的道显明了；这传扬的责任是按着我们的救主上帝的命令交托给我的—
TITUS|1|4|我写信给在共同的信仰上作我真儿子的 提多 。愿恩惠、平安 从父上帝和我们的救主基督耶稣归给你！
TITUS|1|5|我从前把你留在 克里特 ，是要你将那没有办完的事都办妥，又照我所吩咐你的，在各城设立长老。
TITUS|1|6|若有无可指责的人，只作一个妇人的丈夫，儿女也是信主的，没有人告他们放荡，不受约束，就可以设立。
TITUS|1|7|监督既然是上帝的管家，必须无可指责、不自负、不暴躁、不酗酒、不好斗、不贪财；
TITUS|1|8|却要乐意接待外人、好善、克己、正直、圣洁、节制，
TITUS|1|9|坚守合乎教义的可靠之道，就能将健全的教导劝勉人，又能驳倒争辩的人。
TITUS|1|10|因为也有许多人不受约束，说空话欺哄人，尤其是那些奉割礼的人。
TITUS|1|11|这些人的口必须堵住，因为他们贪不义之财，将不该教导的事教导人，败坏人的全家。
TITUS|1|12|克里特 人中有一个本地的先知说：“ 克里特 人常说谎话，是恶兽，贪吃懒做。”
TITUS|1|13|这个见证是真的。为这缘故，你要严厉地责备他们，使他们在信仰上健全。
TITUS|1|14|不要听 犹太 人无稽的传说和背弃真理之人的命令。
TITUS|1|15|在洁净的人，凡物都洁净；在污秽不信的人，什么都不洁净，连心地和天良也都污秽了。
TITUS|1|16|他们宣称认识上帝，却在行为上否认他；他们是可憎恶的，是悖逆的，不配做任何好事。
TITUS|2|1|至于你，你所讲的总要合乎那健全的教导。
TITUS|2|2|劝老年人要有节制、端正、克己，在信心、爱心、耐心上都要健全。
TITUS|2|3|又要劝年长的妇女在操守上恭正，不说谗言，不作酒的奴隶，用善道教导人，
TITUS|2|4|好指教年轻的妇女爱丈夫，爱儿女，
TITUS|2|5|克己，贞洁，理家，善良，顺服自己的丈夫，免得上帝的道被毁谤。
TITUS|2|6|同样，要劝年轻人凡事克己。
TITUS|2|7|你要显出自己是好行为的榜样，在教导上要正直、庄重，
TITUS|2|8|言语健全，无可指责，使那反对的人，因说不出我们有什么不好而自觉羞愧。
TITUS|2|9|要劝仆人顺服自己的主人，凡事讨他的喜悦，不可顶撞他，
TITUS|2|10|不可私窃财物；要凡事显出完美的忠诚，好事事都能荣耀我们救主上帝的教导。
TITUS|2|11|因为，上帝救众人的恩典已经显明出来，
TITUS|2|12|训练我们除去不敬虔的心和世俗的情欲，在今世过克己、正直、敬虔的生活，
TITUS|2|13|等候福乐的盼望，并等候至大的上帝和我们的救主 耶稣基督的荣耀显现。
TITUS|2|14|他为我们的缘故舍己，为了要赎我们脱离一切罪恶，又洁净我们作他自己的子民，热心为善。
TITUS|2|15|这些事你要讲明，要充分运用你的职权劝勉人，责备人。不要让任何人轻看你。
TITUS|3|1|你要提醒众人，叫他们顺服执政的、掌权的，要服从，预备行各样善事。
TITUS|3|2|不要毁谤，不要争吵，要和气，对众人总要显出温柔。
TITUS|3|3|我们从前也是无知、悖逆、受迷惑，作各样私欲和宴乐的奴隶，在恶毒、嫉妒中度日，是可恨的，而且彼此相恨。
TITUS|3|4|但到了我们救主上帝的恩慈和慈爱显明的时候，
TITUS|3|5|他救了我们，并不是因我们自己所行的义，而是照他的怜悯，藉着重生的洗和圣灵的更新。
TITUS|3|6|圣灵就是上帝藉着我们的救主耶稣基督厚厚地浇灌在我们身上的，
TITUS|3|7|好让我们因他的恩得称为义，可以凭着永生的盼望成为后嗣 。
TITUS|3|8|这话是可信的。 我愿你坚持这些事，使那些已信上帝的人留心行善 。这都是美好且对人有益的。
TITUS|3|9|要远避愚拙的辩论、家谱、纷争和因律法而起的争辩，因为这都是虚妄无益的。
TITUS|3|10|分门结党的人，警戒过一两次后就要拒绝跟他来往；
TITUS|3|11|因为你知道这样的人已经背道，常常犯罪，自己定自己的罪了。
TITUS|3|12|我打发 亚提马 或 推基古 到你那里去的时候，你要赶紧往 尼哥坡里 来见我，因为我已经决定在那里过冬。
TITUS|3|13|你要赶紧给 西纳 律师和 亚波罗 送行，让他们没有缺乏。
TITUS|3|14|我们的人也该学习行善，帮助有迫切需要的人，这样才不会不结果子。
TITUS|3|15|跟我同在一起的人都向你问安。请代向在信仰上爱我们的人问安。愿恩惠与你们众人同在！
PHLM|1|1|为基督耶稣被囚的 保罗 ，同弟兄 提摩太 ，写信给我们所亲爱的同工 腓利门 、
PHLM|1|2|亚腓亚 姊妹，和我们的战友 亚基布 ，以及在你家里的教会。
PHLM|1|3|愿恩惠、平安 从我们的父上帝和主耶稣基督归给你们！
PHLM|1|4|我在祷告中记念你的时候，常为你感谢我的上帝，
PHLM|1|5|因听说你对众圣徒的爱心，和你对主耶稣的信心。
PHLM|1|6|愿你与人分享信心的时候，能产生功效，让人知道我们 所行的各样善事都是为基督做的。
PHLM|1|7|弟兄啊，由于你的爱心，我得到极大的快乐和安慰，因为众圣徒的心从你得到舒畅。
PHLM|1|8|虽然我靠着基督能放胆吩咐你做该做的事，
PHLM|1|9|可是像我这上了年纪的 保罗 ，现在又是为基督耶稣被囚的，宁可凭着爱心求你，
PHLM|1|10|就是为我在捆锁中所生的儿子 阿尼西谋 求你。
PHLM|1|11|从前他与你没有益处，但如今与你我都有益处。
PHLM|1|12|我现在打发他回到你那里去，他是我心肝。
PHLM|1|13|我本来有意将他留下，在我为福音所受的捆锁中替你伺候我。
PHLM|1|14|但不知道你的意见，我不愿意这样做，好使你的善行不是出于勉强，而是出于自愿。
PHLM|1|15|他暂时离开你，也许是要让你永远得着他，
PHLM|1|16|不再是奴隶，而是高过奴隶，是亲爱的弟兄；对我确实如此，何况对你呢！无论在肉身或在主里更是如此。
PHLM|1|17|所以，你若以我为同伴，就接纳他，如同接纳我一样。
PHLM|1|18|他若亏负你，或欠你什么，都算在我的账上吧，
PHLM|1|19|我必偿还。这是我— 保罗 亲笔写的。我并不用对你说，甚至你自己也亏欠我呢！
PHLM|1|20|弟兄啊，希望你使我在主里因你得益处，让我的心在基督里得到舒畅。
PHLM|1|21|我写信给你，深信你必顺服，知道你所要做的，必过于我所说的。
PHLM|1|22|此外，还请给我预备住处，因为我盼望藉着你们的祷告，必蒙恩回到你们那里去。
PHLM|1|23|为基督耶稣与我一同坐监的 以巴弗 问候你。
PHLM|1|24|我的同工 马可 、 亚里达古 、 底马 、 路加 也都问候你。
PHLM|1|25|愿 主耶稣基督的恩与你们的灵同在。
HEB|1|1|古时候，上帝藉着众先知多次多方向列祖说话，
HEB|1|2|末世，藉着他儿子向我们说话，又立他为承受万有的，也藉着他创造宇宙。
HEB|1|3|他是上帝荣耀的光辉，是上帝本体的真像，常用他大能的命令托住万有。他洗净了人的罪，就坐在高天至大者的右边。
HEB|1|4|他所承受的名比天使的名更尊贵，所以他远比天使崇高。
HEB|1|5|上帝曾对哪一个天使说过： “你是我的儿子； 我今日生了你”？ 又说过： “我要作他的父； 他要作我的子”呢？
HEB|1|6|再者，上帝引领他长子 进入世界的时候，说： “上帝的使者都要拜他。”
HEB|1|7|关于使者，他说： “上帝以风为使者， 以火焰为仆役。”
HEB|1|8|关于子，他却说： “上帝啊，你的宝座是永永远远的； 你国度的权杖是正直的权杖。
HEB|1|9|你喜爱公义，恨恶罪恶； 所以上帝，就是你的上帝，用喜乐油膏你， 胜过膏你的同伴。”
HEB|1|10|他又说： “主啊，你起初立了地的根基， 天也是你手所造的。
HEB|1|11|天地都会消灭，你却长存； 天地都会像衣服渐渐旧了；
HEB|1|12|你要将天地卷起来，像卷一件外衣， 天地像衣服都会改变。 你却永不改变； 你的年数没有穷尽。”
HEB|1|13|上帝曾对哪一个天使说： “你坐在我的右边， 等我使你的仇敌作你的脚凳”？
HEB|1|14|众天使不都是事奉的灵，奉差遣为那将要承受救恩的人服务的吗？
HEB|2|1|所以，我们必须越发注意所听见的道，免得我们随流失去。
HEB|2|2|既然那藉着天使所传的话是确定的，凡违背不听从的，都受了该受的报应；
HEB|2|3|我们若忽略这么大的救恩，怎能逃避呢？这拯救起先是主亲自讲的，后来是听见的人给我们证实了。
HEB|2|4|上帝又按自己的旨意，更用神迹奇事、百般的异能，和圣灵所给的恩赐，与他们一同作见证。
HEB|2|5|我们所说将来的世界，上帝没有交给天使管辖。
HEB|2|6|但有人在某处证明说： “人算什么，你竟顾念他； 世人算什么，你竟眷顾他。
HEB|2|7|你使他暂时比天使微小 ， 赐他荣耀尊贵为冠冕， 你派他管理你手所造的，
HEB|2|8|使万物都服在他的脚下。” 既然使万物都服他 ，就没有剩下一样不服他的了。只是如今我们还不见万物都服他；
HEB|2|9|惟独见那成为暂时比天使微小的耶稣，因为受了死的痛苦，得了尊贵荣耀为冠冕，好使他因着上帝的恩，为人人经历了死亡。
HEB|2|10|原来那为万物所属、为万物所本的，为要领许多儿子进入荣耀，使救他们的元帅因受苦难而得以完全，本是合宜的。
HEB|2|11|因那使人成圣的，和那些得以成圣的，都是出于一。为这缘故，他称他们为弟兄也不以为耻，
HEB|2|12|说： “我要将你的名传给我的弟兄， 在会众中我要颂扬你。”
HEB|2|13|他又说： “我要依赖他。” 他又说： “看哪！我与上帝所给我的儿女都在这里。”
HEB|2|14|既然儿女同有血肉之躯，他也照样亲自成了血肉之躯，为能藉着死败坏那掌管死权的，就是魔鬼，
HEB|2|15|并要释放那些一生因怕死而作奴隶的人。
HEB|2|16|诚然，他并没有帮助天使，而是帮助了 亚伯拉罕 的后裔。
HEB|2|17|所以，他凡事应当与他的弟兄相同，为要在上帝的事上成为慈悲忠信的大祭司，为百姓的罪献上赎罪祭。
HEB|2|18|既然他自己被试探而受苦，他能帮助被试探的人。
HEB|3|1|同蒙天召的圣洁弟兄啊，要思想我们所宣认为使者、为大祭司的耶稣；
HEB|3|2|他向指派他的尽忠，如同 摩西 向上帝的全 家尽忠一样。
HEB|3|3|他比 摩西 配得更多的荣耀，好像建造房屋的人比房屋更尊荣；
HEB|3|4|因为房屋都必有人建造，但建造万物的是上帝。
HEB|3|5|摩西 作为仆人，向上帝的全家尽忠，为将来要谈论的事作证；
HEB|3|6|但是基督作为儿子，治理上帝的家。我们若坚持因盼望而有的胆量和夸耀，我们就是他的家了。
HEB|3|7|所以，正如圣灵所说： “今日，你们若听他的话，
HEB|3|8|就不可硬着心，像在背叛之时， 就如在旷野受试探之日。
HEB|3|9|在那里，你们的祖宗试探我， 并且观看我的作为，
HEB|3|10|有四十年之久。 所以，我厌烦那世代， 说：他们的心常常迷糊， 竟不知道我的道路！
HEB|3|11|我在怒中起誓： 他们断不可进入我的安息！”
HEB|3|12|弟兄们，你们要谨慎，免得你们中间有人存着邪恶不信的心，离弃了永生的上帝。
HEB|3|13|总要趁着还有今日，天天彼此相劝，免得你们中间有人被罪迷惑，心肠刚硬了。
HEB|3|14|只要我们将起初确实的信心坚持到底，就在基督里有份了。
HEB|3|15|经上说： “今日，你们若听他的话， 就不可硬着心，像在背叛之时。”
HEB|3|16|听见他而又背叛他的是谁呢？岂不是跟着 摩西 从 埃及 出来的众人吗？
HEB|3|17|上帝向谁发怒四十年之久呢？岂不是那些犯罪而陈尸在旷野的人吗？
HEB|3|18|他向谁起誓，不容他们进入他的安息呢？岂不是向那些不信从的人吗？
HEB|3|19|这样看来，他们不能进入安息是因为不信的缘故了。
HEB|4|1|所以，既然进入他安息的应许依旧存在，我们就该存畏惧的心，免得我们 中间有人似乎没有得到安息。
HEB|4|2|因为的确有福音传给我们像传给他们一样；只是所听见的道对他们无益，因为他们没有以信心与所听见的道配合。
HEB|4|3|但我们已经信的人进入安息，正如上帝所说： “我在怒中起誓： 他们断不可进入我的安息！” 其实造物之工，从创世以来已经完成了。
HEB|4|4|论到第七日，有一处说：“到第七日，上帝就歇了他一切工作。”
HEB|4|5|又有一处说：“他们断不可进入我的安息！”
HEB|4|6|既有这安息保留着让一些人进入，那些先前听见福音的人，因不信从而不得进去，
HEB|4|7|所以上帝多年后藉着 大卫 的书，又定了一天—“今日”，如以上所引的说： “今日，你们若听他的话， 就不可硬着心。”
HEB|4|8|若是 约书亚 已使他们享了安息，后来上帝就不会再提别的日子了。
HEB|4|9|这样看来，另有一安息日的安息为上帝的子民保留着。
HEB|4|10|因为那些进入安息的，也是歇了自己的工作，正如上帝歇了他的工作一样。
HEB|4|11|所以，我们务必竭力进入那安息，免得有人学了不顺从而跌倒了。
HEB|4|12|上帝的道是活泼的，是有功效的，比一切两刃的剑更锋利，甚至魂与灵、骨节与骨髓，都能刺入、剖开，连心中的思念和主意都能辨明。
HEB|4|13|被造的，没有一样在他面前不是显露的；万物在他眼前都是赤露敞开的，我们必须向他交账。
HEB|4|14|既然我们有一位伟大、进入高天的大祭司，就是耶稣—上帝的儿子，我们应当持定所宣认的道。
HEB|4|15|因为我们的大祭司并非不能体恤我们的软弱；他也在各方面受过试探，与我们一样，只是他没有犯罪。
HEB|4|16|所以，我们只管坦然无惧地来到施恩的宝座前，为要得怜悯，蒙恩惠，作及时的帮助。
HEB|5|1|凡从人间挑选的大祭司都是奉派替人办理属上帝的事，要为罪献上礼物和祭物 。
HEB|5|2|他能体谅无知和迷失的人，因为他自己也是被软弱所困，
HEB|5|3|因此他理当为百姓和自己的罪献祭。
HEB|5|4|没有人可擅自取得大祭司的尊荣，惟有蒙上帝所选召的才可以，像 亚伦 一样。
HEB|5|5|同样，基督也没有自取作大祭司的荣耀，而是在乎向他说话的那一位，他说： “你是我的儿子， 我今日生了你。”
HEB|5|6|就如又有一处说： “你是照着 麦基洗德 的体系 永远为祭司。”
HEB|5|7|基督在他肉身的日子，曾大声哀哭，流泪祷告，恳求那能救他免死的上帝，就因他的虔诚蒙了应允。
HEB|5|8|他虽然为儿子，还是因所受的苦难学了顺从。
HEB|5|9|既然他得以完全，就为凡顺从他的人成了永远得救的根源，
HEB|5|10|并蒙上帝照着 麦基洗德 的体系宣称他为大祭司。
HEB|5|11|论到这事，我们有好些话要说，可是很难解释，因为你们听不进去。
HEB|5|12|按时间说，你们早该作教师了，谁知还需要有人再将上帝圣言基础的要道教导你们；你们成了那需要吃奶、不能吃干粮的人。
HEB|5|13|凡只能吃奶的，就不熟练仁义的道理，因为他是婴孩。
HEB|5|14|惟独长大成人的才能吃干粮，他们的心窍因练习而灵活，能分辨善恶了。
HEB|6|1|所以，我们应当离开基督道理的基础，竭力进到成熟的地步；不必再立根基，就如懊悔致死的行为、信靠上帝、
HEB|6|2|各样洗礼、按手礼、死人复活，以及永远的审判等的教导。
HEB|6|3|上帝若准许，我们就这样做。
HEB|6|4|论到那些已经蒙了光照、尝过天恩的滋味、又于圣灵有份、并尝过上帝的话的美味，和来世权能的人，若再离弃真道，就不可能使他们重新懊悔了；因为他们亲自把上帝的儿子重钉十字架，公然羞辱他。
HEB|6|5|
HEB|6|6|
HEB|6|7|就如一块田地吸收过屡次下的雨水，生长蔬菜，合乎耕种的人用，就从上帝得福。
HEB|6|8|这块田地若长荆棘和蒺藜，必被废弃，近于诅咒，结局就是焚烧。
HEB|6|9|亲爱的，虽然这样说，我们仍深信你们有更好的情况，更接近救恩。
HEB|6|10|因为上帝并非不公义，竟忘记你们的工作和你们为他的名所显的爱心，就是你们过去和现在伺候圣徒的爱心。
HEB|6|11|我们盼望你们各人都显出同样的热忱，一直到底，好达成所确信的指望。
HEB|6|12|这样你们才不会懒惰，却成为效法那些藉着信和忍耐承受应许的人。
HEB|6|13|当初上帝应许 亚伯拉罕 的时候，因为没有比自己更大的可以指着起誓，就指着自己起誓，
HEB|6|14|说：“我必多多赐福给你；我必使你大大增多。”
HEB|6|15|这样， 亚伯拉罕 因恒心等待而得了所应许的。
HEB|6|16|人都是指着比自己大的起誓，并且以起誓作保证，了结各样的争论。
HEB|6|17|照样，上帝愿意为那承受应许的人更有力地显明他的旨意不可更改，他以起誓作保证。
HEB|6|18|藉这两件不可更改的事—在这些事上，上帝绝不会说谎—我们这些逃往避难所的人能得到强有力的鼓励，去抓住那摆在我们前头的指望。
HEB|6|19|我们有这指望，如同灵魂的锚，又坚固又牢靠，进入幔子后面的至圣所。
HEB|6|20|为我们作先锋的耶稣，既照着 麦基洗德 的体系成了永远的大祭司，已经进入了。
HEB|7|1|这 麦基洗德 就是 撒冷 王，是至高上帝的祭司。他在 亚伯拉罕 打败诸王回来的时候迎接他，并给他祝福。
HEB|7|2|亚伯拉罕 也将自己所得来的一切，取十分之一给他。他头一个名字翻译出来是“公义的王”，他又名“ 撒冷 王”，是和平王的意思。
HEB|7|3|他无父、无母、无族谱、无生之始、无命之终，是与上帝的儿子相似，他永远作祭司。
HEB|7|4|你们想一想，这个人多么伟大啊！连先祖 亚伯拉罕 都拿战利品的十分之一给他。
HEB|7|5|那得祭司职分的 利未 子孙，奉命照例向百姓取十分之一，这百姓是自己的弟兄，虽是从 亚伯拉罕 亲身生的，还是照例取十分之一。
HEB|7|6|惟独 麦基洗德 那不与他们同族谱的，从 亚伯拉罕 收取了十分之一，并且给蒙应许的 亚伯拉罕 祝福。
HEB|7|7|向来位分大的给位分小的祝福，这是无可争议的。
HEB|7|8|在这事上，一方面，收取十分之一的都是必死的人；另一方面，收取十分之一的却是那位被证实是活着的。
HEB|7|9|我们可以说，那接受十分之一的 利未 也是藉着 亚伯拉罕 纳了十分之一，
HEB|7|10|因为 麦基洗德 迎接 亚伯拉罕 的时候， 利未 还在他先祖的身体里面。
HEB|7|11|那么，如果百姓藉着 利未 人的祭司职任能达到完全—因为百姓是在这职分下领受律法的—为什么还需要按照 麦基洗德 的体系另外兴起一位祭司，而不按照 亚伦 的体系呢？
HEB|7|12|既然祭司的职分已更改，律法也需要更改。
HEB|7|13|因为这些话所指的人本属别的支派，那支派里从来没有一人在祭坛前事奉的。
HEB|7|14|很明显地，我们的主是从 犹大 出来的；但关于这支派， 摩西 并没有提到祭司。
HEB|7|15|倘若有另一位像 麦基洗德 的祭司兴起来，我的话就更显而易见了。
HEB|7|16|他成为祭司，并不是照属肉身的条例，而是照无穷 生命的大能。
HEB|7|17|因为有给他作见证的说： “你是照着 麦基洗德 的体系 永远为祭司。”
HEB|7|18|一方面，先前的诫命因软弱无能而废掉了，
HEB|7|19|（律法本来就不能成就什么）；另一方面，一个更好的指望被引进来，靠这指望，我们就可以亲近上帝。
HEB|7|20|再者，耶稣成为祭司，并不是没有上帝的誓言；其他的祭司被指派时并没有这种誓言，
HEB|7|21|只有耶稣是起誓立的，因为那位立他的对他说： “主起了誓， 绝不改变。 你是永远为祭司。”
HEB|7|22|既是起誓立的，耶稣也作了更美之约的中保。
HEB|7|23|一方面，那些成为祭司的数目本来多，是因为受死亡限制不能长久留住。
HEB|7|24|另一方面，这位既是永远留住的，他具有不可更换的祭司职任。
HEB|7|25|所以，凡靠着他进到上帝面前的人，他都能拯救到底，因为他长远活着为他们祈求。
HEB|7|26|这样一位圣洁、无邪恶、无玷污、远离罪人、高过诸天的大祭司，对我们是最合适的；
HEB|7|27|他不像那些大祭司，每日必须先为自己的罪，后为百姓的罪献祭，因为他只一次将自己献上就把这事成全了。
HEB|7|28|律法所立的大祭司本是有弱点的人，但在律法以后，上帝以起誓的话立了儿子为大祭司，成为完全，直到永远。
HEB|8|1|我们所讲的事，其中第一要紧的就是：我们有这样一位大祭司，他已经坐在天上至大者宝座的右边，
HEB|8|2|在圣所，就是在真帐幕里作仆役；这帐幕是主所支搭的，不是人所支搭的。
HEB|8|3|凡大祭司都是为献礼物和祭物设立的，所以这位大祭司也必须有所献上。
HEB|8|4|他若在地上，就不用作祭司，因为已经有照律法献礼物的祭司了。
HEB|8|5|他们所供奉的本是天上之事的样式和影像，正如 摩西 将要造帐幕的时候，上帝警戒他，说：“要谨慎，一切都要照着在山上指示你的样式去做。”
HEB|8|6|如今耶稣已经得了更优越的事奉，正如他作更美之约的中保；这约原是凭更美之应许立的。
HEB|8|7|第一个约若没有瑕疵，就无须寻求第二个约了。
HEB|8|8|所以上帝指责他们说： “主说，看哪，日子将到， 我要与 以色列 家 和 犹大 家另立新的约；
HEB|8|9|不像我拉着他们祖宗的手 领他们出 埃及 地的时候， 与他们所立的约； 因为他们不恒心守我的约， 所以我也不理他们；这是主说的。
HEB|8|10|主又说： 那些日子以后， 我与 以色列 家所立的约是这样： 我要将我的律法放在他们的心思里， 写在他们的心上； 我要作他们的上帝， 他们要作我的子民。
HEB|8|11|他们各人不用教导自己的乡亲和自己的弟兄，说：你要认识主； 因为从最小的到最大的， 他们都要认识我。
HEB|8|12|我要宽恕他们的不义， 绝不再记得他们的罪恶。”
HEB|8|13|既然上帝提到“新的约”，那么第一个约就成为旧的了；而那渐旧渐衰的必然很快消逝了。
HEB|9|1|原来连第一个约都有敬拜的礼仪和属世界的圣幕。
HEB|9|2|因为那预备好了的帐幕，第一层叫圣所，里面有灯台、供桌和供饼。
HEB|9|3|第二层幔子后又有一层帐幕，叫至圣所，
HEB|9|4|有金香坛和四周包金的约柜，柜里有盛吗哪的金罐、 亚伦 那根发过芽的杖和两块约版；
HEB|9|5|柜上面有荣耀的基路伯罩着施恩座。有关这一切我现在不能一一细说。
HEB|9|6|这些物件既如此预备齐了，众祭司就不断地进第一层帐幕行拜上帝的礼。
HEB|9|7|至于第二层帐幕，惟有大祭司一年一次独自进去，没有一次不带着血，为自己献上，也为百姓无意所犯的过错献上。
HEB|9|8|圣灵藉此指明，第一层帐幕仍存在的时候，进入至圣所的路还没有显示。
HEB|9|9|那第一层帐幕是现今时代的一个预表，表示所献的礼物和祭物都不能使敬拜的人在良心上得以完全。
HEB|9|10|这些事只不过是有关饮食和各种洁净的规矩，是属肉体的条例，它的功效是直到新次序的时期来到为止。
HEB|9|11|但现在基督已经来到，作了已实现的美事的大祭司，经过那更大更全备的帐幕，不是人手所造，也不是属于这世界的；
HEB|9|12|他不用山羊和牛犊的血，而是用自己的血，只一次进入至圣所就获得了永远的赎罪。
HEB|9|13|若山羊和公牛的血，以及母牛犊的灰，洒在不洁的人身上，尚且使人成圣，身体洁净，
HEB|9|14|何况基督的血，他藉着永远的灵把自己无瑕疵地献给上帝，更能洗净我们 的良心，除去致死的行为，好事奉那位永生的上帝。
HEB|9|15|为此，基督作了新约的中保；因为他的死，赎了人在第一个约之时所犯的罪过，使蒙召的人能得着所应许永远的产业。
HEB|9|16|凡有遗嘱，必须证实立遗嘱的人已经死了。
HEB|9|17|因为人死了，遗嘱才有效力；立遗嘱的人尚在，遗嘱就不能生效。
HEB|9|18|所以，第一个约也是用血立的。
HEB|9|19|因为 摩西 当日照着律法将各样诫命传给众百姓，就拿朱红色绒和牛膝草，把牛犊、山羊 的血和水洒在书上，又洒在众百姓身上，
HEB|9|20|说：“这血就是上帝与你们立约的凭据。”
HEB|9|21|他又照样把血洒在帐幕和敬拜用的各样器皿上。
HEB|9|22|按着律法，几乎每样东西都是用血洁净的；没有流血，就没有赦罪。
HEB|9|23|这样，照着天上样式做的物件必须用这些礼仪去洁净，但那天上的一切，自然当用更美的祭物去洁净。
HEB|9|24|因为基督并没有进了人手所造的圣所—这不过是真圣所的影像—而是进到天上，如今为我们出现在上帝面前。
HEB|9|25|他也无须多次将自己献上，像大祭司每年带着牛羊的血进入至圣所。
HEB|9|26|如果这样，他从创世以来就必须多次受苦了。但如今，他在今世的末期显现，仅一次把自己献为祭，好除掉罪。
HEB|9|27|按着命定，人人都有一死，死后且有审判。
HEB|9|28|同样，基督既然一次献上，担当了许多人的罪，将来要第二次显现，与罪无关，而是为了拯救热切等候他的人。
HEB|10|1|既然律法只不过是未来美好事物的影子，不是本体的真像，就不能藉着每年常献一样的祭物，使那些进前来的人完全。
HEB|10|2|若不然，献祭的事岂不早已停止了吗？因为敬拜的人仅只一次洁净，良心就不再觉得有罪了。
HEB|10|3|但是这些祭物使人每年都想起罪来，
HEB|10|4|因为公牛和山羊的血不能除罪。
HEB|10|5|所以，基督到世上来的时候，就说： “祭物和礼物不是你所要的， 但你曾给我预备了身体。
HEB|10|6|燔祭和赎罪祭 是你不喜欢的。
HEB|10|7|那时我说： 看哪！我来了，我的事在经卷上已经记载了； 上帝啊！我来为要照你的旨意行。”
HEB|10|8|以上说：“祭物和礼物，以及燔祭和赎罪祭，不是你所要的，也不是你喜欢的。”这都是按着律法献的。
HEB|10|9|他接着说：“看哪！我来了，为要照你的旨意行。”可见他除去在先的，为要立定在后的。
HEB|10|10|我们凭着这旨意，藉着耶稣基督，仅只一次献上他的身体就得以成圣。
HEB|10|11|所有的祭司天天站着事奉上帝，屡次献上一样的祭物，这祭物永不能除罪。
HEB|10|12|但基督献了一次永远有效的赎罪祭，就坐在上帝的右边，
HEB|10|13|从此等候他的仇敌成为他的脚凳。
HEB|10|14|因为他仅只一次献祭，就使那些得以成圣的人永远完全。
HEB|10|15|圣灵也对我们作证，因为他说过：
HEB|10|16|“主说：那些日子以后， 我与他们所立的约是这样的： 我要将我的律法放在他们的心上， 又要写在他们的心思里。”
HEB|10|17|并说： “他们的罪恶和他们的过犯， 我绝不再记得。”
HEB|10|18|这些罪过既已蒙赦免，就不用再为罪献祭了。
HEB|10|19|所以，弟兄们，既然我们靠着耶稣的血得以坦然进入至圣所，
HEB|10|20|是藉着他给我们开了一条又新又活的路，从幔子经过，这幔子就是他的身体。
HEB|10|21|既然我们有一位伟大祭司治理上帝的家，
HEB|10|22|那么，我们该用诚心和充足的信心，同已蒙洁净、无亏的良心，和清水洗净了的身体来亲近上帝。
HEB|10|23|我们要坚守所宣认的指望，毫不动摇，因为应许我们的那位是信实的。
HEB|10|24|我们要彼此相顾，激发爱心，勉励行善；
HEB|10|25|不可停止聚会，好像那些停止惯了的人，倒要彼此劝勉，既然知道那日子临近，就更当如此。
HEB|10|26|如果我们领受真理的知识以后仍故意犯罪，就不再有赎罪的祭物，
HEB|10|27|惟有战战兢兢等候审判和那将吞灭众敌人的烈火了。
HEB|10|28|任何人干犯 摩西 的律法，凭两个或三个证人，尚且必须处死，不得宽赦，
HEB|10|29|更何况践踏上帝儿子的人，他们将那使他成圣之约的血当作不洁净，又亵慢施恩的圣灵的人，你们想，他不该受更严厉的惩罚吗？
HEB|10|30|因为我们知道谁说： “伸冤在我， 我必报应。” 又说： “主要审判他的百姓。”
HEB|10|31|落在永生上帝的手里真是可怕呀！
HEB|10|32|你们要追念往日；你们蒙了光照以后，忍受了许多痛苦的挣扎：
HEB|10|33|一面在众人面前公然被毁谤，遭患难；一面陪伴那些受这样苦难的人。
HEB|10|34|你们同情那些遭监禁的人，也欣然忍受你们的家业被人抢去，因为你们知道自己有更美好更长存的家业。
HEB|10|35|所以，不可丢弃你们无惧的心，存这样的心必得大赏赐。
HEB|10|36|你们必须忍耐，使你们行完了上帝的旨意，可以获得所应许的。
HEB|10|37|因为 “还有一点点时候， 那要来的就来，必不迟延。
HEB|10|38|只是我的义人必因信得生； 他若退缩，我心就不喜欢他。”
HEB|10|39|我们却不是退缩以致沉沦的那等人，而是有信心以致得生命的人。
HEB|11|1|信就是对所盼望之事有把握，对未见之事有确据。
HEB|11|2|古人因着这信获得了赞许。
HEB|11|3|因着信，我们知道这宇宙是藉上帝的话造成的。这样，看得见的是从看不见的造出来的。
HEB|11|4|因着信， 亚伯 献祭给上帝比 该隐 所献的更美，因此获得了赞许为义人，上帝亲自悦纳了他的礼物。他虽然死了，却因这信仍旧在说话。
HEB|11|5|因着信， 以诺 被接去，得以不见死，人也找不着他，因为上帝已经把他接去了；只是他被接去以前，已讨得上帝的喜悦而蒙赞许。
HEB|11|6|没有信，就不能讨上帝的喜悦，因为到上帝面前来的人必须信有上帝，并且信他会赏赐寻求他的人。
HEB|11|7|因着信， 挪亚 既蒙上帝指示他未见的事，动了敬畏的心，造了方舟，使他全家得救。藉此他定了那世代的罪，自己也承受了那从信而来的义。
HEB|11|8|因着信， 亚伯拉罕 蒙召的时候就遵命出去，往将来要承受为基业的地方去；他出去的时候还不知往哪里去。
HEB|11|9|因着信，他就在所应许之地作客，好像在异乡，居住在帐棚里，与蒙同一个应许的 以撒 和 雅各 一样。
HEB|11|10|因为他等候着那座有根基的城，就是上帝所设计和建造的。
HEB|11|11|因着信， 撒拉 自己已过了生育的年龄还能怀孕，因为她认为应许她的那位是可信的 ；
HEB|11|12|所以，从一个仿佛已死的人竟生出子孙，如同天上的星那样众多，海边的沙那样无数。
HEB|11|13|这些人都是存着信心死的，并没有得着所应许的，却从远处观望，且欢喜迎接。他们承认自己在地上是客旅，是寄居的。
HEB|11|14|说这样话的人是表明自己要寻找一个家乡。
HEB|11|15|他们若想念所离开的家乡，还有回去的机会。
HEB|11|16|其实他们所羡慕的是一个更美的，就是在天上的家乡。所以，上帝并不因他们称他为上帝 而觉得羞耻，因为他已经为他们预备了一座城。
HEB|11|17|因着信， 亚伯拉罕 被考验的时候把 以撒 献上，这就是那领受了应许的人甘心把自己独生的儿子献上。
HEB|11|18|论到这儿子，上帝曾说：“从 以撒 生的才要称为你的后裔。”
HEB|11|19|他认为上帝甚至能使人从死人中复活，意味着他得回了他的儿子。
HEB|11|20|因着信， 以撒 指着将来的事给 雅各 、 以扫 祝福。
HEB|11|21|因着信， 雅各 临死的时候给 约瑟 的两个儿子个别祝福，扶着拐杖敬拜上帝。
HEB|11|22|因着信， 约瑟 临终的时候提到 以色列 人将来要出 埃及 ，并为自己的骸骨留下遗言。
HEB|11|23|因着信， 摩西 生下来，他的父母见他是个俊美的孩子，把他藏了三个月，并不怕王的命令。
HEB|11|24|因着信， 摩西 长大了不肯称为法老女儿之子。
HEB|11|25|他宁可和上帝的百姓一同受苦，也不愿在罪中享受片刻的欢乐。
HEB|11|26|他把为弥赛亚受凌辱看得比 埃及 的财物更宝贵，因为他想望所要得的赏赐。
HEB|11|27|因着信，他离开 埃及 ，不怕王的愤怒，因为他恒心忍耐，如同看见那不能看见的上帝。
HEB|11|28|因着信，他设立逾越节，在门上洒血，免得那毁灭者加害 以色列 人的长子。
HEB|11|29|因着信，他们过 红海 如行干地； 埃及 人试着要过去就被淹没了。
HEB|11|30|因着信， 以色列 人围绕 耶利哥城 七日，城墙就倒塌了。
HEB|11|31|因着信，妓女 喇合 曾友善地接待探子，就没有跟那些不顺从的人一同灭亡。
HEB|11|32|我还要说什么呢？若要一一细说 基甸 、 巴拉 、 参孙 、 耶弗他 、 大卫 、 撒母耳 和众先知的事，时间就不够了。
HEB|11|33|他们藉着信，制伏了敌国，行了公义，得了应许，堵住了狮子的口，
HEB|11|34|灭了烈火的威力，在锋利的刀剑下逃生，从软弱变为刚强，争战中显出勇猛，打退外邦的全军。
HEB|11|35|有些妇人得回从死人中复活的亲人。又有人忍受严刑，拒绝被释放，为要得着更美好的复活。
HEB|11|36|又有人忍受戏弄、鞭打、捆锁、监禁、各等的磨炼；
HEB|11|37|他们被石头打死，被锯锯死， 被刀杀，披着绵羊山羊的皮各处奔跑，受贫穷、患难、虐待。
HEB|11|38|这世界配不上他们，他们在旷野、山岭、山洞、地穴，飘流无定。
HEB|11|39|这些人都是因信获得了赞许，却仍未得着所应许的，
HEB|11|40|因为上帝给我们预备了更美好的事，若没有我们，他们就不能达到完全。
HEB|12|1|所以，既然我们有这许多见证人如同云彩围绕着我们，就该卸下各样重担和紧紧缠累的罪，以坚忍的心奔那摆在我们前头的路程，
HEB|12|2|仰望我们信心的创始成终者耶稣，他因那摆在前面的喜乐，轻看羞辱，忍受了十字架的苦难，如今已坐在上帝宝座的右边。
HEB|12|3|你们要仔细想想这位忍受了罪人如此顶撞的耶稣，你们就不致心灰意懒了。
HEB|12|4|你们与罪恶争斗，还没有抵抗到流血的地步。
HEB|12|5|你们又忘了上帝劝你们如同劝儿女的那些话，说： “我儿啊，不可轻看主的管教， 被他责备的时候不可灰心；
HEB|12|6|因为主所爱的，他必管教， 又鞭打他所接纳的每一个孩子。”
HEB|12|7|为了受管教，你们要忍受。上帝待你们如同待儿女。哪有儿女不被父亲管教的呢？
HEB|12|8|管教原是众儿女共同所领受的；你们若不受管教，就是私生子，不是儿女了。
HEB|12|9|再者，我们曾有肉身之父管教我们，我们尚且敬重他，何况灵性之父，我们岂不更当顺服他而得生命吗？
HEB|12|10|肉身之父都是短时间随己意管教我们，惟有灵性之父管教我们是要我们得益处，使我们在他的圣洁上有份。
HEB|12|11|凡管教的事，当时不觉得快乐，反觉得痛苦；后来却为那经过锻鍊的人结出平安的果子，就是义的果子。
HEB|12|12|所以，你们要把下垂的手举起来，发酸的腿挺直；
HEB|12|13|要为自己的脚把道路修直了，使瘸了的腿不再脱臼，反而得到痊愈。
HEB|12|14|你们要追求与众人和睦，并要追求圣洁；人非圣洁不能见主。
HEB|12|15|要谨慎，免得有人失去了上帝的恩典；免得有毒根生出来扰乱你们，因而使许多人沾染污秽，
HEB|12|16|免得有人淫乱，或不敬虔如 以扫 ，他因一点点食物把自己长子的名分卖了。
HEB|12|17|后来你们知道，他想要承受父亲的祝福，竟被拒绝，虽然流着泪苦求，却得不着门路使他父亲回心转意。
HEB|12|18|你们不是来到那可触摸的山，那里有火焰、密云、黑暗、暴风、
HEB|12|19|角声，和说话的声音；当时那些听见这声音的，都求不要再向他们说话，
HEB|12|20|因为他们担当不起所命令他们的话，说：“靠近这山的，即使是走兽，也要用石头打死。”
HEB|12|21|所见的景象极其可怕，以致 摩西 说：“我恐惧战兢。”
HEB|12|22|但是你们是来到 锡安山 ，永生上帝的城，就是天上的 耶路撒冷 ，那里有千千万万的天使，
HEB|12|23|有名字记录在天上众长子的盛会，有审判众人的上帝和成为完全的义人的灵魂，
HEB|12|24|并新约的中保耶稣，以及所洒的血；这血所说的信息比 亚伯 的血所说的更美。
HEB|12|25|你们总要谨慎，不可拒绝那向你们说话的，因为那些拒绝了在地上警戒他们的，尚且不能逃罪，何况我们违背那从天上警戒我们的呢？
HEB|12|26|当时他的声音震动了地，但如今他应许说：“再一次我不单要震动地，还要震动天。”
HEB|12|27|这“再一次”的话是指明被震动的要像受造之物一样被挪去，使那不被震动的能常存。
HEB|12|28|所以，既然我们得了不能被震动的国度，就要感恩，照着上帝所喜悦的，用虔诚、敬畏的心事奉上帝，
HEB|12|29|因为我们的上帝是吞灭的火。
HEB|13|1|你们务要常存弟兄相爱的心。
HEB|13|2|不可忘记用爱心接待旅客，因为曾经有人这样做，在无意中接待了天使。
HEB|13|3|要记念受监禁的人，好像与他们同受监禁；要记念受虐待的人，好像你们也亲身受虐待一样。
HEB|13|4|婚姻，人人都当尊重，共眠的床也不可污秽，因为淫乱和通奸的人，上帝必审判。
HEB|13|5|不可贪爱钱财，要以自己所有的为满足，因为上帝曾说：“我绝不撇下你，也绝不丢弃你。”
HEB|13|6|所以，我们可以勇敢地说： “主是我的帮助， 我必不惧怕。 人能把我怎么样呢？”
HEB|13|7|从前引导你们、传上帝的道给你们的人，你们要记念他们，效法他们的信心，回顾他们为人的结局。
HEB|13|8|耶稣基督昨日、今日，一直到永远，是一样的。
HEB|13|9|你们不要被种种怪异的教训勾引了去，因为人的心靠恩典得坚固才是好的，并不是靠饮食。那在饮食上用心的，从来没有得到益处。
HEB|13|10|我们有一祭坛，上面的祭物是那些在会幕中供职的人无权可吃的。
HEB|13|11|因为牲畜的血被大祭司带入至圣所作赎罪祭，牲畜的体却在营外烧掉。
HEB|13|12|所以，耶稣也在城门外受苦，为要用自己的血使百姓成圣。
HEB|13|13|这样，我们也当走出营外，到他那里去，忍受他所受的凌辱。
HEB|13|14|在这里，我们本没有永存的城，而是在寻求那将要来的城。
HEB|13|15|我们应当藉着耶稣，常常以颂赞为祭献给上帝，这是那宣认他名的人嘴唇所结的果子。
HEB|13|16|只是不可忘记行善和分享，因为这样的祭物是上帝所喜悦的。
HEB|13|17|你们要服从那些引导你们的，并且要顺服，因为他们为你们的灵魂时刻警醒，像在上帝面前交账的人，让他们在交账的时候有喜乐，而不是叹息，叹息就对你们无益了。
HEB|13|18|请你们为我们祷告；因为我们自觉良心无亏，愿意凡事按正道而行。
HEB|13|19|我更求你们为我祷告，使我快些回到你们那里去。
HEB|13|20|但愿赐平安 的上帝，就是那凭永约之血，把群羊的大牧人—我们主耶稣从死人中领出来的上帝，
HEB|13|21|在各样善事上装备你们，使你们遵行他的旨意；又藉着耶稣基督在我们 里面行他所喜悦的事。愿荣耀归给他，直到永永远远 。阿们！
HEB|13|22|弟兄们，我简略地写信给你们，希望你们听我劝勉的话。
HEB|13|23|你们该知道，我们的弟兄 提摩太 已经重获自由了；他若很快就来，我必同他去见你们。
HEB|13|24|请你们向带领你们的诸位和众圣徒问安。从 意大利 来的人也向你们问安。
HEB|13|25|愿恩惠与你们众人同在。
JAS|1|1|上帝和主耶稣基督的仆人 雅各 问候散居在各处的十二个支派的人。
JAS|1|2|我的弟兄们，你们遭受各种试炼时，都要认为是大喜乐，
JAS|1|3|因为知道你们的信心经过考验，就生忍耐。
JAS|1|4|但要让忍耐发挥完全的功用，使你们能又完全又完整，一无所缺。
JAS|1|5|你们中间若有缺少智慧的，该求那厚赐与众人又不斥责人的上帝，上帝必赐给他。
JAS|1|6|只要凭着信心求，一点也不疑惑；因为那疑惑的人，就像海中的波浪被风吹动翻腾。
JAS|1|7|这样的人不要想从主那里得到什么。
JAS|1|8|三心二意的人，在他一切所行的路上都摇摆不定。
JAS|1|9|卑微的弟兄要因高升而夸耀，
JAS|1|10|富足的却要因被降卑而夸耀，因为富足的人要消逝，如同草上的花一样。
JAS|1|11|太阳出来，热风刮起，草就枯干，花也凋谢，它美丽的样子就消失了；那富足的人在他一生的奔波中也要这样衰残。
JAS|1|12|忍受试炼的人有福了，因为他经过考验以后必得生命的冠冕，这是主应许给爱他之人的。
JAS|1|13|人被诱惑，不可说：“我是被上帝诱惑”；因为上帝是不被恶诱惑的，他也不诱惑人。
JAS|1|14|但每一个人被诱惑是因自己的私欲牵引而被诱惑的。
JAS|1|15|私欲既怀了胎，就生出罪来；罪既长成，就生出死来。
JAS|1|16|我亲爱的弟兄们，不要被欺骗了。
JAS|1|17|各样美善的恩泽和各样完美的赏赐都是从上头来的，从众光之父那里降下来的；在他并没有改变，也没有转动的影儿。
JAS|1|18|他按自己的旨意，用真理的道生了我们，使我们在他所造的万物中成为初熟的果子。
JAS|1|19|我亲爱的弟兄们，你们要明白：你们每一个人要快快地听，慢慢地说，慢慢地动怒，
JAS|1|20|因为人的怒气并不能实现上帝的义。
JAS|1|21|所以，你们要除去一切的污秽和累积的恶毒，要存温柔的心领受所栽种的道，就是能救你们灵魂的道。
JAS|1|22|但是，你们要作行道的人，不要只作听道的人，自己欺骗自己。
JAS|1|23|因为只听道而不行道的，就像人对着镜子观看自己本来的面目，
JAS|1|24|注视后，就离开，立刻忘了自己的相貌如何。
JAS|1|25|惟有查看那完美、使人自由的律法，并且时常遵守的，他不是听了就忘，而是切实行出来，这样的人在所行的事上必然蒙福。
JAS|1|26|若有人自以为虔诚，却不勒住自己的舌头，反欺骗自己的心，这人的虔诚是徒然的。
JAS|1|27|在上帝—我们的父面前，清洁没有玷污的虔诚就是看顾在患难中的孤儿寡妇，并且保守自己不沾染世俗。
JAS|2|1|我的弟兄们，你们信奉我们荣耀的主耶稣基督，就不可按着外貌待人。
JAS|2|2|若有一个人戴着金戒指，穿着华丽的衣服，进入你们的会堂，又有一个穷人穿着肮脏的衣服也进去，
JAS|2|3|而你们只看重那穿华丽衣服的人，说：“请坐在这里”，又对那穷人说：“你站在那里”，或“坐在我脚凳旁”；
JAS|2|4|这岂不是你们偏心待人，用恶意评断人吗？
JAS|2|5|我亲爱的弟兄们，请听，上帝岂不是拣选了世上的贫穷人，使他们在信心上富足，并承受他所应许给那些爱他之人的国吗？
JAS|2|6|你们却羞辱贫穷的人。欺压你们，拉你们到公堂去的，不就是这些富有的人吗？
JAS|2|7|毁谤为你们求告时所奉的尊名的，不就是他们吗？
JAS|2|8|经上记着：“要爱邻 如己”，你们若切实守这至尊的律法，你们就做得很好。
JAS|2|9|但你们若按外貌待人就是犯罪，是被律法定为犯法的。
JAS|2|10|因为凡遵守全部律法的，只违背了一条就是违犯了所有的律法。
JAS|2|11|原来那说“不可奸淫”的，也说“不可杀人”。你就是不奸淫，却杀人，也是成为违犯律法的。
JAS|2|12|既然你们要按使人自由的律法受审判，就要照这律法说话行事。
JAS|2|13|因为对那不怜悯人的，他们要受没有怜悯的审判；怜悯胜过审判。
JAS|2|14|我的弟兄们，若有人说自己有信心，却没有行为，有什么益处呢？这信心能救他吗？
JAS|2|15|若是弟兄或是姊妹没有衣服穿，又缺少日用的饮食；
JAS|2|16|你们中间有人对他们说：“平平安安地去吧！愿你们穿得暖，吃得饱”，却不给他们身体所需要的，这有什么益处呢？
JAS|2|17|信心也是这样，若没有行为是死的。
JAS|2|18|但是有人会说：“你有信心，我有行为。”把你没有行为的信心给我看，我就藉着我的行为把我的信心给你看。
JAS|2|19|你信上帝只有一位，你信得很好；连鬼魔也信，且怕得发抖。
JAS|2|20|你这虚浮的人哪，你愿意知道没有行为的信心是没有用的吗？
JAS|2|21|我们的祖宗 亚伯拉罕 把他儿子 以撒 献在坛上，岂不是因行为得称义吗？
JAS|2|22|可见信心是与他的行为相辅并行，而且信心是因着行为才得以成全的。
JAS|2|23|这正应验了经上所说：“ 亚伯拉罕 信了上帝，这就算他为义”；他又得称为上帝的朋友。
JAS|2|24|这样看来，人称义是因着行为，不是单因着信。
JAS|2|25|同样，妓女 喇合 接待使者，又放他们从另一条路出去，不也是因行为称义吗？
JAS|2|26|所以，就如身体没有灵魂是死的，信心没有行为也是死的。
JAS|3|1|我的弟兄们，不要许多人做教师，因为你们知道，我们做教师的要接受更严厉的审判。
JAS|3|2|原来我们在许多事上都有过失；若有人在言语上没有过失，他就是完全的人，也能勒住自己的全身。
JAS|3|3|我们若把嚼环放在马嘴里使它们驯服，就能控制它们的全身。
JAS|3|4|再看船只，虽然甚大，又被强风猛吹，只用小小的舵就随着掌舵的意思转动。
JAS|3|5|同样，舌头是小肢体，却能说大话。 看哪，最小的火能点燃最大的树林。
JAS|3|6|舌头就是火。在我们百体中，舌头是个不义的世界，能玷污全身，也能烧毁生命的轮子，而且是被地狱的火点燃的。
JAS|3|7|各类的走兽、飞禽、爬虫、水族，本来都可以制伏，也已经被人制伏了；
JAS|3|8|惟独舌头没有人能制伏，是永不静止的邪恶，充满了害死人的毒气。
JAS|3|9|我们用舌头颂赞我们的主—我们的天父，又用舌头诅咒照着上帝形像被造的人。
JAS|3|10|颂赞和诅咒从同一个口出来。我的弟兄们，这是不应该的。
JAS|3|11|泉源能从一个出口发出甜苦两样的水吗？
JAS|3|12|我的弟兄们，无花果树能生橄榄吗？葡萄树能结无花果吗？咸水也不能流出甜水来。
JAS|3|13|你们中间谁是有智慧有见识的呢？他就当在智慧的温柔上显出他的善行来。
JAS|3|14|你们心里若怀着恶毒的嫉妒和自私，就不可自夸，不可说谎话抵挡真理。
JAS|3|15|这样的智慧不是从上头下来的，而是属地上的，属情欲的，属鬼魔的。
JAS|3|16|在何处有嫉妒、自私，在何处就有动乱和各样的坏事。
JAS|3|17|惟独从上头来的智慧，先是清洁，后是和平、温良、柔顺，满有怜悯和美善的果子，没有偏私，没有虚伪。
JAS|3|18|正义的果实是为促进和平的人用和平栽种出来的。
JAS|4|1|你们中间的冲突是哪里来的？争执是哪里来的？不是从你们肢体中交战着的私欲来的吗？
JAS|4|2|你们贪恋，得不着就杀人；你们嫉妒，不能得手就起争执和冲突；你们得不着，是因为你们不求。
JAS|4|3|你们求也得不着，是因为你们妄求，为了要浪费在你们的宴乐中。
JAS|4|4|你们这些淫乱的人哪，岂不知道与世俗为友就是与上帝为敌吗？所以，凡想要与世俗为友的，就是与上帝为敌了。
JAS|4|5|经上说：“上帝爱安置在我们里面的灵，爱到嫉妒的地步。” 你们以为这话是徒然的吗？
JAS|4|6|但是他赐更多的恩典，正如经上说： “上帝抵挡骄傲的人， 但赐恩给谦卑的人。”
JAS|4|7|所以，要顺服上帝。要抵挡魔鬼，魔鬼就必逃避你们；
JAS|4|8|要亲近上帝，上帝就必亲近你们。有罪的人哪，要洁净你们的手！心怀二意的人哪，要清洁你们的心！
JAS|4|9|你们要愁苦，悲哀，哭泣；要将欢笑变为悲哀，欢乐变为愁闷。
JAS|4|10|要在主面前谦卑，他就使你们高升。
JAS|4|11|弟兄们，不可彼此诋毁。诋毁弟兄或评断弟兄的人，就是诋毁律法，评断律法；你若评断律法，就不是遵行律法，而是评断者了。
JAS|4|12|立法者和审判者只有一位；他就是那能拯救人也能毁灭人的。你是谁，竟敢评断你的邻舍！
JAS|4|13|注意！有人说：“今天或明天我们要往某城去，在那里住一年，做买卖赚钱。”
JAS|4|14|其实明天如何，你们还不知道。你们的生命是什么呢？你们 原来是一片云雾，出现片刻就不见了。
JAS|4|15|你们倒应当说：“主若愿意，我们就能活着，也可以做这事或那事。”
JAS|4|16|现今你们竟然狂傲自夸；凡这样的自夸都是邪恶的。
JAS|4|17|所以，人若知道该行善而不去行，这就是他的罪了。
JAS|5|1|注意！你们这些富足人哪，要为将要临到你们身上的灾难哭泣、号啕。
JAS|5|2|你们的财物腐烂了，你们的衣服被虫子蛀了。
JAS|5|3|你们的金银都生锈了；这锈要证明你们的不是，又要像火一样吞吃你们的肉。你们在这末世只知道积蓄钱财。
JAS|5|4|工人给你们收割庄稼，你们克扣他们的工钱；这工钱在喊冤，而且收割工人的冤声已经进入万军之主的耳朵了。
JAS|5|5|你们在地上享奢华宴乐，把自己养肥了，等候宰杀的日子。
JAS|5|6|你们定了义人的罪，把他杀害，他没有抵抗你们。
JAS|5|7|所以弟兄们，你们要忍耐，直到主来。看哪，农夫等候着地里宝贵的出产，耐心地等到它得了秋霖春雨。
JAS|5|8|你们也要忍耐，坚固你们的心，因为主来的日子近了。
JAS|5|9|弟兄们，你们不要彼此埋怨，免得受审判。看哪，审判的主站在门口了。
JAS|5|10|弟兄们，你们要把那先前奉主名说话的众先知作能受苦、能忍耐的榜样。
JAS|5|11|看哪，那些忍耐的人，我们称他们是有福的。你们听见过 约伯 的忍耐，也看见主给他的结局，知道主是充满怜悯和慈悲的。
JAS|5|12|我的弟兄们，最要紧的是不可起誓；不可指着天起誓，也不可指着地起誓，任何誓都不可起。你们说话，是，就说是；不是，就说不是，免得你们落在审判之下。
JAS|5|13|你们中间若有人受苦，他该祷告；有人喜乐，他该歌颂。
JAS|5|14|你们中间若有人病了，他该请教会的长老们来为他祷告，奉主的名为他抹油。
JAS|5|15|出于信心的祈祷必能救那病人，主必叫他起来；他若犯了罪，也必蒙赦免。
JAS|5|16|所以，你们要彼此认罪，互相代求，使你们得医治。义人祈祷所发的力量是大有功效的。
JAS|5|17|以利亚 与我们是同样性情的人，他恳切地祈求不要下雨，地上就三年六个月没有下雨。
JAS|5|18|他又祷告，天就降下雨来，地就有了出产。
JAS|5|19|我的弟兄们，你们中间若有人迷失了真理而有人使他回转，
JAS|5|20|这人该知道，使一个罪人从迷途中回转，会从死亡中把他的灵魂救回来，而且遮盖许多的罪。
1PET|1|1|耶稣基督的使徒 彼得 写信给那些被拣选，分散在 本都 、 加拉太 、 加帕多家 、 亚细亚 、 庇推尼 寄居的人，
1PET|1|2|就是照父上帝的预知，藉着圣灵得以成圣，以致顺服耶稣基督，又蒙他血所洒的人。愿恩惠、平安 多多地赐给你们！
1PET|1|3|愿颂赞归于我们主耶稣基督的父上帝！他曾照自己的大怜悯，藉着耶稣基督从死人中复活，重生了我们，使我们有活的盼望，
1PET|1|4|好得到不朽坏、不玷污、不衰残、为你们存留在天上的基业，
1PET|1|5|就是为你们这些藉着信、蒙上帝大能保守的人，能获得他所预备、到末世要显现的救恩。
1PET|1|6|虽然你们必须在百般试炼中暂时忧愁，你们要为此喜乐 ，
1PET|1|7|使你们的信心既被考验，就比那被火试炼仍然能坏的金子更显宝贵，可以在耶稣基督显现的时候得著称赞、荣耀、尊贵。
1PET|1|8|虽然你们没有见过他，却是爱他；如今虽看不见，你们却因信他而有说不出来、满有荣光的喜乐，
1PET|1|9|因为你们 得到信心的效果，就是灵魂的得救。
1PET|1|10|论到这救恩，那预先说你们要得恩典的众先知已经详细地搜索查考过，
1PET|1|11|查考在他们心里的基督的灵预先证明基督受苦难，后来得荣耀，是指什么时候，什么样的情况。
1PET|1|12|他们得了启示，知道他们所服事的不是自己，而是你们。那藉着从天上差来的圣灵传福音给你们的人，现在将这些事传给你们；这些事连天使也都切望察看呢！
1PET|1|13|所以，要准备 好你们的心，谨慎自守，专心盼望耶稣基督显现的时候带给你们的恩惠。
1PET|1|14|作为顺服的儿女，就不要效法从前蒙昧无知的时候那放纵私欲的样子。
1PET|1|15|但那召你们的既是圣洁，你们在一切所行的事上也要圣洁；
1PET|1|16|因为经上记着：“你们要成为圣，因为我是神圣的。”
1PET|1|17|既然你们称那不偏待人、按各人行为审判人的主为父 ，就当存敬畏的心，度你们在世寄居的日子。
1PET|1|18|你们知道，你们得以从你们祖先传下来虚妄的行为中救赎出来，不是靠着会朽坏的金银等物，
1PET|1|19|而是凭着基督的宝血，如同无瑕疵、无玷污的羔羊的血。
1PET|1|20|基督是上帝在创世以前所预知，而在这末世才为你们显现的。
1PET|1|21|你们也因着他而信那使他从死人中复活、又给他荣耀的上帝，好让你们的信心和盼望都在于上帝。
1PET|1|22|既然你们因顺从真理而洁净了自己的心灵，能真诚爱弟兄，就该以清洁的心 彼此切实相爱。
1PET|1|23|你们蒙了重生，不是由于会朽坏的种子，而是由于不会朽坏的种子，是藉着上帝永活常存的道。
1PET|1|24|因为 “凡血肉之躯的尽都如草， 他的一切荣美像草上的花； 草必枯干，花必凋谢，
1PET|1|25|惟有主的道永远常存。” 这话就是传给你们的福音。
1PET|2|1|所以，你们要除去一切的恶毒，一切诡诈、假善、嫉妒，和一切毁谤的话。
1PET|2|2|要爱慕那纯净的灵奶，像初生的婴孩爱慕奶一样，好使你们藉着它成长，以致得救，
1PET|2|3|因为你们已经尝过主恩的滋味。
1PET|2|4|要亲近主，他是活石，虽然被人所丢弃，却是上帝所拣选、所珍贵的。
1PET|2|5|你们作为活石，要被建造成属灵的殿，成为圣洁的祭司，藉着耶稣基督献上蒙上帝悦纳的属灵祭物。
1PET|2|6|因为经上说： “看哪，我把一块石头放在 锡安 — 一块蒙拣选、珍贵的房角石； 信靠他的人必不蒙羞。”
1PET|2|7|所以，这石头在你们信的人是珍贵的；在那不信的人却有话说： “匠人所丢弃的石头 已作了房角的头块石头。”
1PET|2|8|又说： “作了绊脚的石头， 使人跌倒的磐石。” 他们绊跌，因为不顺从这道，这也是预定的。
1PET|2|9|不过，你们是被拣选的一族，是君尊的祭司，是神圣的国度，是属上帝的子民，要使你们宣扬那召你们出黑暗入奇妙光明者的美德。
1PET|2|10|“你们从前不是子民， 现在却成了上帝的子民； 从前未曾蒙怜悯， 现在却蒙了怜悯。”
1PET|2|11|亲爱的，你们是客旅，是寄居的，我劝你们要禁戒肉体的情欲；这情欲是与灵魂争战的。
1PET|2|12|你们在外邦人中要品行端正，好让那些人，虽然毁谤你们是作恶的，会因看见你们的好行为而在鉴察 的日子归荣耀给上帝。
1PET|2|13|你们为主的缘故要顺服人的一切制度，或是在上的君王，
1PET|2|14|或是君王所派惩恶赏善的官员。
1PET|2|15|因为上帝的旨意原是要你们以行善来堵住糊涂无知人的口。
1PET|2|16|虽然你们是自由的，却不可藉着自由遮盖恶毒，总要作上帝的仆人。
1PET|2|17|务要尊重众人；要敬爱教中的弟兄姊妹；要敬畏上帝；要尊敬君王。
1PET|2|18|你们作奴仆的，凡事要存敬畏的心顺服主人；不但顺服善良温和的，就是乖僻的也要顺服。
1PET|2|19|倘若你们为使良心对得起上帝，忍受冤屈的痛苦，这是可赞许的。
1PET|2|20|你们若因犯罪受责打而忍耐，有什么可称赞的呢？但你们若因行善受苦而忍耐，这在上帝看来是可赞许的。
1PET|2|21|你们蒙召就是为此，因为基督也为你们受过苦，给你们留下榜样，为要使你们跟随他的脚踪。
1PET|2|22|“他并没有犯罪， 口里也没有诡诈。”
1PET|2|23|他被辱骂不还口，受害也不说威吓的话，只将自己交托给公义的审判者。
1PET|2|24|他被挂在木头上，亲身担当了我们的罪，使我们既然在罪上死，就得以在义上活。因他受的鞭伤，你们得了医治。
1PET|2|25|你们从前好像迷路的羊，如今却归回你们灵魂的牧人和监督了。
1PET|3|1|同样，你们作妻子的，要顺服自己的丈夫，这样，即使有不信从道理的丈夫，也会因妻子的品行，并非言语，而感化过来，
1PET|3|2|因为看见了你们敬虔纯洁的品行。
1PET|3|3|你们不要藉外表来妆饰自己，如编头发，戴金饰，穿美丽的衣裳等，
1PET|3|4|而要有蕴藏在人内心不衰退的美，以温柔娴静的心妆饰自己；这在上帝面前是极宝贵的。
1PET|3|5|因为古时仰赖上帝的圣洁妇人正是以此为妆饰，顺服自己的丈夫。
1PET|3|6|就如 撒拉 听从 亚伯拉罕 ，称他为主。你们只要行善，不怕任何恐吓，就成为 撒拉 的女儿了。
1PET|3|7|同样，你们作丈夫的，要按情理 跟妻子共同生活，体贴女性是比较软弱的器皿；要尊重她，因为她也与你一同承受生命之恩。这样，你们的祷告就不会受阻碍。
1PET|3|8|总而言之，你们都要同心，彼此体恤，相爱如弟兄，存怜悯和谦卑的心。
1PET|3|9|不要以恶报恶，以辱骂还辱骂，倒要祝福，因为你们正是为此蒙召的，好使你们承受福气。
1PET|3|10|因为经上说： “凡要爱惜生命、 享受好日子的人， 要禁止舌头不出恶言， 嘴唇不说诡诈的话。
1PET|3|11|也要弃恶行善， 寻求和睦，一心追求。
1PET|3|12|因为主的眼看顾义人， 他的耳听他们的祈祷； 但主向行恶的人变脸。”
1PET|3|13|你们若热心行善，有谁会害你们呢？
1PET|3|14|即使你们为义受苦，也是有福的。不要怕人的威吓，也不要惊慌；
1PET|3|15|只要心里奉主基督为圣，尊他为主。有人问你们心中盼望的理由，要随时准备答覆；
1PET|3|16|不过，要以温柔、敬畏的心回答。要存无亏的良心，使你们在何事上被毁谤，就在何事上使那些凌辱你们在基督里有好品行的人自觉羞愧。
1PET|3|17|上帝的旨意若是要你们因行善受苦，这总比因行恶受苦好。
1PET|3|18|因为基督也曾一次为罪受苦 ， 就是义的代替不义的， 为要引领你们 到上帝面前。 在肉体里，他被治死； 但在灵里，他复活了。
1PET|3|19|他藉这灵也曾去向那些在监狱里的灵传道，
1PET|3|20|就是那些从前在 挪亚 预备方舟、上帝容忍等待的时候不信从的人。当时进入方舟，藉着水得救的不多，只有八个人。
1PET|3|21|这水所预表的洗礼，现在藉着耶稣基督的复活拯救你们，不是除掉肉体的污秽，而是向上帝恳求有无亏的良心。
1PET|3|22|耶稣已经到天上去，在上帝的右边，众天使、有权柄的、有权能的都服从了他。
1PET|4|1|既然基督在肉身受苦，你们也该将这样的心志作为兵器，因为在肉身受过苦的已经与罪断绝了，
1PET|4|2|使你们从今以后不再随从人的情欲，只顺从上帝的旨意，在世度余下的光阴。
1PET|4|3|因为你们从前随从外邦人的心意，生活在淫荡、情欲、醉酒、荒宴、狂饮和可憎的偶像崇拜中，时候已经够了。
1PET|4|4|在这些事上，他们见你们不与他们同奔放荡无度的路就以为怪，毁谤你们。
1PET|4|5|他们必须在那位将要审判活人死人的主面前交账。
1PET|4|6|为此，死人也曾有福音传给他们，要使他们的肉体按着人受审判，他们的灵却靠上帝活着。
1PET|4|7|万物的结局近了。所以你们要谨慎自守，要警醒祷告。
1PET|4|8|最要紧的是彼此切实相爱，因为爱能遮掩许多的罪。
1PET|4|9|你们要互相款待，不发怨言。
1PET|4|10|人人要照自己所得的恩赐彼此服事，作上帝各种恩赐的好管家。
1PET|4|11|若有人讲道，他要按着上帝的圣言讲；若有人服事，他要按着上帝所赐的力量服事，好让上帝在凡事上因耶稣基督得荣耀。愿荣耀和权能都归给他，直到永永远远。阿们！
1PET|4|12|亲爱的，有火一般的考验临到你们，不要奇怪，似乎是遭遇非常的事；
1PET|4|13|倒要欢喜，因为你们是与基督一同受苦，使你们在他荣耀显现的时候也可以欢喜快乐。
1PET|4|14|你们若为基督的名受辱骂是有福的，因为荣耀的灵，就是上帝的灵，在你们身上。
1PET|4|15|你们中间，不可有人因为杀人、偷窃、作恶、好管闲事而受苦。
1PET|4|16|若有人因是基督徒而受苦，不要引以为耻，倒要因这名而归荣耀给上帝。
1PET|4|17|因为时候到了，审判要从上帝的家开始；若是先从我们开始，那么，不信从上帝福音的人将有何等的结局呢？
1PET|4|18|“若是义人还仅仅得救， 不虔敬和犯罪的人将有何地可站呢？”
1PET|4|19|所以，照上帝旨意受苦的人要一心为善，将自己的灵魂交给那信实的造物主。
1PET|5|1|所以，我这同作长老，作基督受苦的证人和分享将来所要显现的荣耀的人，勉励在你们中间的长老们：
1PET|5|2|务要牧养在你们当中上帝的群羊，按着上帝的旨意照顾他们 ，不是出于勉强，而是出于甘心；也不是因为贪财，而是出于乐意。
1PET|5|3|不要辖制所托付你们的群羊，而是要作他们的榜样。
1PET|5|4|到了大牧人显现的时候，你们必得到那永不衰残、荣耀的冠冕。
1PET|5|5|同样，你们年轻的，要顺服年长的。你们大家都要以谦卑当衣服穿上，彼此顺服，因为 “上帝抵挡骄傲的人， 但赐恩给谦卑的人。”
1PET|5|6|所以，你们要谦卑服在上帝大能的手下，这样，到了适当的时候，他必使你们升高。
1PET|5|7|你们要将一切的忧虑卸给上帝，因为他顾念你们。
1PET|5|8|务要谨慎，要警醒。因为你们的仇敌魔鬼，如同咆哮的狮子，走来走去，寻找可吞吃的人。
1PET|5|9|你们要用坚固的信心抵挡他，因为知道你们在世上的众弟兄也正在经历这样的苦难。
1PET|5|10|那赐一切恩典的上帝曾在基督 里召了你们，得享他永远的荣耀，在你们暂受苦难之后，必要亲自成全你们，坚固你们，赐力量给你们，建立你们 。
1PET|5|11|愿权能归给他，直到永永远远。阿们！
1PET|5|12|我简单地写了这信，托我所看为忠心的弟兄 西拉 交给你们，劝勉你们，又证明这恩是上帝真实的恩典；你们务要在这恩上站立得住。
1PET|5|13|在 巴比伦 与你们同蒙拣选的教会向你们问安。我儿子 马可 也向你们问安。
1PET|5|14|你们要用爱心彼此亲吻问安。愿平安 归给你们所有在基督里的人！
2PET|1|1|耶稣基督的仆人和使徒 西门．彼得 写信给那因我们的上帝和 救主耶稣基督的义，与我们同得一样宝贵信心的人。
2PET|1|2|愿恩惠、平安 ，因你们认识上帝和我们的主耶稣，多多加给你们！
2PET|1|3|上帝的神能已把一切关乎生命和虔敬的事赐给我们，因我们认识那用自己荣耀和美德召我们的上帝。
2PET|1|4|因此，他已把又宝贵又极大的应许赐给我们，使我们既脱离世上从情欲来的败坏，就得分享上帝的本性。
2PET|1|5|正因这缘故，你们要分外地努力。有了信心，又要加上德行；有了德行，又要加上知识；
2PET|1|6|有了知识，又要加上节制；有了节制，又要加上忍耐；有了忍耐，又要加上虔敬；
2PET|1|7|有了虔敬，又要加上爱弟兄的心；有了爱弟兄的心，又要加上爱众人的心。
2PET|1|8|你们有了这几样，再继续增长，就必使你们在认识我们的主耶稣基督上，不至于懒散和不结果子了。
2PET|1|9|没有这几样的人就是瞎眼，是短视，忘了他过去的罪已经得了洁净。
2PET|1|10|所以，弟兄们，要更加努力，使你们的蒙召和被选坚定不移。你们实行这几样，就永不失脚。
2PET|1|11|这样，必叫你们丰丰富富地得以进入我们主－救主耶稣基督永远的国度。
2PET|1|12|虽然你们已经知道这些事，并且在你们已有的真道上得到坚固，我还是要常常提醒你们这些事。
2PET|1|13|我认为趁我还在这帐棚的时候，应该激发你们的记忆，
2PET|1|14|因为知道我脱离这帐棚的时候快到了，正如我们的主耶稣基督所指示我的。
2PET|1|15|我也要尽心竭力，使你们在我去世以后时常记念这些事。
2PET|1|16|我们从前把我们主耶稣基督的大能和他来临的事告诉你们，并不是随从一些捏造出来的无稽传说，我们是曾经亲眼见过他的威荣的人。
2PET|1|17|他从父上帝得尊贵荣耀的时候，从至高无上的荣耀有声音出来，对他说：“这是我的爱子，我所喜悦的。”
2PET|1|18|我们同他在圣山的时候，亲自听见这声音从天上出来。
2PET|1|19|我们有先知更确实的信息，你们要好好地留意这信息，如同留意照耀在暗处的明灯，直等到天亮，晨星在你们心里升起的时候。
2PET|1|20|第一要紧的，你们要知道，经上所有的预言是不可随私意解释的，
2PET|1|21|因为预言从来没有出于人意的，而是人被圣灵感动说出上帝的话来。
2PET|2|1|从前在民间有假先知起来；同样，将来在你们中间也会有假教师，偷偷地引进使人灭亡的异端。他们甚至不认买他们的主人，自取迅速灭亡。
2PET|2|2|许多人会随从他们淫荡的行为，以致真理之道因他们的缘故被毁谤。
2PET|2|3|他们因贪婪，要用捏造的言语在你们身上取得利益。他们的惩罚，自古以来并不迟延；他们的灭亡也必迅速来到。
2PET|2|4|既然上帝没有宽容犯了罪的天使，反而把他们丢在地狱里，囚禁在幽暗中等候审判；
2PET|2|5|既然上帝也没有宽容上古的世界，曾叫洪水临到那不敬虔的世界，只保护了报公义信息的 挪亚 一家八口；
2PET|2|6|既然上帝判决了 所多玛 和 蛾摩拉 ，将二城倾覆 ，焚烧成灰，作为后世不敬虔人的鉴戒，
2PET|2|7|只搭救了那常为恶人的淫荡忧伤的义人 罗得 —
2PET|2|8|因为那义人住在他们当中，他正义的心因天天看见和听见他们不法的事而伤痛；
2PET|2|9|那么，主知道搭救敬虔的人脱离试炼，把不义的人留在惩罚之下等候审判的日子，
2PET|2|10|尤其那些随从肉体、放纵污秽的情欲、藐视主的权威的人更是如此。 他们胆大任性，无惧地毁谤众尊荣者；
2PET|2|11|就是天使，虽然力量权能更大，在对他们宣告从主来的审判的时候还不用毁谤的话 。
2PET|2|12|但这些人好像没有理性的牲畜，生来就是要被捉拿宰杀的。他们毁谤自己所不知道的事，正在败坏人的时候，自己也遭遇败坏，
2PET|2|13|为所行的不义受不义的工钱。他们喜爱白昼狂欢，他们已被玷污，又有瑕疵，正与你们一同欢宴，以自己的诡诈为乐。
2PET|2|14|他们满眼是淫色，是止不住的罪，引诱心不坚定的人，心中习惯了贪婪，正是被诅咒的种类。
2PET|2|15|他们离弃了正路，走入歧途，随从 比珥 的儿子 巴兰 的路； 巴兰 就是那贪爱不义的工钱的人，
2PET|2|16|他却为自己的过犯受了责备，而那不能说话的驴以人的声音阻止了先知的狂妄。
2PET|2|17|这些人是无水的泉源，是狂风催逼的雾气，有漆黑的幽暗为他们存留。
2PET|2|18|他们说虚妄夸大的话，用肉体的情欲和淫荡的事引诱那些刚脱离错谬生活的人。
2PET|2|19|他们应许人自由，自己却作了腐败的奴隶，因为人被谁制伏就是谁的奴隶。
2PET|2|20|倘若他们因认识我们的主和救主耶稣基督而得以脱离世上的污秽，后来又被污秽缠住，被制伏，他们末后的景况就比先前更不好了。
2PET|2|21|他们知道义路，竟背弃了传授给他们那神圣的诫命，倒不如不知道为妙。
2PET|2|22|俗语说得好，这话正印证在他们身上了： “狗转过来吃自己所吐的；” 又说： “猪洗净了，又回到烂泥里打滚。”
2PET|3|1|亲爱的，我现在写给你们的是第二封信。在这两封信里，我都提醒你们，激发你们真诚的心，
2PET|3|2|要你们记得圣先知预先所说的话和主—救主的命令，就是使徒所传给你们的。
2PET|3|3|第一要紧的，你们要知道，在末世必有好讥诮的人随从自己的私欲出来讥诮，
2PET|3|4|说：“他要来临的应许在哪里呢？因为从列祖长眠以来，万物与起初创造的时候仍是一样啊！”
2PET|3|5|他们故意忘记这事，就是从太古凭上帝的话有了天，并由水而出和藉着水而成的地；
2PET|3|6|藉着水，当时的世界被水淹没而消灭了。
2PET|3|7|但现在的天地还是凭着上帝的话存留，直留到不敬虔之人受审判遭沉沦的日子，用火焚烧。
2PET|3|8|亲爱的，有一件事你们不可忘记，就是：主看一日如千年，千年如一日。
2PET|3|9|主没有迟延他的应许，就如有人以为他是迟延，其实他是宽容你们，不愿一人沉沦，而是人人都来悔改。
2PET|3|10|但主的日子要像贼一样来到；那日，天必在轰然一声中消失，天体都要被烈火熔化，地和地上的万物都要烧尽 。
2PET|3|11|既然这一切都要如此消失，你们 处世为人必须圣洁敬虔，
2PET|3|12|等候并催促上帝的日子来到。因为在那日，天要被火烧而消灭，天体都要被烈火熔化。
2PET|3|13|但照他的应许，我们等候新天新地，其中有正义常住。
2PET|3|14|所以，亲爱的，既然你们等候这些事，就要竭力使自己没有玷污，无可指责，在主前和睦；
2PET|3|15|并且要以我们主的容忍作为你们得救的机会，就如我们所亲爱的弟兄 保罗 ，照着所赐给他的智慧写信给你们。
2PET|3|16|他一切的信上都谈到这事。信中有些难明白的，那无学问、不坚定的人加以曲解，如曲解别的经书一样，自取灭亡。
2PET|3|17|所以，亲爱的，既然你们预先知道这事，就当防备，免得被恶人的错谬诱惑，从自己稳定的立场上坠落。
2PET|3|18|你们倒要在我们的主和救主耶稣基督的恩典和知识上有长进。愿荣耀归给他，从今直到永远之日。阿们！
1JOHN|1|1|论到从起初原有的生命之道，就是我们所听见、所看见、亲眼看过、亲手摸过的－
1JOHN|1|2|这生命已经显现出来，我们看见了，现在又作见证，把原与父同在，并且向我们显现过的那永远的生命传扬给你们－
1JOHN|1|3|我们把所看见、所听见的传扬给你们，为要使你们也与我们有团契，而我们的团契是与父和他儿子耶稣基督所共有的。
1JOHN|1|4|我们把这些事写给你们，使我们 的喜乐得以满足。
1JOHN|1|5|上帝就是光，在他毫无黑暗；这是我们从主所听见，又报给你们的信息。
1JOHN|1|6|我们若说，我们与上帝有团契，却仍在黑暗里行走，就是说谎话，不实行真理了。
1JOHN|1|7|我们若在光明中行走，如同上帝在光明中，就彼此有团契，他儿子耶稣的血就洗净我们一切的罪。
1JOHN|1|8|我们若说自己没有罪，就是欺骗自己，真理就不在我们里面了。
1JOHN|1|9|我们若认自己的罪，上帝是信实的，是公义的，必要赦免我们的罪，洗净我们一切的不义。
1JOHN|1|10|我们若说自己没有犯过罪，就是把上帝当作说谎的，他的道就不在我们里面了。
1JOHN|2|1|我的孩子们哪，我把这些话写给你们，是要你们不犯罪。若有人犯罪，在父那里我们有一位中保，就是那义者耶稣基督。
1JOHN|2|2|他为我们的罪作了赎罪祭，不单是为我们的罪，也是为普天下人的罪。
1JOHN|2|3|我们若遵守上帝的命令，就知道我们确实认识他。
1JOHN|2|4|人若说“我认识他”，却不遵守他的命令，就是说谎话的，真理就不在他里面了。
1JOHN|2|5|凡遵守他的道的，爱上帝的心确实地在他里面达到完全了。由此我们知道我们是在他里面。
1JOHN|2|6|凡说自己住在他里面的，就该照着他所行的去行。
1JOHN|2|7|亲爱的，我写给你们的不是一条新命令，而是你们从起初所受的旧命令；这旧命令就是你们所听过的道。
1JOHN|2|8|然而，我写给你们的是一条新命令，在基督里是真实的，在你们也是真实的，因为黑暗渐渐消逝，真光已经在照耀。
1JOHN|2|9|人若说自己在光明中，却恨他的弟兄，他到如今还是在黑暗里。
1JOHN|2|10|那爱弟兄的，就是住在光明中，他不会使人失足犯罪 。
1JOHN|2|11|惟独那恨弟兄的，是在黑暗里，也在黑暗里行走，不知道往哪里去，因为黑暗使他的眼睛瞎了。
1JOHN|2|12|孩子们哪，我写信给你们， 因为你们的罪藉着基督的名得了赦免。
1JOHN|2|13|父老们啊，我写信给你们， 因为你们认识从起初就有的那一位。 青年们哪，我写信给你们， 因为你们胜过了那恶者。
1JOHN|2|14|孩子们哪，我曾写信给你们， 因为你们认识父。 父老们啊，我曾写信给你们， 因为你们认识从起初就有的那一位。 青年们哪，我曾写信给你们， 因为你们刚强， 上帝的道常存在你们心里， 你们也胜过了那恶者。
1JOHN|2|15|不要爱世界和世界上的东西，若有人爱世界，爱父的心就不在他里面了。
1JOHN|2|16|因为凡世界上的东西，好比肉体的情欲、眼目的情欲和今生的骄傲，都不是从父来的，而是从世界来的。
1JOHN|2|17|这世界和世上的情欲都要消逝，惟独那遵行上帝旨意的人永远常存。
1JOHN|2|18|孩子们哪，如今是末世的时光了。你们曾听过那敌基督者要来，现在有好些敌基督者已经出来了；由此我们就知道，如今是末世的时光了。
1JOHN|2|19|他们从我们中间出去，却不是属我们的，若是属我们的，就必仍旧与我们同在。他们出去，这就显明他们都不是属我们的。
1JOHN|2|20|你们从那圣者受了恩膏，并且你们大家都知道 。
1JOHN|2|21|我写信给你们，不是因你们不认识真理，而是因你们认识，并且知道一切虚谎都不是从真理出来的。
1JOHN|2|22|谁是说谎话的呢？不就是那不认耶稣为基督的吗？那不认父与子的，这个人就是敌基督的。
1JOHN|2|23|凡不认子的，就没有父；宣认子的，连父也有了。
1JOHN|2|24|论到你们，务要将那从起初所听见的常存在心里；若将从起初所听见的存在心里，你们就会住在子里面，也会住在父里面。
1JOHN|2|25|基督所应许我们的就是永生。
1JOHN|2|26|我将这些话写给你们，是论到那些迷惑你们的人说的。
1JOHN|2|27|至于你们，你们从基督所受的恩膏常存在你们心里，并不用人教导你们，自有他的恩膏在凡事上教导你们。这恩膏是真的，不是假的，你们要按这恩膏的教导住在他里面。
1JOHN|2|28|孩子们哪，你们要住在基督里面。这样，他若显现，我们就可以坦然无惧；当他来临的时候，在他面前不至于惭愧。
1JOHN|2|29|你们若知道他是公义的，就知道凡行公义的人都是他所生的。
1JOHN|3|1|你们看父赐给我们的是何等的慈爱，让我们得以称为上帝的儿女；我们也真是他的儿女。世人不认识我们 的理由，是因他们未曾认识父。
1JOHN|3|2|亲爱的，我们现在是上帝的儿女，将来如何还未显明。我们所知道的是：基督显现的时候，我们会像他，因为我们将见到他的本相。
1JOHN|3|3|凡对他有这指望的，就洁净自己，像他是洁净的一样。
1JOHN|3|4|凡犯罪的，就是做违背律法的事；违背律法就是罪。
1JOHN|3|5|你们知道，基督曾显现是要除掉罪 ；在他并没有罪。
1JOHN|3|6|凡住在他里面的，不犯罪；凡犯罪的，未曾看见他，也未曾认识他。
1JOHN|3|7|孩子们哪，不要让人迷惑了你们；行义的才是义人，正如基督是义的。
1JOHN|3|8|犯罪的是出于魔鬼，因为魔鬼从起初就犯罪。上帝的儿子显现出来，是为了要毁灭魔鬼的作为。
1JOHN|3|9|凡从上帝生的，不犯罪，因上帝的道 存在他里面，他也不能犯罪，因为他是由上帝所生的。
1JOHN|3|10|这就显明谁是上帝的儿女，谁是魔鬼的儿女了。凡不行义的，不是出于上帝，不爱他弟兄的，也是如此。
1JOHN|3|11|我们要彼此相爱。这就是你们从起初所听到的信息。
1JOHN|3|12|不要像 该隐 ；他是属那邪恶者，杀了自己的弟弟。为什么杀了他呢？因为自己的行为是邪恶的，而弟弟的行为是正直的。
1JOHN|3|13|弟兄们，世人若恨你们，不要惊讶。
1JOHN|3|14|我们知道，我们已经出死入生了，因为我们爱弟兄。没有爱心的，仍住在死中。
1JOHN|3|15|凡恨自己弟兄的，就是杀人的；你们知道，凡杀人的，没有永生住在他里面。
1JOHN|3|16|基督为我们舍命，我们从此就知道何为爱；我们也当为弟兄舍命。
1JOHN|3|17|凡有世上财物的，看见弟兄缺乏，却关闭了恻隐的心，上帝的爱怎能住在他里面呢？
1JOHN|3|18|孩子们哪，我们相爱，不要只在言语或舌头上，总要以行为和真诚表现出来。
1JOHN|3|19|从这一点，我们会知道，我们是出于真理的，并且我们在上帝面前可以安心，
1JOHN|3|20|即使我们的心责备自己，上帝比我们的心大，他知道一切。
1JOHN|3|21|亲爱的，我们的心若不责备我们，在上帝面前就可以坦然无惧了。
1JOHN|3|22|我们一切所求的，就从他得着，因为我们遵守他的命令，行他所喜悦的事。
1JOHN|3|23|上帝的命令就是：我们要信他儿子耶稣基督的名，并且照他所赐给我们的命令彼此相爱。
1JOHN|3|24|遵守上帝命令的，住在上帝里面，而上帝也住在他里面。从这一点，我们知道上帝住在我们里面，这是由于他所赐给我们的圣灵。
1JOHN|4|1|亲爱的，一切的灵不可都信，总要察验那些灵是否出于上帝，因为有许多假先知已经来到世上。
1JOHN|4|2|凡宣认耶稣基督是成了肉身而来的灵就是出于上帝的，由此你们可以认出上帝的灵来；
1JOHN|4|3|凡不宣认耶稣的灵，不是出于上帝。这是那敌基督者的灵；你们从前听见他要来，现在他已经在世上了。
1JOHN|4|4|孩子们哪，你们是属上帝的，并且胜过了假先知，因为那在你们里面的比那在世界上的更大。
1JOHN|4|5|他们是属世界的，所以讲论世界的事，而世人也听从他们。
1JOHN|4|6|我们是属上帝的，认识上帝的就听从我们；不属上帝的就不听从我们。从此我们可以认出真理的灵和错谬的灵来。
1JOHN|4|7|亲爱的，我们要彼此相爱，因为爱是从上帝来的。凡有爱的都是由上帝而生，并且认识上帝。
1JOHN|4|8|没有爱的就不认识上帝，因为上帝就是爱。
1JOHN|4|9|上帝差他独一的儿子到世上来，使我们藉着他得生命；由此，上帝对我们的爱就显明了。
1JOHN|4|10|不是我们爱上帝，而是上帝爱我们，差他的儿子为我们的罪作了赎罪祭；这就是爱。
1JOHN|4|11|亲爱的，既然上帝这样爱我们，我们也要彼此相爱。
1JOHN|4|12|从来没有人见过上帝，我们若彼此相爱，上帝就住在我们里面，他的爱在我们里面得以完满了。
1JOHN|4|13|因为上帝将他的灵赐给我们，由此我们知道我们是住在他里面，而他也住在我们里面。
1JOHN|4|14|父差子作世人的救主，这是我们所看见并且作见证的。
1JOHN|4|15|凡宣认耶稣为上帝儿子的，上帝就住在他里面，而他也住在上帝里面。
1JOHN|4|16|我们知道并且深信上帝是爱我们的。 上帝就是爱，住在爱里面的就是住在上帝里面；上帝也住在他里面。
1JOHN|4|17|由此，爱在我们里面得以完满：我们可以在审判的日子坦然无惧，因为基督如何，我们在这世上也如何。
1JOHN|4|18|在爱里没有惧怕；完满的爱把惧怕驱逐出去，因为惧怕里含着惩罚，惧怕的人在爱里尚未得到完满。
1JOHN|4|19|我们爱，因为上帝先爱我们。
1JOHN|4|20|人若说“我爱上帝”，却恨他的弟兄，就是说谎了；不爱他看得见的弟兄，就不能爱看不见的上帝 。
1JOHN|4|21|爱上帝的，也要爱弟兄；这是我们从上帝所受的命令。
1JOHN|5|1|凡信耶稣是基督的，都是从上帝生的；凡爱生他之上帝的，也必爱从上帝生的 。
1JOHN|5|2|我们爱上帝，又实行 他的命令，由此就知道我们爱上帝的儿女了。
1JOHN|5|3|我们遵守上帝的命令，这就是爱他了，而且他的命令并不是难守的。
1JOHN|5|4|因为凡从上帝生的就胜过世界；使我们胜过世界的就是我们的信心。
1JOHN|5|5|胜过世界的是谁呢？不就是那信耶稣是上帝儿子的吗？
1JOHN|5|6|这藉着水和血而来的，就是耶稣基督，不是单用水，而是用水又用血，并且有圣灵作见证，因为圣灵就是真理。
1JOHN|5|7|作见证的有三：
1JOHN|5|8|就是圣灵、水与血，这三样也都是一致的。
1JOHN|5|9|既然我们领受人的见证，上帝的见证更该领受 了，因为上帝的见证是为他儿子作的。
1JOHN|5|10|信上帝儿子的，就有这见证在他心里；不信上帝的，就是把上帝当作说谎的，因为不信上帝为他儿子作的见证。
1JOHN|5|11|这见证就是：上帝赐给我们永生，而这永生是在他儿子里面的。
1JOHN|5|12|那有上帝儿子的，就有生命；没有上帝儿子的，就没有生命。
1JOHN|5|13|我把这些话写给你们信奉上帝儿子之名的人，要让你们知道自己有永生。
1JOHN|5|14|我们若照着上帝的旨意祈求，他就垂听我们；这就是我们对他所存坦然无惧的心。
1JOHN|5|15|既然我们知道他听我们一切所求的，就知道我们所求于他的，无不得着。
1JOHN|5|16|人若看见弟兄犯了不至于死的罪，就要为他祈求，上帝必将生命赐给他—有些人犯的罪是不至于死的；有的是至于死的罪，我不是说要为这罪祈求。
1JOHN|5|17|一切不义的事都是罪，但也有不至于死的罪。
1JOHN|5|18|我们知道，凡从上帝生的，必不犯罪；从上帝生的那一位，必保守他，那邪恶者无法加害于他。
1JOHN|5|19|我们知道，我们是属上帝的，而全世界都伏在那邪恶者的权势之下。
1JOHN|5|20|我们知道，上帝的儿子已经来到，并且将悟性赐给我们，使我们认识那位真实者，我们也在那位真实者里面，就是在他儿子耶稣基督里面。这是真神，也是永生。
1JOHN|5|21|孩子们哪，你们要远避偶像。
2JOHN|1|1|我作长老的写信给蒙拣选的夫人 和她的儿女，就是我真心所爱的；不但我爱，也是一切认识真理的人所爱的，
2JOHN|1|2|这是因为真理住在我们里面，也必与我们同在直到永远。
2JOHN|1|3|愿恩惠、怜悯、平安 从父上帝和他儿子耶稣基督，在真理和爱中必与我们同在。
2JOHN|1|4|我非常欢喜见你的儿女，有照我们从父所受之命令遵行真理的。
2JOHN|1|5|夫人哪，我现在请求你，我们大家要彼此相爱。我写给你的，并不是一条新命令，而是我们从起初就有的。
2JOHN|1|6|这就是爱，就是照他的命令行事；这就是命令，你们要照这命令行，正如你们从起初所听见的。
2JOHN|1|7|有许多迷惑人的已经来到世上，他们不宣认耶稣基督是成了肉身来的；这样的人是迷惑人的，是敌基督的。
2JOHN|1|8|你们要小心，不要失去你们 所完成的工作，而要得到充足的赏赐。
2JOHN|1|9|凡越过基督的教导而不持守的，就没有上帝；凡持守这教导的，就有父又有子。
2JOHN|1|10|若有人到你们那里而不传这教导，不要接他到家里，也不要向他问安；
2JOHN|1|11|因为向他问安的，就在他的恶行上有份。
2JOHN|1|12|我还有许多事要写给你们，却不愿意用纸用墨，但盼望到你们那里，与你们面对面谈论，使我们的喜乐得以满足。
2JOHN|1|13|你那蒙拣选的姊妹的儿女向你问安。
3JOHN|1|1|我作长老的写信给亲爱的 该犹 ，就是我真心所爱的。
3JOHN|1|2|亲爱的，我愿你事事安宁，身体健康，正如你的心神安宁一样。
3JOHN|1|3|我非常欢喜，有弟兄到这里来，证实你对真理的忠诚，就是你按着真理而行。
3JOHN|1|4|我听见我的儿女按真理而行，我的欢喜没有比这个更大的。
3JOHN|1|5|亲爱的，你对弟兄，特别是对作客旅的弟兄所做的都是忠诚的。
3JOHN|1|6|他们在教会面前证实了你的爱；你若以对得起上帝的方式，为他们送行就好了；
3JOHN|1|7|因为他们是为基督的名 出外，并没有从未信的人接受什么。
3JOHN|1|8|所以，我们应当接待这样的人，好让我们与他们在真理上成为同工。
3JOHN|1|9|我曾写过一些东西给教会，但他们中间那好作领袖的 丢特腓 不接纳我们。
3JOHN|1|10|为此，我若去，要提起他所做的事，就是他用恶言攻击我们，还不满足，他自己不接纳弟兄，有人愿意接纳，他还阻止，并且把接纳弟兄的人赶出教会。
3JOHN|1|11|亲爱的，不要效法恶，只要效法善。行善的人属乎上帝；行恶的人未曾见过上帝。
3JOHN|1|12|低米丢 行善，有众人给他作见证，又有真理给他作见证，就是我们也给他作见证，你知道我们的见证是真的。
3JOHN|1|13|我还有许多事要写给你，却不愿意用笔墨来写给你，
3JOHN|1|14|但盼望很快见到你，我们好面对面谈论。
3JOHN|1|15|愿你平安！朋友们都向你问安。请你替我按著名字一一向朋友们问安。
JUDE|1|1|耶稣基督的仆人、 雅各 的兄弟 犹大 ，写信给那些被召、在父上帝里蒙爱、为耶稣基督保守的人。
JUDE|1|2|愿怜悯、平安 、慈爱多多加给你们！
JUDE|1|3|亲爱的，我一直很迫切地想要写信给你们，论到我们同享的救恩，但我觉得有必要现在就写信劝你们，要为从前一次交付给圣徒的真道竭力奋斗。
JUDE|1|4|因为有些人偷偷地进来，就是早就被判定受惩罚的不虔诚的人，他们把我们上帝的恩典变为放纵情欲的机会，并且不认独一的主宰—我们的主耶稣基督。
JUDE|1|5|这一切的事，你们虽然知道，我却仍要提醒你们：从前主 只一次就 救了他的百姓出 埃及 地，后来却把那些不信的灭绝了。
JUDE|1|6|至于那些不守本位、离开自己住处的天使，主用锁链把他们永远拘留在黑暗里，等候大日子的审判。
JUDE|1|7|同样， 所多玛 、 蛾摩拉 和周围城镇的人也跟着他们一样犯淫乱，随从逆性的情欲，以致遭受永不熄灭之火的惩罚，作为众人的鉴戒。
JUDE|1|8|照样，这些做梦的人也污秽身体，轻慢掌权者，毁谤众尊荣者。
JUDE|1|9|天使长 米迦勒 为 摩西 的尸首与魔鬼争辩的时候，尚且不敢用毁谤的话谴责他，只说：“主责备你吧！”
JUDE|1|10|但这些人毁谤他们所不知道的。他们与那些没有理性的牲畜一样，只做本性所知道的事，败坏了自己。
JUDE|1|11|他们有祸了！因为他们走 该隐 的道路，又为财利往 巴兰 的错谬里直奔，并在 可拉 的背叛中灭亡了。
JUDE|1|12|这样的人是你们爱筵上的污点 ；他们无所惧怕地同你们宴乐，仿佛牧人只顾喂饱自己。他们是无雨的浮云，被风飘荡；是秋天没有果子的树，死而又死，连根被拔出来；
JUDE|1|13|是海里的狂浪，涌出自己可耻的沫子来；是流荡的星，有漆黑的幽暗永远为他们保留着。
JUDE|1|14|亚当 的七世孙 以诺 曾预言这些人说：“看哪，主带着他的千万圣者来临，
JUDE|1|15|要审判众人，证实一切不敬虔的人所妄行一切不敬虔的事，又证实不敬虔的罪人所说顶撞他的刚愎的话。”
JUDE|1|16|这些人喜出怨言，责怪他人，随从自己的情欲而行，口说夸大的话，为自己的利益谄媚人。
JUDE|1|17|亲爱的，至于你们，要记得我们主耶稣基督的使徒从前所说的话。
JUDE|1|18|他们曾对你们说过，末世必有好嘲弄的人随从自己不敬虔的私欲而行。
JUDE|1|19|这就是那些好结党分派、属乎血气、没有圣灵的人。
JUDE|1|20|亲爱的，至于你们，要在至圣的真道上造就自己，藉着圣灵祷告，
JUDE|1|21|保守自己常在上帝的爱中，仰望我们主耶稣基督的怜悯，进入永生。
JUDE|1|22|有些人心中犹疑 ，你们要怜悯 他们；
JUDE|1|23|有些人你们要从火中抢出来，搭救他们 ；有些人你们要存惧怕的心怜悯他们，连那被情欲污染的衣服也要厌恶。
JUDE|1|24|愿那能保守你们不失脚，使你们无瑕无疵、欢欢喜喜站在他荣耀之前的、
JUDE|1|25|我们的救主独一的上帝，藉着我们的主耶稣基督，得享荣耀、威严、能力、权柄，从万古以前，到现今，直到永永远远。阿们！
REV|1|1|耶稣基督的启示，就是上帝赐给他，要他将必须快要发生的事指示他的众仆人。他差遣使者指明给他的仆人 约翰 ，
REV|1|2|约翰 就将上帝的道和耶稣基督的见证，凡自己所看见的，都见证出来。
REV|1|3|诵读这书上预言的，和那些听见又遵守其中所记载的，都是有福的，因为时候近了。
REV|1|4|约翰 写信给 亚细亚 的七个教会。愿那位今在、昔在、以后永在的上帝，与他宝座前的七灵，和那忠信的见证者、从死人中复活的首生者 、世上君王的元首耶稣基督，赐恩惠和平安 给你们。 他爱我们，用自己的血使我们从罪中得释放 ，
REV|1|5|
REV|1|6|又使我们成为国度，作他父上帝的祭司。愿荣耀、权能归给他，直到永永远远 。阿们！
REV|1|7|“看哪，他驾云降临； 众目都要看见他， 连刺他的人也要看见他； 地上的万族要因他哀哭。” 这是真实的。阿们！
REV|1|8|主上帝说：“我是阿拉法，我是俄梅戛 ，是今在、昔在、以后永在的全能者。”
REV|1|9|我— 约翰 就是你们的弟兄，在耶稣里和你们一同在患难、国度、忍耐里有份的，为上帝的道，并为给耶稣作的见证，曾在那名叫 拔摩 的海岛上。
REV|1|10|有一主日我被圣灵感动，听见在我后面有大声音如吹号，
REV|1|11|说：“把你所看见的写在书上，寄给 以弗所 、 士每拿 、 别迦摩 、 推雅推喇 、 撒狄 、 非拉铁非 、 老底嘉 那七个教会。”
REV|1|12|我转过身来要看看是谁的声音在跟我说话。我一转过来，看见了七个金灯台；
REV|1|13|在灯台中间有一位好像人子的，身穿垂到脚的长袍，胸间束着金带。
REV|1|14|他的头与发皆白，如白羊毛，如雪；他的眼睛好像火焰，
REV|1|15|双脚好像在炉中锻鍊得发亮的铜，声音好像众水的声音。
REV|1|16|他右手拿着七颗星，从他口中吐出一把两刃的利剑，面貌好像烈日放光。
REV|1|17|我看见了他，就仆倒在他脚前，像死人一样。他用右手按着我说：“不要怕。我是首先的，是末后的，
REV|1|18|又是永活的。我曾死过，看哪，我是活着的，直到永永远远；并且我拿着死亡和阴间的钥匙。
REV|1|19|所以，你要把所看见的事、现在的事和以后将发生的事，都写下来。
REV|1|20|至于你所看见、在我右手中的七颗星和那七个金灯台的奥秘就是：七颗星是七个教会的使者，七个灯台是七个教会。”
REV|2|1|“你要写信给 以弗所 教会的使者，说：‘那右手拿着七颗星，在七个金灯台中间行走的这样说：
REV|2|2|我知道你的行为、劳碌、忍耐，也知道你不容忍恶人。你也曾察验那自称为使徒却不是使徒的，看出他们是假的。
REV|2|3|你能忍耐，曾为我的名劳苦而不困倦。
REV|2|4|然而，有一件事我要责备你，就是你把起初的爱心抛弃了。
REV|2|5|所以你要回想你是从哪里坠落的，并且要悔改，做起初所做的工作。你若不悔改，我要到你那里去，把你的灯台从原处挪去。
REV|2|6|然而你还有一件可取的事，就是你恨恶 尼哥拉 派的行为，这种行为也是我所恨恶的。
REV|2|7|凡有耳朵的都应当听圣灵向众教会所说的话。得胜的，我必将上帝乐园中生命树的果子赐给他吃。’”
REV|2|8|“你要写信给 士每拿 教会的使者，说：‘那首先的、末后的，死过又活了的这样说：
REV|2|9|我知道你的患难和贫穷—其实你却是富足的，也知道那自称是 犹太 人的所说毁谤的话，其实他们不是 犹太 人，而是撒但会堂的人。
REV|2|10|你将要受的苦，你不用怕。看哪！魔鬼要把你们中间几个人下在监里，使你们受考验，你们要遭受苦难十日。你务要至死忠心，我就赐给你那生命的冠冕。
REV|2|11|凡有耳朵的都应当听圣灵向众教会所说的话。得胜的必不受第二次死的害。’”
REV|2|12|“你要写信给 别迦摩 教会的使者，说：‘那有两刃利剑的这样说：
REV|2|13|我知道你的居所，就是有撒但座位之处；当我忠心的见证人 安提帕 在你们中间，在撒但所住的地方被杀之时，你还坚守我的名，没有否认对我的信仰。
REV|2|14|然而，有几件事我要责备你，就是在你那里有人服从了 巴兰 的教训；这 巴兰 曾教唆 巴勒 将绊脚石放在 以色列 人面前，使他们吃祭过偶像之物，并且犯淫乱。
REV|2|15|同样，你那里也有人服从了 尼哥拉 派的教训。
REV|2|16|所以，你当悔改；若不悔改，我很快就到你那里来，用我口中的剑攻击他们。
REV|2|17|凡有耳朵的都应当听圣灵向众教会所说的话。得胜的，我必将那隐藏的吗哪赐给他，并赐他一块白石，石上写着新的名字，除了那领受的以外，没有人认识。’”
REV|2|18|“你要写信给 推雅推喇 教会的使者，说：‘上帝的儿子，那位眼睛如火焰、双脚像发亮的铜的这样说：
REV|2|19|我知道你的行为：爱心、信心、勤劳、忍耐；又知道你末后所行的善事比起初所行的更多。
REV|2|20|然而，有一件事我要责备你，就是你容忍那自称是先知的妇人 耶洗别 教唆我的仆人，引诱他们犯淫乱，吃祭过偶像之物。
REV|2|21|我曾给她悔改的机会，她却不肯悔改她的淫行。
REV|2|22|看吧，我要使她病倒在床上。那些与她犯奸淫的人若不悔改他们的行为，我也要使他们同受大患难。
REV|2|23|我又要杀死她的儿女，众教会就知道，我是那察看人肺腑心肠的，我要照你们的行为报应各人。
REV|2|24|至于你们其余的 推雅推喇 人，就是一切不随从这教训，不明白他们所谓撒但深奥之理的人，我告诉你们，我不会再把别的担子放在你们身上。
REV|2|25|你们只要持守那已经有的，直到我来。
REV|2|26|那得胜又遵守我命令到底的， 我要赐给他权柄制伏列国；
REV|2|27|他必用铁杖管辖他们， 如同打碎陶器，
REV|2|28|像我也从我父领受了权柄一样。我又要把晨星赐给他。
REV|2|29|凡有耳朵的都应当听圣灵向众教会所说的话。’”
REV|3|1|“你要写信给 撒狄 教会的使者，说：‘那有上帝的七灵和七颗星的这样说：我知道你的行为，就是名义上你是活的，实际上你是死的。
REV|3|2|你要警醒，坚固那些剩下、快要死的，因为我发现你的行为，在我上帝面前没有一样是完全的。
REV|3|3|所以，要记得你所领受和听见的；要遵守，并要悔改。你若不警醒，我必如贼一样来到；我几时来到你那里，你绝不会知道。
REV|3|4|然而，在 撒狄 你还有几位是未曾污秽自己衣服的，他们会穿白衣与我同行，因为他们是配穿的。
REV|3|5|得胜的必这样穿白衣，我也不从生命册上涂去他的名；我要在我父面前，和我父的众使者面前，宣认他的名。
REV|3|6|凡有耳朵的都应当听圣灵向众教会所说的话。’”
REV|3|7|“你要写信给 非拉铁非 教会的使者，说： ‘那神圣、真实的， 拿着 大卫 的钥匙， 开了就没有人能关， 关了就没有人能开的这样说：
REV|3|8|我知道你的行为。看哪，我在你面前给你一个敞开的门，是没有人能关的。我知道你有一点力量，也遵守我的道，没有否认我的名。
REV|3|9|那属撒但会堂的，自称是 犹太 人，其实不是 犹太 人，而是说谎话的，我要使他们来到你脚前下拜，使他们知道我已经爱你了。
REV|3|10|因为你遵守了我坚忍的道，我也必在普天下人受试炼的时候保守你免受试炼。
REV|3|11|我必快来，你要持守你所有的，免得人夺去你的冠冕。
REV|3|12|得胜的，我要使他在我上帝的殿中作柱子，他必不再从那里出去。我又要把我上帝的名和我上帝城的名—从天上我上帝那里降下来的新 耶路撒冷 ，和我的新名，都写在他上面。
REV|3|13|凡有耳朵的都应当听圣灵向众教会所说的话。’”
REV|3|14|“你要写信给 老底嘉 教会的使者，说：‘那位阿们、诚信真实的见证者、上帝创造的根源这样说：
REV|3|15|我知道你的行为，你也不冷也不热；我巴不得你或冷或热。
REV|3|16|既然你如温水，也不冷也不热，我要从我口中把你吐出去。
REV|3|17|你说：我是富足的，已经发了财，一样都不缺，却不知道你是困苦、可怜、贫穷、瞎眼、赤身的。
REV|3|18|我劝你向我买从火中锻鍊出来的金子，使你富足；又买白衣穿上，使你赤身的羞耻不露出来；又买眼药抹你的眼睛，使你能看见。
REV|3|19|凡我所疼爱的，我就责备管教。所以，你要发热心，也要悔改。
REV|3|20|看哪，我站在门外叩门，若有听见我声音而开门的，我要进到他那里去，我与他，他与我一起吃饭。
REV|3|21|得胜的，我要赐他在我宝座上与我同坐，就如我得了胜，在我父的宝座上与他同坐一般。
REV|3|22|凡有耳朵的都应当听圣灵向众教会所说的话。’”
REV|4|1|这些事以后，我观看，看见天上有一道门开着。我头一次听见的那好像吹号的声音对我说：“你上这里来，我要把此后必须发生的事指示你。”
REV|4|2|我立刻被圣灵感动，见有一个宝座安置在天上，有一位坐在宝座上。
REV|4|3|那坐着的，看来好像碧玉和红宝石；又有彩虹围着宝座，光彩好像绿宝石。
REV|4|4|宝座的周围又有二十四个座位，上面坐着二十四位长老，身穿白衣，头上戴着金冠冕。
REV|4|5|有闪电、声音、雷轰从宝座中发出。在宝座前点着七支火炬，就是上帝的七灵。
REV|4|6|宝座前有一个如同水晶的玻璃海。 宝座的周围，四边有四个活物，遍体前后都长满了眼睛。
REV|4|7|第一个活物像狮子，第二个像牛犊，第三个的脸像人脸，第四个像飞鹰。
REV|4|8|四个活物各有六个翅膀，遍体内外都长满了眼睛。他们昼夜不住地说： “圣哉！圣哉！圣哉！ 主—全能的上帝； 昔在、今在、以后永在！”
REV|4|9|每逢四活物将荣耀、尊贵、感谢归给那坐在宝座上、活到永永远远者的时候，
REV|4|10|二十四位长老就俯伏敬拜坐在宝座上活到永永远远的那一位，又把他们的冠冕放在宝座前，说：
REV|4|11|“我们的主，我们的上帝， 你配得荣耀、尊贵、权柄， 因为你创造了万物， 万物因你的旨意被创造而存在。”
REV|5|1|我看见坐在宝座那位的右手中有书卷，正反面都写着字，用七个印密封着。
REV|5|2|我又看见一位大力的天使大声宣告说：“有谁配展开那书卷，揭开那七个印呢？”
REV|5|3|在天上、地上、地底下，没有人能展开、能阅览那书卷。
REV|5|4|因为没有人配展开、阅览那书卷，我就大哭。
REV|5|5|长老中有一位对我说：“不要哭。看哪， 犹大 支派中的狮子， 大卫 的根，他已得胜，能展开那书卷，揭开那七个印。”
REV|5|6|我又看见宝座和四个活物，以及长老之中有羔羊站着，像是被杀的，有七个角七只眼睛，就是上帝的七 灵，奉差遣往普天下去的。
REV|5|7|这羔羊前来，从坐在宝座上那位的右手中拿了书卷。
REV|5|8|他一拿了书卷，四活物和二十四位长老就俯伏在羔羊面前，各拿着琴和盛满了香的金炉；这香就是众圣徒的祈祷。
REV|5|9|他们唱新歌，说： “你配拿书卷， 配揭开它的七印； 因为你曾被杀，用自己的血 从各支派、各语言、各民族、各邦国中买了人来，使他们归于上帝，
REV|5|10|又使他们成为国民和祭司，归于我们的上帝； 他们将在地上执掌王权。”
REV|5|11|我又观看，我听见宝座和活物及长老的周围有许多天使的声音；他们的数目有千千万万，
REV|5|12|大声说： “被杀的羔羊配得 权能、丰富、智慧、力量、 尊贵、荣耀、颂赞。
REV|5|13|我又听见在天上、地上、地底下、沧海里和天地间一切所有被造之物，都说： “愿颂赞、尊贵、荣耀、权势， 都归给坐在宝座上的那位和羔羊， 直到永永远远！”
REV|5|14|四活物就说：“阿们！”众长老也俯伏敬拜。
REV|6|1|我看见羔羊揭开七个印中第一个印的时候，听见四活物中的一个活物，声音如雷，说：“你来！”
REV|6|2|我就观看，看见一匹白马，骑在马上的拿着弓，并有冠冕赐给他。他出来征服，胜而又胜。
REV|6|3|羔羊揭开第二个印的时候，我听见第二个活物说：“你来！”
REV|6|4|就另有一匹马出来，是红色的；有权柄赐给了那骑马的，要从地上夺去太平，使人彼此相杀；他又接受了一把大刀。
REV|6|5|羔羊揭开第三个印的时候，我听见第三个活物说：“你来！”我就观看，看见一匹黑马；骑在马上的，手里拿着天平。
REV|6|6|我听见在四个活物中似乎有声音说：“一个银币买一升麦子，一个银币买三升大麦；油和酒不可糟蹋。”
REV|6|7|羔羊揭开第四个印的时候，我听见第四个活物说：“你来！”
REV|6|8|我就观看，看见一匹灰色马；骑在马上的，名字叫作“死”，阴间也随着他；有权柄赐给他们，可以用刀剑、饥荒、瘟疫、野兽，杀害地上四分之一的人。
REV|6|9|羔羊揭开第五个印的时候，我看见在祭坛底下有曾为上帝的道，并为作见证而被杀的人的灵魂，
REV|6|10|大声喊着说：“神圣真实的主宰啊，你不审判住在地上的人，为我们所流的血伸冤，要到几时呢？”
REV|6|11|于是有白袍赐给他们各人；又有话吩咐他们还要歇息片刻，等到与他们同作仆人的，和他们的弟兄，像他们一样被杀的人的数目凑足的时候。
REV|6|12|羔羊揭开第六个印的时候，我看见地大震动，太阳变黑像粗麻布，整个月亮变红像血，
REV|6|13|天上的星辰坠落在地上，如同无花果树被大风摇动，落下未熟的果子一样。
REV|6|14|天就裂开，好像书卷被卷起来；山岭海岛都被移动离开原位。
REV|6|15|地上的君王、臣宰、将军、富户、壮士，和一切为奴的、自主的，都藏在山洞和岩石穴里，
REV|6|16|向山和岩石说：“倒在我们身上吧！把我们藏起来，躲避坐宝座者的脸面和羔羊的愤怒；
REV|6|17|因为他们遭愤怒的大日子到了，谁能站得住呢？”
REV|7|1|此后，我看见四位天使站在地的四角，执掌地上四方的风，使风不吹在地上、海上和各种树上。
REV|7|2|我又看见另有一位天使从日出之地上来，拿着永生上帝的印。他向那得到权柄能伤害地和海的四位天使大声喊着，
REV|7|3|说：“你们不可伤害地、海和树林，等我们在我们上帝众仆人的额上盖了印。”
REV|7|4|我听见 以色列 人各支派中受印的数目有十四万四千；
REV|7|5|犹大 支派中受印的有一万二千； 吕便 支派中有一万二千； 迦得 支派中有一万二千；
REV|7|6|亚设 支派中有一万二千； 拿弗他利 支派中有一万二千； 玛拿西 支派中有一万二千；
REV|7|7|西缅 支派中有一万二千； 利未 支派中有一万二千； 以萨迦 支派中有一万二千；
REV|7|8|西布伦 支派中有一万二千； 约瑟 支派中有一万二千； 便雅悯 支派中受印的有一万二千。
REV|7|9|此后，我观看，看见有许多人，没有人能计算，是从各邦国、各支派、各民族、各语言来的，站在宝座和羔羊面前，身穿白衣，手拿棕树枝，
REV|7|10|大声喊着说： “愿救恩归于坐在宝座上我们的上帝， 也归于羔羊！”
REV|7|11|众天使都站在宝座和众长老，以及四个活物的周围，俯伏在宝座前，敬拜上帝，
REV|7|12|说： “阿们！颂赞、荣耀、智慧、 感谢、尊贵、权能、 力量都归于我们的上帝， 直到永永远远。阿们！”
REV|7|13|长老中有一位回应我说：“这些穿白衣的是谁？是从哪里来的？”
REV|7|14|我对他说：“我主啊，你是知道的。”他向我说：“这些人是从大患难中出来的，他们曾用羔羊的血把衣裳洗得洁白。
REV|7|15|所以，他们在上帝宝座前， 昼夜在他殿中事奉他； 那坐在宝座上的要用帐幕覆庇他们。
REV|7|16|他们不再饥，不再渴； 太阳必不伤害他们， 任何炎热也不伤害他们，
REV|7|17|因为宝座中的羔羊必牧养他们， 领他们到生命水的泉源； 上帝必擦去他们一切的眼泪。”
REV|8|1|羔羊揭开第七个印的时候，天上寂静约有半小时。
REV|8|2|我看见那站在上帝面前的七位天使，有七枝号赐给他们。
REV|8|3|另有一位天使拿着金香炉来，站在祭坛旁边；有许多香赐给他，要和众圣徒的祈祷一同献在宝座前的金坛上。
REV|8|4|那香的烟和众圣徒的祈祷从天使的手中一同升到上帝面前。
REV|8|5|天使拿着香炉，盛满了坛上的火，倒在地上；就有雷轰、响声、闪电、地震。
REV|8|6|拿着七枝号筒的七位天使预备好要吹号。
REV|8|7|第一位天使吹号，就有冰雹和火搀着血扔在地上；地的三分之一和树的三分之一被烧掉了，一切的青草也被烧掉了。
REV|8|8|第二位天使吹号，就有像火烧着的大山扔在海中；海的三分之一变成血，
REV|8|9|海中有生命的被造之物死了三分之一，船只也毁坏了三分之一。
REV|8|10|第三位天使吹号，就有烧着的大星好像火把从天上坠下来，落在江河的三分之一和众水的泉源上。
REV|8|11|这星名叫“苦艾”；众水的三分之一变为苦艾，许多人因水变苦而死了。
REV|8|12|第四位天使吹号，太阳的三分之一、月亮的三分之一、星辰的三分之一都被击打，以致日月星的三分之一变黑了，白昼的三分之一没有光，黑夜也是这样。
REV|8|13|我观看，听见一只在空中飞的鹰大声说：“祸哉！祸哉！祸哉！地上的居民哪，其余的三位天使快要吹号了！”
REV|9|1|第五位天使吹号，我就看见一颗星从天上坠落到地上；有无底坑的钥匙赐给它。
REV|9|2|它开了无底坑，就有烟从坑里往上冒，好像大火炉的烟；太阳和天空都因这烟昏暗了。
REV|9|3|有蝗虫从烟中出来，飞到地上，有权柄赐给它们，好像地上的蝎子有权柄一样。
REV|9|4|它们奉命不可伤害地上的草、各样绿色植物和各种树木，惟独可伤害额上没有上帝印记的人；
REV|9|5|但是不许蝗虫害死他们，只可使他们受痛苦五个月；这痛苦就像人被蝎子螫了的痛苦一样。
REV|9|6|在那些日子，人求死，却死不了；想死，死却避开他们。
REV|9|7|蝗虫的形状好像预备上阵的战马一样，头上戴的好像金冠冕，脸面好像男人的脸面，
REV|9|8|头发像女人的头发，牙齿像狮子的牙齿；
REV|9|9|它们胸前有甲，好像铁甲；又有翅膀的响声，好像许多车马奔跑上阵的声音。
REV|9|10|它们有尾巴像蝎子，长着毒刺，尾巴上的毒刺有能力伤害人五个月。
REV|9|11|它们有无底坑的使者作它们的王，按着 希伯来 话名叫 亚巴顿 ， 希腊 话名话叫 亚玻伦 。
REV|9|12|第一样灾祸过去了；看哪，还有两样灾祸要来。
REV|9|13|第六位天使吹号，我听见有声音从上帝面前金坛的四 角发出来，
REV|9|14|吩咐那吹号的第六位天使，说：“把那捆绑在 幼发拉底 大河的四个使者释放了。”
REV|9|15|那四个使者就被释放；他们原是预备好，在特定的年、月、日、时，要杀人类的三分之一。
REV|9|16|骑兵有二亿；他们的数目我听见了。
REV|9|17|我在异象中看见那些马和骑马的：骑马的穿着火红、紫玛瑙及硫磺色的胸甲；马的头好像狮子的头，有火、有烟、有硫磺从马的口中喷出来。
REV|9|18|从马的口中所喷出来的火、烟和硫磺这三样灾害杀了人类的三分之一。
REV|9|19|马的能力在于它们的口和尾巴；它们的尾巴像蛇，有头，用头来伤害人。
REV|9|20|其余未曾被这些灾难所杀的人仍旧不为自己手所做的悔改，还是去拜鬼魔和那些不能看、不能听、不能走，用金、银、铜、木、石所造的偶像。
REV|9|21|他们也不为自己所犯的那些凶杀、邪术、淫乱、偷窃的事悔改。
REV|10|1|我又看见另一位大力的天使从天降下，披着云彩，头上有彩虹，脸面像太阳，两脚像火柱。
REV|10|2|他手里拿着展开的小书卷。他右脚踏海，左脚踏地，
REV|10|3|大声呼喊，好像狮子吼叫。呼喊完了，就有七个雷发出声音。
REV|10|4|七个雷发声后，我正要写出来，就听见从天上有声音说：“七个雷所说的，你要封上，不可写出来。”
REV|10|5|我所看见的那踏海踏地的天使向天举起右手，
REV|10|6|指着创造天和天上之物、地和地上之物、海和海中之物、直活到永永远远的那位起誓，说：“不再有时日了 。”
REV|10|7|但在第七位天使要吹号的日子，上帝的奥秘就要成全了，正如上帝向他仆人众先知所宣告的。
REV|10|8|我先前从天上所听见的那声音又吩咐我说：“你去，把那踏海踏地之天使手中展开的小书卷拿过来。”
REV|10|9|我就走到天使那里，对他说，请他把小书卷给我。他对我说：“你拿去，把它吃光。它会使你肚子发苦，然而在你口中会甘甜如蜜。”
REV|10|10|于是我从天使手中把小书卷接过来，把它吃光了，在我口中果然甘甜如蜜，吃了以后，我肚子觉得发苦。
REV|10|11|天使们对我说：“你必须指着许多民族、邦国、语言、君王再说预言。”
REV|11|1|有一根芦苇，像丈量的杖，赐给我；且有话说：“起来！将上帝的殿和祭坛，以及在殿中礼拜的人，都量一量。
REV|11|2|只是殿外的院子不用量，因为这是要给外邦人的；他们将践踏圣城四十二个月。
REV|11|3|“我要赐权柄给我那两个见证人，穿着粗麻衣说预言一千二百六十天。”
REV|11|4|他们就是那站在世界之主面前的两棵橄榄树和两个灯台。
REV|11|5|若有人想要害他们，就有火从他们口中喷出来，烧灭仇敌；凡想要害他们的都必须这样被杀。
REV|11|6|这二人有权柄关闭天空，使他们说预言的日子不下雨；又有权柄使水变为血，并且能随时随意用各样的灾害击打大地世界。
REV|11|7|他们作完见证的时候，那从无底坑里上来的兽要跟他们交战，并且得胜，把他们杀了。
REV|11|8|他们的尸首将倒在大城的街道上；这城按着灵意叫 所多玛 ，又叫 埃及 ，就是他们的主钉十字架的地方。
REV|11|9|从各民族、支派、语言、邦国中有人观看他们的尸首三天半，又不许人把尸首安放在坟墓里。
REV|11|10|住在地上的人会因他们而欢喜快乐，互相馈送礼物，因为这两位先知曾使住在地上的人受痛苦。
REV|11|11|过了这三天半，有生命的气息从上帝那里进入他们里面，他们就站起来；看见他们的人都大大惧怕。
REV|11|12|两位先知听见有大声音从天上对他们说：“上这里来。”他们就驾着云上了天，他们的仇敌也看见了。
REV|11|13|正在那时候，地大震动，城倒塌了十分之一；因地震而死的有七千人，其余的都恐惧，归荣耀给天上的上帝。
REV|11|14|第二样灾祸过去了；看哪，第三样灾祸快到了。
REV|11|15|第七位天使吹号，天上就有大声音说： “世上的国已成了我们的主和他所立的基督的国了。 他要作王直到永永远远！”
REV|11|16|在上帝面前，坐在自己座位上的二十四位长老都俯伏在地上敬拜上帝，
REV|11|17|说： “今在昔在的主—全能的上帝啊， 我们感谢你！ 因你执掌大权作王了。
REV|11|18|外邦发怒， 你的愤怒临到了。 审判死人的时候也到了； 你的仆人众先知、众圣徒及敬畏你名的人， 连大带小得赏赐的时候到了； 你毁灭那些毁灭大地者的时候也到了。”
REV|11|19|于是，上帝天上的圣所开了，在他圣所中，他的约柜出现了；随后有闪电、响声、雷轰、地震、大冰雹。
REV|12|1|天上出现了一个大兆头：有一个妇人身披太阳，脚踏月亮，头戴十二颗星的冠冕；
REV|12|2|她怀了孕，在生产的阵痛中疼痛地喊叫。
REV|12|3|天上又出现了另一个兆头：有一条大红龙 ，有七个头十个角；七个头上戴着七个冠冕。
REV|12|4|它的尾巴拖拉着天上星辰的三分之一，把它们摔在地上。然后龙站在那将要生产的妇人面前，等她生产后要吞吃她的孩子。
REV|12|5|妇人生了一个男孩子，就是将来要用铁杖管辖 万国的；她的孩子被提到上帝和他宝座那里去。
REV|12|6|妇人就逃到旷野，在那里有上帝给她预备的地方，使她在那里被供养一千二百六十天。
REV|12|7|天上发生了争战。 米迦勒 同他的使者与龙作战，龙同它的使者也起来应战，
REV|12|8|它们都打败了，天上再也没有它们的地方。
REV|12|9|大龙就是那古蛇，名叫魔鬼，又叫撒但，是迷惑普天下的；它被摔在地上，它的使者也一同被摔下去。
REV|12|10|我听见在天上有大声音说： “我上帝的救恩、能力、国度， 和他所立的基督的权柄现在都来到了。 因为那个在我们上帝面前、 昼夜控告我们弟兄的， 已经被摔下去了。
REV|12|11|弟兄胜过那条龙是因羔羊的血， 和因自己所见证的道。 虽然至于死，他们也不惜自己的性命。
REV|12|12|所以，诸天和住在其中的， 你们都快乐吧！ 只是地和海有祸了！ 因为魔鬼知道自己的时候不多， 就气愤愤地下到你们那里去了。”
REV|12|13|龙见自己被摔在地上，就迫害那生男孩子的妇人。
REV|12|14|于是有大鹰的两个翅膀赐给妇人，让她能飞到旷野，到自己的地方，躲避那蛇。她在那里受供养一载二载半载。
REV|12|15|蛇在妇人背后，从口中喷出水来，像河一样，要将妇人冲走。
REV|12|16|地却帮助了妇人，开口吞了从龙口喷出来的水。
REV|12|17|于是龙向妇人发怒，去与她其余的儿女作战，就是与那些遵守上帝命令 、为耶稣作见证的 。
REV|12|18|那时龙站在海边沙滩上。
REV|13|1|我又看见一只兽从海里上来，有十个角七个头；在十个角上戴着十个冠冕，七个头上有亵渎的名号。
REV|13|2|我所看见的兽，形状像豹，脚像熊的脚，口像狮子的口。那条龙将自己的能力、座位和大权柄都给了它。
REV|13|3|我看见兽的七个头中，有一个似乎受了致命伤，那伤却医好了。全地的人都很惊讶，跟从了那只兽。
REV|13|4|他们都拜那条龙，因为它把自己的权柄给了兽；又拜那只兽，说：“谁能比这只兽，谁能与它交战呢？”
REV|13|5|龙又赐给那只兽说夸大亵渎话的口，又赐给它权柄可以任意行事四十二个月。
REV|13|6|那兽就开口向上帝说亵渎的话，亵渎上帝的名和他的帐幕，就是那些住在天上的。
REV|13|7|它又被准许与圣徒作战，并且得胜，也赐给它权柄，可以制伏各支派、各民族、各语言、各邦国。
REV|13|8|凡住在地上、名字从创世以来没有记在被杀羔羊的生命册上的人都要拜它。
REV|13|9|凡有耳朵的都听吧！
REV|13|10|该被掳掠的，必被掳掠； 该被刀杀的，必被刀杀。 在此，圣徒要有耐心和信心。
REV|13|11|我又看见另一只兽从地里上来。它有两个角如同羔羊，说话好像龙。
REV|13|12|它在第一只兽面前施行第一只兽所有的权柄，并且使地和住在地上的人拜那致命伤被医好了的第一只兽。
REV|13|13|这只兽又行大奇事，甚至在人面前使火从天降在地上。
REV|13|14|它得了权柄在第一只兽面前能行奇事，迷惑住在地上的人，告诉他们要为那受过刀伤还活着的兽造个像。
REV|13|15|又有权柄赐给它，让那只兽的像有生气，并且能说话，又使所有不拜兽像的人都被杀害。
REV|13|16|它又使众人，无论大小、贫富，自主的、为奴的，都在右手上，或是在额上，打一个印记；
REV|13|17|这样，除了那有印记，有兽的名或有兽名数字的，都不得买或卖。
REV|13|18|在此，要有智慧：让有悟性的人解开兽的数目吧，因为这是一个人的数字，那数字是六百六十六。
REV|14|1|我又观看，看见羔羊站在 锡安山 ，和他在一起的有十四万四千人，都有他的名和他父亲的名写在额上。
REV|14|2|我听见从天上有声音，像众水的声音和大雷的声音，我所听见的声音好像琴师所弹的琴声。
REV|14|3|他们在宝座前，和在四活物及众长老前唱新歌，除了从地上买来的那十四万四千人以外，没有人能学这歌。
REV|14|4|这些人未曾沾染妇女，他们原是童身。羔羊无论往哪里去，他们都跟随他。他们是从人间买来的，作为初熟的果子归给上帝和羔羊。
REV|14|5|在他们口中找不出谎言，他们是没有瑕疵的。
REV|14|6|我又看见另一位天使在空中飞翔，有永远的福音要传给住在地上的人，就是各邦国、各支派、各语言、各民族。
REV|14|7|他大声说：“要敬畏上帝，把荣耀归给他，因为他施行审判的时候已经到了。要敬拜那创造天、地、海和水源的主。”
REV|14|8|另有第二位天使接着说：“倾覆了！那曾叫列国喝淫乱、烈怒之酒的大 巴比伦 倾覆了！”
REV|14|9|另有第三位天使接着他们，大声说：“若有人拜那只兽和兽像，在额上或在手上受了印记，
REV|14|10|他也必喝上帝烈怒的酒；这酒是斟在上帝愤怒的杯中的纯酒。他要在圣天使和羔羊面前，在火与硫磺之中受痛苦。
REV|14|11|使他们受痛苦的烟往上冒，直到永永远远。那些拜兽和兽像，受了它名字的印记的人，昼夜不得安宁。”
REV|14|12|在此，遵守上帝命令 和坚信耶稣真道的圣徒要有耐心。
REV|14|13|我听见从天上有声音说：“你要写下：从今以后，在主里死去的人有福了。”圣灵说：“是的，他们要从自己的劳苦中得安息，因为工作的成果永随着他们。”
REV|14|14|我又观看，看见有一片白云，云上坐着一位好像是人子的，头上戴着金冠冕，手里拿着锋利的镰刀。
REV|14|15|另有一位天使从圣所出来，向那坐在云上的大声喊着：“伸出你的镰刀来收割吧，因为收割的时候已经到了，地上的庄稼已经熟透了。”
REV|14|16|于是那坐在云上的把镰刀向地上挥去，地上的庄稼就收割了。
REV|14|17|另有一位天使从天上的圣所出来，他也拿着锋利的镰刀。
REV|14|18|另有一位天使从祭坛出来，是有权柄管火的，向那拿着锋利镰刀的大声喊着说：“伸出锋利的镰刀来，收取地上葡萄树的果子，因为葡萄熟透了。”
REV|14|19|那天使就把镰刀向地上挥去，收取了地上的葡萄，扔进上帝愤怒的大醡酒池里。
REV|14|20|那醡酒池在城外被踹踏，有血从醡酒池里流出来，涨到马的嚼环那么高，约有一千六百斯他迪 那么远。
REV|15|1|我看见在天上有另一兆头，大而且奇，就是七位天使掌管末了的七种灾难，因为上帝的烈怒在这七种灾难中发尽了。
REV|15|2|我看见仿佛有搀杂火的玻璃海；又看见那些胜了那兽和兽像，以及它名字的数字的人，都站在玻璃海上，拿着上帝的竖琴。
REV|15|3|他们唱上帝仆人 摩西 的歌和羔羊的歌，说： “主—全能的上帝啊， 你的作为又伟大又奇妙！ 万国之王啊， 你的道路又公义又真实！
REV|15|4|主啊，谁敢不敬畏你， 不把荣耀归于你的名？ 因为只有你是神圣的。 万民都要来， 在你面前敬拜， 因你公义的作为已经彰显了。”
REV|15|5|此后，我看见在天上那存放法柜的圣所开了。
REV|15|6|那掌管七种灾难的七位天使从圣所出来，穿着洁白明亮的细麻衣 ，胸间束着金带。
REV|15|7|四个活物中，有一个把盛满了活到永永远远之上帝烈怒的七个金碗给了那七位天使。
REV|15|8|圣所中充满了上帝的荣耀和权能而来的烟。没有人能进入圣所，直等到那七位天使降完了七种灾难。
REV|16|1|我听见有大声音从圣所里出来，向那七位天使说：“你们去，把盛着上帝烈怒的七碗倾倒在地上。”
REV|16|2|第一位天使去，把碗倾倒在地上，就有又臭又毒的疮生在那些有兽的印记和拜兽像的人身上。
REV|16|3|第二位天使把碗倾倒在海里，海就变成像死人的血一样，海里所有的活物都死了。
REV|16|4|第三位天使把碗倾倒在河流和水源里，水就变成血了。
REV|16|5|我听见掌管众水的天使说： “昔在、今在的圣者啊， 你做的判断公义；
REV|16|6|因他们曾流过圣徒与先知的血， 现在你给他们血喝， 这是他们该受的。”
REV|16|7|我又听见祭坛中有声音说： “是的，主—全能的上帝啊， 你的判断又真实又公义！”
REV|16|8|第四位天使把碗倾倒在太阳上，使太阳可用火烤人。
REV|16|9|人被炎热所烤，就亵渎那有权掌管这些灾难的上帝的名，他们没有悔改，也没有把荣耀归给上帝。
REV|16|10|第五位天使把碗倾倒在兽的座位上，兽的国就变成黑暗。人因疼痛而咬自己的舌头；
REV|16|11|又因所受的疼痛和生的疮，就亵渎天上的上帝，也没有为他们的行为悔改。
REV|16|12|第六位天使把碗倾倒在大 幼发拉底河 上，河水就干了，为要给从日出之地所来的众王预备道路。
REV|16|13|我又看见三个污秽的灵，好像青蛙，从龙的口、兽的口和假先知的口中出来。
REV|16|14|他们本是鬼魔的灵，施行奇事，到普天下众王那里去，召集他们在全能者上帝的大日子作战。
REV|16|15|看哪，我来像贼一样。那警醒、穿着衣服的人有福了；他不至于赤身而行，给人看见他的羞耻。
REV|16|16|于是，那三个鬼魔把众王聚集在 希伯来 话叫作 哈米吉多顿 的地方。
REV|16|17|第七位天使把碗倾倒在空中，就有大声音从圣所的宝座上出来，说：“成了！”
REV|16|18|又有闪电、响声、雷轰、大地震，自从地上有人以来没有这样大、这样厉害的地震。
REV|16|19|那大城裂为三段，列国的城也都倒塌了。上帝记起了大 巴比伦城 ，把那盛自己烈怒的酒杯递给她。
REV|16|20|各海岛都逃避了，众山也不见了。
REV|16|21|又有大冰雹从天掉落在人身上，每一个约重一他连得，以致人因冰雹的灾难而亵渎上帝，因为那灾难太大了。
REV|17|1|拿着七个碗的七位天使中，有一位前来对我说：“来，我要让你看那坐在众水之上的大淫妇所要受的惩罚；
REV|17|2|地上的君王都曾与她行淫，住在地上的人也喝醉了她淫乱的酒。”
REV|17|3|我在圣灵感动下，被天使带到旷野去，我看见一个女人骑在朱红色的兽上；那只兽有七个头十个角，遍体有亵渎的名号。
REV|17|4|那女人穿着紫色和朱红色的衣服，用金子、宝石、珍珠作妆饰，手拿着金杯，杯中盛满了可憎之物和她淫乱的污秽。
REV|17|5|在她额上写着奥秘的名字，说：“大 巴比伦 ，世上的淫妇和一切可憎之物的母。”
REV|17|6|我又看见那女人喝醉了圣徒的血和为耶稣作见证的人的血。 我看见她，非常诧异。
REV|17|7|天使对我说：“你为什么诧异呢？我要把这女人和驮着她那七头十角的兽的奥秘告诉你。
REV|17|8|你曾看见的兽，以前有，现在没有，将来要从无底坑里上来，又归于沉沦。凡住在地上、名字从创世以来没有记在生命册上的人看见那只兽都要诧异，因为它以前有，现在没有，以后再有。
REV|17|9|在此要有智慧的心思：那七个头就是女人所坐的七座山；他们又是七个王，
REV|17|10|五个已经倒了，一个还在，一个还没有来到；他来的时候必须只暂时停留。
REV|17|11|那以前有、现在没有的兽就是第八个，他也和那七个同列，正归于沉沦。
REV|17|12|你曾看见的那十个角就是十个王；他们还没有得到国度，但他们要和那只兽同得权柄作王一个时辰。
REV|17|13|他们同心把自己的能力权柄交给那只兽。
REV|17|14|他们将与羔羊作战，羔羊必胜过他们，因为羔羊是万主之主、万王之王，而同羔羊在一起的是蒙召、被选、忠心的人。”
REV|17|15|天使又对我说：“你所看见那淫妇坐的众水，就是许多民族、人民、邦国、语言。
REV|17|16|你所看见的那十个角与兽必恨这淫妇，他们要使她孤独赤身，又要吃她的肉，用火将她烧尽。
REV|17|17|因为上帝使诸王同心执行他的旨意，把他们自己的国交给那只兽，直等到上帝的话都应验了。
REV|17|18|你所看见的那女人就是管辖地上众王的大城。”
REV|18|1|此后，我看见另一位有大权柄的天使从天降下，地由于他的荣耀而发光。
REV|18|2|他以强而有力的声音喊着说： “倾覆了！大 巴比伦 倾覆了！ 她成了鬼魔的住处， 各样污秽之灵的巢穴， 各样污秽之鸟的窝， 各样污秽可憎之兽的出没处 。
REV|18|3|因为列国都喝了她淫乱大怒的酒 ； 地上的君王和她行淫； 地上的商人因她极度奢华而发了财。”
REV|18|4|我又听见另一个声音从天上说： “我的民哪，从那城出来吧！ 免得和她在罪上有份， 受她所受的灾殃；
REV|18|5|因她的罪恶滔天， 上帝已经记得她的不义。
REV|18|6|她怎样待人，也要怎样待她， 按她所行的加倍地报应她； 用她调酒的杯加倍调给她喝。
REV|18|7|她怎样荣耀自己，怎样奢华， 也要使她照样痛苦悲哀。 因她心里说： ‘我坐了皇后的位， 并不是寡妇， 绝不至于悲哀。’
REV|18|8|所以在一天之内，她的灾殃要一齐来到， 就是死亡、悲哀、饥荒。 她将被火烧尽， 因为审判她的主上帝大有能力。”
REV|18|9|地上的君王，与她行淫、一同奢华的，看见烧她的烟，就必为她哭泣哀号；
REV|18|10|因怕她的痛苦，就远远地站着，说： “祸哉，祸哉，这大城！ 坚固的 巴比伦城 啊！ 一时之间，你的审判要来到了。”
REV|18|11|地上的商人也都为她哭泣悲哀，因为没有人再买他们的货物了；
REV|18|12|这货物就是金、银、宝石、珍珠、细麻布、丝绸、紫色和朱红色衣料、各样香木、各样象牙的器皿、各样极宝贵的木头和铜、铁、大理石的器皿，
REV|18|13|和肉桂、豆蔻、香料、香膏、乳香、酒、油、细面、麦子、牛、羊、马、马车，以及奴隶、人口。
REV|18|14|“你所贪爱的果子离开了你； 你一切的珍馐美味和华美的物件 都从你那里毁灭， 绝对见不到了。”
REV|18|15|贩卖这些货物、藉着她发财的商人，因怕她的痛苦，就远远地站着哭泣悲哀，
REV|18|16|说： “祸哉，祸哉，这大城！ 她穿着细麻、 紫色、朱红色的衣服， 用金子、宝石、珍珠为妆饰。
REV|18|17|一时之间，这么多的财富就归于无有了。” 所有的船长和到处航海的，水手以及所有靠海为业的，都远远地站着，
REV|18|18|看见烧她的烟，就喊着说：“有哪一个城能跟这大城比呢？”
REV|18|19|于是他们把灰尘撒在头上，哭泣悲哀地喊着说： “祸哉，祸哉，这大城！ 凡有船在海中的， 都因她的珍宝成了富足。 她在一时之间就成为荒芜。
REV|18|20|天哪，众圣徒、众使徒、众先知啊！ 你们都要因她欢喜， 因为上帝已经在她身上为你们伸了冤。”
REV|18|21|有一位大力的天使举起一块石头，好像大磨石，扔在海里，说： “ 巴比伦 大城 也必这样猛力地被扔下去， 绝对见不到了。
REV|18|22|弹琴、歌唱、 吹笛、吹号的声音， 在你中间绝对听不见了； 各行手艺的技工 在你中间绝对见不到了； 推磨的声音 在你中间绝对听不见了；
REV|18|23|灯台的光 在你中间绝对不再照耀了； 新郎和新娘的声音 在你中间绝对听不见了。 你的商人原来是地上的显要； 万国也被你的邪术迷惑了。
REV|18|24|先知、圣徒和地上一切被杀的人的血都在这城里找到了。”
REV|19|1|此后，我听见好像有一大群人在天上大声说： “哈利路亚 ！ 救恩、荣耀、权能都属于我们的上帝。
REV|19|2|他的判断又真实又公义； 因他判断了那大淫妇， 她用淫行败坏了世界。 上帝为他的仆人伸冤， 向淫妇讨流仆人血的罪。”
REV|19|3|他们又一次说： “哈利路亚！ 烧淫妇的烟往上冒，直到永永远远。”
REV|19|4|那二十四位长老和四活物就俯伏敬拜坐在宝座上的上帝，说： “阿们。哈利路亚！”
REV|19|5|接着，有声音从宝座出来说： “上帝的众仆人哪， 凡敬畏他的， 无论大小， 都要赞美我们的上帝！”
REV|19|6|我听见好像一大群人的声音，像众水的声音，像大雷的声音，说： “哈利路亚！ 因为主─我们的上帝 、 全能者，作王了。
REV|19|7|我们要欢喜快乐， 将荣耀归给他； 因为羔羊的婚期到了， 他的新娘也自己预备好了，
REV|19|8|她蒙恩得穿明亮洁白的细麻衣： 这细麻衣就是圣徒们的义行。”
REV|19|9|天使对我说：“你要写下来：凡被请赴羔羊婚宴的人有福了！”他又对我说：“这些都是上帝真实的话。”
REV|19|10|我就俯伏在他脚前要拜他。他对我说：“千万不可！我和你，以及那些为耶稣作见证的弟兄同是仆人。你要敬拜上帝。”因为那些为耶稣作见证的人有预言的灵。
REV|19|11|后来我看见天开了。有一匹白马，骑在马上的称为 “诚信”、“真实”，他审判和争战都凭着公义。
REV|19|12|他的眼睛如 火焰，头上戴着许多冠冕；他身上写着一个名字，除了他自己没有人知道。
REV|19|13|他穿着浸过血的衣服；他的名称为“上帝之道”。
REV|19|14|众天军都骑着白马，穿着又白又洁净的细麻衣跟随他。
REV|19|15|有利剑从他口中出来，用来击打列国。他要用铁杖管辖 他们，并且要踹全能上帝烈怒的醡酒池。
REV|19|16|在他衣服和大腿上写着“万王之王，万主之主”的名号。
REV|19|17|我又看见一位天使站在太阳中，向天空一切的飞鸟大声喊着说：“你们聚集来赴上帝的大宴席，
REV|19|18|为要吃君王的肉、将军的肉、壮士的肉、马和骑士的肉、一切自主的和为奴的，以及尊贵的和卑贱的肉。”
REV|19|19|我又看见那兽和地上的君王，和他们的军队都聚集，要与白马骑士和他的军队作战。
REV|19|20|那兽被擒拿了；那在兽面前曾行奇事、迷惑了接受兽的印记和拜兽像的人的假先知，也与兽同被擒拿。他们两个就活生生地被扔进烧着硫磺的火湖里，
REV|19|21|其余的人被白马骑士口中吐出来的剑杀了；所有的飞鸟都吃饱了他们的肉。
REV|20|1|我又看见一位天使从天降下，手里拿着无底坑的钥匙和一条大铁链。
REV|20|2|他抓住那龙，那古蛇，就是魔鬼、撒但，把它捆绑了一千年，
REV|20|3|扔在无底坑里，把无底坑关闭，用印封上，使它不再迷惑列国，等到那一千年满了。这些事以后，它必须暂时被释放。
REV|20|4|我又看见一些宝座，坐在上面的有审判的权柄赐给他们。我又看见那些因为给耶稣作见证，并为上帝之道被斩首的人的灵魂，和没有拜过那兽与兽像、也没有在额上和手上打过它印记的人的灵魂。他们都复活了，与基督一同作王一千年。
REV|20|5|这是头一次的复活。其余的死人还没有复活，直等那一千年满了。
REV|20|6|在头一次复活有份的有福了，圣洁了！第二次的死在他们身上没有权柄，但他们要作上帝和基督的祭司，也要与基督一同作王一千年。
REV|20|7|那一千年满了，撒但会从监牢里被释放，
REV|20|8|出来要迷惑地上四方的列国，就是 歌革 和 玛各 ，使他们聚集争战。他们的人数多如海沙。
REV|20|9|他们上来布满了全地，围住圣徒的营与蒙爱的城，就有火从天降下，烧灭了他们。
REV|20|10|那迷惑他们的魔鬼被扔进硫磺的火湖里，就是那兽和假先知所在的地方，他们会昼夜受折磨，直到永永远远。
REV|20|11|我又看见一个白色的大宝座和那坐在上面的；天和地都从他面前逃避，再也找不到它们的位置了。
REV|20|12|我又看见死了的人，无论大小，都站在宝座前。案卷都展开了，并另有一卷展开，就是生命册。死了的人都凭着这些案卷所记载的，照他们所行的受审判。
REV|20|13|于是海交出其中的死人，死亡和阴间也交出其中的死人；他们都照各人所行的受审判。
REV|20|14|死亡和阴间也被扔进火湖里，这火湖就是第二次的死。
REV|20|15|凡名字没有记在生命册上的人，就被扔进火湖里。
REV|21|1|我又看见一个新天新地，因为先前的天和先前的地已经过去了，海也不再有了。
REV|21|2|我又看见圣城，新 耶路撒冷 由上帝那里，从天而降，预备好了，就如新娘打扮整齐，等候丈夫。
REV|21|3|我听见有大声音从宝座出来，说： “看哪，上帝的帐幕在人间！ 他要和他们同住， 他们要作他的子民。 上帝要亲自与他们同在。
REV|21|4|上帝要擦去他们一切的眼泪； 不再有死亡， 也不再有悲哀、哭号、痛苦， 因为先前的事都过去了。”
REV|21|5|那位坐在宝座上的说：“看哪，我把一切都更新了！”他又说：“你要写下来，因为这些话是可信靠的，是真实的。”
REV|21|6|他又对我说：“成了！我是阿拉法，我是俄梅戛；我是开始，我是终结。我要把生命的泉水白白赐给那口渴的人喝。
REV|21|7|得胜的要承受这些为业；我要作他的上帝，他要作我的儿子。
REV|21|8|至于胆怯的、不信的、可憎的、杀人的、淫乱的、行邪术的、拜偶像的和一切说谎话的人，他们将在烧着硫磺的火湖里有份；这是第二次的死。”
REV|21|9|拿着七个金碗、盛满末后七种灾祸的七位天使中，有一位来对我说：“你来，我要给你看新娘，就是羔羊的妻子。”
REV|21|10|我在圣灵感动下，天使带我到一座高大的山，给我看由上帝那里、从天而降的圣城 耶路撒冷 ，
REV|21|11|这城有上帝的荣耀，它光辉如同极贵的宝石，好像碧玉，明如水晶。
REV|21|12|它有高大的墙，有十二个门，门上有十二位天使，门上又写着 以色列 人十二个支派的名字 。
REV|21|13|东边有三个门，北边有三个门，南边有三个门，西边有三个门。
REV|21|14|城墙有十二个根基，根基上有羔羊十二使徒的名字。
REV|21|15|那对我说话的天使拿着金的芦苇当尺，要量那城、城门和城墙。
REV|21|16|城是四方的，长宽一样。天使用芦苇量那城，共有一万二千斯他迪，长、宽、高都是一样。
REV|21|17|他又量了城墙，按着人的尺寸，就是天使的尺寸，共有一百四十四肘。
REV|21|18|墙是碧玉造的；城是纯金的，如同明净的玻璃。
REV|21|19|城墙的根基是用各样宝石修饰的：第一个根基是碧玉，第二是蓝宝石，第三是绿玛瑙，第四是绿宝石，
REV|21|20|第五是红玛瑙，第六是红宝石，第七是黄璧玺，第八是水苍玉，第九是红璧玺，第十是翡翠，第十一是紫玛瑙，第十二是紫晶。
REV|21|21|十二个门是十二颗珍珠；每一个门是一颗珍珠造的。城内的街道是纯金的，好像透明的玻璃。
REV|21|22|我没有看见城内有殿，因主—全能者上帝和羔羊就是城的殿。
REV|21|23|那城内不用日月光照，因为有上帝的荣耀光照，又有羔羊为城的灯。
REV|21|24|列国要藉着城的光行走；地上的君王要把自己的荣耀带给那城。
REV|21|25|城门白昼总不关闭，在那里没有黑夜。
REV|21|26|人要将列国的荣耀尊贵带给那城。
REV|21|27|凡不洁净的，和那行可憎与虚谎之事的人，都不得进那城，只有名字写在羔羊生命册上的才得进去。
REV|22|1|天使又让我看一道生命水的河，明亮如水晶，从上帝和羔羊的宝座流出来，
REV|22|2|经过城内街道的中央；在河的两边有生命树，结十二样 的果子，每月都结果子；树上的叶子可作医治万民之用。
REV|22|3|以后不再有任何诅咒。在城里将有上帝和羔羊的宝座。他的仆人都要事奉他，
REV|22|4|也要见他的面。他的名字将写在他们的额上。
REV|22|5|不再有黑夜；他们也不需要灯光或日光，因为主上帝要光照他们。他们要作王，直到永永远远。
REV|22|6|天使又对我说：“这些话是可信靠的，是真实的。主，就是赐灵感给众先知的上帝，差遣他的使者，要将必须快要发生的事指示他的众仆人。”
REV|22|7|“看哪，我必快来！凡遵守这书上预言的有福了。”
REV|22|8|这些事是我－ 约翰 所听见所看见的。当我听见看见时，就俯伏在指示我的天使脚前要拜他。
REV|22|9|他对我说：“千万不可！我与你和你的弟兄众先知，以及那些守这书上的话的人，同是作仆人。你要敬拜上帝。”
REV|22|10|他又对我说：“不可封了这书上的预言，因为时候近了。
REV|22|11|不义的，让他仍旧不义；污秽的，让他仍旧污秽；为义的，让他仍旧为义；圣洁的，让他仍旧圣洁。”
REV|22|12|“看哪，我必快来！赏罚在我，要照每个人所行的报应他。
REV|22|13|我是阿拉法，我是俄梅戛；我是首先的，我是末后的；我是开始，我是终结。”
REV|22|14|那些洗净自己衣服的有福了！他们可得权柄到生命树那里，也能从门进城。
REV|22|15|城外有犬类、行邪术的、淫乱的、杀人的、拜偶像的，以及所有喜爱和行虚谎的人。
REV|22|16|“我－耶稣差遣我的使者，为了众教会向你们证明这些事。我是 大卫 的根，是他的后裔；我是明亮的晨星。”
REV|22|17|圣灵和新娘都说：“来！”听见的人也要说：“来！”口渴的人也要来，愿意的人都可以白白取生命的水喝。
REV|22|18|我警告一切听见这书上预言的人：若有人在这预言上加添什么，上帝必将记在这书上的灾祸加在他身上。
REV|22|19|这书上的预言，若有人删去什么，上帝必从这书上所记的生命树和圣城删去他的份。
REV|22|20|证明这些事的说：“是的，我必快来！”阿们！主耶稣啊，我愿你来！
REV|22|21|愿主耶稣的恩惠与众圣徒同在。阿们！
