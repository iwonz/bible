2CHR|1|1|confortatus est ergo Salomon filius David in regno suo et Dominus erat cum eo et magnificavit eum in excelsum
2CHR|1|2|praecepitque Salomon universo Israheli tribunis et centurionibus et ducibus et iudicibus omnis Israhel et principibus familiarum
2CHR|1|3|et abiit cum universa multitudine in excelsum Gabaon ubi erat tabernaculum foederis Dei quod fecit Moses famulus Dei in solitudine
2CHR|1|4|arcam autem Dei adduxerat David de Cariathiarim in locum quem paraverat ei et ubi fixerat illi tabernaculum hoc est in Hierusalem
2CHR|1|5|altare quoque aeneum quod fabricatus fuerat Beselehel filius Uri filii Ur ibi erat coram tabernaculo Domini quod et requisivit Salomon et omnis ecclesia
2CHR|1|6|ascenditque Salomon ad altare aeneum coram tabernaculo foederis Domini et obtulit in eo mille hostias
2CHR|1|7|ecce autem in ipsa nocte apparuit ei Deus dicens postula quod vis ut dem tibi
2CHR|1|8|dixitque Salomon Deo tu fecisti cum David patre meo misericordiam magnam et constituisti me regem pro eo
2CHR|1|9|nunc igitur Domine Deus impleatur sermo tuus quem pollicitus es David patri meo tu enim fecisti me regem super populum tuum multum qui tam innumerabilis est quam pulvis terrae
2CHR|1|10|da mihi sapientiam et intellegentiam ut egrediar coram populo tuo et ingrediar quis enim potest hunc populum tuum digne qui tam grandis est iudicare
2CHR|1|11|dixit autem Deus ad Salomonem quia hoc magis placuit cordi tuo et non postulasti divitias et substantiam et gloriam neque animas eorum qui te oderunt sed nec dies vitae plurimos petisti autem sapientiam et scientiam ut iudicare possis populum meum super quem constitui te regem
2CHR|1|12|sapientia et scientia data sunt tibi divitias autem et substantiam et gloriam dabo tibi ita ut nullus in regibus nec ante te nec post te fuerit similis tui
2CHR|1|13|venit ergo Salomon ab excelso Gabaon in Hierusalem coram tabernaculo foederis et regnavit super Israhel
2CHR|1|14|congregavitque sibi currus et equites et facti sunt ei mille quadringenti currus et duodecim milia equitum et fecit eos esse in urbibus quadrigarum et cum rege in Hierusalem
2CHR|1|15|praebuitque rex argentum et aurum in Hierusalem quasi lapides et cedros quasi sycomoros quae nascuntur in campestribus multitudine magna
2CHR|1|16|adducebantur autem ei et equi de Aegypto et de Coa a negotiatoribus regis qui ibant et coemebant pretio
2CHR|1|17|quadrigam equorum sescentis argenteis et equum centum quinquaginta similiter de universis regnis Cettheorum et a regibus Syriae emptio celebrabatur
2CHR|2|1|decrevit autem Salomon aedificare domum nomini Domini et palatium sibi
2CHR|2|2|et numeravit septuaginta milia virorum portantium umeris et octoginta milia qui caederent lapides in montibus praepositosque eorum tria milia sescentos
2CHR|2|3|misit quoque ad Hiram regem Tyri dicens sicut egisti cum David patre meo et misisti ei ligna cedrina ut aedificaret sibi domum in qua et habitavit
2CHR|2|4|sic fac mecum ut aedificem domum nomini Domini Dei mei et consecrem eam ad adolendum incensum coram illo et fumiganda aromata et ad propositionem panum sempiternam et holocaustomata mane et vespere sabbatis quoque et neomeniis et sollemnitatibus Domini Dei nostri in sempiternum quae mandata sunt Israheli
2CHR|2|5|domus autem quam aedificare cupio magna est magnus est enim Deus noster super omnes deos
2CHR|2|6|quis ergo poterit praevalere ut aedificet ei dignam domum si caelum et caeli caelorum capere eum non queunt quantus ego sum ut possim ei aedificare domum sed ad hoc tantum ut adoleatur incensum coram illo
2CHR|2|7|mitte igitur mihi virum eruditum qui noverit operari in auro et argento aere ferro purpura coccino et hyacintho et qui sciat scalpere celata cum his artificibus quos mecum habeo in Iudaea et in Hierusalem quos praeparavit David pater meus
2CHR|2|8|sed et ligna cedrina mitte mihi et arceuthina et pinea de Libano scio enim quod servi tui noverint caedere ligna de Libano et erunt servi mei cum servis tuis
2CHR|2|9|ut parentur mihi ligna plurima domus enim quam cupio aedificare magna est nimis et inclita
2CHR|2|10|praeterea operariis qui caesuri sunt ligna servis tuis dabo in cibaria tritici choros viginti milia et hordei choros totidem olei quoque sata viginti milia
2CHR|2|11|dixit autem Hiram rex Tyri per litteras quas miserat Salomoni quia dilexit Dominus populum suum idcirco te regnare fecit super eum
2CHR|2|12|et addidit dicens benedictus Dominus Deus Israhel qui fecit caelum et terram qui dedit David regi filium sapientem et eruditum et sensatum atque prudentem ut aedificaret domum Domino et palatium sibi
2CHR|2|13|misi ergo tibi virum prudentem et scientissimum Hiram patrem meum
2CHR|2|14|filium mulieris de filiabus Dan cuius pater Tyrius fuit qui noverit operari in auro et argento et aere et ferro et marmore et lignis in purpura quoque et hyacintho et bysso et coccino et qui sciat celare omnem scalpturam et adinvenire prudenter quodcumque in opere necessarium est cum artificibus tuis et cum artificibus domini mei David patris tui
2CHR|2|15|triticum ergo et hordeum et oleum et vinum quae pollicitus es domine mi mitte servis tuis
2CHR|2|16|nos autem caedemus ligna de Libano quot necessaria habueris et adplicabimus ea ratibus per mare in Ioppe tuum erit transferre ea in Hierusalem
2CHR|2|17|numeravit igitur Salomon omnes viros proselytos qui erant in terra Israhel post dinumerationem quam dinumeravit David pater eius et inventi sunt centum quinquaginta milia et tria milia sescenti
2CHR|2|18|fecitque ex eis septuaginta milia qui umeris onera portarent et octoginta milia qui lapides in montibus caederent tria milia autem et sescentos praepositos operum populi
2CHR|3|1|et coepit Salomon aedificare domum Domini in Hierusalem in monte Moria qui demonstratus fuerat David patri eius in loco quem paraverat David in area Ornan Iebusei
2CHR|3|2|coepit autem aedificare mense secundo anno quarto regni sui
2CHR|3|3|et haec sunt fundamenta quae iecit Salomon ut aedificaret domum Dei longitudinis cubitos in mensura prima sexaginta latitudinis cubitos viginti
2CHR|3|4|porticum vero ante frontem quae tendebatur in longum iuxta mensuram latitudinis domus cubitorum viginti porro altitudo centum viginti cubitorum erat et deauravit eam intrinsecus auro mundissimo
2CHR|3|5|domum quoque maiorem texit tabulis ligneis abiegnis et lamminas auri obrizi adfixit per totum scalpsitque in ea palmas et quasi catenulas se invicem conplectentes
2CHR|3|6|stravit quoque pavimentum templi pretiosissimo marmore decore multo
2CHR|3|7|porro aurum erat probatissimum de cuius lamminis texit domum et trabes eius et postes et parietes et ostia et celavit cherubin in parietibus
2CHR|3|8|fecit quoque domum sancti sanctorum longitudinem iuxta latitudinem domus cubitorum viginti et latitudinem similiter viginti cubitorum et lamminis aureis texit eam quasi talentis sescentis
2CHR|3|9|sed et clavos fecit aureos ita ut singuli clavi siclos quinquagenos adpenderent cenacula quoque texit auro
2CHR|3|10|fecit etiam in domo sancti sanctorum cherubin duo opere statuario et texit eos auro
2CHR|3|11|alae cherubin viginti cubitis extendebantur ita ut una ala haberet cubitos quinque et tangeret parietem domus et altera quinque cubitos habens alam tangeret alterius cherub
2CHR|3|12|similiter cherub alterius ala quinque habebat cubitos et tangebat parietem et ala eius altera quinque cubitorum alam cherub alterius contingebat
2CHR|3|13|igitur alae utriusque cherubin expansae erant et extendebantur per cubitos viginti ipsi autem stabant erectis pedibus et facies eorum versae erant ad exteriorem domum
2CHR|3|14|fecit quoque velum ex hyacintho purpura coccino et bysso et intexuit ei cherubin
2CHR|3|15|ante fores etiam templi duas columnas quae triginta et quinque cubitos habebant altitudinis porro capita earum quinque cubitorum
2CHR|3|16|necnon et quasi catenulas in oraculo et superposuit eas capitibus columnarum malagranata etiam centum quae catenulis interposuit
2CHR|3|17|ipsas quoque columnas posuit in vestibulo templi unam a dextris et alteram a sinistris eam quae a dextris erat vocavit Iachin et quae ad levam Booz
2CHR|4|1|fecit quoque altare aeneum viginti cubitorum longitudinis et viginti cubitorum latitudinis et decem cubitorum altitudinis
2CHR|4|2|mare etiam fusile decem cubitis a labio usque ad labium rotundum per circuitum quinque cubitos habebat altitudinis et funiculus triginta cubitorum ambiebat gyrum eius
2CHR|4|3|similitudo quoque boum erat subter illud et decem cubitis quaedam extrinsecus celaturae quasi duobus versibus alvum maris circuibant boves autem erant fusiles
2CHR|4|4|et ipsum mare super duodecim boves inpositum erat quorum tres respiciebant aquilonem et alii tres occidentem porro tres alii meridiem et tres qui reliqui erant orientem mare habentes superpositum posteriora autem boum erant intrinsecus sub mari
2CHR|4|5|porro vastitas eius habebat mensuram palmi et labium illius erat quasi labium calicis vel repandi lilii capiebatque mensurae tria milia metretas
2CHR|4|6|fecit quoque concas decem et posuit quinque a dextris et quinque a sinistris ut lavarent in eis omnia quae in holocaustum oblaturi erant porro in mari sacerdotes lavabantur
2CHR|4|7|fecit autem et candelabra aurea decem secundum speciem qua iussa erant fieri et posuit ea in templo quinque a dextris et quinque a sinistris
2CHR|4|8|necnon et mensas decem posuitque eas in templo quinque a dextris et quinque a sinistris fialas quoque aureas centum
2CHR|4|9|fecit etiam atrium sacerdotum et basilicam grandem et ostia in basilica quae texit aere
2CHR|4|10|porro mare posuit in latere dextro contra orientem ad meridiem
2CHR|4|11|fecit autem Hiram lebetas quoque et creagras et fialas et conplevit omne opus regis in domo Dei
2CHR|4|12|hoc est columnas duas et epistylia et capita et quasi quaedam retiacula quae capita tegerent super epistylia
2CHR|4|13|malagranata quoque quadringenta et retiacula duo ita ut bini ordines malagranatorum singulis retiaculis iungerentur quae protegerent epistylia et capita columnarum
2CHR|4|14|bases etiam fecit et concas quas superposuit basibus
2CHR|4|15|mare unum bovesque duodecim sub mari
2CHR|4|16|et lebetas et creagras et fialas omnia vasa fecit Salomoni Hiram pater eius in domo Domini ex aere mundissimo
2CHR|4|17|in regione Iordanis fudit ea rex in argillosa terra inter Socchoth et Saredatha
2CHR|4|18|erat autem multitudo vasorum innumerabilis ita ut ignoraretur pondus aeris
2CHR|4|19|fecitque Salomon omnia vasa domus Dei et altare aureum et mensas et super eas panes propositionis
2CHR|4|20|candelabra quoque cum lucernis suis ut lucerent ante oraculum iuxta ritum ex auro purissimo
2CHR|4|21|et florentia quaedam et lucernas et forcipes aureos omnia de auro mundissimo facta sunt
2CHR|4|22|thymiamateria quoque et turibula et fialas et mortariola ex auro purissimo et ostia celavit templi interioris id est in sancto sanctorum et ostia templi forinsecus aurea sicque conpletum est omne opus quod fecit Salomon in domo Domini
2CHR|5|1|intulit igitur Salomon omnia quae voverat David pater suus argentum et aurum et universa vasa posuit in thesauris domus Dei
2CHR|5|2|post quae congregavit maiores natu Israhel et cunctos principes tribuum et capita familiarum de filiis Israhel in Hierusalem ut adducerent arcam foederis Domini de civitate David quae est Sion
2CHR|5|3|venerunt igitur ad regem omnes viri Israhel in die sollemni mensis septimi
2CHR|5|4|cumque venissent cuncti seniorum Israhel portaverunt Levitae arcam
2CHR|5|5|et intulerunt eam et omnem paraturam tabernaculi porro vasa sanctuarii quae erant in tabernaculo portaverunt sacerdotes cum Levitis
2CHR|5|6|rex autem Salomon et universus coetus Israhel et omnes qui fuerant congregati ante arcam immolabant arietes et boves absque ullo numero tanta enim erat multitudo victimarum
2CHR|5|7|et intulerunt sacerdotes arcam foederis Domini in locum suum id est ad oraculum templi in sancta sanctorum subter alas cherubin
2CHR|5|8|ita ut cherubin expanderent alas suas super locum in quo posita erat arca et ipsam arcam tegerent cum vectibus eius
2CHR|5|9|vectium autem quibus portabatur arca quia paululum longiores erant capita parebant ante oraculum si vero quis paululum fuisset extrinsecus eos videre non poterat fuit itaque arca ibi usque in praesentem diem
2CHR|5|10|nihilque erat aliud in arca nisi duae tabulae quas posuerat Moses in Horeb quando legem dedit Dominus filiis Israhel egredientibus ex Aegypto
2CHR|5|11|egressis autem sacerdotibus de sanctuario omnes enim sacerdotes qui ibi potuerant inveniri sanctificati sunt nec adhuc illo tempore vices et ministeriorum ordo inter eos divisus erat
2CHR|5|12|tam Levitae quam cantores id est et qui sub Asaph erant et qui sub Heman et qui sub Idithun filii et fratres eorum vestiti byssinis cymbalis et psalteriis et citharis concrepabant stantes ad orientalem plagam altaris cumque eis sacerdotes centum viginti canentes tubis
2CHR|5|13|igitur cunctis pariter et tubis et voce et cymbalis et organis et diversi generis musicorum concinentibus et vocem in sublime tollentibus longe sonitus audiebatur ita ut cum Dominum laudare coepissent et dicere confitemini Domino quoniam bonus quoniam in aeternum misericordia eius impleretur domus Domini nube
2CHR|5|14|nec possent sacerdotes stare et ministrare propter caliginem conpleverat enim gloria Domini domum Dei
2CHR|6|1|tunc Salomon ait Dominus pollicitus est ut habitaret in caligine
2CHR|6|2|ego autem aedificavi domum nomini eius ut habitaret ibi in perpetuum
2CHR|6|3|et convertit faciem suam et benedixit universae multitudini Israhel nam omnis turba stabat intenta et ait
2CHR|6|4|benedictus Dominus Deus Israhel qui quod locutus est David patri meo opere conplevit dicens
2CHR|6|5|a die qua eduxi populum meum de terra Aegypti non elegi civitatem de cunctis tribubus Israhel ut aedificaretur in ea domus nomini meo neque elegi quemquam alium virum ut esset dux in populo meo Israhel
2CHR|6|6|sed elegi Hierusalem ut sit nomen meum in ea et elegi David ut constituerem eum super populum meum Israhel
2CHR|6|7|cumque fuisset voluntatis David patris mei ut aedificaret domum nomini Domini Dei Israhel
2CHR|6|8|dixit Dominus ad eum quia haec fuit voluntas tua ut aedificares domum nomini meo bene quidem fecisti habere huiuscemodi voluntatem
2CHR|6|9|sed non tu aedificabis domum verum filius tuus qui egredietur de lumbis tuis ipse aedificabit domum nomini meo
2CHR|6|10|conplevit ergo Dominus sermonem suum quem locutus fuerat et ego surrexi pro David patre meo et sedi super thronum Israhel sicut locutus est Dominus et aedificavi domum nomini Domini Dei Israhel
2CHR|6|11|et posui in ea arcam in qua est pactum Domini quod pepigit cum filiis Israhel
2CHR|6|12|stetit ergo coram altare Domini ex adverso universae multitudinis Israhel et extendit manus suas
2CHR|6|13|siquidem fecerat Salomon basem aeneam et posuerat eam in medio basilicae habentem quinque cubitos longitudinis et quinque cubitos latitudinis et tres cubitos in altum stetitque super eam et deinceps flexis genibus contra universam multitudinem Israhel et palmis in caelum levatis
2CHR|6|14|ait Domine Deus Israhel non est similis tui Deus in caelo et in terra qui custodis pactum et misericordiam cum servis tuis qui ambulant coram te in toto corde suo
2CHR|6|15|qui praestitisti servo tuo David patri meo quaecumque locutus fueras ei et quae ore promiseras opere conplesti sicut et praesens tempus probat
2CHR|6|16|nunc ergo Domine Deus Israhel imple servo tuo patri meo David quaecumque locutus es dicens non deficiet ex te vir coram me qui sedeat super thronum Israhel ita tamen si custodierint filii tui vias suas et ambulaverint in lege mea sicut et tu ambulasti coram me
2CHR|6|17|et nunc Domine Deus Israhel firmetur sermo tuus quem locutus es servo tuo David
2CHR|6|18|ergone credibile est ut habitet Deus cum hominibus super terram si caelum et caeli caelorum non te capiunt quanto magis domus ista quam aedificavi
2CHR|6|19|sed ad hoc tantum facta est ut respicias orationem servi tui et obsecrationem eius Domine Deus meus audias et preces quas fundit famulus tuus coram te
2CHR|6|20|ut aperias oculos tuos super domum istam diebus et noctibus super locum in quo pollicitus es ut invocaretur nomen tuum
2CHR|6|21|et exaudires orationem quam servus tuus orat in eo exaudi preces famuli tui et populi tui Israhel quicumque oraverit in loco isto et exaudi de habitaculo tuo id est de caelis et propitiare
2CHR|6|22|si peccaverit quispiam in proximum suum et iurare contra eum paratus venerit seque maledicto constrinxerit coram altari in domo ista
2CHR|6|23|tu audies de caelo et facies iudicium servorum tuorum ita ut reddas iniquo viam suam in caput proprium et ulciscaris iustum retribuens ei secundum iustitiam suam
2CHR|6|24|si superatus fuerit populus tuus Israhel ab inimicis peccabunt enim tibi et conversi egerint paenitentiam et obsecraverint nomen tuum et fuerint deprecati in loco isto
2CHR|6|25|tu exaudi de caelo et propitiare peccato populi tui Israhel et reduc eos in terram quam dedisti eis et patribus eorum
2CHR|6|26|si clauso caelo pluvia non fluxerit propter peccata populi et deprecati te fuerint in loco isto et confessi nomini tuo et conversi a peccatis suis cum eos adflixeris
2CHR|6|27|exaudi de caelo Domine et dimitte peccata servis tuis et populi tui Israhel et doce eos viam bonam per quam ingrediantur et da pluviam terrae quam dedisti populo tuo ad possidendum
2CHR|6|28|fames si orta fuerit in terra et pestilentia erugo et aurugo et lucusta et brucus et hostes vastatis regionibus portas obsederint civitatis omnisque plaga et infirmitas presserit
2CHR|6|29|si quis de populo tuo Israhel fuerit deprecatus cognoscens plagam et infirmitatem suam et expanderit manus suas in domo hac
2CHR|6|30|tu exaudi de caelo de sublimi scilicet habitaculo tuo et propitiare et redde unicuique secundum vias suas quas nosti eum habere in corde suo tu enim solus nosti corda filiorum hominum
2CHR|6|31|ut timeant te et ambulent in viis tuis cunctis diebus quibus vivunt super faciem terrae quam dedisti patribus nostris
2CHR|6|32|externum quoque qui non est de populo tuo Israhel si venerit de terra longinqua propter nomen tuum magnum et propter manum tuam robustam et brachium tuum extentum et adoraverit in loco isto
2CHR|6|33|tu exaudies de caelo firmissimo habitaculo tuo et facies cuncta pro quibus invocaverit te ille peregrinus ut sciant omnes populi terrae nomen tuum et timeant te sicut populus tuus Israhel et cognoscant quia nomen tuum invocatum est super domum hanc quam aedificavi
2CHR|6|34|si egressus fuerit populus tuus ad bellum contra adversarios suos per viam in qua miseris eos adorabunt te contra viam in qua civitas haec est quam elegisti et domus quam aedificavi nomini tuo
2CHR|6|35|ut exaudias de caelo preces eorum et obsecrationem et ulciscaris
2CHR|6|36|si autem et peccaverint tibi neque enim est homo qui non peccet et iratus fueris eis et tradideris hostibus et captivos eos duxerint in terram longinquam vel certe quae iuxta est
2CHR|6|37|et conversi corde suo in terra ad quam captivi ducti fuerant egerint paenitentiam et deprecati te fuerint in terra captivitatis suae dicentes peccavimus inique fecimus iniuste egimus
2CHR|6|38|et reversi fuerint ad te in toto corde suo et in tota anima sua in terra captivitatis suae ad quam ducti sunt adorabunt te contra viam terrae suae quam dedisti patribus eorum et urbis quam elegisti et domus quam aedificavi nomini tuo
2CHR|6|39|ut exaudias de caelo hoc est de firmo habitaculo tuo preces eorum et facias iudicium et dimittas populo tuo quamvis peccatori
2CHR|6|40|tu es enim Deus meus aperiantur quaeso oculi tui et aures tuae intentae sint ad orationem quae fit in loco isto
2CHR|6|41|nunc igitur consurge Domine Deus in requiem tuam tu et arca fortitudinis tuae sacerdotes tui Domine Deus induantur salute et sancti tui laetentur in bonis
2CHR|6|42|Domine Deus ne averseris faciem christi tui memento misericordiarum David servi tui
2CHR|7|1|cumque conplesset Salomon fundens preces ignis descendit de caelo et devoravit holocausta et victimas et maiestas Domini implevit domum
2CHR|7|2|nec poterant sacerdotes ingredi templum Domini eo quod implesset maiestas Domini templum Domini
2CHR|7|3|sed et omnes filii Israhel videbant descendentem ignem et gloriam Domini super domum et corruentes proni in terram super pavimentum stratum lapide adoraverunt et laudaverunt Dominum quoniam bonus quoniam in aeternum misericordia eius
2CHR|7|4|rex autem et omnis populus immolabant victimas coram Domino
2CHR|7|5|mactavit igitur rex Salomon hostias boum viginti duo milia arietum centum viginti milia et dedicavit domum Dei rex et universus populus
2CHR|7|6|sacerdotes autem stabant in officiis suis et Levitae in organis carminum Domini quae fecit David rex ad laudandum Dominum quoniam in aeternum misericordia eius hymnos David canentes per manus suas porro sacerdotes canebant tubis ante eos cunctusque Israhel stabat
2CHR|7|7|sanctificavit quoque Salomon medium atrii ante templum Domini obtulerat enim ibi holocausta et adipes pacificorum quia altare aeneum quod fecerat non poterat sustinere holocausta et sacrificia et adipes
2CHR|7|8|fecit ergo Salomon sollemnitatem in tempore illo septem diebus et omnis Israhel cum eo ecclesia magna valde ab introitu Emath usque ad torrentem Aegypti
2CHR|7|9|fecitque die octavo collectam eo quod dedicasset altare septem diebus et sollemnitatem celebrasset diebus septem
2CHR|7|10|igitur in die vicesimo tertio mensis septimi dimisit populos ad tabernacula sua laetantes atque gaudentes super bono quod fecerat Dominus David et Salomoni et Israhel populo suo
2CHR|7|11|conplevitque Salomon domum Domini et domum regis et omnia quae disposuerat in corde suo ut faceret in domo Domini et in domo sua et prosperatus est
2CHR|7|12|apparuit autem ei Dominus nocte et ait audivi orationem tuam et elegi locum istum mihi in domum sacrificii
2CHR|7|13|si clausero caelum et pluvia non fluxerit et mandavero et praecepero lucustae ut devoret terram et misero pestilentiam in populum meum
2CHR|7|14|conversus autem populus meus super quos invocatum est nomen meum deprecatus me fuerit et exquisierit faciem meam et egerit paenitentiam a viis suis pessimis et ego exaudiam de caelo et propitius ero peccatis eorum et sanabo terram eorum
2CHR|7|15|oculi quoque mei erunt aperti et aures meae erectae ad orationem eius qui in loco isto oraverit
2CHR|7|16|elegi enim et sanctificavi locum istum ut sit nomen meum ibi in sempiternum et permaneant oculi mei et cor meum ibi cunctis diebus
2CHR|7|17|tu quoque si ambulaveris coram me sicut ambulavit David pater tuus et feceris iuxta omnia quae praecepi tibi et iustitias meas iudiciaque servaveris
2CHR|7|18|suscitabo thronum regni tui sicut pollicitus sum David patri tuo dicens non auferetur de stirpe tua vir qui sit princeps in Israhel
2CHR|7|19|si autem aversi fueritis et dereliqueritis iustitias meas et praecepta mea quae proposui vobis et abeuntes servieritis diis alienis et adoraveritis eos
2CHR|7|20|evellam vos de terra mea quam dedi vobis et domum hanc quam sanctificavi nomini meo proiciam a facie mea et tradam eam in parabolam et in exemplum cunctis populis
2CHR|7|21|et domus ista erit in proverbium universis transeuntibus et dicent stupentes quare fecit Dominus sic terrae huic et domui huic
2CHR|7|22|respondebuntque quia dereliquerunt Dominum Deum patrum suorum qui eduxit eos de terra Aegypti et adprehenderunt deos alienos et adoraverunt eos atque coluerunt idcirco venerunt super eos universa haec mala
2CHR|8|1|expletis autem viginti annis postquam aedificavit Salomon domum Domini et domum suam
2CHR|8|2|civitates quas dederat Hiram Salomoni aedificavit et habitare ibi fecit filios Israhel
2CHR|8|3|abiit quoque in Emath Suba et obtinuit eam
2CHR|8|4|et aedificavit Palmyram in deserto et alias civitates munitissimas aedificavit in Emath
2CHR|8|5|extruxitque Bethoron superiorem et Bethoron inferiorem civitates muratas habentes portas et vectes et seras
2CHR|8|6|Baalath etiam et omnes urbes firmissimas quae fuerunt Salomonis cunctasque urbes quadrigarum et urbes equitum omnia quae voluit Salomon atque disposuit aedificavit in Hierusalem et in Libano et in universa terra potestatis suae
2CHR|8|7|omnem populum qui derelictus fuerat de Hettheis et Amorreis et Ferezeis et Eveis et Iebuseis qui non erant de stirpe Israhel
2CHR|8|8|de filiis eorum et de posteris quos non interfecerant filii Israhel subiugavit Salomon in tributarios usque in diem hanc
2CHR|8|9|porro de filiis Israhel non posuit ut servirent operibus regis ipsi enim erant viri bellatores et duces primi et principes quadrigarum et equitum eius
2CHR|8|10|omnes autem principes exercitus regis Salomonis fuerunt ducenti quinquaginta qui erudiebant populum
2CHR|8|11|filiam vero Pharaonis transtulit de civitate David in domum quam aedificaverat ei dixit enim non habitabit uxor mea in domo David regis Israhel eo quod sanctificata sit quia ingressa est eam arca Domini
2CHR|8|12|tunc obtulit Salomon holocausta Domino super altare Domini quod extruxerat ante porticum
2CHR|8|13|ut per singulos dies offerretur in eo iuxta praeceptum Mosi in sabbatis et in kalendis et in festis diebus ter per annum id est in sollemnitate azymorum et in sollemnitate ebdomadarum et in sollemnitate tabernaculorum
2CHR|8|14|et constituit iuxta dispositionem David patris sui officia sacerdotum in ministeriis suis et Levitas in ordine suo ut laudarent et ministrarent coram sacerdotibus iuxta ritum uniuscuiusque diei et ianitores in divisionibus suis per portam et portam sic enim praeceperat David homo Dei
2CHR|8|15|nec praetergressi sunt de mandatis regis tam sacerdotes quam Levitae ex omnibus quae praeceperat et in custodiis thesaurorum
2CHR|8|16|omnes inpensas praeparatas habuit Salomon ex eo die quo fundavit domum Domini usque in diem quo perfecit eam
2CHR|8|17|tunc abiit Salomon in Hesiongaber et in Ahilath ad oram maris Rubri quae est in terra Edom
2CHR|8|18|misit autem ei Hiram per manum servorum suorum naves et nautas gnaros maris et abierunt cum servis Salomonis in Ophir tuleruntque inde quadringenta quinquaginta talenta auri et adtulerunt ad regem Salomonem
2CHR|9|1|regina quoque Saba cum audisset famam Salomonis venit ut temptaret eum enigmatibus in Hierusalem cum magnis opibus et camelis qui portabant aromata et auri plurimum gemmasque pretiosas cumque venisset ad Salomonem locuta est ei quaecumque erant in corde suo
2CHR|9|2|et exposuit ei Salomon omnia quae proposuerat nec quicquam fuit quod ei non perspicuum fecerit
2CHR|9|3|quod postquam vidit sapientiam scilicet Salomonis et domum quam aedificaverat
2CHR|9|4|necnon cibaria mensae eius et habitacula servorum et officia ministrorum eius et vestimenta eorum pincernas quoque et vestes eorum et victimas quas immolabat in domo Domini non erat prae stupore ultra in ea spiritus
2CHR|9|5|dixitque ad regem verus sermo quem audieram in terra mea de virtutibus et sapientia tua
2CHR|9|6|non credebam narrantibus donec ipsa venissem et vidissent oculi mei et probassem vix medietatem mihi sapientiae tuae fuisse narratam vicisti famam virtutibus tuis
2CHR|9|7|beati viri tui et beati servi tui hii qui adsistunt coram te in omni tempore et audiunt sapientiam tuam
2CHR|9|8|sit Dominus Deus tuus benedictus qui voluit te ordinare super thronum suum regem Domini Dei tui quia diligit Deus Israhel et vult servare eum in aeternum idcirco posuit te super eum regem ut facias iudicia atque iustitiam
2CHR|9|9|dedit autem regi centum viginti talenta auri et aromata multa nimis et gemmas pretiosissimas non fuerunt aromata talia ut haec quae dedit regina Saba regi Salomoni
2CHR|9|10|sed et servi Hiram cum servis Salomonis adtulerunt aurum de Ophir et ligna thyina et gemmas pretiosissimas
2CHR|9|11|de quibus fecit rex de lignis scilicet thyinis gradus in domo Domini et in domo regia citharas quoque et psalteria cantoribus numquam visa sunt in terra Iuda ligna talia
2CHR|9|12|rex autem Salomon dedit reginae Saba cuncta quae voluit et quae postulavit multo plura quam adtulerat ad eum quae reversa abiit in terram suam cum servis suis
2CHR|9|13|erat autem pondus auri quod adferebatur Salomoni per annos singulos sescenta sexaginta sex talenta auri
2CHR|9|14|excepta ea summa quam legati diversarum gentium et negotiatores adferre consueverant omnesque reges Arabiae et satrapae terrarum qui conportabant aurum et argentum Salomoni
2CHR|9|15|fecit igitur rex Salomon ducentas hastas aureas de summa sescentorum aureorum qui in hastis singulis expendebantur
2CHR|9|16|trecenta quoque scuta aurea trecentorum aureorum quibus tegebantur scuta singula posuitque ea rex in armamentario quod erat consitum nemore
2CHR|9|17|fecit quoque rex solium eburneum grande et vestivit illud auro mundissimo
2CHR|9|18|sexque gradus quibus ascendebatur ad solium et scabillum aureum et brachiola duo altrinsecus et duos leones stantes iuxta brachiola
2CHR|9|19|sed et alios duodecim leunculos stantes super sex gradus ex utraque parte non fuit tale solium in universis regnis
2CHR|9|20|omnia quoque vasa convivii regis erant aurea et vasa domus saltus Libani ex auro purissimo argentum enim in diebus illis pro nihilo reputabatur
2CHR|9|21|siquidem naves regis ibant in Tharsis cum servis Hiram semel in annis tribus et deferebant inde aurum et argentum et ebur et simias et pavos
2CHR|9|22|magnificatus est igitur Salomon super omnes reges terrae divitiis et gloria
2CHR|9|23|omnesque reges terrarum desiderabant faciem videre Salomonis ut audirent sapientiam quam dederat Deus in corde eius
2CHR|9|24|et deferebant ei munera vasa argentea et aurea et vestes et arma et aromata equos et mulos per singulos annos
2CHR|9|25|habuit quoque Salomon quadraginta milia equorum in stabulis et curruum equitumque duodecim milia constituitque eos in urbibus quadrigarum et ubi erat rex in Hierusalem
2CHR|9|26|exercuit etiam potestatem super cunctos reges a fluvio Eufraten usque ad terram Philisthinorum id est usque ad terminos Aegypti
2CHR|9|27|tantamque copiam praebuit argenti in Hierusalem quasi lapidum et cedrorum tantam multitudinem velut sycaminorum quae gignuntur in campestribus
2CHR|9|28|adducebantur autem ei equi de Aegypto cunctisque regionibus
2CHR|9|29|reliqua vero operum Salomonis priorum et novissimorum scripta sunt in verbis Nathan prophetae et in libris Ahiae Silonitis in visione quoque Iaddo videntis contra Hieroboam filium Nabath
2CHR|9|30|regnavit autem Salomon in Hierusalem super omnem Israhel quadraginta annis
2CHR|9|31|dormivitque cum patribus suis et sepelierunt eum in civitate David regnavitque pro eo Roboam filius eius
2CHR|10|1|profectus est autem Roboam in Sychem illuc enim cunctus Israhel convenerat ut constituerent eum regem
2CHR|10|2|quod cum audisset Hieroboam filius Nabath qui erat in Aegypto fugerat quippe illuc ante Salomonem statim reversus est
2CHR|10|3|vocaveruntque eum et venit cum universo Israhel et locuti sunt ad Roboam dicentes
2CHR|10|4|pater tuus durissimo iugo nos pressit tu leviora impera patre tuo qui nobis gravem inposuit servitutem et paululum de onere subleva ut serviamus tibi
2CHR|10|5|qui ait post tres dies revertimini ad me cumque abisset populus
2CHR|10|6|iniit consilium cum senibus qui steterant coram patre eius Salomone dum adviveret dicens quid datis consilii ut respondeam populo
2CHR|10|7|qui dixerunt ei si placueris populo huic et lenieris eos verbis clementibus servient tibi omni tempore
2CHR|10|8|at ille reliquit consilium senum et cum iuvenibus tractare coepit qui cum eo nutriti fuerant et erant in comitatu illius
2CHR|10|9|dixitque ad eos quid vobis videtur vel respondere quid debeo populo huic qui dixit mihi subleva iugum quod inposuit nobis pater tuus
2CHR|10|10|at illi responderunt ut iuvenes et nutriti cum eo in deliciis atque dixerunt sic loqueris populo qui dixit tibi pater tuus adgravavit iugum nostrum tu subleva et sic respondebis eis minimus digitus meus grossior est lumbis patris mei
2CHR|10|11|pater meus inposuit vobis iugum grave et ego maius pondus adponam pater meus cecidit vos flagellis ego vero caedam scorpionibus
2CHR|10|12|venit ergo Hieroboam et universus populus ad Roboam die tertio sicut praeceperat eis
2CHR|10|13|responditque rex dura derelicto consilio seniorum
2CHR|10|14|locutusque est iuxta iuvenum voluntatem pater meus grave vobis inposuit iugum quod ego gravius faciam pater meus cecidit vos flagellis ego vero caedam scorpionibus
2CHR|10|15|et non adquievit populi precibus erat enim voluntatis Dei ut conpleretur sermo eius quem locutus fuerat per manum Ahiae Silonitis ad Hieroboam filium Nabath
2CHR|10|16|populus autem universus rege duriora dicente sic locutus est ad eum non est nobis pars in David neque hereditas in filio Isai revertere in tabernacula tua Israhel tu autem pasce domum tuam David et abiit Israhel in tabernacula sua
2CHR|10|17|super filios autem Israhel qui habitabant in civitatibus Iuda regnavit Roboam
2CHR|10|18|misitque rex Roboam Aduram qui praeerat tributis et lapidaverunt eum filii Israhel et mortuus est porro rex Roboam currum festinavit ascendere et fugit in Hierusalem
2CHR|10|19|recessitque Israhel a domo David usque ad diem hanc
2CHR|11|1|venit autem Roboam in Hierusalem et convocavit universam domum Iuda et Beniamin in centum octoginta milibus electorum atque bellantium ut dimicaret contra Israhel et converteret ad se regnum suum
2CHR|11|2|factusque est sermo Domini ad Semeiam hominem Dei dicens
2CHR|11|3|loquere ad Roboam filium Salomonis regem Iuda et ad universum Israhel qui est in Iuda et Beniamin
2CHR|11|4|haec dicit Dominus non ascendetis neque pugnabitis contra fratres vestros revertatur unusquisque in domum suam quia mea hoc gestum est voluntate qui cum audissent sermonem Domini reversi sunt nec perrexerunt contra Hieroboam
2CHR|11|5|habitavit autem Roboam in Hierusalem et aedificavit civitates muratas in Iuda
2CHR|11|6|extruxitque Bethleem et Aetham et Thecue
2CHR|11|7|Bethsur quoque et Soccho et Odollam
2CHR|11|8|necnon Geth et Maresa et Ziph
2CHR|11|9|sed et Aduram et Lachis et Azecha
2CHR|11|10|Saraa quoque et Ahilon et Hebron quae erant in Iuda et Beniamin civitates munitissimas
2CHR|11|11|cumque clausisset eas muris posuit in eis principes ciborumque horrea hoc est olei et vini
2CHR|11|12|sed et in singulis urbibus fecit armamentaria scutorum et hastarum firmavitque eas multa diligentia et imperavit super Iudam et Beniamin
2CHR|11|13|sacerdotes autem et Levitae qui erant in universo Israhel venerunt ad eum de cunctis sedibus suis
2CHR|11|14|relinquentes suburbana et possessiones suas et transeuntes ad Iudam et Hierusalem eo quod abiecisset eos Hieroboam et posteri eius ne sacerdotio Domini fungerentur
2CHR|11|15|qui constituit sibi sacerdotes excelsorum et daemonum vitulorumque quos fecerat
2CHR|11|16|sed et de cunctis tribubus Israhel quicumque dederant cor suum ut quaererent Dominum Deum Israhel venerunt Hierusalem ad immolandas victimas Domino Deo patrum suorum
2CHR|11|17|et roboraverunt regnum Iuda et confirmaverunt Roboam filium Salomonis per tres annos ambulaverunt enim in viis David et Salomonis annis tantum tribus
2CHR|11|18|duxit autem Roboam uxorem Maalath filiam Hierimuth filii David Abiail quoque filiam Heliab filii Isai
2CHR|11|19|quae peperit ei filios Ieus et Somoriam et Zoom
2CHR|11|20|post hanc quoque accepit Maacha filiam Absalom quae peperit ei Abia et Ethai et Ziza et Salumith
2CHR|11|21|amavit autem Roboam Maacha filiam Absalom super omnes uxores suas et concubinas nam uxores decem et octo duxerat concubinasque sexaginta et genuit viginti octo filios et sexaginta filias
2CHR|11|22|constituit vero in capite Abiam filium Maacha ducem super fratres suos ipsum enim regem facere cogitabat
2CHR|11|23|qui sapientior fuit et potentior super omnes filios eius et in cunctis finibus Iuda et Beniamin et in universis civitatibus muratis praebuitque eis escas plurimas et multas petivit uxores
2CHR|12|1|cumque roboratum fuisset regnum Roboam et confortatum dereliquit legem Domini et omnis Israhel cum eo
2CHR|12|2|anno autem quinto regni Roboam ascendit Sesac rex Aegypti in Hierusalem quia peccaverunt Domino
2CHR|12|3|cum mille ducentis curribus et sexaginta milibus equitum nec erat numerus vulgi quod venerat cum eo ex Aegypto Lybies scilicet et Trogoditae et Aethiopes
2CHR|12|4|cepitque civitates munitissimas in Iuda et venit usque Hierusalem
2CHR|12|5|Semeias autem propheta ingressus est ad Roboam et principes Iuda qui congregati fuerant in Hierusalem fugientes Sesac dixitque ad eos haec dicit Dominus vos reliquistis me et ego reliqui vos in manu Sesac
2CHR|12|6|consternatique principes Israhel et rex dixerunt iustus est Dominus
2CHR|12|7|cumque vidisset Dominus quod humiliati essent factus est sermo Domini ad Semeiam dicens quia humiliati sunt non disperdam eos daboque eis pauxillum auxilii et non stillabit furor meus super Hierusalem per manum Sesac
2CHR|12|8|verumtamen servient ei ut sciant distantiam servitutis meae et servitutis regni terrarum
2CHR|12|9|recessit itaque Sesac rex Aegypti ab Hierusalem sublatis thesauris domus Domini et domus regis omniaque secum tulit et clypeos aureos quos fecerat Salomon
2CHR|12|10|pro quibus fecit rex aeneos et tradidit illos principibus scutariorum qui custodiebant vestibulum palatii
2CHR|12|11|cumque introiret rex domum Domini veniebant scutarii et tollebant eos iterumque referebant ad armamentarium suum
2CHR|12|12|verumtamen quia humiliati sunt aversa est ab eis ira Domini nec deleti sunt penitus siquidem et in Iuda inventa sunt opera bona
2CHR|12|13|confortatus est igitur rex Roboam in Hierusalem atque regnavit quadraginta autem et unius anni erat cum regnare coepisset et decem septemque annis regnavit in Hierusalem urbe quam elegit Dominus ut confirmaret nomen suum ibi de cunctis tribubus Israhel nomenque matris eius Naama Ammanitis
2CHR|12|14|fecit autem malum et non praeparavit cor suum ut quaereret Dominum
2CHR|12|15|opera vero Roboam prima et novissima scripta sunt in libris Semeiae prophetae et Addo videntis et diligenter exposita pugnaveruntque adversum se Roboam et Hieroboam cunctis diebus
2CHR|12|16|et dormivit Roboam cum patribus suis sepultusque est in civitate David et regnavit Abia filius eius pro eo
2CHR|13|1|anno octavodecimo regis Hieroboam regnavit Abia super Iudam
2CHR|13|2|tribus annis regnavit in Hierusalem nomenque matris eius Michaia filia Urihel de Gabaa et erat bellum inter Abia et Hieroboam
2CHR|13|3|cumque inisset Abia certamen et haberet bellicosissimos viros et electorum quadringenta milia Hieroboam instruxit e contra aciem octingenta milia virorum qui et ipsi electi erant et ad bella fortissimi
2CHR|13|4|stetit igitur Abia super montem Someron qui erat in Ephraim et ait audi Hieroboam et omnis Israhel
2CHR|13|5|num ignoratis quod Dominus Deus Israhel dederit regnum David super Israhel in sempiternum ipsi et filiis eius pactum salis
2CHR|13|6|et surrexit Hieroboam filius Nabath servus Salomonis filii David et rebellavit contra dominum suum
2CHR|13|7|congregatique sunt ad eum viri vanissimi et filii Belial et praevaluerunt contra Roboam filium Salomonis porro Roboam erat rudis et corde pavido nec potuit resistere eis
2CHR|13|8|nunc ergo vos dicitis quod resistere possitis regno Domini quod possidet per filios David habetisque grandem populi multitudinem atque vitulos aureos quos fecit vobis Hieroboam in deos
2CHR|13|9|et eiecistis sacerdotes Domini filios Aaron atque Levitas et fecistis vobis sacerdotes sicut omnes populi terrarum quicumque venerit et initiaverit manum suam in tauro in bubus et in arietibus septem fit sacerdos eorum qui non sunt dii
2CHR|13|10|noster autem Dominus Deus est quem non relinquimus sacerdotesque ministrant Domino de filiis Aaron et Levitae sunt in ordine suo
2CHR|13|11|holocausta quoque offerunt Domino per singulos dies mane et vespere et thymiama iuxta legis praecepta confectum et proponuntur panes in mensa mundissima estque apud nos candelabrum aureum et lucernae eius ut accendantur semper ad vesperam nos quippe custodimus praecepta Domini Dei nostri quem vos reliquistis
2CHR|13|12|ergo in exercitu nostro dux Deus est et sacerdotes eius qui clangunt tubis et resonant contra vos filii Israhel nolite pugnare contra Dominum Deum patrum vestrorum quia non vobis expedit
2CHR|13|13|haec illo loquente Hieroboam retro moliebatur insidias cumque ex adverso hostium staret ignorantem Iudam suo ambiebat exercitu
2CHR|13|14|respiciensque Iudas vidit instare bellum ex adverso et post tergum et clamavit ad Dominum ac sacerdotes tubis canere coeperunt
2CHR|13|15|omnesque viri Iuda vociferati sunt et ecce illis clamantibus perterruit Deus Hieroboam et omnem Israhel qui stabat ex adverso Abia et Iuda
2CHR|13|16|fugeruntque filii Israhel Iudam et tradidit eos Deus in manu eorum
2CHR|13|17|percussit ergo eos Abia et populus eius plaga magna et corruerunt vulnerati ex Israhel quingenta milia virorum fortium
2CHR|13|18|humiliatique sunt filii Israhel in tempore illo et vehementissime confortati filii Iuda eo quod sperassent in Domino Deo patrum suorum
2CHR|13|19|persecutus est autem Abia fugientem Hieroboam et cepit civitates eius Bethel et filias eius et Hiesena cum filiabus suis Ephron quoque et filias eius
2CHR|13|20|nec valuit ultra resistere Hieroboam in diebus Abia quem percussit Dominus et mortuus est
2CHR|13|21|igitur Abia confortato imperio suo accepit uxores quattuordecim procreavitque viginti duos filios et sedecim filias
2CHR|13|22|reliqua autem sermonum Abia viarumque et operum eius scripta sunt diligentissime in libro prophetae Addo
2CHR|14|1|dormivit autem Abia cum patribus suis et sepelierunt eum in civitate David regnavitque Asa filius eius pro eo in cuius diebus quievit terra annis decem
2CHR|14|2|fecit autem Asa quod bonum et placitum erat in conspectu Dei sui et subvertit altaria peregrini cultus et excelsa
2CHR|14|3|et confregit statuas lucosque succidit
2CHR|14|4|ac praecepit Iudae ut quaereret Dominum Deum patrum suorum et faceret legem et universa mandata
2CHR|14|5|et abstulit e cunctis urbibus Iuda aras et fana et regnavit in pace
2CHR|14|6|aedificavit quoque urbes munitas in Iuda quia quietus erat et nulla temporibus eius bella surrexerant pacem Domino largiente
2CHR|14|7|dixit autem Iudae aedificemus civitates istas et vallemus muris et roboremus turribus et portis et seris donec a bellis quieta sunt omnia eo quod quaesierimus Dominum Deum patrum nostrorum et dederit nobis pacem per gyrum aedificaverunt igitur et nullum in extruendo inpedimentum fuit
2CHR|14|8|habuit autem Asa in exercitu suo portantium scuta et hastas de Iuda trecenta milia de Beniamin vero scutariorum et sagittariorum ducenta octoginta milia omnes isti viri fortissimi
2CHR|14|9|egressus est autem contra eos Zara Aethiops cum exercitu decies centena milia et curribus trecentis et venit usque Maresa
2CHR|14|10|porro Asa perrexit obviam et instruxit aciem ad bellum in valle Sephata quae est iuxta Maresa
2CHR|14|11|et invocavit Dominum Deum et ait Domine non est apud te ulla distantia utrum in paucis auxilieris an in pluribus adiuva nos Domine Deus noster in te enim et in tuo nomine habentes fiduciam venimus contra hanc multitudinem Domine Deus noster tu es non praevaleat contra te homo
2CHR|14|12|exterruit itaque Dominus Aethiopas coram Asa et Iuda fugeruntque Aethiopes
2CHR|14|13|et persecutus est eos Asa et populus qui cum eo erat usque Gerar et ruerunt Aethiopes usque ad internicionem quia Domino caedente contriti sunt et exercitu illius proeliante tulerunt ergo spolia multa
2CHR|14|14|et percusserunt omnes civitates per circuitum Gerare grandis quippe cunctos terror invaserat et diripuerunt urbes et multam praedam asportaverunt
2CHR|14|15|sed et caulas ovium destruentes tulerunt pecorum infinitam multitudinem et camelorum reversique sunt Hierusalem
2CHR|15|1|Azarias autem filius Oded facto in se spiritu Dei
2CHR|15|2|egressus est in occursum Asa et dixit ei audite me Asa et omnis Iuda et Beniamin Dominus vobiscum quia fuistis cum eo si quaesieritis eum invenietis si autem dereliqueritis derelinquet vos
2CHR|15|3|transibunt autem multi dies in Israhel absque Deo vero et absque sacerdote doctore et absque lege
2CHR|15|4|cumque reversi fuerint in angustia sua ad Dominum Deum Israhel et quaesierint eum repperient
2CHR|15|5|in tempore illo non erit pax egredienti et ingredienti sed terrores undique in cunctis habitatoribus terrarum
2CHR|15|6|pugnabit enim gens contra gentem et civitas contra civitatem quia Dominus conturbabit eos in omni angustia
2CHR|15|7|vos ergo confortamini et non dissolvantur manus vestrae erit enim merces operi vestro
2CHR|15|8|quod cum audisset Asa verba scilicet et prophetiam Oded prophetae confortatus est et abstulit idola de omni terra Iuda et Beniamin et ex urbibus quas ceperat montis Ephraim et dedicavit altare Domini quod erat ante porticum Domini
2CHR|15|9|congregavitque universum Iuda et Beniamin et advenas cum eis de Ephraim et de Manasse et de Symeon plures enim ad eum confugerant ex Israhel videntes quod Dominus Deus illius esset cum eo
2CHR|15|10|cumque venissent Hierusalem mense tertio anno quintodecimo regni Asa
2CHR|15|11|immolaverunt Domino in die illa de manubiis et praeda quam adduxerant boves septingentos et arietes septem milia
2CHR|15|12|et intravit ex more ad corroborandum foedus ut quaererent Dominum Deum patrum suorum in toto corde et in tota anima sua
2CHR|15|13|si quis autem inquit non quaesierit Dominum Deum Israhel moriatur a minimo usque ad maximum a viro usque ad mulierem
2CHR|15|14|iuraveruntque Domino voce magna in iubilo et in clangore tubae et in sonitu bucinarum
2CHR|15|15|omnes qui erant in Iuda cum execratione in omni enim corde suo iuraverunt et in tota voluntate quaesierunt eum et invenerunt praestititque eis Dominus requiem per circuitum
2CHR|15|16|sed et Maacham matrem Asa regis ex augusto deposuit imperio eo quod fecisset in luco simulacrum Priapi quod omne contrivit et in frusta comminuens conbusit in torrente Cedron
2CHR|15|17|excelsa autem derelicta sunt in Israhel attamen cor Asa erat perfectum cunctis diebus eius
2CHR|15|18|ea quae voverat pater suus et ipse intulit in domum Domini argentum et aurum vasorumque diversam supellectilem
2CHR|15|19|bellum vero non fuit usque ad tricesimum quintum annum regni Asa
2CHR|16|1|anno autem tricesimo sexto regni eius ascendit Baasa rex Israhel in Iudam et muro circumdabat Rama ut nullus tute posset egredi et ingredi de regno Asa
2CHR|16|2|protulit ergo Asa argentum et aurum de thesauris domus Domini et de thesauris regis misitque ad Benadad regem Syriae qui habitabat in Damasco dicens
2CHR|16|3|foedus inter me et te est pater quoque meus et pater tuus habuere concordiam quam ob rem misi tibi argentum et aurum ut rupto foedere quod habes cum Baasa rege Israhel facias eum a me recedere
2CHR|16|4|quo conperto Benadad misit principes exercituum suorum ad urbes Israhel qui percusserunt Ahion et Dan et Abelmaim et universas urbes muratas Nepthalim
2CHR|16|5|quod cum audisset Baasa desivit aedificare Rama et intermisit opus suum
2CHR|16|6|porro Asa rex adsumpsit universum Iudam et tulerunt lapides Rama et ligna quae aedificationi praeparaverat Baasa aedificavitque ex eis Gabaa et Maspha
2CHR|16|7|in tempore illo venit Anani propheta ad Asam regem Iuda et dixit ei quia habuisti fiduciam in rege Syriae et non in Domino Deo tuo idcirco evasit Syriae regis exercitus de manu tua
2CHR|16|8|nonne Aethiopes et Lybies multo plures erant quadrigis et equitibus et multitudine nimia quos cum Domino credidisses tradidit in manu tua
2CHR|16|9|oculi enim eius contemplantur universam terram et praebent fortitudinem his qui corde perfecto credunt in eum stulte igitur egisti et propter hoc ex praesenti tempore contra te bella consurgent
2CHR|16|10|iratusque Asa adversus videntem iussit eum mitti in nervum valde quippe super hoc fuerat indignatus et interfecit de populo in tempore illo plurimos
2CHR|16|11|opera autem Asa prima et novissima scripta sunt in libro regum Iuda et Israhel
2CHR|16|12|aegrotavit etiam Asa anno tricesimo nono regni sui dolore pedum vehementissimo et nec in infirmitate sua quaesivit Dominum sed magis in medicorum arte confisus est
2CHR|16|13|dormivitque cum patribus suis et mortuus est anno quadragesimo primo regni sui
2CHR|16|14|et sepelierunt eum in sepulchro suo quod foderat sibi in civitate David posueruntque eum super lectulum suum plenum aromatibus et unguentis meretriciis quae erant pigmentariorum arte confecta et conbuserunt super eum ambitione nimia
2CHR|17|1|regnavit autem Iosaphat filius eius pro eo et invaluit contra Israhel
2CHR|17|2|constituitque militum numeros in cunctis urbibus Iudae quae erant vallatae muris praesidiaque disposuit in terra Iuda et in civitatibus Ephraim quas ceperat Asa pater eius
2CHR|17|3|et fuit Dominus cum Iosaphat quia ambulavit in viis David patris sui primis et non speravit in Baalim
2CHR|17|4|sed in Deo patris sui et perrexit in praeceptis illius et non iuxta peccata Israhel
2CHR|17|5|confirmavitque Dominus regnum in manu eius et dedit omnis Iuda munera Iosaphat factaeque sunt ei infinitae divitiae et multa gloria
2CHR|17|6|cumque sumpsisset cor eius audaciam propter vias Domini etiam excelsa et lucos de Iuda abstulit
2CHR|17|7|tertio autem anno regni sui misit de principibus suis Benail et Obdiam et Zacchariam et Nathanahel et Micheam ut docerent in civitatibus Iuda
2CHR|17|8|et cum eis Levitas Semeiam et Nathaniam et Zabadiam Asahel quoque et Semiramoth et Ionathan Adoniam et Tobiam et Tobadoniam Levitas et cum eis Elisama et Ioram sacerdotes
2CHR|17|9|docebantque in Iuda habentes librum legis Domini et circuibant cunctas urbes Iuda atque erudiebant populum
2CHR|17|10|itaque factus est pavor Domini super omnia regna terrarum quae erant per gyrum Iuda nec audebant bellare contra Iosaphat
2CHR|17|11|sed et Philisthei Iosaphat munera deferebant et vectigal argenti Arabes quoque adducebant pecora arietum septem milia septingentos et hircos totidem
2CHR|17|12|crevit ergo Iosaphat et magnificatus est usque in sublime atque aedificavit in Iuda domos ad instar turrium urbesque muratas
2CHR|17|13|et multa opera patravit in urbibus Iuda viri quoque bellatores et robusti erant in Hierusalem
2CHR|17|14|quorum iste numerus per domos atque familias singulorum in Iuda principes exercitus Ednas dux et cum eo robustissimorum trecenta milia
2CHR|17|15|post hunc Iohanan princeps et cum eo ducenta octoginta milia
2CHR|17|16|post istum quoque Amasias filius Zechri consecratus Domino et cum eo ducenta milia virorum fortium
2CHR|17|17|hunc sequebatur robustus ad proelia Heliada et cum eo tenentium arcum et clypeum ducenta milia
2CHR|17|18|post istum etiam Iozabath et cum eo centum octoginta milia expeditorum militum
2CHR|17|19|hii omnes erant ad manum regis exceptis aliis quos posuerat in urbibus muratis et in universo Iuda
2CHR|18|1|fuit ergo Iosaphat dives et inclitus multum et adfinitate coniunctus est Ahab
2CHR|18|2|descenditque post annos ad eum in Samariam ad cuius adventum mactavit Ahab arietes et boves plurimos et populo qui venerat cum eo persuasitque illi ut ascenderet in Ramoth Galaad
2CHR|18|3|dixitque Ahab rex Israhel ad Iosaphat regem Iuda veni mecum in Ramoth Galaad cui ille respondit ut ego et tu sicut populus tuus sic et populus meus tecumque erimus in bello
2CHR|18|4|dixitque Iosaphat ad regem Israhel consule obsecro inpraesentiarum sermonem Domini
2CHR|18|5|congregavitque rex Israhel prophetarum quadringentos viros et dixit ad eos in Ramoth Galaad ad bellandum ire debemus an quiescere at illi ascende inquiunt et tradet Deus in manu regis
2CHR|18|6|dixitque Iosaphat numquid non est hic prophetes Domini ut ab illo etiam requiramus
2CHR|18|7|et ait rex Israhel ad Iosaphat est vir unus a quo possumus quaerere Domini voluntatem sed ego odi eum quia non prophetat mihi bonum sed malum omni tempore est autem Micheas filius Iembla dixitque Iosaphat ne loquaris rex hoc modo
2CHR|18|8|vocavit ergo rex Israhel unum de eunuchis et dixit ei voca cito Micheam filium Iembla
2CHR|18|9|porro rex Israhel et Iosaphat rex Iuda uterque sedebant in solio suo vestiti cultu regio sedebant autem in area iuxta portam Samariae omnesque prophetae vaticinabantur coram eis
2CHR|18|10|Sedecias vero filius Chanana fecit sibi cornua ferrea et ait haec dicit Dominus his ventilabis Syriam donec conteras eam
2CHR|18|11|omnesque prophetae similiter prophetabant atque dicebant ascende in Ramoth Galaad et prosperaberis et tradet eos Dominus in manu regis
2CHR|18|12|nuntius autem qui ierat ad vocandum Micheam ait illi en verba omnium prophetarum uno ore bona regi adnuntiant quaeso ergo te ut et sermo tuus ab eis non dissentiat loquarisque prospera
2CHR|18|13|cui respondit Micheas vivit Dominus quia quodcumque dixerit Deus meus hoc loquar
2CHR|18|14|venit ergo ad regem cui rex ait Michea ire debemus in Ramoth Galaad ad bellandum an quiescere cui ille respondit ascendite cuncta enim prospera evenient et tradentur hostes in manus vestras
2CHR|18|15|dixitque rex iterum atque iterum te adiuro ut non mihi loquaris nisi quod verum est in nomine Domini
2CHR|18|16|at ille ait vidi universum Israhel dispersum in montibus sicut oves absque pastore et dixit Dominus non habent isti dominos revertatur unusquisque ad domum suam in pace
2CHR|18|17|et ait rex Israhel ad Iosaphat nonne dixi tibi quod non prophetaret iste mihi quicquam boni sed ea quae mala sunt
2CHR|18|18|at ille idcirco ait audite verbum Domini vidi Dominum sedentem in solio suo et omnem exercitum caeli adsistentem ei a dextris et sinistris
2CHR|18|19|et dixit Dominus quis decipiet Ahab regem Israhel ut ascendat et corruat in Ramoth Galaad cumque diceret unus hoc modo et alter alio
2CHR|18|20|processit spiritus et stetit coram Domino et ait ego decipiam eum cui Dominus in quo inquit decipies
2CHR|18|21|at ille respondit egrediar et ero spiritus mendax in ore omnium prophetarum eius dixitque Dominus decipies et praevalebis egredere et fac ita
2CHR|18|22|nunc igitur ecce dedit Dominus spiritum mendacii in ore omnium prophetarum tuorum et Dominus locutus est de te mala
2CHR|18|23|accessit autem Sedecias filius Chanana et percussit Micheae maxillam et ait per quam viam transivit spiritus Domini a me ut loqueretur tibi
2CHR|18|24|dixitque Micheas tu ipse videbis in die illo quando ingressus fueris cubiculum de cubiculo ut abscondaris
2CHR|18|25|praecepit autem rex Israhel dicens tollite Micheam et ducite eum ad Amon principem civitatis et ad Ioas filium Ammelech
2CHR|18|26|et dicetis haec dicit rex mittite hunc in carcerem et date ei panis modicum et aquae pauxillum donec revertar in pace
2CHR|18|27|dixitque Micheas si reversus fueris in pace non est locutus Dominus in me et ait audite populi omnes
2CHR|18|28|igitur ascenderunt rex Israhel et Iosaphat rex Iuda in Ramoth Galaad
2CHR|18|29|dixitque rex Israhel ad Iosaphat mutabo habitum et sic ad pugnandum vadam tu autem induere vestibus tuis mutatoque rex Israhel habitu venit ad bellum
2CHR|18|30|rex autem Syriae praeceperat ducibus equitatus sui dicens ne pugnetis contra minimum aut contra maximum nisi contra solum regem Israhel
2CHR|18|31|itaque cum vidissent principes equitatus Iosaphat dixerunt rex Israhel iste est et circumdederunt eum dimicantes at ille clamavit ad Dominum et auxiliatus est ei atque avertit eos ab illo
2CHR|18|32|cum enim vidissent duces equitatus quod non esset rex Israhel reliquerunt eum
2CHR|18|33|accidit autem ut unus e populo sagittam in incertum iaceret et percuteret regem Israhel inter cervicem et scapulas at ille aurigae suo ait converte manum tuam et educ me de acie quia vulneratus sum
2CHR|18|34|et finita est pugna in die illo porro rex Israhel stabat in curru suo contra Syros usque ad vesperam et mortuus est occidente sole
2CHR|19|1|reversus est autem Iosaphat rex Iuda domum suam pacifice in Hierusalem
2CHR|19|2|cui occurrit Hieu filius Anani videns et ait ad eum impio praebes auxilium et his qui oderunt Dominum amicitia iungeris et idcirco iram quidem Domini merebaris
2CHR|19|3|sed bona opera inventa sunt in te eo quod abstuleris lucos de terra Iuda et praeparaveris cor tuum ut requireres Dominum
2CHR|19|4|habitavit ergo Iosaphat in Hierusalem rursumque egressus est ad populum de Bersabee usque ad montem Ephraim et revocavit eos ad Dominum Deum patrum suorum
2CHR|19|5|constituitque iudices terrae in cunctis civitatibus Iuda munitis per singula loca
2CHR|19|6|et praecipiens iudicibus videte ait quid faciatis non enim hominis exercetis iudicium sed Domini et quodcumque iudicaveritis in vos redundabit
2CHR|19|7|sit timor Domini vobiscum et cum diligentia cuncta facite non est enim apud Dominum Deum nostrum iniquitas nec personarum acceptio nec cupido munerum
2CHR|19|8|in Hierusalem quoque constituit Iosaphat Levitas et sacerdotes et principes familiarum ex Israhel ut iudicium et causam Domini iudicarent habitatoribus eius
2CHR|19|9|praecepitque eis dicens sic agetis in timore Dei fideliter et corde perfecto
2CHR|19|10|omnem causam quae venerit ad vos fratrum vestrorum qui habitant in urbibus suis inter cognationem et cognationem ubicumque quaestio est de lege de mandato de caerimoniis de iustificationibus ostendite eis ut non peccent in Dominum et ne veniat ira super vos et super fratres vestros sic ergo agetis et non peccabitis
2CHR|19|11|Amarias autem sacerdos et pontifex vester in his quae ad Dominum pertinent praesidebit porro Zabadias filius Ismahel qui est dux in domo Iuda super ea opera erit quae ad regis officium pertinent habetisque magistros Levitas coram vobis confortamini et agite diligenter et erit Dominus cum bonis
2CHR|20|1|post haec congregati sunt filii Moab et filii Ammon et cum eis de Ammanitis ad Iosaphat ut pugnarent contra eum
2CHR|20|2|veneruntque nuntii et indicaverunt Iosaphat dicentes venit contra te multitudo magna de his locis quae trans mare sunt et de Syria et ecce consistunt in Asasonthamar quae est Engaddi
2CHR|20|3|Iosaphat autem timore perterritus totum se contulit ad rogandum Dominum et praedicavit ieiunium universo Iuda
2CHR|20|4|congregatusque Iudas ad precandum Dominum sed et omnes de urbibus suis venerunt ad obsecrandum eum
2CHR|20|5|cumque stetisset Iosaphat in medio coetu Iudae et Hierusalem in domo Domini ante atrium novum
2CHR|20|6|ait Domine Deus patrum nostrorum tu es Deus in caelo et dominaris cunctis regnis gentium in manu tua est fortitudo et potentia nec quisquam tibi potest resistere
2CHR|20|7|nonne tu Deus noster interfecisti omnes habitatores terrae huius coram populo tuo Israhel et dedisti eam semini Abraham amici tui in sempiternum
2CHR|20|8|habitaveruntque in ea et extruxerunt in illa sanctuarium nomini tuo dicentes
2CHR|20|9|si inruerint super nos mala gladius iudicii pestilentia et fames stabimus coram domo hac in conspectu tuo in qua invocatum est nomen tuum et clamabimus ad te in tribulationibus nostris et exaudies salvosque facies
2CHR|20|10|nunc igitur ecce filii Ammon et Moab et mons Seir per quos non concessisti Israheli ut transirent quando egrediebantur de Aegypto sed declinaverunt ab eis et non interfecerunt illos
2CHR|20|11|e contrario agunt et nituntur eicere nos de possessione quam tradidisti nobis
2CHR|20|12|Deus noster ergo non iudicabis eos in nobis quidem non tanta est fortitudo ut possimus huic multitudini resistere quae inruit super nos sed cum ignoremus quid agere debeamus hoc solum habemus residui ut oculos nostros dirigamus ad te
2CHR|20|13|omnis vero Iuda stabat coram Domino cum parvulis et uxoribus et liberis suis
2CHR|20|14|erat autem Hiazihel filius Zacchariae filii Banaiae filii Hiehihel filii Mathaniae Levites de filiis Asaph super quem factus est spiritus Domini in medio turbae
2CHR|20|15|et ait adtendite omnis Iuda et qui habitatis Hierusalem et tu rex Iosaphat haec dicit Dominus vobis nolite timere nec paveatis hanc multitudinem non est enim vestra pugna sed Dei
2CHR|20|16|cras descendetis contra eos ascensuri enim sunt per clivum nomine Sis et invenietis illos in summitate torrentis qui est contra solitudinem Hieruhel
2CHR|20|17|non eritis vos qui dimicabitis sed tantummodo confidenter state et videbitis auxilium Domini super vos o Iuda et Hierusalem nolite timere nec paveatis cras egredimini contra eos et Dominus erit vobiscum
2CHR|20|18|Iosaphat ergo et Iuda et omnes habitatores Hierusalem ceciderunt proni in terram coram Domino et adoraverunt eum
2CHR|20|19|porro Levitae de filiis Caath et de filiis Core laudabant Dominum Deum Israhel voce magna in excelsum
2CHR|20|20|cumque mane surrexissent egressi sunt per desertum Thecuae profectisque eis stans Iosaphat in medio eorum dixit audite me Iuda et omnes habitatores Hierusalem credite in Domino Deo vestro et securi eritis credite prophetis eius et cuncta evenient prospera
2CHR|20|21|deditque consilium populo et statuit cantores Domini ut laudarent eum in turmis suis et antecederent exercitum ac voce consona dicerent confitemini Domino quoniam in aeternum misericordia eius
2CHR|20|22|cumque coepissent laudes canere vertit Dominus insidias eorum in semet ipsos filiorum scilicet Ammon et Moab et montis Seir qui egressi fuerant ut pugnarent contra Iudam et percussi sunt
2CHR|20|23|namque filii Ammon et Moab consurrexerunt adversum habitatores montis Seir ut interficerent et delerent eos cumque hoc opere perpetrassent etiam in semet ipsos versi mutuis concidere vulneribus
2CHR|20|24|porro Iudas cum venisset ad speculam quae respicit solitudinem vidit procul omnem late regionem plenam cadaveribus nec superesse quemquam qui necem potuisset evadere
2CHR|20|25|venit ergo Iosaphat et omnis populus cum eo ad detrahenda spolia mortuorum inveneruntque inter cadavera variam supellectilem vestes quoque et vasa pretiosissima et diripuerunt ita ut omnia portare non possent nec per tres dies spolia auferre pro praedae magnitudine
2CHR|20|26|die autem quarto congregati sunt in valle Benedictionis etenim quoniam ibi benedixerant Domino vocaverunt locum illum vallis Benedictionis usque in praesentem diem
2CHR|20|27|reversusque est omnis vir Iuda et habitatores Hierusalem et Iosaphat ante eos in Hierusalem cum laetitia magna eo quod dedisset eis Dominus gaudium de inimicis suis
2CHR|20|28|ingressique sunt Hierusalem cum psalteriis et citharis et tubis in domum Domini
2CHR|20|29|inruit autem pavor Domini super universa regna terrarum cum audissent quod pugnasset Dominus contra inimicos Israhel
2CHR|20|30|quievitque regnum Iosaphat et praebuit ei Deus pacem per circuitum
2CHR|20|31|regnavit igitur Iosaphat super Iudam et erat triginta quinque annorum cum regnare coepisset viginti autem et quinque annis regnavit in Hierusalem nomen matris eius Azuba filia Selachi
2CHR|20|32|et ambulavit in via patris sui Asa nec declinavit ab ea faciens quae placita erant coram Domino
2CHR|20|33|verumtamen excelsa non abstulit et adhuc populus non direxerat cor suum ad Dominum Deum patrum suorum
2CHR|20|34|reliqua autem gestorum Iosaphat priorum et novissimorum scripta sunt in verbis Hieu filii Anani quae digessit in libro regum Israhel
2CHR|20|35|post haec iniit amicitias Iosaphat rex Iuda cum Ochozia rege Israhel cuius opera fuerunt impiissima
2CHR|20|36|et particeps fuit ut facerent naves quae irent in Tharsis feceruntque classem in Asiongaber
2CHR|20|37|prophetavit autem Eliezer filius Dodoau de Maresa ad Iosaphat dicens quia habuisti foedus cum Ochozia percussit Dominus opera tua contritaeque sunt naves nec potuerunt ire in Tharsis
2CHR|21|1|dormivit autem Iosaphat cum patribus suis et sepultus est cum eis in civitate David regnavitque Ioram filius eius pro eo
2CHR|21|2|qui habuit fratres filios Iosaphat Azariam et Hiahihel et Zacchariam et Azariam et Michahel et Saphatiam omnes hii filii Iosaphat regis Israhel
2CHR|21|3|deditque eis pater suus multa munera argenti et auri et pensitationes cum civitatibus munitissimis in Iuda regnum autem tradidit Ioram eo quod esset primogenitus
2CHR|21|4|surrexit ergo Ioram super regnum patris sui cumque se confirmasset occidit omnes fratres suos gladio et quosdam de principibus Israhel
2CHR|21|5|triginta duo annorum erat Ioram cum regnare coepisset et octo annis regnavit in Hierusalem
2CHR|21|6|ambulavitque in viis regum Israhel sicut egerat domus Ahab filia quippe Ahab erat uxor eius et fecit malum in conspectu Domini
2CHR|21|7|noluit autem Dominus disperdere domum David propter pactum quod inierat cum eo et quia promiserat ut daret illi lucernam et filiis eius omni tempore
2CHR|21|8|in diebus illis rebellavit Edom ne esset subditus Iudae et constituit sibi regem
2CHR|21|9|cumque transisset Ioram cum principibus suis et cuncto equitatu qui erat secum surrexit nocte et percussit Edom qui se circumdederat et omnes duces equitatus eius
2CHR|21|10|attamen rebellavit Edom ne esset sub dicione Iuda usque ad hanc diem eo tempore et Lobna recessit ne esset sub manu illius dereliquerat enim Dominum Deum patrum suorum
2CHR|21|11|insuper et excelsa fabricatus est in urbibus Iuda et fornicari fecit habitatores Hierusalem et praevaricari Iudam
2CHR|21|12|adlatae sunt autem ei litterae ab Helia propheta in quibus scriptum erat haec dicit Dominus Deus David patris tui quoniam non ambulasti in viis Iosaphat patris tui et in viis Asa regis Iuda
2CHR|21|13|sed incessisti per iter regum Israhel et fornicari fecisti Iudam et habitatores Hierusalem imitatus fornicationem domus Ahab insuper et fratres tuos domum patris tui meliores te occidisti
2CHR|21|14|ecce Dominus percutiet te plaga magna cum populo tuo et filiis et uxoribus tuis universaque substantia tua
2CHR|21|15|tu autem aegrotabis pessimo languore uteri donec egrediantur vitalia tua paulatim per dies singulos
2CHR|21|16|suscitavit ergo Dominus contra Ioram spiritum Philisthinorum et Arabum qui confines sunt Aethiopibus
2CHR|21|17|et ascenderunt in terram Iuda et vastaverunt eam diripueruntque cunctam substantiam quae inventa est in domo regis insuper et filios eius et uxores nec remansit ei filius nisi Ioachaz qui minimus natu erat
2CHR|21|18|et super haec omnia percussit eum Dominus alvi languore insanabili
2CHR|21|19|cumque diei succederet dies et temporum spatia volverentur duorum annorum expletus est circulus et sic longa consumptus tabe ita ut egereret etiam viscera sua languore pariter et vita caruit mortuusque est in infirmitate pessima et non fecit ei populus secundum morem conbustionis exequias sicut fecerat maioribus eius
2CHR|21|20|triginta duum annorum fuit cum regnare coepisset et octo annis regnavit in Hierusalem ambulavitque non recte et sepelierunt eum in civitate David verumtamen non in sepulchro regum
2CHR|22|1|constituerunt autem habitatores Hierusalem Ochoziam filium eius minimum regem pro eo omnes enim maiores natu qui ante eum fuerant interfecerant latrones Arabum qui inruerant in castra regnavitque Ochozias filius Ioram regis Iuda
2CHR|22|2|filius quadraginta duo annorum erat Ochozias cum regnare coepisset et uno anno regnavit in Hierusalem nomen matris eius Otholia filia Amri
2CHR|22|3|sed et ipse ingressus est per vias domus Ahab mater enim eius inpulit eum ut impie ageret
2CHR|22|4|fecit igitur malum in conspectu Domini sicut domus Ahab ipsi enim fuerunt ei consiliarii post mortem patris sui in interitum eius
2CHR|22|5|ambulavitque in consiliis eorum et perrexit cum Ioram filio Ahab rege Israhel in bellum contra Azahel regem Syriae in Ramoth Galaad vulneraveruntque Syri Ioram
2CHR|22|6|qui reversus est ut curaretur in Hiezrahel multas enim plagas acceperat in supradicto certamine igitur Azarias filius Ioram rex Iuda descendit ut inviseret Ioram filium Ahab in Hiezrahel aegrotantem
2CHR|22|7|voluntatis quippe fuit Dei adversum Ochoziam ut veniret ad Ioram et cum venisset egrederetur cum eo adversum Hieu filium Namsi quem unxit Dominus ut deleret domum Ahab
2CHR|22|8|cum ergo subverteret Hieu domum Ahab invenit principes Iuda et filios fratrum Ochoziae qui ministrabant ei et interfecit illos
2CHR|22|9|ipsumque perquirens Ochoziam conprehendit latentem in Samaria adductumque ad se occidit et sepelierunt eum eo quod esset filius Iosaphat qui quaesierat Dominum in toto corde suo nec erat ultra spes aliqua ut de stirpe regnaret Ochoziae
2CHR|22|10|siquidem Otholia mater eius videns quod mortuus esset filius suus surrexit et interfecit omnem stirpem regiam domus Ioram
2CHR|22|11|porro Iosabeth filia regis tulit Ioas filium Ochoziae et furata est eum de medio filiorum regis cum interficerentur absconditque cum nutrice sua in cubiculo lectulorum Iosabeth autem quae absconderat eum erat filia regis Ioram uxor Ioiadae pontificis soror Ochoziae et idcirco Otholia non interfecit eum
2CHR|22|12|fuit ergo cum eis in domo Dei absconditus sex annis quibus regnavit Otholia super terram
2CHR|23|1|anno autem septimo confortatus Ioiadae adsumpsit centuriones Azariam videlicet filium Hieroam et Ismahel filium Iohanan Azariam quoque filium Oded et Maasiam filium Adaiae et Elisaphat filium Zechri et iniit cum eis foedus
2CHR|23|2|qui circumeuntes Iudam congregaverunt Levitas de cunctis urbibus Iuda et principes familiarum Israhel veneruntque in Hierusalem
2CHR|23|3|iniit igitur omnis multitudo pactum in domo Domini cum rege dixitque ad eos Ioiadae ecce filius regis regnabit sicut locutus est Dominus super filios David
2CHR|23|4|iste est ergo sermo quem facietis
2CHR|23|5|tertia pars vestrum qui veniunt ad sabbatum sacerdotum et Levitarum et ianitorum erit in portis tertia vero pars ad domum regis et tertia in porta quae appellatur Fundamenti omne vero reliquum vulgus sit in atriis domus Domini
2CHR|23|6|nec quisquam alius ingrediatur domum Domini nisi sacerdotes et qui ministrant de Levitis ipsi tantummodo ingrediantur quia sanctificati sunt et omne reliquum vulgus observet custodias Domini
2CHR|23|7|Levitae autem circumdent regem habentes singuli arma sua et si quis alius ingressus fuerit templum interficiatur sintque cum rege et intrante et egrediente
2CHR|23|8|fecerunt igitur Levitae et universus Iuda iuxta omnia quae praeceperat Ioiadae pontifex et adsumpserunt singuli viros qui sub se erant et veniebant per ordinem sabbati cum his qui iam impleverant sabbatum et egressuri erant siquidem Ioiadae pontifex non dimiserat abire turmas quae sibi per singulas ebdomadas succedere consueverant
2CHR|23|9|deditque Ioiadae sacerdos centurionibus lanceas clypeosque et peltas regis David quas consecraverat in domo Domini
2CHR|23|10|constituitque omnem populum tenentium pugiones a parte templi dextra usque ad partem templi sinistram coram altari et templo per circuitum regis
2CHR|23|11|et eduxerunt filium regis et inposuerunt ei diadema dederuntque in manu eius tenendam legem et constituerunt eum regem unxit quoque illum Ioiadae pontifex et filii eius inprecatique sunt atque dixerunt vivat rex
2CHR|23|12|quod cum audisset Otholia vocem scilicet currentium atque laudantium regem ingressa est ad populum in templum Domini
2CHR|23|13|cumque vidisset regem stantem super gradum in introitu et principes turmasque circa eum omnem quoque populum terrae gaudentem atque clangentem tubis et diversi generis organis concinentem vocemque laudantium scidit vestimenta sua et ait insidiae insidiae
2CHR|23|14|egressus autem Ioiadae pontifex ad centuriones et principes exercitus dixit eis educite illam extra septa templi et interficiatur foris gladio praecepitque sacerdos ne occideretur in domo Domini
2CHR|23|15|et inposuerunt cervicibus eius manus cumque intrasset portam Equorum domus regis interfecerunt eam ibi
2CHR|23|16|pepigit autem Ioiadae foedus inter se universumque populum et regem ut esset populus Domini
2CHR|23|17|itaque ingressus est omnis populus domum Baal et destruxerunt eam et altaria ac simulacra illius confregerunt Matthan quoque sacerdotem Baal interfecerunt ante aras
2CHR|23|18|constituit autem Ioiadae praepositos in domo Domini et sub manibus sacerdotum ac Levitarum quos distribuit David in domo Domini ut offerrent holocausta Domino sicut scriptum est in lege Mosi in gaudio et canticis iuxta dispositionem David
2CHR|23|19|constituit quoque ianitores in portis domus Domini ut non ingrederetur eam inmundus in omni re
2CHR|23|20|adsumpsitque centuriones et fortissimos viros ac principes populi et omne vulgus terrae et fecerunt descendere regem de domo Domini et introire per medium portae superioris in domum regis et conlocaverunt eum in solio regali
2CHR|23|21|laetatusque est omnis populus terrae et urbs quievit porro Otholia interfecta est gladio
2CHR|24|1|septem annorum erat Ioas cum regnare coepisset et quadraginta annis regnavit in Hierusalem nomen matris eius Sebia de Bersabee
2CHR|24|2|fecitque quod bonum est coram Domino cunctis diebus Ioiadae sacerdotis
2CHR|24|3|accepit autem ei Ioiadae uxores duas e quibus genuit filios et filias
2CHR|24|4|post quae placuit Ioas ut instauraret domum Domini
2CHR|24|5|congregavitque sacerdotes et Levitas et dixit eis egredimini ad civitates Iuda et colligite de universo Israhel pecuniam ad sarta tecta templi Dei vestri per singulos annos festinatoque hoc facite porro Levitae egere neglegentius
2CHR|24|6|vocavitque rex Ioiadae principem et dixit ei quare non tibi fuit curae ut cogeres Levitas inferre de Iuda et de Hierusalem pecuniam quae constituta est a Mose servo Domini ut inferret eam omnis multitudo Israhel in tabernaculum testimonii
2CHR|24|7|Otholia enim impiissima et filii eius destruxerunt domum Domini et de universis quae sanctificata fuerant templo Domini ornaverunt fanum Baalim
2CHR|24|8|praecepit ergo rex et fecerunt arcam posueruntque eam iuxta portam domus Domini forinsecus
2CHR|24|9|et praedicatum est in Iuda et Hierusalem ut deferrent singuli pretium Domino quod constituit Moses servus Dei super omnem Israhel in deserto
2CHR|24|10|laetatique sunt cuncti principes et omnis populus et ingressi contulerunt in arcam Domini atque miserunt ita ut impleretur
2CHR|24|11|cumque tempus esset ut deferrent arcam coram rege per manus Levitarum videbant enim multam pecuniam ingrediebatur scriba regis et quem primus sacerdos constituerat effundebantque pecuniam quae erat in arca porro arcam reportabant ad locum suum sicque faciebant per singulos dies et congregata est infinita pecunia
2CHR|24|12|quam dederunt rex et Ioiada his qui praeerant operibus domus Domini at illi conducebant ex ea caesores lapidum et artifices operum singulorum ut instaurarent domum Domini fabros quoque ferri et aeris ut quod cadere coeperat fulciretur
2CHR|24|13|egeruntque hii qui operabantur industrie et obducebatur parietum cicatrix per manus eorum ac suscitaverunt domum Domini in statum pristinum et firme eam stare fecerunt
2CHR|24|14|cumque conplessent omnia opera detulerunt coram rege et Ioiadae reliquam partem pecuniae de qua facta sunt vasa templi in ministerium et ad holocausta fialae quoque et cetera vasa aurea et argentea et offerebantur holocausta in domo Domini iugiter cunctis diebus Ioiadae
2CHR|24|15|senuit autem Ioiadae plenus dierum et mortuus est cum centum triginta esset annorum
2CHR|24|16|sepelieruntque eum in civitate David cum regibus eo quod fecisset bonum cum Israhel et cum domo eius
2CHR|24|17|postquam autem obiit Ioiada ingressi sunt principes Iuda et adoraverunt regem qui delinitus obsequiis eorum adquievit eis
2CHR|24|18|et dereliquerunt templum Domini Dei patrum suorum servieruntque lucis et sculptilibus et facta est ira contra Iudam et Hierusalem propter hoc peccatum
2CHR|24|19|mittebatque eis prophetas ut reverterentur ad Dominum quos protestantes illi audire nolebant
2CHR|24|20|spiritus itaque Dei induit Zacchariam filium Ioiadae sacerdotem et stetit in conspectu populi et dixit eis haec dicit Dominus quare transgredimini praeceptum Domini quod vobis non proderit et dereliquistis Dominum ut derelinqueret vos
2CHR|24|21|qui congregati adversus eum miserunt lapides iuxta regis imperium in atrio domus Domini
2CHR|24|22|et non est recordatus Ioas rex misericordiae quam fecerat Ioiadae pater illius secum sed interfecit filium eius qui cum moreretur ait videat Dominus et requirat
2CHR|24|23|cumque evolutus esset annus ascendit contra eum exercitus Syriae venitque in Iudam et Hierusalem et interfecit cunctos principes populi atque universam praedam miserunt regi Damascum
2CHR|24|24|et certe cum permodicus venisset numerus Syrorum tradidit Dominus manibus eorum infinitam multitudinem eo quod reliquissent Dominum Deum patrum suorum in Ioas quoque ignominiosa exercuere iudicia
2CHR|24|25|et abeuntes dimiserunt eum in languoribus magnis surrexerunt autem contra eum servi sui in ultionem sanguinis filii Ioiadae sacerdotis et occiderunt eum in lectulo suo et mortuus est sepelieruntque eum in civitate David sed non in sepulchris regum
2CHR|24|26|insidiati vero sunt ei Zabath filius Semath Ammanitidis et Iozabath filius Semarith Moabitidis
2CHR|24|27|porro filii eius ac summa pecuniae quae adunata fuerat sub eo et instauratio domus Dei scripta sunt diligentius in libro regum regnavitque Amasias filius eius pro eo
2CHR|25|1|viginti quinque annorum erat Amasias cum regnare coepisset et viginti novem annis regnavit in Hierusalem nomen matris eius Ioaden de Hierusalem
2CHR|25|2|fecitque bonum in conspectu Domini verumtamen non in corde perfecto
2CHR|25|3|cumque roboratum sibi videret imperium iugulavit servos qui occiderant regem patrem suum
2CHR|25|4|sed filios eorum non interfecit sicut scriptum est in libro legis Mosi ubi praecepit Dominus dicens non occidentur patres pro filiis neque filii pro patribus suis sed unusquisque in suo peccato morietur
2CHR|25|5|congregavit igitur Amasias Iudam et constituit eos per familias tribunosque et centuriones in universo Iuda et Beniamin et recensuit a viginti annis sursum invenitque triginta milia iuvenum qui egrederentur ad pugnam et tenerent hastam et clypeum
2CHR|25|6|mercede quoque conduxit de Israhel centum milia robustorum centum talentis argenti
2CHR|25|7|venit autem homo Dei ad illum et ait o rex ne egrediatur tecum exercitus Israhel non est enim Dominus cum Israhel et cunctis filiis Ephraim
2CHR|25|8|quod si putas in robore exercitus bella consistere superari te faciet Deus ab hostibus Dei quippe est et adiuvare et in fugam vertere
2CHR|25|9|dixitque Amasias ad hominem Dei quid ergo fiet de centum talentis quae dedi militibus Israhel et respondit ei homo Dei habet Dominus unde tibi dare possit multo his plura
2CHR|25|10|separavit itaque Amasias exercitum qui venerat ad eum ex Ephraim ut reverteretur in locum suum at illi contra Iudam vehementer irati reversi sunt in regionem suam
2CHR|25|11|porro Amasias confidenter eduxit populum suum et abiit in vallem Salinarum percussitque filios Seir decem milia
2CHR|25|12|et alia decem milia virorum ceperunt filii Iuda et adduxerunt ad praeruptum cuiusdam petrae praecipitaveruntque eos de summo in praeceps qui universi crepuerunt
2CHR|25|13|at ille exercitus quem remiserat Amasias ne secum iret ad proelium diffusus est in civitatibus Iuda a Samaria usque Bethoron et interfectis tribus milibus diripuit praedam magnam
2CHR|25|14|Amasias vero post caedem Idumeorum et adlatos deos filiorum Seir statuit illos in deos sibi et adorabat eos et illis adolebat incensum
2CHR|25|15|quam ob rem iratus Dominus contra Amasiam misit ad illum prophetam qui diceret ei cur adorasti deos qui non liberaverunt populum suum de manu tua
2CHR|25|16|cumque haec ille loqueretur respondit ei num consiliarius regis es quiesce ne interficiam te discedensque propheta scio inquit quod cogitaverit Dominus occidere te qui et fecisti hoc malum et insuper non adquievisti consilio meo
2CHR|25|17|igitur Amasias rex Iuda inito pessimo consilio misit ad Ioas filium Ioachaz filii Hieu regem Israhel dicens veni videamus nos mutuo
2CHR|25|18|at ille remisit nuntium dicens carduus qui est in Libano misit ad cedrum Libani dicens da filiam tuam filio meo uxorem et ecce bestiae quae erant in silva Libani transierunt et conculcaverunt carduum
2CHR|25|19|dixisti percussi Edom et idcirco erigitur cor tuum in superbiam sede in domo tua cur malum adversum te provocas ut cadas et tu et Iudas tecum
2CHR|25|20|noluit audire Amasias eo quod Domini esset voluntas ut traderetur in manibus hostium propter deos Edom
2CHR|25|21|ascendit igitur Ioas rex Israhel et mutuos sibi praebuere conspectus Amasias autem rex Iuda erat in Bethsames Iudae
2CHR|25|22|corruitque Iudas coram Israhel et fugit in tabernacula sua
2CHR|25|23|porro Amasiam regem Iuda filium Ioas filii Ioachaz cepit Ioas rex Israhel in Bethsames et adduxit in Hierusalem destruxitque murum eius a porta Ephraim usque ad portam Anguli quadringentis cubitis
2CHR|25|24|omne quoque aurum et argentum et universa vasa quae reppererat in domo Dei et apud Obededom in thesauris etiam domus regiae necnon et filios obsidum reduxit Samariam
2CHR|25|25|vixit autem Amasias filius Ioas rex Iuda postquam mortuus est Ioas filius Ioachaz rex Israhel quindecim annis
2CHR|25|26|reliqua vero sermonum Amasiae priorum et novissimorum scripta sunt in libro regum Iuda et Israhel
2CHR|25|27|qui postquam recessit a Domino tetenderunt ei insidias in Hierusalem cumque fugisset Lachis miserunt et interfecerunt eum ibi
2CHR|25|28|reportantesque super equos sepelierunt eum cum patribus suis in civitate David
2CHR|26|1|omnis autem populus Iuda filium eius Oziam annorum sedecim constituit regem pro patre suo Amasia
2CHR|26|2|ipse aedificavit Ahilath et restituit eam dicioni Iudae postquam dormivit rex cum patribus suis
2CHR|26|3|sedecim annorum erat Ozias cum regnare coepisset et quinquaginta duobus annis regnavit in Hierusalem nomen matris eius Hiechelia de Hierusalem
2CHR|26|4|fecitque quod erat rectum in oculis Domini iuxta omnia quae fecerat Amasias pater eius
2CHR|26|5|et exquisivit Deum in diebus Zacchariae intellegentis et videntis Deum cumque requireret Dominum direxit eum in omnibus
2CHR|26|6|denique egressus est et pugnavit contra Philisthim et destruxit murum Geth et murum Iabniae murumque Azoti aedificavit quoque oppida in Azoto et in Philisthim
2CHR|26|7|et adiuvit eum Deus contra Philisthim et contra Arabas qui habitabant in Gurbaal et contra Ammanitas
2CHR|26|8|pendebantque Ammanitae munera Oziae et divulgatum est nomen eius usque ad introitum Aegypti propter crebras victorias
2CHR|26|9|aedificavitque Ozias turres in Hierusalem super portam Anguli et super portam Vallis et reliquas in eodem muri latere firmavitque eas
2CHR|26|10|extruxit etiam turres in solitudine et fodit cisternas plurimas eo quod haberet multa pecora tam in campestribus quam in heremi vastitate vineas quoque habuit et vinitores in montibus et in Carmelo erat quippe homo agriculturae deditus
2CHR|26|11|fuit autem exercitus bellatorum eius qui procedebant ad proelia sub manu Hiehihel scribae Maasiaeque doctoris et sub manu Ananiae qui erat de ducibus regis
2CHR|26|12|omnisque numerus principum per familias virorum fortium duum milium sescentorum
2CHR|26|13|et sub eis universus exercitus trecentorum et septem milium quingentorum qui erant apti ad bella et pro rege contra adversarios dimicabant
2CHR|26|14|praeparavit quoque eis Ozias id est cuncto exercitui clypeos et hastas et galeas et loricas arcusque et fundas ad iaciendos lapides
2CHR|26|15|et fecit in Hierusalem diversi generis machinas quas in turribus conlocavit et in angulis murorum ut mitterent sagittas et saxa grandia egressumque est nomen eius procul eo quod auxiliaretur ei Dominus et corroborasset illum
2CHR|26|16|sed cum roboratus esset elevatum est cor eius in interitum suum et neglexit Dominum Deum suum ingressusque templum Domini adolere voluit incensum super altare thymiamatis
2CHR|26|17|statimque ingressus post eum Azarias sacerdos et cum eo sacerdotes Domini octoginta viri fortissimi
2CHR|26|18|restiterunt regi atque dixerunt non est tui officii Ozia ut adoleas incensum Domino sed sacerdotum hoc est filiorum Aaron qui consecrati sunt ad huiuscemodi ministerium egredere de sanctuario ne contempseris quia non reputabitur tibi in gloriam hoc a Domino Deo
2CHR|26|19|iratusque est Ozias et tenens in manu turibulum ut adoleret incensum minabatur sacerdotibus statimque orta est lepra in fronte eius coram sacerdotibus in domo Domini super altare thymiamatis
2CHR|26|20|cumque respexisset eum Azarias pontifex et omnes reliqui sacerdotes viderunt lepram in fronte eius et festinato expulerunt eum sed et ipse perterritus adceleravit egredi eo quod sensisset ilico plagam Domini
2CHR|26|21|fuit igitur Ozias rex leprosus usque ad diem mortis suae et habitavit in domo separata plenus lepra ob quam et eiectus fuerat de domo Domini porro Ioatham filius eius rexit domum regis et iudicabat populum terrae
2CHR|26|22|reliqua autem sermonum Oziae priorum et novissimorum scripsit Esaias filius Amos propheta
2CHR|26|23|dormivitque Ozias cum patribus suis et sepelierunt eum in agro regalium sepulchrorum eo quod esset leprosus regnavitque Ioatham filius eius pro eo
2CHR|27|1|viginti quinque annorum erat Ioatham cum regnare coepisset et sedecim annis regnavit in Hierusalem nomen matris eius Hierusa filia Sadoc
2CHR|27|2|fecitque quod rectum erat coram Domino iuxta omnia quae fecerat Ozias pater suus excepto quod non est ingressus templum Domini et adhuc populus delinquebat
2CHR|27|3|ipse aedificavit portam domus Domini Excelsam et in muro Ophel multa construxit
2CHR|27|4|urbes quoque aedificavit in montibus Iuda et in saltibus castella et turres
2CHR|27|5|ipse pugnavit contra regem filiorum Ammon et vicit eos dederuntque ei filii Ammon in tempore illo centum talenta argenti et decem milia choros tritici ac totidem choros hordei haec ei praebuerunt filii Ammon in anno secundo et tertio
2CHR|27|6|corroboratusque est Ioatham eo quod direxisset vias suas coram Domino Deo suo
2CHR|27|7|reliqua autem sermonum Ioatham et omnes pugnae eius et opera scripta sunt in libro regum Israhel et Iuda
2CHR|27|8|viginti quinque annorum erat cum regnare coepisset et sedecim annis regnavit in Hierusalem
2CHR|27|9|dormivitque Ioatham cum patribus suis et sepelierunt eum in civitate David et regnavit Achaz filius eius pro eo
2CHR|28|1|viginti annorum erat Achaz cum regnare coepisset et sedecim annis regnavit in Hierusalem non fecit rectum in conspectu Domini sicut David pater eius
2CHR|28|2|sed ambulavit in viis regum Israhel insuper et statuas fudit Baalim
2CHR|28|3|ipse est qui adolevit incensum in valle Benennon et lustravit filios suos in igne iuxta ritum gentium quas interfecit Dominus in adventu filiorum Israhel
2CHR|28|4|sacrificabat quoque et thymiama succendebat in excelsis et in collibus et sub omni ligno frondoso
2CHR|28|5|tradiditque eum Dominus Deus eius in manu regis Syriae qui percussit eum magnamque praedam de eius cepit imperio et adduxit in Damascum manibus quoque regis Israhel traditus est et percussus plaga grandi
2CHR|28|6|occiditque Phacee filius Romeliae de Iuda centum viginti milia in die uno omnes viros bellatores eo quod reliquissent Dominum Deum patrum suorum
2CHR|28|7|eodem tempore occidit Zechri vir potens ex Ephraim Masiam filium regis et Ezricam ducem domus eius Helcanam quoque secundum a rege
2CHR|28|8|ceperuntque filii Israhel de fratribus suis ducenta milia mulierum puerorum et puellarum et infinitam praedam pertuleruntque eam in Samariam
2CHR|28|9|ea tempestate erat ibi propheta Domini nomine Oded qui egressus obviam exercitui venientium in Samariam dixit eis ecce iratus Dominus Deus patrum vestrorum contra Iudam tradidit eos manibus vestris et occidistis illos atrociter ita ut caelum pertingeret vestra crudelitas
2CHR|28|10|insuper filios Iuda et Hierusalem vultis vobis subicere in servos et ancillas quod nequaquam facto opus est peccatis enim super hoc Domino Deo vestro
2CHR|28|11|sed audite consilium meum et reducite captivos quos adduxistis de fratribus vestris quia magnus furor Domini inminet vobis
2CHR|28|12|steterunt itaque viri de principibus filiorum Ephraim Azarias filius Iohanan Barachias filius Mosollamoth Hiezechias filius Sellum et Amasa filius Adali contra eos qui veniebant de proelio
2CHR|28|13|et dixerunt eis non introducetis huc captivos ne peccemus Domino quare vultis adicere super peccata nostra et vetera cumulare delicta grande quippe peccatum est et ira furoris Domini inminet super Israhel
2CHR|28|14|dimiseruntque viri bellatores praedam et universa quae ceperant coram principibus et omni multitudine
2CHR|28|15|steteruntque viri quos supra memoravimus et adprehendentes captivos omnesque qui nudi erant vestierunt de spoliis cumque vestissent eos et calciassent et refecissent cibo ac potu unxissent quoque propter laborem et adhibuissent eis curam quicumque ambulare non poterant et erant inbecillo corpore inposuerunt eos iumentis et adduxerunt Hierichum civitatem Palmarum ad fratres eorum ipsique reversi sunt Samariam
2CHR|28|16|tempore illo misit rex Achaz ad regem Assyriorum auxilium postulans
2CHR|28|17|veneruntque Idumei et percusserunt multos ex Iuda et ceperunt praedam magnam
2CHR|28|18|Philisthim quoque diffusi sunt per urbes campestres et ad meridiem Iuda ceperuntque Bethsames et Ahilon et Gaderoth Soccho quoque et Thamnam et Gamzo cum viculis suis et habitaverunt in eis
2CHR|28|19|humiliaverat enim Dominus Iudam propter Achaz regem Iuda eo quod nudasset eum auxilio et contemptui habuisset Dominum
2CHR|28|20|adduxitque contra eum Thaglathphalnasar regem Assyriorum qui et adflixit eum et nullo resistente vastavit
2CHR|28|21|igitur Achaz spoliata domo Domini et domo regum et principum dedit regi Assyriorum munera et tamen nihil ei profuit
2CHR|28|22|insuper et in tempore angustiae suae auxit contemptum in Dominum ipse per se rex Achaz
2CHR|28|23|immolavit diis Damasci victimas percussoribus suis et dixit dii regum Syriae auxiliantur eis quos ego placabo hostiis et aderunt mihi cum e contrario ipsi fuerint ruina eius et universo Israhel
2CHR|28|24|direptis itaque Achaz omnibus vasis domus Dei atque confractis clusit ianuas templi Dei et fecit sibi altaria in universis angulis Hierusalem
2CHR|28|25|in omnibus quoque urbibus Iuda extruxit aras ad cremandum tus atque ad iracundiam provocavit Dominum Deum patrum suorum
2CHR|28|26|reliqua autem sermonum eius et omnium operum priorum et novissimorum scripta sunt in libro regum Iuda et Israhel
2CHR|28|27|dormivitque Achaz cum patribus suis et sepelierunt eum in civitate Hierusalem neque enim receperunt eum in sepulchra regum Israhel regnavitque Ezechias filius eius pro eo
2CHR|29|1|igitur Ezechias regnare coepit cum viginti quinque esset annorum et viginti novem annis regnavit in Hierusalem nomen matris eius Abia filia Zacchariae
2CHR|29|2|fecitque quod erat placitum in conspectu Domini iuxta omnia quae fecerat David pater eius
2CHR|29|3|ipse anno et mense primo regni sui aperuit valvas domus Domini et instauravit eas
2CHR|29|4|adduxitque sacerdotes atque Levitas et congregavit eos in plateam orientalem
2CHR|29|5|dixitque ad eos audite me Levitae et sanctificamini mundate domum Domini Dei patrum vestrorum auferte omnem inmunditiam de sanctuario
2CHR|29|6|peccaverunt patres nostri et fecerunt malum in conspectu Domini Dei nostri derelinquentes eum averterunt facies suas a tabernaculo Domini et praebuerunt dorsum
2CHR|29|7|cluserunt ostia quae erant in porticu et extinxerunt lucernas incensumque non adoleverunt et holocausta non obtulerunt in sanctuario Deo Israhel
2CHR|29|8|concitatus est itaque furor Domini super Iudam et Hierusalem tradiditque eos in commotionem et in interitum et in sibilum sicut ipsi cernitis oculis vestris
2CHR|29|9|en corruerunt patres nostri gladiis filii nostri et filiae nostrae et coniuges captivae ductae sunt propter hoc scelus
2CHR|29|10|nunc igitur placet mihi ut ineamus foedus cum Domino Deo Israhel et avertat a nobis furorem irae suae
2CHR|29|11|filii mi nolite neglegere vos elegit Dominus ut stetis coram eo et ministretis illi colatis eum et cremetis incensum
2CHR|29|12|surrexerunt ergo Levitae Maath filius Amasiae et Iohel filius Azariae de filiis Caath porro de filiis Merari Cis filius Abdai et Azarias filius Iallelel de filiis autem Gersom Ioha filius Zemma et Eden filius Ioaha
2CHR|29|13|at vero de filiis Elisaphan Samri et Iahihel de filiis quoque Asaph Zaccharias et Mathanias
2CHR|29|14|necnon de filiis Heman Iahihel et Semei sed et de filiis Idithun Semeias et Ozihel
2CHR|29|15|congregaveruntque fratres suos et sanctificati sunt et ingressi iuxta mandatum regis et imperium Domini ut expiarent domum Dei
2CHR|29|16|sacerdotes quoque ingressi templum Domini ut sanctificarent illud extulerunt omnem inmunditiam quam intro reppererant in vestibulum domus Domini quam tulerunt Levitae et asportaverunt ad torrentem Cedron foras
2CHR|29|17|coeperunt autem prima die mensis primi mundare et in die octava eiusdem mensis ingressi sunt porticum templi Domini expiaveruntque templum diebus octo et in die sextadecima mensis eiusdem quod coeperant impleverunt
2CHR|29|18|ingressi quoque sunt ad Ezechiam regem et dixerunt ei sanctificavimus omnem domum Domini et altare holocaustoseos vasaque eius necnon et mensam propositionis cum omnibus vasis suis
2CHR|29|19|cunctamque templi supellectilem quam polluerat rex Achaz in regno suo postquam praevaricatus est et ecce exposita sunt omnia coram altari Domini
2CHR|29|20|consurgensque diluculo Ezechias rex adunavit omnes principes civitatis et ascendit domum Domini
2CHR|29|21|obtuleruntque simul tauros septem arietes septem agnos septem et hircos septem pro peccato pro regno pro sanctuario pro Iuda dixit quoque sacerdotibus filiis Aaron ut offerrent super altare Domini
2CHR|29|22|mactaverunt igitur tauros et susceperunt sacerdotes sanguinem et fuderunt illud super altare mactaverunt etiam arietes et illorum sanguinem super altare fuderunt immolaverunt agnos et fuderunt super altare sanguinem
2CHR|29|23|adplicaverunt hircos pro peccato coram rege et universa multitudine inposueruntque manus suas super eos
2CHR|29|24|et immolaverunt illos sacerdotes et asperserunt sanguinem eorum altari pro piaculo universi Israhelis pro omni quippe Israhel praeceperat rex ut holocaustum fieret et pro peccato
2CHR|29|25|constituit quoque Levitas in domo Domini cum cymbalis et psalteriis et citharis secundum dispositionem David et Gad videntis regis et Nathan prophetae siquidem Domini praeceptum fuit per manum prophetarum eius
2CHR|29|26|steteruntque Levitae tenentes organa David et sacerdotes tubas
2CHR|29|27|et iussit Ezechias ut offerrent holocaustum super altare cumque offerrentur holocausta coeperunt laudes canere Domino et clangere tubis atque in diversis organis quae David rex Israhel reppererat concrepare
2CHR|29|28|omni autem turba adorante cantores et hii qui tenebant tubas erant in officio suo donec conpleretur holocaustum
2CHR|29|29|cumque finita esset oblatio incurvatus est rex et omnes qui erant cum eo et adoraverunt
2CHR|29|30|praecepitque Ezechias et principes Levitis ut laudarent Dominum sermonibus David et Asaph videntis qui laudaverunt eum magna laetitia et curvato genu adoraverunt
2CHR|29|31|Ezechias autem etiam haec addidit implestis manus vestras Domino accedite et offerte victimas et laudes in domo Domini obtulit ergo universa multitudo hostias et laudes et holocausta mente devota
2CHR|29|32|porro numerus holocaustorum quae obtulit multitudo hic fuit tauros septuaginta arietes centum agnos ducentos
2CHR|29|33|sanctificaveruntque Domino boves sescentos et oves tria milia
2CHR|29|34|sacerdotes vero pauci erant nec poterant sufficere ut pelles holocaustorum detraherent unde et Levitae fratres eorum adiuverunt eos donec impleretur opus et sanctificarentur antistites Levitae quippe faciliori ritu sanctificantur quam sacerdotes
2CHR|29|35|fuerunt igitur holocausta plurima adipes pacificorum et libamina holocaustorum et conpletus est cultus domus Domini
2CHR|29|36|laetatusque est Ezechias et omnis populus eo quod ministerium Domini esset expletum de repente quippe hoc fieri placuerat
2CHR|30|1|misit quoque Ezechias ad omnem Israhel et Iudam scripsitque epistulas ad Ephraim et Manassem ut venirent ad domum Domini in Hierusalem et facerent phase Domino Deo Israhel
2CHR|30|2|inito ergo consilio regis et principum et universi coetus Hierusalem decreverunt ut facerent phase mense secundo
2CHR|30|3|non enim occurrerant facere in tempore suo quia sacerdotes qui possent sufficere sanctificati non fuerant et populus necdum congregatus erat in Hierusalem
2CHR|30|4|placuitque sermo regi et omni multitudini
2CHR|30|5|et decreverunt ut mitterent nuntios in universum Israhel de Bersabee usque Dan ut venirent et facerent phase Domino Deo Israhel in Hierusalem multi enim non fecerant sicut lege praescriptum est
2CHR|30|6|perrexeruntque cursores cum epistulis ex regis imperio et principum eius in universum Israhel et Iudam iuxta quod rex iusserat praedicantes filii Israhel revertimini ad Dominum Deum Abraham et Isaac et Israhel et revertetur ad reliquias quae effugerunt manum regis Assyriorum
2CHR|30|7|nolite fieri sicut patres vestri et fratres qui recesserunt a Domino Deo patrum suorum et tradidit eos in interitum ut ipsi cernitis
2CHR|30|8|nolite indurare cervices vestras sicut patres vestri tradite manus Domino et venite ad sanctuarium eius quod sanctificavit in aeternum servite Domino Deo patrum vestrorum et avertetur a vobis ira furoris eius
2CHR|30|9|si enim vos reversi fueritis ad Dominum fratres vestri et filii habebunt misericordiam coram dominis suis qui illos duxere captivos et revertentur in terram hanc pius enim et clemens est Dominus Deus vester et non avertet faciem suam a vobis si reversi fueritis ad eum
2CHR|30|10|igitur cursores pergebant velociter de civitate in civitatem per terram Ephraim et Manasse usque Zabulon illis inridentibus et subsannantibus eos
2CHR|30|11|attamen quidam viri ex Aser et Manasse et Zabulon adquiescentes consilio venerunt Hierusalem
2CHR|30|12|in Iuda vero facta est manus Domini ut daret eis cor unum et facerent iuxta praeceptum regis et principum verbum Domini
2CHR|30|13|congregatique sunt in Hierusalem populi multi ut facerent sollemnitatem azymorum in mense secundo
2CHR|30|14|et surgentes destruxerunt altaria quae erant in Hierusalem atque universa in quibus idolis adolebatur incensum subvertentes proiecerunt in torrentem Cedron
2CHR|30|15|immolaverunt autem phase quartadecima die mensis secundi sacerdotes quoque atque Levitae tandem sanctificati obtulerunt holocausta in domo Domini
2CHR|30|16|steteruntque in ordine suo iuxta dispositionem et legem Mosi hominis Dei sacerdotes vero suscipiebant effundendum sanguinem de manibus Levitarum
2CHR|30|17|eo quod multa turba sanctificata non esset et idcirco Levitae immolarent phase his qui non occurrerant sanctificari Domino
2CHR|30|18|magna etiam pars populi de Ephraim et Manasse et Isachar et Zabulon quae sanctificata non fuerat comedit phase non iuxta quod scriptum est et oravit pro eis Ezechias dicens Dominus bonus propitiabitur
2CHR|30|19|cunctis qui in toto corde requirunt Dominum Deum patrum suorum et non inputabit eis quod minus sanctificati sunt
2CHR|30|20|quem exaudivit Dominus et placatus est populo
2CHR|30|21|feceruntque filii Israhel qui inventi sunt in Hierusalem sollemnitatem azymorum septem diebus in laetitia magna laudantes Dominum per singulos dies Levitae quoque et sacerdotes per organa quae suo officio congruebant
2CHR|30|22|et locutus est Ezechias ad cor omnium Levitarum qui habebant intellegentiam bonam super Domino et comederunt septem diebus sollemnitatis immolantes victimas pacificorum et laudantes Dominum Deum patrum suorum
2CHR|30|23|placuitque universae multitudini ut celebrarent etiam alios dies septem quod et fecerunt cum ingenti gaudio
2CHR|30|24|Ezechias enim rex Iuda praebuerat multitudini mille tauros et septem milia ovium principes vero dederant populo tauros mille et oves decem milia sanctificata ergo est sacerdotum plurima multitudo
2CHR|30|25|et hilaritate perfusa omnis turba Iuda tam sacerdotum et Levitarum quam universae frequentiae quae venerat ex Israhel proselytorum quoque de terra Israhel et habitantium in Iuda
2CHR|30|26|factaque est grandis celebritas in Hierusalem qualis a diebus Salomonis filii David regis Israhel in ea urbe non fuerat
2CHR|30|27|surrexerunt autem sacerdotes atque Levitae benedicentes populo et exaudita est vox eorum pervenitque oratio in habitaculum sanctum caeli
2CHR|31|1|cumque haec fuissent rite celebrata egressus est omnis Israhel qui inventus fuerat in urbibus Iuda et fregerunt simulacra succideruntque lucos demoliti sunt excelsa et altaria destruxerunt non solum de universo Iuda et Beniamin sed de Ephraim quoque et Manasse donec penitus everterent reversique sunt omnes filii Israhel in possessiones et civitates suas
2CHR|31|2|Ezechias vero constituit turmas sacerdotales et leviticas per divisiones suas unumquemque in officio proprio tam sacerdotum videlicet quam Levitarum ad holocausta et pacifica ut ministrarent et confiterentur canerentque in portis castrorum Domini
2CHR|31|3|pars autem regis erat ut de propria eius substantia offerretur holocaustum mane semper et vespere sabbatis quoque et kalendis et sollemnitatibus ceteris sicut scriptum est in lege Mosi
2CHR|31|4|praecepit etiam populo habitantium Hierusalem ut darent partes sacerdotibus et Levitis et possent vacare legi Domini
2CHR|31|5|quod cum percrebruisset in auribus multitudinis plurimas obtulere primitias filii Israhel frumenti vini et olei mellis quoque et omnium quae gignit humus decimas obtulerunt
2CHR|31|6|sed et filii Israhel et Iuda qui habitabant in urbibus Iuda obtulerunt decimas boum et ovium decimasque sanctorum quae voverant Domino Deo suo atque universa portantes fecerunt acervos plurimos
2CHR|31|7|mense tertio coeperunt acervorum iacere fundamenta et mense septimo conpleverunt eos
2CHR|31|8|cumque ingressi fuissent Ezechias et principes eius viderunt acervos et benedixerunt Domino ac populo Israhel
2CHR|31|9|interrogavitque Ezechias sacerdotes et Levitas cur ita iacerent acervi
2CHR|31|10|respondit illi Azarias sacerdos primus de stirpe Sadoc dicens ex quo coeperunt offerri primitiae in domo Domini comedimus et saturati sumus remanseruntque plurima eo quod benedixerit Dominus populo suo reliquiarum autem copia est ista quam cernis
2CHR|31|11|praecepit igitur Ezechias ut praepararent horrea in domo Domini quod cum fecissent
2CHR|31|12|intulerunt tam primitias quam decimas et quaecumque voverant fideliter fuit autem praefectus eorum Chonenias Levita et Semei frater eius secundus
2CHR|31|13|post quem Ieihel et Azazias et Naath et Asahel et Ierimoth Iozabath quoque et Helihel et Iesmachias et Maath et Banaias praepositi sub manibus Choneniae et Semei fratris eius ex imperio Ezechiae regis et Azariae pontificis domus Domini ad quos omnia pertinebant
2CHR|31|14|Core vero filius Iemna Levites et ianitor orientalis portae praepositus erat his quae sponte offerebantur Domino primitiisque et consecratis in sancta sanctorum
2CHR|31|15|et sub cura eius Eden et Meniamin Hiesue et Sameias Amarias quoque et Sechenias in civitatibus sacerdotum ut fideliter distribuerent fratribus suis partes minoribus atque maioribus
2CHR|31|16|exceptis maribus ab annis tribus et supra cunctis qui ingrediebantur templum Domini et quicquid per dies singulos conducebat in ministerio atque observationibus iuxta divisiones suas
2CHR|31|17|sacerdotibus per familias et Levitis a vicesimo anno et supra per ordines et turmas suas
2CHR|31|18|universaeque multitudini tam uxoribus quam liberis eorum utriusque sexus fideliter cibi de his quae sanctificata fuerant praebebantur
2CHR|31|19|sed et filiorum Aaron per agros et suburbana urbium singularum dispositi erant viri qui partes distribuerent universo sexui masculino de sacerdotibus et Levitis
2CHR|31|20|fecit ergo Ezechias universa quae diximus in omni Iuda operatusque est bonum et rectum et verum coram Domino Deo suo
2CHR|31|21|in universa cultura ministerii domus Domini iuxta legem et caerimonias volens requirere Deum suum in toto corde suo fecitque et prosperatus est
2CHR|32|1|post quae et huiuscemodi veritatem venit Sennacherib rex Assyriorum et ingressus Iudam obsedit civitates munitas volens eas capere
2CHR|32|2|quod cum vidisset Ezechias venisse scilicet Sennacherib et totum belli impetum verti contra Hierusalem
2CHR|32|3|inito cum principibus consilio virisque fortissimis ut obturarent capita fontium quae erant extra urbem et hoc omnium decernente sententia
2CHR|32|4|congregavit plurimam multitudinem et obturaverunt cunctos fontes et rivum qui fluebat in medio terrae dicentes ne veniant reges Assyriorum et inveniant aquarum abundantiam
2CHR|32|5|aedificavit quoque agens industrie omnem murum qui fuerat dissipatus et extruxit turres desuper et forinsecus alterum murum instauravitque Mello in civitate David et fecit universi generis armaturam et clypeos
2CHR|32|6|constituitque principes bellatorum in exercitu et convocavit universos in platea portae civitatis ac locutus est ad cor eorum dicens
2CHR|32|7|viriliter agite et confortamini nolite timere nec paveatis regem Assyriorum et universam multitudinem quae est cum eo multo enim plures nobiscum sunt quam cum illo
2CHR|32|8|cum illo est brachium carneum nobiscum Dominus Deus noster qui auxiliator est noster pugnatque pro nobis confortatusque est populus huiuscemodi verbis Ezechiae regis Iuda
2CHR|32|9|quae postquam gesta sunt misit Sennacherib rex Assyriorum servos suos Hierusalem ipse enim cum universo exercitu obsidebat Lachis ad Ezechiam regem Iuda et ad omnem populum qui erat in urbe dicens
2CHR|32|10|haec dicit Sennacherib rex Assyriorum in quo habentes fiduciam sedetis obsessi in Hierusalem
2CHR|32|11|num Ezechias decipit vos ut tradat morti in fame et siti adfirmans quod Dominus Deus vester liberet vos de manu regis Assyriorum
2CHR|32|12|numquid non iste est Ezechias qui destruxit excelsa illius et altaria et praecepit Iudae et Hierusalem dicens coram altari uno adorabitis et in ipso conburetis incensum
2CHR|32|13|an ignoratis quae ego fecerim et patres mei cunctis terrarum populis numquid praevaluerunt dii gentium omniumque terrarum liberare regionem suam de manu mea
2CHR|32|14|quis est de universis diis gentium quas vastaverunt patres mei qui potuerit eruere populum suum de manu mea ut possit etiam Deus vester eruere vos de hac manu
2CHR|32|15|non vos ergo decipiat Ezechias nec vana persuasione deludat neque credatis ei si enim nullus potuit deus cunctarum gentium atque regnorum liberare populum suum de manu mea et de manu patrum meorum consequenter nec Deus vester poterit eruere vos de hac manu
2CHR|32|16|sed et alia multa locuti sunt servi eius contra Dominum Deum et contra Ezechiam servum eius
2CHR|32|17|epistulas quoque scripsit plenas blasphemiae in Dominum Deum Israhel et locutus est adversus eum sicut dii gentium ceterarum non potuerunt liberare populos suos de manu mea sic et Deus Ezechiae eruere non poterit populum suum de manu ista
2CHR|32|18|insuper et clamore magno lingua iudaica contra populum qui sedebat in muris Hierusalem personabat ut terreret eos et caperet civitatem
2CHR|32|19|locutusque est contra Deum Hierusalem sicut adversum deos populorum terrae opera manuum hominum
2CHR|32|20|oraverunt igitur Ezechias rex et Esaias filius Amos prophetes adversum hanc blasphemiam ac vociferati sunt usque in caelum
2CHR|32|21|et misit Dominus angelum qui percussit omnem virum robustum et bellatorem et principem exercitus regis Assyriorum reversusque est cum ignominia in terram suam cumque ingressus esset domum dei sui filii qui egressi fuerant de utero eius interfecerunt eum gladio
2CHR|32|22|salvavitque Dominus Ezechiam et habitatores Hierusalem de manu Sennacherib regis Assyriorum et de manu omnium et praestitit ei quietem per circuitum
2CHR|32|23|multi etiam deferebant hostias et sacrificia Domino Hierusalem et munera Ezechiae regi Iuda qui exaltatus est post haec coram cunctis gentibus
2CHR|32|24|in diebus illis aegrotavit Ezechias usque ad mortem et oravit Dominum exaudivitque eum et dedit ei signum
2CHR|32|25|sed non iuxta beneficia quae acceperat retribuit quia elevatum est cor eius et facta est contra eum ira et contra Iudam ac Hierusalem
2CHR|32|26|humiliatusque est postea eo quod exaltatum fuisset cor eius tam ipse quam habitatores Hierusalem et idcirco non venit super eos ira Domini in diebus Ezechiae
2CHR|32|27|fuit autem Ezechias dives et inclitus valde et thesauros sibi plurimos congregavit argenti auri et lapidis pretiosi aromatum et armorum universi generis et vasorum magni pretii
2CHR|32|28|apothecas quoque frumenti vini et olei et praesepia omnium iumentorum caulasque pecoribus
2CHR|32|29|et urbes exaedificavit habebat quippe greges ovium et armentorum innumerabiles eo quod dedisset ei Dominus substantiam multam nimis
2CHR|32|30|ipse est Ezechias qui obturavit superiorem fontem aquarum Gion et avertit eas subter ad occidentem urbis David in omnibus operibus suis fecit prospere quae voluit
2CHR|32|31|attamen in legatione principum Babylonis qui missi fuerant ad eum ut interrogarent de portento quod acciderat super terram dereliquit eum Deus ut temptaretur et nota fierent omnia quae erant in corde eius
2CHR|32|32|reliqua autem sermonum Ezechiae et misericordiarum eius scripta sunt in visione Esaiae filii Amos prophetae et in libro regum Iuda et Israhel
2CHR|32|33|dormivitque Ezechias cum patribus suis et sepelierunt eum supra sepulchra filiorum David et celebravit eius exequias universus Iuda et omnes habitatores Hierusalem regnavitque Manasses filius eius pro eo
2CHR|33|1|duodecim annorum erat Manasses cum regnare coepisset et quinquaginta quinque annis regnavit in Hierusalem
2CHR|33|2|fecit autem malum coram Domino iuxta abominationes gentium quas subvertit Dominus coram filiis Israhel
2CHR|33|3|et conversus instauravit excelsa quae demolitus fuerat Ezechias pater eius construxitque aras Baalim et fecit lucos et adoravit omnem militiam caeli et coluit eam
2CHR|33|4|aedificavit quoque altaria in domo Domini de qua dixerat Dominus in Hierusalem erit nomen meum in aeternum
2CHR|33|5|aedificavit autem ea cuncto exercitui caeli in duobus atriis domus Domini
2CHR|33|6|transireque fecit filios suos per ignem in valle Benennon observabat somnia sectabatur auguria maleficis artibus inserviebat habebat secum magos et incantatores multaque mala operatus est coram Domino ut inritaret eum
2CHR|33|7|sculptile quoque et conflatile signum posuit in domo Domini de qua locutus est Dominus ad David et ad Salomonem filium eius dicens in domo hac et in Hierusalem quam elegi de cunctis tribubus Israhel ponam nomen meum in sempiternum
2CHR|33|8|et movere non faciam pedem Israhel de terra quam tradidi patribus eorum ita dumtaxat si custodierint facere quae praecepi eis cunctamque legem et caerimonias atque iudicia per manum Mosi
2CHR|33|9|igitur Manasses seduxit Iudam et habitatores Hierusalem ut facerent malum super omnes gentes quas subverterat Dominus a facie filiorum Israhel
2CHR|33|10|locutusque est Dominus ad eum et ad populum illius et adtendere noluerunt
2CHR|33|11|idcirco superinduxit eis principes exercitus regis Assyriorum ceperuntque Manassen et vinctum catenis atque conpedibus duxerunt Babylonem
2CHR|33|12|qui postquam coangustatus est oravit Dominum Deum suum et egit paenitentiam valde coram Deo patrum suorum
2CHR|33|13|deprecatusque est eum et obsecravit intente et exaudivit orationem eius reduxitque eum Hierusalem in regnum suum et cognovit Manasses quod Dominus ipse esset Deus
2CHR|33|14|post haec aedificavit murum extra civitatem David ad occidentem Gion in convalle ab introitu portae Piscium per circuitum usque ad Ophel et exaltavit illum vehementer constituitque principes exercitus in cunctis civitatibus Iuda munitis
2CHR|33|15|et abstulit deos alienos et simulacrum de domo Domini aras quoque quas fecerat in monte domus Domini et in Hierusalem et proiecit omnia extra urbem
2CHR|33|16|porro instauravit altare Domini et immolavit super illud victimas et pacifica et laudem praecepitque Iudae ut serviret Domino Deo Israhel
2CHR|33|17|attamen adhuc populus immolabat in excelsis Domino Deo suo
2CHR|33|18|reliqua autem gestorum Manasse et obsecratio eius ad Deum suum verba quoque videntium qui loquebantur ad eum in nomine Domini Dei Israhel continentur in sermonibus regum Israhel
2CHR|33|19|oratio quoque eius et exauditio et cuncta peccata atque contemptus loca etiam in quibus aedificavit excelsa et fecit lucos et statuas antequam ageret paenitentiam scripta sunt in sermonibus Ozai
2CHR|33|20|dormivit ergo Manasses cum patribus suis et sepelierunt eum in domo sua regnavitque pro eo filius eius Amon
2CHR|33|21|viginti duo annorum erat Amon cum regnare coepisset et duobus annis regnavit in Hierusalem
2CHR|33|22|fecitque malum in conspectu Domini sicut fecerat Manasses pater eius et cunctis idolis quae Manasses fuerat fabricatus immolavit atque servivit
2CHR|33|23|et non est reveritus faciem Domini sicut reveritus est Manasses pater eius et multo maiora deliquit
2CHR|33|24|cumque coniurassent adversus eum servi sui interfecerunt eum in domo sua
2CHR|33|25|porro reliqua populi multitudo caesis his qui Amon percusserant constituit regem Iosiam filium eius pro eo
2CHR|34|1|octo annorum erat Iosias cum regnare coepisset et triginta et uno annis regnavit in Hierusalem
2CHR|34|2|fecitque quod erat rectum in conspectu Domini et ambulavit in viis David patris sui non declinavit neque ad dexteram neque ad sinistram
2CHR|34|3|octavo autem anno regni sui cum adhuc esset puer coepit quaerere Deum patris sui David et duodecimo anno postquam coeperat mundavit Iudam et Hierusalem ab excelsis et lucis simulacrisque et sculptilibus
2CHR|34|4|destruxeruntque coram eo aras Baalim et simulacra quae superposita fuerant demoliti sunt lucos etiam et sculptilia succidit atque comminuit et super tumulos eorum qui eis immolare consueverant fragmenta dispersit
2CHR|34|5|ossa praeterea sacerdotum conbusit in altaribus idolorum mundavitque Iudam et Hierusalem
2CHR|34|6|sed et in urbibus Manasse et Ephraim et Symeon usque Nepthalim cuncta subvertit
2CHR|34|7|cumque altaria dissipasset et lucos et sculptilia contrivisset in frusta cunctaque delubra demolitus esset de universa terra Israhel reversus est Hierusalem
2CHR|34|8|igitur anno octavodecimo regni sui mundata iam terra et templo Domini misit Saphan filium Eseliae et Maasiam principem civitatis et Ioha filium Ioachaz a commentariis ut instaurarent domum Domini Dei sui
2CHR|34|9|qui venerunt ad Helciam sacerdotem magnum acceptamque ab eo pecuniam quae inlata fuerat in domum Domini et quam congregaverant Levitae ianitores de Manasse et Ephraim et universis reliquiis Israhel ab omni quoque Iuda et Beniamin et habitatoribus Hierusalem
2CHR|34|10|tradiderunt in manibus eorum qui praeerant operariis in domo Domini ut instaurarent templum et infirma quaeque sarcirent
2CHR|34|11|at illi dederunt eam artificibus et cementariis ut emerent lapides de lapidicinis et ligna ad commissuras aedificii et ad contignationem domorum quas destruxerant reges Iuda
2CHR|34|12|qui fideliter cuncta faciebant erant autem praepositi operantium Iaath et Abdias de filiis Merari Zaccharias et Mosollam de filiis Caath qui urguebant opus omnes Levitae scientes organis canere
2CHR|34|13|super eos vero qui ad varios usus onera portabant erant scribae et magistri de Levitis ianitores
2CHR|34|14|cumque efferrent pecuniam quae inlata fuerat in templum Domini repperit Helcias sacerdos librum legis Domini per manum Mosi
2CHR|34|15|et ait ad Saphan scribam librum legis inveni in domo Domini et tradidit ei
2CHR|34|16|at ille intulit volumen ad regem et nuntiavit ei dicens omnia quae dedisti in manu servorum tuorum ecce conplentur
2CHR|34|17|argentum quod reppertum est in domo Domini conflaverunt datumque est praefectis artificum et diversa opera fabricantium
2CHR|34|18|praeterea tradidit mihi Helcias sacerdos hunc librum quem cum rege praesente recitasset
2CHR|34|19|audissetque ille verba legis scidit vestimenta sua
2CHR|34|20|et praecepit Helciae et Ahicam filio Saphan et Abdon filio Micha Saphan quoque scribae et Asaiae servo regis dicens
2CHR|34|21|ite et orate Dominum pro me et pro reliquiis Israhel et Iuda super universis sermonibus libri istius qui reppertus est magnus enim furor Domini stillavit super nos eo quod non custodierint patres nostri verba Domini ut facerent omnia quae scripta sunt in isto volumine
2CHR|34|22|abiit igitur Helcias et hii qui simul a rege missi fuerant ad Holdan propheten uxorem Sellum filii Thecuath filii Hasra custodis vestium quae habitabat Hierusalem in secunda et locuti sunt ei verba quae supra narravimus
2CHR|34|23|at illa respondit eis haec dicit Dominus Deus Israhel dicite viro qui misit vos ad me
2CHR|34|24|haec dicit Dominus ecce ego inducam mala super locum istum et super habitatores eius cunctaque maledicta quae scripta sunt in libro hoc quem legerunt coram rege Iuda
2CHR|34|25|quia dereliquerunt me et sacrificaverunt diis alienis ut me ad iracundiam provocarent in cunctis operibus manuum suarum idcirco stillavit furor meus super locum istum et non extinguetur
2CHR|34|26|ad regem autem Iuda qui misit vos pro Domino deprecando sic loquimini haec dicit Dominus Deus Israhel quoniam audisti verba voluminis
2CHR|34|27|atque emollitum est cor tuum et humiliatus es in conspectu Dei super his quae dicta sunt contra locum hunc et habitatores Hierusalem reveritusque faciem meam scidisti vestimenta tua et flevisti coram me ego quoque exaudivi te dicit Dominus
2CHR|34|28|iam enim colligam te ad patres tuos et infereris in sepulchrum tuum in pace nec videbunt oculi tui omne malum quod ego inducturus sum super locum istum et super habitatores eius rettulerunt itaque regi cuncta quae dixerat
2CHR|34|29|at ille convocatis universis maioribus natu Iuda et Hierusalem
2CHR|34|30|ascendit domum Domini unaque omnes viri Iuda et habitatores Hierusalem sacerdotes et Levitae et cunctus populus a minimo usque ad maximum quibus audientibus in domo Domini legit rex omnia verba voluminis
2CHR|34|31|et stans in tribunali suo percussit foedus coram Domino ut ambularet post eum et custodiret praecepta et testimonia et iustificationes eius in toto corde suo et in tota anima sua faceretque quae scripta sunt in volumine illo quem legerat
2CHR|34|32|adiuravit quoque super hoc omnes qui repperti fuerant in Hierusalem et Beniamin et fecerunt habitatores Hierusalem iuxta pactum Domini Dei patrum suorum
2CHR|34|33|abstulit ergo Iosias cunctas abominationes de universis regionibus filiorum Israhel et fecit omnes qui residui erant in Israhel servire Domino Deo suo cunctis diebus eius non recesserunt a Domino Deo patrum suorum
2CHR|35|1|fecit autem Iosias in Hierusalem phase Domino quod immolatum est quartadecima die mensis primi
2CHR|35|2|et constituit sacerdotes in officiis suis hortatusque est eos ut ministrarent in domo Domini
2CHR|35|3|Levitis quoque ad quorum eruditionem omnis Israhel sanctificabatur Domino locutus est ponite arcam in sanctuario templi quod aedificavit Salomon filius David rex Israhel nequaquam enim eam ultra portabitis nunc autem ministrate Domino Deo vestro et populo eius Israhel
2CHR|35|4|et praeparate vos per domos et cognationes vestras in divisionibus singulorum sicut praecepit David rex Israhel et descripsit Salomon filius eius
2CHR|35|5|ministrate in sanctuario per familias turmasque leviticas
2CHR|35|6|et sanctificati immolate phase fratres etiam vestros ut possint iuxta verba quae locutus est Dominus in manu Mosi facere praeparate
2CHR|35|7|dedit praeterea Iosias omni populo qui ibi fuerat inventus in sollemnitatem phase agnos et hedos de gregibus et reliqui pecoris triginta milia boumque tria milia haec de regis universa substantia
2CHR|35|8|duces quoque eius sponte quod voluerant obtulerunt tam populo quam sacerdotibus et Levitis porro Helcias et Zaccharias et Iehihel principes domus Domini dederunt sacerdotibus ad faciendum phase pecora commixtim duo milia sescenta et boves trecentos
2CHR|35|9|Chonenias autem Semeias etiam et Nathanahel fratres eius necnon Asabias et Iahihel et Iozabath principes Levitarum dederunt ceteris Levitis ad celebrandum phase quinque milia pecorum et boves quingentos
2CHR|35|10|praeparatumque est ministerium et steterunt sacerdotes in officio suo Levitae quoque in turmis iuxta regis imperium
2CHR|35|11|et immolatum est phase asperseruntque sacerdotes manu sua sanguinem et Levitae detraxerunt pelles holocaustorum
2CHR|35|12|et separaverunt ea ut darent per domos et familias singulorum et offerrentur Domino sicut scriptum est in libro Mosi de bubus quoque fecere similiter
2CHR|35|13|et assaverunt phase super ignem iuxta quod lege praeceptum est pacificas vero hostias coxerunt in lebetis et caccabis et ollis et festinato distribuerunt universae plebi
2CHR|35|14|sibi autem et sacerdotibus postea paraverunt nam in oblatione holocaustorum et adipum usque ad noctem sacerdotes fuerant occupati unde Levitae et sibi et sacerdotibus filiis Aaron paraverunt novissimis
2CHR|35|15|porro cantores filii Asaph stabant in ordine suo iuxta praeceptum David et Asaph et Heman et Idithun prophetarum regis ianitores vero per portas singulas observabant ita ut ne puncto quidem discederent a ministerio quam ob rem et fratres eorum Levitae paraverunt eis cibos
2CHR|35|16|omnis igitur cultura Domini rite conpleta est in die illa ut facerent phase et offerrent holocausta super altare Domini iuxta praeceptum regis Iosiae
2CHR|35|17|feceruntque filii Israhel qui repperti fuerant ibi phase in tempore illo et sollemnitatem azymorum septem diebus
2CHR|35|18|non fuit phase simile huic in Israhel a diebus Samuhelis prophetae sed nec quisquam de cunctis regibus Israhel fecit phase sicut Iosias sacerdotibus et Levitis et omni Iuda et Israhel qui reppertus fuerat et habitantibus in Hierusalem
2CHR|35|19|octavodecimo anno regni Iosiae hoc phase celebratum est
2CHR|35|20|postquam instauraverat Iosias templum ascendit Nechao rex Aegypti ad pugnandum in Charchamis iuxta Eufraten et processit in occursum eius Iosias
2CHR|35|21|at ille missis ad eum nuntiis ait quid mihi et tibi est rex Iuda non adversum te hodie venio sed contra aliam pugno domum ad quam me Deus festinato ire praecepit desine adversum Deum facere qui mecum est ne interficiat te
2CHR|35|22|noluit Iosias reverti sed praeparavit contra eum bellum nec adquievit sermonibus Nechao ex ore Dei verum perrexit ut dimicaret in campo Mageddo
2CHR|35|23|ibique vulneratus a sagittariis dixit pueris suis educite me de proelio quia oppido vulneratus sum
2CHR|35|24|qui transtulerunt eum de curru in alterum currum qui sequebatur eum more regio et asportaverunt in Hierusalem mortuusque est et sepultus in mausoleo patrum suorum et universus Iuda et Hierusalem luxerunt eum
2CHR|35|25|Hieremias maxime cuius omnes cantores atque cantrices usque in praesentem diem lamentationes super Iosia replicant et quasi lex obtinuit in Israhel ecce scriptum fertur in Lamentationibus
2CHR|35|26|reliqua autem sermonum Iosiae et misericordiarum eius quae lege praecepta sunt Domini
2CHR|35|27|opera quoque illius prima et novissima scripta sunt in libro regum Israhel et Iuda
2CHR|36|1|tulit ergo populus terrae Ioachaz filium Iosiae et constituit regem pro patre suo in Hierusalem
2CHR|36|2|viginti trium annorum erat Ioachaz cum regnare coepisset et tribus mensibus regnavit in Hierusalem
2CHR|36|3|amovit autem eum rex Aegypti cum venisset Hierusalem et condemnavit terram centum talentis argenti et talento auri
2CHR|36|4|constituitque regem pro eo Eliacim fratrem eius super Iudam et Hierusalem et vertit nomen eius Ioacim ipsum vero Ioachaz tulit secum et adduxit in Aegyptum
2CHR|36|5|viginti quinque annorum erat Ioacim cum regnare coepisset et undecim annis regnavit in Hierusalem fecitque malum coram Domino Deo suo
2CHR|36|6|contra hunc ascendit Nabuchodonosor rex Chaldeorum et vinctum catenis duxit in Babylonem
2CHR|36|7|ad quam et vasa Domini transtulit et posuit ea in templo suo
2CHR|36|8|reliqua autem verborum Ioacim et abominationum eius quas operatus est et quae inventa sunt in eo continentur in libro regum Israhel et Iuda regnavitque Ioachin filius eius pro eo
2CHR|36|9|octo annorum erat Ioachin cum regnare coepisset et tribus mensibus ac decem diebus regnavit in Hierusalem fecitque malum in conspectu Domini
2CHR|36|10|cumque anni circulus volveretur misit Nabuchodonosor rex qui et adduxerunt eum in Babylonem asportatis simul pretiosissimis vasis domus Domini regem vero constituit Sedeciam fratrem eius super Iudam et Hierusalem
2CHR|36|11|viginti et unius anni erat Sedecias cum regnare coepisset et undecim annis regnavit in Hierusalem
2CHR|36|12|fecitque malum in oculis Domini Dei sui nec erubuit faciem Hieremiae prophetae loquentis ad se ex ore Domini
2CHR|36|13|a rege quoque Nabuchodonosor recessit qui adiuraverat eum per Deum et induravit cervicem suam et cor ut non reverteretur ad Dominum Deum Israhel
2CHR|36|14|sed et universi principes sacerdotum et populus praevaricati sunt inique iuxta universas abominationes gentium et polluerunt domum Domini quam sanctificaverat sibi in Hierusalem
2CHR|36|15|mittebat autem Dominus Deus patrum suorum ad illos per manum nuntiorum suorum de nocte consurgens et cotidie commonens eo quod parceret populo et habitaculo suo
2CHR|36|16|at illi subsannabant nuntios Dei et parvipendebant sermones eius inludebantque prophetis donec ascenderet furor Domini in populum eius et esset nulla curatio
2CHR|36|17|adduxit enim super eos regem Chaldeorum et interfecit iuvenes eorum gladio in domo sanctuarii sui non est misertus adulescentis et virginis et senis nec decrepiti quidem sed omnes tradidit manibus eius
2CHR|36|18|universaque vasa domus Domini tam maiora quam minora et thesauros templi et regis et principum transtulit in Babylonem
2CHR|36|19|incenderunt hostes domum Dei destruxerunt murum Hierusalem universas turres conbuserunt et quicquid pretiosum fuerat demoliti sunt
2CHR|36|20|si quis evaserat gladium ductus in Babylonem servivit regi et filiis eius donec imperaret rex Persarum
2CHR|36|21|et conpleretur sermo Domini ex ore Hieremiae et celebraret terra sabbata sua cunctis enim diebus desolationis egit sabbatum usque dum conplerentur septuaginta anni
2CHR|36|22|anno autem primo Cyri regis Persarum ad explendum sermonem Domini quem locutus fuerat per os Hieremiae suscitavit Dominus spiritum Cyri regis Persarum qui iussit praedicari in universo regno suo etiam per scripturam dicens
2CHR|36|23|haec dicit Cyrus rex Persarum omnia regna terrae dedit mihi Dominus Deus caeli et ipse praecepit mihi ut aedificarem ei domum in Hierusalem quae est in Iudaea quis ex vobis est in omni populo eius sit Dominus Deus suus cum eo et ascendat
