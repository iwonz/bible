HOS|1|1|The word of the LORD that came unto Hosea, the son of Beeri, in the days of Uzziah, Jotham, Ahaz, and Hezekiah, kings of Judah, and in the days of Jeroboam the son of Joash, king of Israel.
HOS|1|2|The beginning of the word of the LORD by Hosea. And the LORD said to Hosea, Go, take unto thee a wife of whoredoms and children of whoredoms: for the land hath committed great whoredom, departing from the LORD.
HOS|1|3|So he went and took Gomer the daughter of Diblaim; which conceived, and bare him a son.
HOS|1|4|And the LORD said unto him, Call his name Jezreel; for yet a little while, and I will avenge the blood of Jezreel upon the house of Jehu, and will cause to cease the kingdom of the house of Israel.
HOS|1|5|And it shall come to pass at that day, that I will break the bow of Israel, in the valley of Jezreel.
HOS|1|6|And she conceived again, and bare a daughter. And God said unto him, Call her name Loruhamah: for I will no more have mercy upon the house of Israel; but I will utterly take them away.
HOS|1|7|But I will have mercy upon the house of Judah, and will save them by the LORD their God, and will not save them by bow, nor by sword, nor by battle, by horses, nor by horsemen.
HOS|1|8|Now when she had weaned Loruhamah, she conceived, and bare a son.
HOS|1|9|Then said God, Call his name Loammi: for ye are not my people, and I will not be your God.
HOS|1|10|Yet the number of the children of Israel shall be as the sand of the sea, which cannot be measured nor numbered; and it shall come to pass, that in the place where it was said unto them, Ye are not my people, there it shall be said unto them, Ye are the sons of the living God.
HOS|1|11|Then shall the children of Judah and the children of Israel be gathered together, and appoint themselves one head, and they shall come up out of the land: for great shall be the day of Jezreel.
HOS|2|1|Say ye unto your brethren, Ammi; and to your sisters, Ruhamah.
HOS|2|2|Plead with your mother, plead: for she is not my wife, neither am I her husband: let her therefore put away her whoredoms out of her sight, and her adulteries from between her breasts;
HOS|2|3|Lest I strip her naked, and set her as in the day that she was born, and make her as a wilderness, and set her like a dry land, and slay her with thirst.
HOS|2|4|And I will not have mercy upon her children; for they be the children of whoredoms.
HOS|2|5|For their mother hath played the harlot: she that conceived them hath done shamefully: for she said, I will go after my lovers, that give me my bread and my water, my wool and my flax, mine oil and my drink.
HOS|2|6|Therefore, behold, I will hedge up thy way with thorns, and make a wall, that she shall not find her paths.
HOS|2|7|And she shall follow after her lovers, but she shall not overtake them; and she shall seek them, but shall not find them: then shall she say, I will go and return to my first husband; for then was it better with me than now.
HOS|2|8|For she did not know that I gave her corn, and wine, and oil, and multiplied her silver and gold, which they prepared for Baal.
HOS|2|9|Therefore will I return, and take away my corn in the time thereof, and my wine in the season thereof, and will recover my wool and my flax given to cover her nakedness.
HOS|2|10|And now will I discover her lewdness in the sight of her lovers, and none shall deliver her out of mine hand.
HOS|2|11|I will also cause all her mirth to cease, her feast days, her new moons, and her sabbaths, and all her solemn feasts.
HOS|2|12|And I will destroy her vines and her fig trees, whereof she hath said, These are my rewards that my lovers have given me: and I will make them a forest, and the beasts of the field shall eat them.
HOS|2|13|And I will visit upon her the days of Baalim, wherein she burned incense to them, and she decked herself with her earrings and her jewels, and she went after her lovers, and forgat me, saith the LORD.
HOS|2|14|Therefore, behold, I will allure her, and bring her into the wilderness, and speak comfortably unto her.
HOS|2|15|And I will give her her vineyards from thence, and the valley of Achor for a door of hope: and she shall sing there, as in the days of her youth, and as in the day when she came up out of the land of Egypt.
HOS|2|16|And it shall be at that day, saith the LORD, that thou shalt call me Ishi; and shalt call me no more Baali.
HOS|2|17|For I will take away the names of Baalim out of her mouth, and they shall no more be remembered by their name.
HOS|2|18|And in that day will I make a covenant for them with the beasts of the field and with the fowls of heaven, and with the creeping things of the ground: and I will break the bow and the sword and the battle out of the earth, and will make them to lie down safely.
HOS|2|19|And I will betroth thee unto me for ever; yea, I will betroth thee unto me in righteousness, and in judgment, and in lovingkindness, and in mercies.
HOS|2|20|I will even betroth thee unto me in faithfulness: and thou shalt know the LORD.
HOS|2|21|And it shall come to pass in that day, I will hear, saith the LORD, I will hear the heavens, and they shall hear the earth;
HOS|2|22|And the earth shall hear the corn, and the wine, and the oil; and they shall hear Jezreel.
HOS|2|23|And I will sow her unto me in the earth; and I will have mercy upon her that had not obtained mercy; and I will say to them which were not my people, Thou art my people; and they shall say, Thou art my God.
HOS|3|1|Then said the LORD unto me, Go yet, love a woman beloved of her friend, yet an adulteress, according to the love of the LORD toward the children of Israel, who look to other gods, and love flagons of wine.
HOS|3|2|So I bought her to me for fifteen pieces of silver, and for an homer of barley, and an half homer of barley:
HOS|3|3|And I said unto her, Thou shalt abide for me many days; thou shalt not play the harlot, and thou shalt not be for another man: so will I also be for thee.
HOS|3|4|For the children of Israel shall abide many days without a king, and without a prince, and without a sacrifice, and without an image, and without an ephod, and without teraphim:
HOS|3|5|Afterward shall the children of Israel return, and seek the LORD their God, and David their king; and shall fear the LORD and his goodness in the latter days.
HOS|4|1|Hear the word of the LORD, ye children of Israel: for the LORD hath a controversy with the inhabitants of the land, because there is no truth, nor mercy, nor knowledge of God in the land.
HOS|4|2|By swearing, and lying, and killing, and stealing, and committing adultery, they break out, and blood toucheth blood.
HOS|4|3|Therefore shall the land mourn, and every one that dwelleth therein shall languish, with the beasts of the field, and with the fowls of heaven; yea, the fishes of the sea also shall be taken away.
HOS|4|4|Yet let no man strive, nor reprove another: for thy people are as they that strive with the priest.
HOS|4|5|Therefore shalt thou fall in the day, and the prophet also shall fall with thee in the night, and I will destroy thy mother.
HOS|4|6|My people are destroyed for lack of knowledge: because thou hast rejected knowledge, I will also reject thee, that thou shalt be no priest to me: seeing thou hast forgotten the law of thy God, I will also forget thy children.
HOS|4|7|As they were increased, so they sinned against me: therefore will I change their glory into shame.
HOS|4|8|They eat up the sin of my people, and they set their heart on their iniquity.
HOS|4|9|And there shall be, like people, like priest: and I will punish them for their ways, and reward them their doings.
HOS|4|10|For they shall eat, and not have enough: they shall commit whoredom, and shall not increase: because they have left off to take heed to the LORD.
HOS|4|11|Whoredom and wine and new wine take away the heart.
HOS|4|12|My people ask counsel at their stocks, and their staff declareth unto them: for the spirit of whoredoms hath caused them to err, and they have gone a whoring from under their God.
HOS|4|13|They sacrifice upon the tops of the mountains, and burn incense upon the hills, under oaks and poplars and elms, because the shadow thereof is good: therefore your daughters shall commit whoredom, and your spouses shall commit adultery.
HOS|4|14|I will not punish your daughters when they commit whoredom, nor your spouses when they commit adultery: for themselves are separated with whores, and they sacrifice with harlots: therefore the people that doth not understand shall fall.
HOS|4|15|Though thou, Israel, play the harlot, yet let not Judah offend; and come not ye unto Gilgal, neither go ye up to Bethaven, nor swear, The LORD liveth.
HOS|4|16|For Israel slideth back as a backsliding heifer: now the LORD will feed them as a lamb in a large place.
HOS|4|17|Ephraim is joined to idols: let him alone.
HOS|4|18|Their drink is sour: they have committed whoredom continually: her rulers with shame do love, Give ye.
HOS|4|19|The wind hath bound her up in her wings, and they shall be ashamed because of their sacrifices.
HOS|5|1|Hear ye this, O priests; and hearken, ye house of Israel; and give ye ear, O house of the king; for judgment is toward you, because ye have been a snare on Mizpah, and a net spread upon Tabor.
HOS|5|2|And the revolters are profound to make slaughter, though I have been a rebuker of them all.
HOS|5|3|I know Ephraim, and Israel is not hid from me: for now, O Ephraim, thou committest whoredom, and Israel is defiled.
HOS|5|4|They will not frame their doings to turn unto their God: for the spirit of whoredoms is in the midst of them, and they have not known the LORD.
HOS|5|5|And the pride of Israel doth testify to his face: therefore shall Israel and Ephraim fall in their iniquity: Judah also shall fall with them.
HOS|5|6|They shall go with their flocks and with their herds to seek the LORD; but they shall not find him; he hath withdrawn himself from them.
HOS|5|7|They have dealt treacherously against the LORD: for they have begotten strange children: now shall a month devour them with their portions.
HOS|5|8|Blow ye the cornet in Gibeah, and the trumpet in Ramah: cry aloud at Bethaven, after thee, O Benjamin.
HOS|5|9|Ephraim shall be desolate in the day of rebuke: among the tribes of Israel have I made known that which shall surely be.
HOS|5|10|The princes of Judah were like them that remove the bound: therefore I will pour out my wrath upon them like water.
HOS|5|11|Ephraim is oppressed and broken in judgment, because he willingly walked after the commandment.
HOS|5|12|Therefore will I be unto Ephraim as a moth, and to the house of Judah as rottenness.
HOS|5|13|When Ephraim saw his sickness, and Judah saw his wound, then went Ephraim to the Assyrian, and sent to king Jareb: yet could he not heal you, nor cure you of your wound.
HOS|5|14|For I will be unto Ephraim as a lion, and as a young lion to the house of Judah: I, even I, will tear and go away; I will take away, and none shall rescue him.
HOS|5|15|I will go and return to my place, till they acknowledge their offence, and seek my face: in their affliction they will seek me early.
HOS|6|1|Come, and let us return unto the LORD: for he hath torn, and he will heal us; he hath smitten, and he will bind us up.
HOS|6|2|After two days will he revive us: in the third day he will raise us up, and we shall live in his sight.
HOS|6|3|Then shall we know, if we follow on to know the LORD: his going forth is prepared as the morning; and he shall come unto us as the rain, as the latter and former rain unto the earth.
HOS|6|4|O Ephraim, what shall I do unto thee? O Judah, what shall I do unto thee? for your goodness is as a morning cloud, and as the early dew it goeth away.
HOS|6|5|Therefore have I hewed them by the prophets; I have slain them by the words of my mouth: and thy judgments are as the light that goeth forth.
HOS|6|6|For I desired mercy, and not sacrifice; and the knowledge of God more than burnt offerings.
HOS|6|7|But they like men have transgressed the covenant: there have they dealt treacherously against me.
HOS|6|8|Gilead is a city of them that work iniquity, and is polluted with blood.
HOS|6|9|And as troops of robbers wait for a man, so the company of priests murder in the way by consent: for they commit lewdness.
HOS|6|10|I have seen an horrible thing in the house of Israel: there is the whoredom of Ephraim, Israel is defiled.
HOS|6|11|Also, O Judah, he hath set an harvest for thee, when I returned the captivity of my people.
HOS|7|1|When I would have healed Israel, then the iniquity of Ephraim was discovered, and the wickedness of Samaria: for they commit falsehood; and the thief cometh in, and the troop of robbers spoileth without.
HOS|7|2|And they consider not in their hearts that I remember all their wickedness: now their own doings have beset them about; they are before my face.
HOS|7|3|They make the king glad with their wickedness, and the princes with their lies.
HOS|7|4|They are all adulterers, as an oven heated by the baker, who ceaseth from raising after he hath kneaded the dough, until it be leavened.
HOS|7|5|In the day of our king the princes have made him sick with bottles of wine; he stretched out his hand with scorners.
HOS|7|6|For they have made ready their heart like an oven, whiles they lie in wait: their baker sleepeth all the night; in the morning it burneth as a flaming fire.
HOS|7|7|They are all hot as an oven, and have devoured their judges; all their kings are fallen: there is none among them that calleth unto me.
HOS|7|8|Ephraim, he hath mixed himself among the people; Ephraim is a cake not turned.
HOS|7|9|Strangers have devoured his strength, and he knoweth it not: yea, gray hairs are here and there upon him, yet he knoweth not.
HOS|7|10|And the pride of Israel testifieth to his face: and they do not return to the LORD their God, nor seek him for all this.
HOS|7|11|Ephraim also is like a silly dove without heart: they call to Egypt, they go to Assyria.
HOS|7|12|When they shall go, I will spread my net upon them; I will bring them down as the fowls of the heaven; I will chastise them, as their congregation hath heard.
HOS|7|13|Woe unto them! for they have fled from me: destruction unto them! because they have transgressed against me: though I have redeemed them, yet they have spoken lies against me.
HOS|7|14|And they have not cried unto me with their heart, when they howled upon their beds: they assemble themselves for corn and wine, and they rebel against me.
HOS|7|15|Though I have bound and strengthened their arms, yet do they imagine mischief against me.
HOS|7|16|They return, but not to the most High: they are like a deceitful bow: their princes shall fall by the sword for the rage of their tongue: this shall be their derision in the land of Egypt.
HOS|8|1|Set the trumpet to thy mouth. He shall come as an eagle against the house of the LORD, because they have transgressed my covenant, and trespassed against my law.
HOS|8|2|Israel shall cry unto me, My God, we know thee.
HOS|8|3|Israel hath cast off the thing that is good: the enemy shall pursue him.
HOS|8|4|They have set up kings, but not by me: they have made princes, and I knew it not: of their silver and their gold have they made them idols, that they may be cut off.
HOS|8|5|Thy calf, O Samaria, hath cast thee off; mine anger is kindled against them: how long will it be ere they attain to innocency?
HOS|8|6|For from Israel was it also: the workman made it; therefore it is not God: but the calf of Samaria shall be broken in pieces.
HOS|8|7|For they have sown the wind, and they shall reap the whirlwind: it hath no stalk; the bud shall yield no meal: if so be it yield, the strangers shall swallow it up.
HOS|8|8|Israel is swallowed up: now shall they be among the Gentiles as a vessel wherein is no pleasure.
HOS|8|9|For they are gone up to Assyria, a wild ass alone by himself: Ephraim hath hired lovers.
HOS|8|10|Yea, though they have hired among the nations, now will I gather them, and they shall sorrow a little for the burden of the king of princes.
HOS|8|11|Because Ephraim hath made many altars to sin, altars shall be unto him to sin.
HOS|8|12|I have written to him the great things of my law, but they were counted as a strange thing.
HOS|8|13|They sacrifice flesh for the sacrifices of mine offerings, and eat it; but the LORD accepteth them not; now will he remember their iniquity, and visit their sins: they shall return to Egypt.
HOS|8|14|For Israel hath forgotten his Maker, and buildeth temples; and Judah hath multiplied fenced cities: but I will send a fire upon his cities, and it shall devour the palaces thereof.
HOS|9|1|Rejoice not, O Israel, for joy, as other people: for thou hast gone a whoring from thy God, thou hast loved a reward upon every cornfloor.
HOS|9|2|The floor and the winepress shall not feed them, and the new wine shall fail in her.
HOS|9|3|They shall not dwell in the LORD's land; but Ephraim shall return to Egypt, and they shall eat unclean things in Assyria.
HOS|9|4|They shall not offer wine offerings to the LORD, neither shall they be pleasing unto him: their sacrifices shall be unto them as the bread of mourners; all that eat thereof shall be polluted: for their bread for their soul shall not come into the house of the LORD.
HOS|9|5|What will ye do in the solemn day, and in the day of the feast of the LORD?
HOS|9|6|For, lo, they are gone because of destruction: Egypt shall gather them up, Memphis shall bury them: the pleasant places for their silver, nettles shall possess them: thorns shall be in their tabernacles.
HOS|9|7|The days of visitation are come, the days of recompence are come; Israel shall know it: the prophet is a fool, the spiritual man is mad, for the multitude of thine iniquity, and the great hatred.
HOS|9|8|The watchman of Ephraim was with my God: but the prophet is a snare of a fowler in all his ways, and hatred in the house of his God.
HOS|9|9|They have deeply corrupted themselves, as in the days of Gibeah: therefore he will remember their iniquity, he will visit their sins.
HOS|9|10|I found Israel like grapes in the wilderness; I saw your fathers as the firstripe in the fig tree at her first time: but they went to Baalpeor, and separated themselves unto that shame; and their abominations were according as they loved.
HOS|9|11|As for Ephraim, their glory shall fly away like a bird, from the birth, and from the womb, and from the conception.
HOS|9|12|Though they bring up their children, yet will I bereave them, that there shall not be a man left: yea, woe also to them when I depart from them!
HOS|9|13|Ephraim, as I saw Tyrus, is planted in a pleasant place: but Ephraim shall bring forth his children to the murderer.
HOS|9|14|Give them, O LORD: what wilt thou give? give them a miscarrying womb and dry breasts.
HOS|9|15|All their wickedness is in Gilgal: for there I hated them: for the wickedness of their doings I will drive them out of mine house, I will love them no more: all their princes are revolters.
HOS|9|16|Ephraim is smitten, their root is dried up, they shall bear no fruit: yea, though they bring forth, yet will I slay even the beloved fruit of their womb.
HOS|9|17|My God will cast them away, because they did not hearken unto him: and they shall be wanderers among the nations.
HOS|10|1|Israel is an empty vine, he bringeth forth fruit unto himself: according to the multitude of his fruit he hath increased the altars; according to the goodness of his land they have made goodly images.
HOS|10|2|Their heart is divided; now shall they be found faulty: he shall break down their altars, he shall spoil their images.
HOS|10|3|For now they shall say, We have no king, because we feared not the LORD; what then should a king do to us?
HOS|10|4|They have spoken words, swearing falsely in making a covenant: thus judgment springeth up as hemlock in the furrows of the field.
HOS|10|5|The inhabitants of Samaria shall fear because of the calves of Bethaven: for the people thereof shall mourn over it, and the priests thereof that rejoiced on it, for the glory thereof, because it is departed from it.
HOS|10|6|It shall be also carried unto Assyria for a present to king Jareb: Ephraim shall receive shame, and Israel shall be ashamed of his own counsel.
HOS|10|7|As for Samaria, her king is cut off as the foam upon the water.
HOS|10|8|The high places also of Aven, the sin of Israel, shall be destroyed: the thorn and the thistle shall come up on their altars; and they shall say to the mountains, Cover us; and to the hills, Fall on us.
HOS|10|9|O Israel, thou hast sinned from the days of Gibeah: there they stood: the battle in Gibeah against the children of iniquity did not overtake them.
HOS|10|10|It is in my desire that I should chastise them; and the people shall be gathered against them, when they shall bind themselves in their two furrows.
HOS|10|11|And Ephraim is as an heifer that is taught, and loveth to tread out the corn; but I passed over upon her fair neck: I will make Ephraim to ride; Judah shall plow, and Jacob shall break his clods.
HOS|10|12|Sow to yourselves in righteousness, reap in mercy; break up your fallow ground: for it is time to seek the LORD, till he come and rain righteousness upon you.
HOS|10|13|Ye have plowed wickedness, ye have reaped iniquity; ye have eaten the fruit of lies: because thou didst trust in thy way, in the multitude of thy mighty men.
HOS|10|14|Therefore shall a tumult arise among thy people, and all thy fortresses shall be spoiled, as Shalman spoiled Betharbel in the day of battle: the mother was dashed in pieces upon her children.
HOS|10|15|So shall Bethel do unto you because of your great wickedness: in a morning shall the king of Israel utterly be cut off.
HOS|11|1|When Israel was a child, then I loved him, and called my son out of Egypt.
HOS|11|2|As they called them, so they went from them: they sacrificed unto Baalim, and burned incense to graven images.
HOS|11|3|I taught Ephraim also to go, taking them by their arms; but they knew not that I healed them.
HOS|11|4|I drew them with cords of a man, with bands of love: and I was to them as they that take off the yoke on their jaws, and I laid meat unto them.
HOS|11|5|He shall not return into the land of Egypt, and the Assyrian shall be his king, because they refused to return.
HOS|11|6|And the sword shall abide on his cities, and shall consume his branches, and devour them, because of their own counsels.
HOS|11|7|And my people are bent to backsliding from me: though they called them to the most High, none at all would exalt him.
HOS|11|8|How shall I give thee up, Ephraim? how shall I deliver thee, Israel? how shall I make thee as Admah? how shall I set thee as Zeboim? mine heart is turned within me, my repentings are kindled together.
HOS|11|9|I will not execute the fierceness of mine anger, I will not return to destroy Ephraim: for I am God, and not man; the Holy One in the midst of thee: and I will not enter into the city.
HOS|11|10|They shall walk after the LORD: he shall roar like a lion: when he shall roar, then the children shall tremble from the west.
HOS|11|11|They shall tremble as a bird out of Egypt, and as a dove out of the land of Assyria: and I will place them in their houses, saith the LORD.
HOS|11|12|Ephraim compasseth me about with lies, and the house of Israel with deceit: but Judah yet ruleth with God, and is faithful with the saints.
HOS|12|1|Ephraim feedeth on wind, and followeth after the east wind: he daily increaseth lies and desolation; and they do make a covenant with the Assyrians, and oil is carried into Egypt.
HOS|12|2|The LORD hath also a controversy with Judah, and will punish Jacob according to his ways; according to his doings will he recompense him.
HOS|12|3|He took his brother by the heel in the womb, and by his strength he had power with God:
HOS|12|4|Yea, he had power over the angel, and prevailed: he wept, and made supplication unto him: he found him in Bethel, and there he spake with us;
HOS|12|5|Even the LORD God of hosts; the LORD is his memorial.
HOS|12|6|Therefore turn thou to thy God: keep mercy and judgment and wait on thy God continually.
HOS|12|7|He is a merchant, the balances of deceit are in his hand: he loveth to oppress.
HOS|12|8|And Ephraim said, Yet I am become rich, I have found me out substance: in all my labours they shall find none iniquity in me that were sin.
HOS|12|9|And I that am the LORD thy God from the land of Egypt will yet make thee to dwell in tabernacles, as in the days of the solemn feast.
HOS|12|10|I have also spoken by the prophets, and I have multiplied visions, and used similitudes, by the ministry of the prophets.
HOS|12|11|Is there iniquity in Gilead? surely they are vanity: they sacrifice bullocks in Gilgal; yea, their altars are as heaps in the furrows of the fields.
HOS|12|12|And Jacob fled into the country of Syria, and Israel served for a wife, and for a wife he kept sheep.
HOS|12|13|And by a prophet the LORD brought Israel out of Egypt, and by a prophet was he preserved.
HOS|12|14|Ephraim provoked him to anger most bitterly: therefore shall he leave his blood upon him, and his reproach shall his LORD return unto him.
HOS|13|1|When Ephraim spake trembling, he exalted himself in Israel; but when he offended in Baal, he died.
HOS|13|2|And now they sin more and more, and have made them molten images of their silver, and idols according to their own understanding, all of it the work of the craftsmen: they say of them, Let the men that sacrifice kiss the calves.
HOS|13|3|Therefore they shall be as the morning cloud and as the early dew that passeth away, as the chaff that is driven with the whirlwind out of the floor, and as the smoke out of the chimney.
HOS|13|4|Yet I am the LORD thy God from the land of Egypt, and thou shalt know no god but me: for there is no saviour beside me.
HOS|13|5|I did know thee in the wilderness, in the land of great drought.
HOS|13|6|According to their pasture, so were they filled; they were filled, and their heart was exalted; therefore have they forgotten me.
HOS|13|7|Therefore I will be unto them as a lion: as a leopard by the way will I observe them:
HOS|13|8|I will meet them as a bear that is bereaved of her whelps, and will rend the caul of their heart, and there will I devour them like a lion: the wild beast shall tear them.
HOS|13|9|O Israel, thou hast destroyed thyself; but in me is thine help.
HOS|13|10|I will be thy king: where is any other that may save thee in all thy cities? and thy judges of whom thou saidst, Give me a king and princes?
HOS|13|11|I gave thee a king in mine anger, and took him away in my wrath.
HOS|13|12|The iniquity of Ephraim is bound up; his sin is hid.
HOS|13|13|The sorrows of a travailing woman shall come upon him: he is an unwise son; for he should not stay long in the place of the breaking forth of children.
HOS|13|14|I will ransom them from the power of the grave; I will redeem them from death: O death, I will be thy plagues; O grave, I will be thy destruction: repentance shall be hid from mine eyes.
HOS|13|15|Though he be fruitful among his brethren, an east wind shall come, the wind of the LORD shall come up from the wilderness, and his spring shall become dry, and his fountain shall be dried up: he shall spoil the treasure of all pleasant vessels.
HOS|13|16|Samaria shall become desolate; for she hath rebelled against her God: they shall fall by the sword: their infants shall be dashed in pieces, and their women with child shall be ripped up.
HOS|14|1|O israel, return unto the LORD thy God; for thou hast fallen by thine iniquity.
HOS|14|2|Take with you words, and turn to the LORD: say unto him, Take away all iniquity, and receive us graciously: so will we render the calves of our lips.
HOS|14|3|Asshur shall not save us; we will not ride upon horses: neither will we say any more to the work of our hands, Ye are our gods: for in thee the fatherless findeth mercy.
HOS|14|4|I will heal their backsliding, I will love them freely: for mine anger is turned away from him.
HOS|14|5|I will be as the dew unto Israel: he shall grow as the lily, and cast forth his roots as Lebanon.
HOS|14|6|His branches shall spread, and his beauty shall be as the olive tree, and his smell as Lebanon.
HOS|14|7|They that dwell under his shadow shall return; they shall revive as the corn, and grow as the vine: the scent thereof shall be as the wine of Lebanon.
HOS|14|8|Ephraim shall say, What have I to do any more with idols? I have heard him, and observed him: I am like a green fir tree. From me is thy fruit found.
HOS|14|9|Who is wise, and he shall understand these things? prudent, and he shall know them? for the ways of the LORD are right, and the just shall walk in them: but the transgressors shall fall therein.
