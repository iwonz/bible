COL|1|1|Paulus apostolus Christi Iesu per voluntatem Dei et Timotheus frater
COL|1|2|his qui sunt Colossis sanctis et fidelibus fratribus in Christo Iesu gratia vobis et pax a Deo Patre nostro
COL|1|3|gratias agimus Deo et Patri Domini nostri Iesu Christi semper pro vobis orantes
COL|1|4|audientes fidem vestram in Christo Iesu et dilectionem quam habetis in sanctos omnes
COL|1|5|propter spem quae reposita est vobis in caelis quam audistis in verbo veritatis evangelii
COL|1|6|quod pervenit ad vos sicut et in universo mundo est et fructificat et crescit sicut in vobis ex ea die qua audistis et cognovistis gratiam Dei in veritate
COL|1|7|sicut didicistis ab Epaphra carissimo conservo nostro qui est fidelis pro vobis minister Christi Iesu
COL|1|8|qui etiam manifestavit nobis dilectionem vestram in Spiritu
COL|1|9|ideo et nos ex qua die audivimus non cessamus pro vobis orantes et postulantes ut impleamini agnitione voluntatis eius in omni sapientia et intellectu spiritali
COL|1|10|ut ambuletis digne Deo per omnia placentes in omni opere bono fructificantes et crescentes in scientia Dei
COL|1|11|in omni virtute confortati secundum potentiam claritatis eius in omni patientia et longanimitate cum gaudio
COL|1|12|gratias agentes Patri qui dignos nos fecit in partem sortis sanctorum in lumine
COL|1|13|qui eripuit nos de potestate tenebrarum et transtulit in regnum Filii dilectionis suae
COL|1|14|in quo habemus redemptionem remissionem peccatorum
COL|1|15|qui est imago Dei invisibilis primogenitus omnis creaturae
COL|1|16|quia in ipso condita sunt universa in caelis et in terra visibilia et invisibilia sive throni sive dominationes sive principatus sive potestates omnia per ipsum et in ipso creata sunt
COL|1|17|et ipse est ante omnes et omnia in ipso constant
COL|1|18|et ipse est caput corporis ecclesiae qui est principium primogenitus ex mortuis ut sit in omnibus ipse primatum tenens
COL|1|19|quia in ipso conplacuit omnem plenitudinem habitare
COL|1|20|et per eum reconciliare omnia in ipsum pacificans per sanguinem crucis eius sive quae in terris sive quae in caelis sunt
COL|1|21|et vos cum essetis aliquando alienati et inimici sensu in operibus malis
COL|1|22|nunc autem reconciliavit in corpore carnis eius per mortem exhibere vos sanctos et inmaculatos et inreprehensibiles coram ipso
COL|1|23|si tamen permanetis in fide fundati et stabiles et inmobiles ab spe evangelii quod audistis quod praedicatum est in universa creatura quae sub caelo est cuius factus sum ego Paulus minister
COL|1|24|qui nunc gaudeo in passionibus pro vobis et adimpleo ea quae desunt passionum Christi in carne mea pro corpore eius quod est ecclesia
COL|1|25|cuius factus sum ego minister secundum dispensationem Dei quae data est mihi in vos ut impleam verbum Dei
COL|1|26|mysterium quod absconditum fuit a saeculis et generationibus nunc autem manifestatum est sanctis eius
COL|1|27|quibus voluit Deus notas facere divitias gloriae sacramenti huius in gentibus quod est Christus in vobis spes gloriae
COL|1|28|quem nos adnuntiamus corripientes omnem hominem et docentes omnem hominem in omni sapientia ut exhibeamus omnem hominem perfectum in Christo Iesu
COL|1|29|in quo et laboro certando secundum operationem eius quam operatur in me in virtute
COL|2|1|volo enim vos scire qualem sollicitudinem habeam pro vobis et pro his qui sunt Laodiciae et quicumque non viderunt faciem meam in carne
COL|2|2|ut consolentur corda ipsorum instructi in caritate et in omnes divitias plenitudinis intellectus in agnitionem mysterii Dei Patris Christi Iesu
COL|2|3|in quo sunt omnes thesauri sapientiae et scientiae absconditi
COL|2|4|hoc autem dico ut nemo vos decipiat in subtilitate sermonum
COL|2|5|nam et si corpore absens sum sed spiritu vobiscum sum gaudens et videns ordinem vestrum et firmamentum eius quae in Christo est fidei vestrae
COL|2|6|sicut ergo accepistis Christum Iesum Dominum in ipso ambulate
COL|2|7|radicati et superaedificati in ipso et confirmati fide sicut et didicistis abundantes in gratiarum actione
COL|2|8|videte ne quis vos decipiat per philosophiam et inanem fallaciam secundum traditionem hominum secundum elementa mundi et non secundum Christum
COL|2|9|quia in ipso inhabitat omnis plenitudo divinitatis corporaliter
COL|2|10|et estis in illo repleti qui est caput omnis principatus et potestatis
COL|2|11|in quo et circumcisi estis circumcisione non manufacta in expoliatione corporis carnis in circumcisione Christi
COL|2|12|consepulti ei in baptismo in quo et resurrexistis per fidem operationis Dei qui suscitavit illum a mortuis
COL|2|13|et vos cum mortui essetis in delictis et praeputio carnis vestrae convivificavit cum illo donans vobis omnia delicta
COL|2|14|delens quod adversum nos erat chirografum decretis quod erat contrarium nobis et ipsum tulit de medio adfigens illud cruci
COL|2|15|expolians principatus et potestates traduxit palam triumphans illos in semet ipso
COL|2|16|nemo ergo vos iudicet in cibo aut in potu aut in parte diei festi aut neomeniae aut sabbatorum
COL|2|17|quae sunt umbra futurorum corpus autem Christi
COL|2|18|nemo vos seducat volens in humilitate et religione angelorum quae non vidit ambulans frustra inflatus sensu carnis suae
COL|2|19|et non tenens caput ex quo totum corpus per nexus et coniunctiones subministratum et constructum crescit in augmentum Dei
COL|2|20|si mortui estis cum Christo ab elementis mundi quid adhuc tamquam viventes in mundo decernitis
COL|2|21|ne tetigeris neque gustaveris neque contrectaveris
COL|2|22|quae sunt omnia in interitu ipso usu secundum praecepta et doctrinas hominum
COL|2|23|quae sunt rationem quidem habentia sapientiae in superstitione et humilitate et ad non parcendum corpori non in honore aliquo ad saturitatem carnis
COL|3|1|igitur si conresurrexistis Christo quae sursum sunt quaerite ubi Christus est in dextera Dei sedens
COL|3|2|quae sursum sunt sapite non quae supra terram
COL|3|3|mortui enim estis et vita vestra abscondita est cum Christo in Deo
COL|3|4|cum Christus apparuerit vita vestra tunc et vos apparebitis cum ipso in gloria
COL|3|5|mortificate ergo membra vestra quae sunt super terram fornicationem inmunditiam libidinem concupiscentiam malam et avaritiam quae est simulacrorum servitus
COL|3|6|propter quae venit ira Dei super filios incredulitatis
COL|3|7|in quibus et vos ambulastis aliquando cum viveretis in illis
COL|3|8|nunc autem deponite et vos omnia iram indignationem malitiam blasphemiam turpem sermonem de ore vestro
COL|3|9|nolite mentiri invicem expoliantes vos veterem hominem cum actibus eius
COL|3|10|et induentes novum eum qui renovatur in agnitionem secundum imaginem eius qui creavit eum
COL|3|11|ubi non est gentilis et Iudaeus circumcisio et praeputium barbarus et Scytha servus et liber sed omnia et in omnibus Christus
COL|3|12|induite vos ergo sicut electi Dei sancti et dilecti viscera misericordiae benignitatem humilitatem modestiam patientiam
COL|3|13|subportantes invicem et donantes vobis ipsis si quis adversus aliquem habet querellam sicut et Dominus donavit vobis ita et vos
COL|3|14|super omnia autem haec caritatem quod est vinculum perfectionis
COL|3|15|et pax Christi exultet in cordibus vestris in qua et vocati estis in uno corpore et grati estote
COL|3|16|verbum Christi habitet in vobis abundanter in omni sapientia docentes et commonentes vosmet ipsos psalmis hymnis canticis spiritalibus in gratia cantantes in cordibus vestris Deo
COL|3|17|omne quodcumque facitis in verbo aut in opere omnia in nomine Domini Iesu gratias agentes Deo et Patri per ipsum
COL|3|18|mulieres subditae estote viris sicut oportet in Domino
COL|3|19|viri diligite uxores et nolite amari esse ad illas
COL|3|20|filii oboedite parentibus per omnia hoc enim placitum est in Domino
COL|3|21|patres nolite ad indignationem provocare filios vestros ut non pusillo animo fiant
COL|3|22|servi oboedite per omnia dominis carnalibus non ad oculum servientes quasi hominibus placentes sed in simplicitate cordis timentes Dominum
COL|3|23|quodcumque facitis ex animo operamini sicut Domino et non hominibus
COL|3|24|scientes quod a Domino accipietis retributionem hereditatis Domino Christo servite
COL|3|25|qui enim iniuriam facit recipiet id quod inique gessit et non est personarum acceptio
COL|4|1|domini quod iustum est et aequum servis praestate scientes quoniam et vos Dominum habetis in caelo
COL|4|2|orationi instate vigilantes in ea in gratiarum actione
COL|4|3|orantes simul et pro nobis ut Deus aperiat nobis ostium sermonis ad loquendum mysterium Christi propter quod etiam vinctus sum
COL|4|4|ut manifestem illud ita ut oportet me loqui
COL|4|5|in sapientia ambulate ad eos qui foris sunt tempus redimentes
COL|4|6|sermo vester semper in gratia sale sit conditus ut sciatis quomodo oporteat vos unicuique respondere
COL|4|7|quae circa me sunt omnia vobis nota faciet Tychicus carissimus frater et fidelis minister et conservus in Domino
COL|4|8|quem misi ad vos ad hoc ipsum ut cognoscat quae circa vos sunt et consoletur corda vestra
COL|4|9|cum Onesimo carissimo et fideli fratre qui est ex vobis omnia quae hic aguntur nota facient vobis
COL|4|10|salutat vos Aristarchus concaptivus meus et Marcus consobrinus Barnabae de quo accepistis mandata si venerit ad vos excipite illum
COL|4|11|et Iesus qui dicitur Iustus qui sunt ex circumcisione hii soli sunt adiutores in regno Dei qui mihi fuerunt solacio
COL|4|12|salutat vos Epaphras qui ex vobis est servus Christi Iesu semper sollicitus pro vobis in orationibus ut stetis perfecti et pleni in omni voluntate Dei
COL|4|13|testimonium enim illi perhibeo quod habet multum laborem pro vobis et pro his qui sunt Laodiciae et qui Hierapoli
COL|4|14|salutat vos Lucas medicus carissimus et Demas
COL|4|15|salutate fratres qui sunt Laodiciae et Nympham et quae in domo eius est ecclesiam
COL|4|16|et cum lecta fuerit apud vos epistula facite ut et in Laodicensium ecclesia legatur et eam quae Laodicensium est vos legatis
COL|4|17|et dicite Archippo vide ministerium quod accepisti in Domino ut illud impleas
COL|4|18|salutatio mea manu Pauli memores estote vinculorum meorum gratia vobiscum amen
