2THESS|1|1|Paulus et Silvanus et Timotheus ecclesiae Thessalonicensium in Deo Patre nostro et Domino Iesu Christo
2THESS|1|2|gratia vobis et pax a Deo Patre nostro et Domino Iesu Christo
2THESS|1|3|gratias agere debemus Deo semper pro vobis fratres ita ut dignum est quoniam supercrescit fides vestra et abundat caritas uniuscuiusque omnium vestrum in invicem
2THESS|1|4|ita ut et nos ipsi in vobis gloriemur in ecclesiis Dei pro patientia vestra et fide in omnibus persecutionibus vestris et tribulationibus quas sustinetis
2THESS|1|5|in exemplum iusti iudicii Dei ut digni habeamini regno Dei pro quo et patimini
2THESS|1|6|si tamen iustum est apud Deum retribuere tribulationem his qui vos tribulant
2THESS|1|7|et vobis qui tribulamini requiem nobiscum in revelatione Domini Iesu de caelo cum angelis virtutis eius
2THESS|1|8|in flamma ignis dantis vindictam his qui non noverunt Deum et qui non oboediunt evangelio Domini nostri Iesu
2THESS|1|9|qui poenas dabunt in interitu aeternas a facie Domini et a gloria virtutis eius
2THESS|1|10|cum venerit glorificari in sanctis suis et admirabilis fieri in omnibus qui crediderunt quia creditum est testimonium nostrum super vos in die illo
2THESS|1|11|in quo etiam oramus semper pro vobis ut dignetur vos vocatione sua Deus et impleat omnem voluntatem bonitatis et opus fidei in virtute
2THESS|1|12|ut clarificetur nomen Domini nostri Iesu Christi in vobis et vos in illo secundum gratiam Dei nostri et Domini Iesu Christi
2THESS|2|1|rogamus autem vos fratres per adventum Domini nostri Iesu Christi et nostrae congregationis in ipsum
2THESS|2|2|ut non cito moveamini a sensu neque terreamini neque per spiritum neque per sermonem neque per epistulam tamquam per nos quasi instet dies Domini
2THESS|2|3|ne quis vos seducat ullo modo quoniam nisi venerit discessio primum et revelatus fuerit homo peccati filius perditionis
2THESS|2|4|qui adversatur et extollitur supra omne quod dicitur Deus aut quod colitur ita ut in templo Dei sedeat ostendens se quia sit Deus
2THESS|2|5|non retinetis quod cum adhuc essem apud vos haec dicebam vobis
2THESS|2|6|et nunc quid detineat scitis ut reveletur in suo tempore
2THESS|2|7|nam mysterium iam operatur iniquitatis tantum ut qui tenet nunc donec de medio fiat
2THESS|2|8|et tunc revelabitur ille iniquus quem Dominus Iesus interficiet spiritu oris sui et destruet inlustratione adventus sui
2THESS|2|9|eum cuius est adventus secundum operationem Satanae in omni virtute et signis et prodigiis mendacibus
2THESS|2|10|et in omni seductione iniquitatis his qui pereunt eo quod caritatem veritatis non receperunt ut salvi fierent
2THESS|2|11|ideo mittit illis Deus operationem erroris ut credant mendacio
2THESS|2|12|ut iudicentur omnes qui non crediderunt veritati sed consenserunt iniquitati
2THESS|2|13|nos autem debemus gratias agere Deo semper pro vobis fratres dilecti a Deo quod elegerit nos Deus primitias in salutem in sanctificatione Spiritus et fide veritatis
2THESS|2|14|ad quod et vocavit vos per evangelium nostrum in adquisitionem gloriae Domini nostri Iesu Christi
2THESS|2|15|itaque fratres state et tenete traditiones quas didicistis sive per sermonem sive per epistulam nostram
2THESS|2|16|ipse autem Dominus noster Iesus Christus et Deus et Pater noster qui dilexit nos et dedit consolationem aeternam et spem bonam in gratia
2THESS|2|17|exhortetur corda vestra et confirmet in omni opere et sermone bono
2THESS|3|1|de cetero fratres orate pro nobis ut sermo Domini currat et clarificetur sicut et apud vos
2THESS|3|2|et ut liberemur ab inportunis et malis hominibus non enim omnium est fides
2THESS|3|3|fidelis autem Dominus est qui confirmabit vos et custodiet a malo
2THESS|3|4|confidimus autem de vobis in Domino quoniam quae praecipimus et facitis et facietis
2THESS|3|5|Dominus autem dirigat corda vestra in caritate Dei et patientia Christi
2THESS|3|6|denuntiamus autem vobis fratres in nomine Domini nostri Iesu Christi ut subtrahatis vos ab omni fratre ambulante inordinate et non secundum traditionem quam acceperunt a nobis
2THESS|3|7|ipsi enim scitis quemadmodum oporteat imitari nos quoniam non inquieti fuimus inter vos
2THESS|3|8|neque gratis panem manducavimus ab aliquo sed in labore et fatigatione nocte et die operantes ne quem vestrum gravaremus
2THESS|3|9|non quasi non habuerimus potestatem sed ut nosmet ipsos formam daremus vobis ad imitandum nos
2THESS|3|10|nam et cum essemus apud vos hoc denuntiabamus vobis quoniam si quis non vult operari nec manducet
2THESS|3|11|audimus enim inter vos quosdam ambulare inquiete nihil operantes sed curiose agentes
2THESS|3|12|his autem qui eiusmodi sunt denuntiamus et obsecramus in Domino Iesu Christo ut cum silentio operantes suum panem manducent
2THESS|3|13|vos autem fratres nolite deficere benefacientes
2THESS|3|14|quod si quis non oboedit verbo nostro per epistulam hunc notate et non commisceamini cum illo ut confundatur
2THESS|3|15|et nolite quasi inimicum existimare sed corripite ut fratrem
2THESS|3|16|ipse autem Dominus pacis det vobis pacem sempiternam in omni loco Dominus cum omnibus vobis
2THESS|3|17|salutatio mea manu Pauli quod est signum in omni epistula ita scribo
2THESS|3|18|gratia Domini nostri Iesu Christi cum omnibus vobis amen
