MARK|1|1|The beginning of the gospel of Jesus Christ, the Son of God.
MARK|1|2|As it is written in Isaiah the prophet, "Behold, I send my messenger before your face, who will prepare your way,
MARK|1|3|the voice of one crying in the wilderness: Prepare the way of the Lord, make his paths straight."
MARK|1|4|John appeared, baptizing in the wilderness and proclaiming a baptism of repentance for the forgiveness of sins.
MARK|1|5|And all the country of Judea and all Jerusalem were going out to him and were being baptized by him in the river Jordan, confessing their sins.
MARK|1|6|Now John was clothed with camel's hair and wore a leather belt around his waist and ate locusts and wild honey.
MARK|1|7|And he preached, saying, "After me comes he who is mightier than I, the strap of whose sandals I am not worthy to stoop down and untie.
MARK|1|8|I have baptized you with water, but he will baptize you with the Holy Spirit."
MARK|1|9|In those days Jesus came from Nazareth of Galilee and was baptized by John in the Jordan.
MARK|1|10|And when he came up out of the water, immediately he saw the heavens opening and the Spirit descending on him like a dove.
MARK|1|11|And a voice came from heaven, "You are my beloved Son; with you I am well pleased."
MARK|1|12|The Spirit immediately drove him out into the wilderness.
MARK|1|13|And he was in the wilderness forty days, being tempted by Satan. And he was with the wild animals, and the angels were ministering to him.
MARK|1|14|Now after John was arrested, Jesus came into Galilee, proclaiming the gospel of God,
MARK|1|15|and saying, "The time is fulfilled, and the kingdom of God is at hand; repent and believe in the gospel."
MARK|1|16|Passing alongside the Sea of Galilee, he saw Simon and Andrew the brother of Simon casting a net into the sea, for they were fishermen.
MARK|1|17|And Jesus said to them, "Follow me, and I will make you become fishers of men."
MARK|1|18|And immediately they left their nets and followed him.
MARK|1|19|And going on a little farther, he saw James the son of Zebedee and John his brother, who were in their boat mending the nets.
MARK|1|20|And immediately he called them, and they left their father Zebedee in the boat with the hired servants and followed him.
MARK|1|21|And they went into Capernaum, and immediately on the Sabbath he entered the synagogue and was teaching.
MARK|1|22|And they were astonished at his teaching, for he taught them as one who had authority, and not as the scribes.
MARK|1|23|And immediately there was in their synagogue a man with an unclean spirit. And he cried out,
MARK|1|24|"What have you to do with us, Jesus of Nazareth? Have you come to destroy us? I know who you are- the Holy One of God."
MARK|1|25|But Jesus rebuked him, saying, "Be silent, and come out of him!"
MARK|1|26|And the unclean spirit, convulsing him and crying out with a loud voice, came out of him.
MARK|1|27|And they were all amazed, so that they questioned among themselves, saying, "What is this? A new teaching with authority! He commands even the unclean spirits, and they obey him."
MARK|1|28|And at once his fame spread everywhere throughout all the surrounding region of Galilee.
MARK|1|29|And immediately he left the synagogue and entered the house of Simon and Andrew, with James and John.
MARK|1|30|Now Simon's mother-in-law lay ill with a fever, and immediately they told him about her.
MARK|1|31|And he came and took her by the hand and lifted her up, and the fever left her, and she began to serve them.
MARK|1|32|That evening at sundown they brought to him all who were sick or oppressed by demons.
MARK|1|33|And the whole city was gathered together at the door.
MARK|1|34|And he healed many who were sick with various diseases, and cast out many demons. And he would not permit the demons to speak, because they knew him.
MARK|1|35|And rising very early in the morning, while it was still dark, he departed and went out to a desolate place, and there he prayed.
MARK|1|36|And Simon and those who were with him searched for him,
MARK|1|37|and they found him and said to him, "Everyone is looking for you."
MARK|1|38|And he said to them, "Let us go on to the next towns, that I may preach there also, for that is why I came out."
MARK|1|39|And he went throughout all Galilee, preaching in their synagogues and casting out demons.
MARK|1|40|And a leper came to him, imploring him, and kneeling said to him, "If you will, you can make me clean."
MARK|1|41|Moved with pity, he stretched out his hand and touched him and said to him, "I will; be clean."
MARK|1|42|And immediately the leprosy left him, and he was made clean.
MARK|1|43|And Jesus sternly charged him and sent him away at once,
MARK|1|44|and said to him, "See that you say nothing to anyone, but go, show yourself to the priest and offer for your cleansing what Moses commanded, for a proof to them."
MARK|1|45|But he went out and began to talk freely about it, and to spread the news, so that Jesus could no longer openly enter a town, but was out in desolate places, and people were coming to him from every quarter.
MARK|2|1|And when he returned to Capernaum after some days, it was reported that he was at home.
MARK|2|2|And many were gathered together, so that there was no more room, not even at the door. And he was preaching the word to them.
MARK|2|3|And they came, bringing to him a paralytic carried by four men.
MARK|2|4|And when they could not get near him because of the crowd, they removed the roof above him, and when they had made an opening, they let down the bed on which the paralytic lay.
MARK|2|5|And when Jesus saw their faith, he said to the paralytic, "My son, your sins are forgiven."
MARK|2|6|Now some of the scribes were sitting there, questioning in their hearts,
MARK|2|7|"Why does this man speak like that? He is blaspheming! Who can forgive sins but God alone?"
MARK|2|8|And immediately Jesus, perceiving in his spirit that they thus questioned within themselves, said to them, "Why do you question these things in your hearts?
MARK|2|9|Which is easier, to say to the paralytic, 'Your sins are forgiven,' or to say, 'Rise, take up your bed and walk'?
MARK|2|10|But that you may know that the Son of Man has authority on earth to forgive sins"- he said to the paralytic-
MARK|2|11|"I say to you, rise, pick up your bed, and go home."
MARK|2|12|And he rose and immediately picked up his bed and went out before them all, so that they were all amazed and glorified God, saying, "We never saw anything like this!"
MARK|2|13|He went out again beside the sea, and all the crowd was coming to him, and he was teaching them.
MARK|2|14|And as he passed by, he saw Levi the son of Alphaeus sitting at the tax booth, and he said to him, "Follow me." And he rose and followed him.
MARK|2|15|And as he reclined at table in his house, many tax collectors and sinners were reclining with Jesus and his disciples, for there were many who followed him.
MARK|2|16|And the scribes of the Pharisees, when they saw that he was eating with sinners and tax collectors, said to his disciples, "Why does he eat with tax collectors and sinners?"
MARK|2|17|And when Jesus heard it, he said to them, "Those who are well have no need of a physician, but those who are sick. I came not to call the righteous, but sinners."
MARK|2|18|Now John's disciples and the Pharisees were fasting. And people came and said to him, "Why do John's disciples and the disciples of the Pharisees fast, but your disciples do not fast?"
MARK|2|19|And Jesus said to them, "Can the wedding guests fast while the bridegroom is with them? As long as they have the bridegroom with them, they cannot fast.
MARK|2|20|The days will come when the bridegroom is taken away from them, and then they will fast in that day.
MARK|2|21|No one sews a piece of unshrunk cloth on an old garment. If he does, the patch tears away from it, the new from the old, and a worse tear is made.
MARK|2|22|And no one puts new wine into old wineskins. If he does, the wine will burst the skins- and the wine is destroyed, and so are the skins. But new wine is for fresh wineskins."
MARK|2|23|One Sabbath he was going through the grainfields, and as they made their way, his disciples began to pluck heads of grain.
MARK|2|24|And the Pharisees were saying to him, "Look, why are they doing what is not lawful on the Sabbath?"
MARK|2|25|And he said to them, "Have you never read what David did, when he was in need and was hungry, he and those who were with him:
MARK|2|26|how he entered the house of God, in the time of Abiathar the high priest, and ate the bread of the Presence, which it is not lawful for any but the priests to eat, and also gave it to those who were with him?"
MARK|2|27|And he said to them, "The Sabbath was made for man, not man for the Sabbath.
MARK|2|28|So the Son of Man is lord even of the Sabbath."
MARK|3|1|Again he entered the synagogue, and a man was there with a withered hand.
MARK|3|2|And they watched Jesus, to see whether he would heal him on the Sabbath, so that they might accuse him.
MARK|3|3|And he said to the man with the withered hand, "Come here."
MARK|3|4|And he said to them, "Is it lawful on the Sabbath to do good or to do harm, to save life or to kill?" But they were silent.
MARK|3|5|And he looked around at them with anger, grieved at their hardness of heart, and said to the man, "Stretch out your hand." He stretched it out, and his hand was restored.
MARK|3|6|The Pharisees went out and immediately held counsel with the Herodians against him, how to destroy him.
MARK|3|7|Jesus withdrew with his disciples to the sea, and a great crowd followed, from Galilee and Judea
MARK|3|8|and Jerusalem and Idumea and from beyond the Jordan and from around Tyre and Sidon. When the great crowd heard all that he was doing, they came to him.
MARK|3|9|And he told his disciples to have a boat ready for him because of the crowd, lest they crush him,
MARK|3|10|for he had healed many, so that all who had diseases pressed around him to touch him.
MARK|3|11|And whenever the unclean spirits saw him, they fell down before him and cried out, "You are the Son of God."
MARK|3|12|And he strictly ordered them not to make him known.
MARK|3|13|And he went up on the mountain and called to him those whom he desired, and they came to him.
MARK|3|14|And he appointed twelve (whom he also named apostles) so that they might be with him and he might send them out to preach
MARK|3|15|and have authority to cast out demons.
MARK|3|16|He appointed the twelve: Simon (to whom he gave the name Peter);
MARK|3|17|James the son of Zebedee and John the brother of James (to whom he gave the name Boanerges, that is, Sons of Thunder);
MARK|3|18|Andrew, and Philip, and Bartholomew, and Matthew, and Thomas, and James the son of Alphaeus, and Thaddaeus, and Simon the Cananaean,
MARK|3|19|and Judas Iscariot, who betrayed him.
MARK|3|20|Then he went home, and the crowd gathered again, so that they could not even eat.
MARK|3|21|And when his family heard it, they went out to seize him, for they were saying, "He is out of his mind."
MARK|3|22|And the scribes who came down from Jerusalem were saying, "He is possessed by Beelzebul," and "by the prince of demons he casts out the demons."
MARK|3|23|And he called them to him and said to them in parables, "How can Satan cast out Satan?
MARK|3|24|If a kingdom is divided against itself, that kingdom cannot stand.
MARK|3|25|And if a house is divided against itself, that house will not be able to stand.
MARK|3|26|And if Satan has risen up against himself and is divided, he cannot stand, but is coming to an end.
MARK|3|27|But no one can enter a strong man's house and plunder his goods, unless he first binds the strong man. Then indeed he may plunder his house.
MARK|3|28|"Truly, I say to you, all sins will be forgiven the children of man, and whatever blasphemies they utter,
MARK|3|29|but whoever blasphemes against the Holy Spirit never has forgiveness, but is guilty of an eternal sin"-
MARK|3|30|for they had said, "He has an unclean spirit."
MARK|3|31|And his mother and his brothers came, and standing outside they sent to him and called him.
MARK|3|32|And a crowd was sitting around him, and they said to him, "Your mother and your brothers are outside, seeking you."
MARK|3|33|And he answered them, "Who are my mother and my brothers?"
MARK|3|34|And looking about at those who sat around him, he said, "Here are my mother and my brothers!
MARK|3|35|Whoever does the will of God, he is my brother and sister and mother."
MARK|4|1|Again he began to teach beside the sea. And a very large crowd gathered about him, so that he got into a boat and sat in it on the sea, and the whole crowd was beside the sea on the land.
MARK|4|2|And he was teaching them many things in parables, and in his teaching he said to them:
MARK|4|3|"Listen! A sower went out to sow.
MARK|4|4|And as he sowed, some seed fell along the path, and the birds came and devoured it.
MARK|4|5|Other seed fell on rocky ground, where it did not have much soil, and immediately it sprang up, since it had no depth of soil.
MARK|4|6|And when the sun rose it was scorched, and since it had no root, it withered away.
MARK|4|7|Other seed fell among thorns, and the thorns grew up and choked it, and it yielded no grain.
MARK|4|8|And other seeds fell into good soil and produced grain, growing up and increasing and yielding thirtyfold and sixtyfold and a hundredfold."
MARK|4|9|And he said, "He who has ears to hear, let him hear."
MARK|4|10|And when he was alone, those around him with the twelve asked him about the parables.
MARK|4|11|And he said to them, "To you has been given the secret of the kingdom of God, but for those outside everything is in parables,
MARK|4|12|so that "they may indeed see but not perceive, and may indeed hear but not understand, lest they should turn and be forgiven."
MARK|4|13|And he said to them, "Do you not understand this parable? How then will you understand all the parables?
MARK|4|14|The sower sows the word.
MARK|4|15|And these are the ones along the path, where the word is sown: when they hear, Satan immediately comes and takes away the word that is sown in them.
MARK|4|16|And these are the ones sown on rocky ground: the ones who, when they hear the word, immediately receive it with joy.
MARK|4|17|And they have no root in themselves, but endure for a while. Then, when tribulation or persecution arises on account of the word, immediately they fall away.
MARK|4|18|And others are the ones sown among thorns. They are those who hear the word,
MARK|4|19|but the cares of the world and the deceitfulness of riches and the desires for other things enter in and choke the word, and it proves unfruitful.
MARK|4|20|But those that were sown on the good soil are the ones who hear the word and accept it and bear fruit, thirtyfold and sixtyfold and a hundredfold."
MARK|4|21|And he said to them, "Is a lamp brought in to be put under a basket, or under a bed, and not on a stand?
MARK|4|22|For nothing is hidden except to be made manifest; nor is anything secret except to come to light.
MARK|4|23|If anyone has ears to hear, let him hear."
MARK|4|24|And he said to them, "Pay attention to what you hear: with the measure you use, it will be measured to you, and still more will be added to you.
MARK|4|25|For to the one who has, more will be given, and from the one who has not, even what he has will be taken away."
MARK|4|26|And he said, "The kingdom of God is as if a man should scatter seed on the ground.
MARK|4|27|He sleeps and rises night and day, and the seed sprouts and grows; he knows not how.
MARK|4|28|The earth produces by itself, first the blade, then the ear, then the full grain in the ear.
MARK|4|29|But when the grain is ripe, at once he puts in the sickle, because the harvest has come."
MARK|4|30|And he said, "With what can we compare the kingdom of God, or what parable shall we use for it?
MARK|4|31|It is like a grain of mustard seed, which, when sown on the ground, is the smallest of all the seeds on earth,
MARK|4|32|yet when it is sown it grows up and becomes larger than all the garden plants and puts out large branches, so that the birds of the air can make nests in its shade."
MARK|4|33|With many such parables he spoke the word to them, as they were able to hear it.
MARK|4|34|He did not speak to them without a parable, but privately to his own disciples he explained everything.
MARK|4|35|On that day, when evening had come, he said to them, "Let us go across to the other side."
MARK|4|36|And leaving the crowd, they took him with them in the boat, just as he was. And other boats were with him.
MARK|4|37|And a great windstorm arose, and the waves were breaking into the boat, so that the boat was already filling.
MARK|4|38|But he was in the stern, asleep on the cushion. And they woke him and said to him, "Teacher, do you not care that we are perishing?"
MARK|4|39|And he awoke and rebuked the wind and said to the sea, "Peace! Be still!" And the wind ceased, and there was a great calm.
MARK|4|40|He said to them, "Why are you so afraid? Have you still no faith?"
MARK|4|41|And they were filled with great fear and said to one another, "Who then is this, that even wind and sea obey him?"
MARK|5|1|They came to the other side of the sea, to the country of the Gerasenes.
MARK|5|2|And when Jesus had stepped out of the boat, immediately there met him out of the tombs a man with an unclean spirit.
MARK|5|3|He lived among the tombs. And no one could bind him anymore, not even with a chain,
MARK|5|4|for he had often been bound with shackles and chains, but he wrenched the chains apart, and he broke the shackles in pieces. No one had the strength to subdue him.
MARK|5|5|Night and day among the tombs and on the mountains he was always crying out and bruising himself with stones.
MARK|5|6|And when he saw Jesus from afar, he ran and fell down before him.
MARK|5|7|And crying out with a loud voice, he said, "What have you to do with me, Jesus, Son of the Most High God? I adjure you by God, do not torment me."
MARK|5|8|For he was saying to him, "Come out of the man, you unclean spirit!"
MARK|5|9|And Jesus asked him, "What is your name?" He replied, "My name is Legion, for we are many."
MARK|5|10|And he begged him earnestly not to send them out of the country.
MARK|5|11|Now a great herd of pigs was feeding there on the hillside,
MARK|5|12|and they begged him, saying, "Send us to the pigs; let us enter them."
MARK|5|13|So he gave them permission. And the unclean spirits came out, and entered the pigs, and the herd, numbering about two thousand, rushed down the steep bank into the sea and were drowned in the sea.
MARK|5|14|The herdsmen fled and told it in the city and in the country. And people came to see what it was that had happened.
MARK|5|15|And they came to Jesus and saw the demon-possessed man, the one who had had the legion, sitting there, clothed and in his right mind, and they were afraid.
MARK|5|16|And those who had seen it described to them what had happened to the demon-possessed man and to the pigs.
MARK|5|17|And they began to beg Jesus to depart from their region.
MARK|5|18|As he was getting into the boat, the man who had been possessed with demons begged him that he might be with him.
MARK|5|19|And he did not permit him but said to him, "Go home to your friends and tell them how much the Lord has done for you, and how he has had mercy on you."
MARK|5|20|And he went away and began to proclaim in the Decapolis how much Jesus had done for him, and everyone marveled.
MARK|5|21|And when Jesus had crossed again in the boat to the other side, a great crowd gathered about him, and he was beside the sea.
MARK|5|22|Then came one of the rulers of the synagogue, Jairus by name, and seeing him, he fell at his feet
MARK|5|23|and implored him earnestly, saying, "My little daughter is at the point of death. Come and lay your hands on her, so that she may be made well and live."
MARK|5|24|And he went with him. And a great crowd followed him and thronged about him.
MARK|5|25|And there was a woman who had had a discharge of blood for twelve years,
MARK|5|26|and who had suffered much under many physicians, and had spent all that she had, and was no better but rather grew worse.
MARK|5|27|She had heard the reports about Jesus and came up behind him in the crowd and touched his garment.
MARK|5|28|For she said, "If I touch even his garments, I will be made well."
MARK|5|29|And immediately the flow of blood dried up, and she felt in her body that she was healed of her disease.
MARK|5|30|And Jesus, perceiving in himself that power had gone out from him, immediately turned about in the crowd and said, "Who touched my garments?"
MARK|5|31|And his disciples said to him, "You see the crowd pressing around you, and yet you say, 'Who touched me?'"
MARK|5|32|And he looked around to see who had done it.
MARK|5|33|But the woman, knowing what had happened to her, came in fear and trembling and fell down before him and told him the whole truth.
MARK|5|34|And he said to her, "Daughter, your faith has made you well; go in peace, and be healed of your disease."
MARK|5|35|While he was still speaking, there came from the ruler's house some who said, "Your daughter is dead. Why trouble the Teacher any further?"
MARK|5|36|But overhearing what they said, Jesus said to the ruler of the synagogue, "Do not fear, only believe."
MARK|5|37|And he allowed no one to follow him except Peter and James and John the brother of James.
MARK|5|38|They came to the house of the ruler of the synagogue, and Jesus saw a commotion, people weeping and wailing loudly.
MARK|5|39|And when he had entered, he said to them, "Why are you making a commotion and weeping? The child is not dead but sleeping."
MARK|5|40|And they laughed at him. But he put them all outside and took the child's father and mother and those who were with him and went in where the child was.
MARK|5|41|Taking her by the hand he said to her, "Talitha cumi," which means, "Little girl, I say to you, arise."
MARK|5|42|And immediately the girl got up and began walking (for she was twelve years of age), and they were immediately overcome with amazement.
MARK|5|43|And he strictly charged them that no one should know this, and told them to give her something to eat.
MARK|6|1|He went away from there and came to his hometown, and his disciples followed him.
MARK|6|2|And on the Sabbath he began to teach in the synagogue, and many who heard him were astonished, saying, "Where did this man get these things? What is the wisdom given to him? How are such mighty works done by his hands?
MARK|6|3|Is not this the carpenter, the son of Mary and brother of James and Joses and Judas and Simon? And are not his sisters here with us?" And they took offense at him.
MARK|6|4|And Jesus said to them, "A prophet is not without honor, except in his hometown and among his relatives and in his own household."
MARK|6|5|And he could do no mighty work there, except that he laid his hands on a few sick people and healed them.
MARK|6|6|And he marveled because of their unbelief. And he went about among the villages teaching.
MARK|6|7|And he called the twelve and began to send them out two by two, and gave them authority over the unclean spirits.
MARK|6|8|He charged them to take nothing for their journey except a staff- no bread, no bag, no money in their belts-
MARK|6|9|but to wear sandals and not put on two tunics.
MARK|6|10|And he said to them, "Whenever you enter a house, stay there until you depart from there.
MARK|6|11|And if any place will not receive you and they will not listen to you, when you leave, shake off the dust that is on your feet as a testimony against them."
MARK|6|12|So they went out and proclaimed that people should repent.
MARK|6|13|And they cast out many demons and anointed with oil many who were sick and healed them.
MARK|6|14|King Herod heard of it, for Jesus' name had become known. Some said, "John the Baptist has been raised from the dead. That is why these miraculous powers are at work in him."
MARK|6|15|But others said, "He is Elijah." And others said, "He is a prophet, like one of the prophets of old."
MARK|6|16|But when Herod heard of it, he said, "John, whom I beheaded, has been raised."
MARK|6|17|For it was Herod who had sent and seized John and bound him in prison for the sake of Herodias, his brother Philip's wife, because he had married her.
MARK|6|18|For John had been saying to Herod, "It is not lawful for you to have your brother's wife."
MARK|6|19|And Herodias had a grudge against him and wanted to put him to death. But she could not,
MARK|6|20|for Herod feared John, knowing that he was a righteous and holy man, and he kept him safe. When he heard him, he was greatly perplexed, and yet he heard him gladly.
MARK|6|21|But an opportunity came when Herod on his birthday gave a banquet for his nobles and military commanders and the leading men of Galilee.
MARK|6|22|For when Herodias's daughter came in and danced, she pleased Herod and his guests. And the king said to the girl, "Ask me for whatever you wish, and I will give it to you."
MARK|6|23|And he vowed to her, "Whatever you ask me, I will give you, up to half of my kingdom."
MARK|6|24|And she went out and said to her mother, "For what should I ask?" And she said, "The head of John the Baptist."
MARK|6|25|And she came in immediately with haste to the king and asked, saying, "I want you to give me at once the head of John the Baptist on a platter."
MARK|6|26|And the king was exceedingly sorry, but because of his oaths and his guests he did not want to break his word to her.
MARK|6|27|And immediately the king sent an executioner with orders to bring John's head. He went and beheaded him in the prison
MARK|6|28|and brought his head on a platter and gave it to the girl, and the girl gave it to her mother.
MARK|6|29|When his disciples heard of it, they came and took his body and laid it in a tomb.
MARK|6|30|The apostles returned to Jesus and told him all that they had done and taught.
MARK|6|31|And he said to them, "Come away by yourselves to a desolate place and rest a while." For many were coming and going, and they had no leisure even to eat.
MARK|6|32|And they went away in the boat to a desolate place by themselves.
MARK|6|33|Now many saw them going and recognized them, and they ran there on foot from all the towns and got there ahead of them.
MARK|6|34|When he went ashore he saw a great crowd, and he had compassion on them, because they were like sheep without a shepherd. And he began to teach them many things.
MARK|6|35|And when it grew late, his disciples came to him and said, "This is a desolate place, and the hour is now late.
MARK|6|36|Send them away to go into the surrounding countryside and villages and buy themselves something to eat."
MARK|6|37|But he answered them, "You give them something to eat." And they said to him, "Shall we go and buy two hundred denarii worth of bread and give it to them to eat?"
MARK|6|38|And he said to them, "How many loaves do you have? Go and see." And when they had found out, they said, "Five, and two fish."
MARK|6|39|Then he commanded them all to sit down in groups on the green grass.
MARK|6|40|So they sat down in groups, by hundreds and by fifties.
MARK|6|41|And taking the five loaves and the two fish he looked up to heaven and said a blessing and broke the loaves and gave them to the disciples to set before the people. And he divided the two fish among them all.
MARK|6|42|And they all ate and were satisfied.
MARK|6|43|And they took up twelve baskets full of broken pieces and of the fish.
MARK|6|44|And those who ate the loaves were five thousand men.
MARK|6|45|Immediately he made his disciples get into the boat and go before him to the other side, to Bethsaida, while he dismissed the crowd.
MARK|6|46|And after he had taken leave of them, he went up on the mountain to pray.
MARK|6|47|And when evening came, the boat was out on the sea, and he was alone on the land.
MARK|6|48|And he saw that they were making headway painfully, for the wind was against them. And about the fourth watch of the night he came to them, walking on the sea. He meant to pass by them,
MARK|6|49|but when they saw him walking on the sea they thought it was a ghost, and cried out,
MARK|6|50|for they all saw him and were terrified. But immediately he spoke to them and said, "Take heart; it is I. Do not be afraid."
MARK|6|51|And he got into the boat with them, and the wind ceased. And they were utterly astounded,
MARK|6|52|for they did not understand about the loaves, but their hearts were hardened.
MARK|6|53|When they had crossed over, they came to land at Gennesaret and moored to the shore.
MARK|6|54|And when they got out of the boat, the people immediately recognized him
MARK|6|55|and ran about the whole region and began to bring the sick people on their beds to wherever they heard he was.
MARK|6|56|And wherever he came, in villages, cities, or countryside, they laid the sick in the marketplaces and implored him that they might touch even the fringe of his garment. And as many as touched it were made well.
MARK|7|1|Now when the Pharisees gathered to him, with some of the scribes who had come from Jerusalem,
MARK|7|2|they saw that some of his disciples ate with hands that were defiled, that is, unwashed.
MARK|7|3|(For the Pharisees and all the Jews do not eat unless they wash their hands, holding to the tradition of the elders,
MARK|7|4|and when they come from the marketplace, they do not eat unless they wash. And there are many other traditions that they observe, such as the washing of cups and pots and copper vessels and dining couches.)
MARK|7|5|And the Pharisees and the scribes asked him, "Why do your disciples not walk according to the tradition of the elders, but eat with defiled hands?"
MARK|7|6|And he said to them, "Well did Isaiah prophesy of you hypocrites, as it is written, "' This people honors me with their lips, but their heart is far from me;
MARK|7|7|in vain do they worship me, teaching as doctrines the commandments of men.'
MARK|7|8|You leave the commandment of God and hold to the tradition of men."
MARK|7|9|And he said to them, "You have a fine way of rejecting the commandment of God in order to establish your tradition!
MARK|7|10|For Moses said, 'Honor your father and your mother'; and, 'Whoever reviles father or mother must surely die.'
MARK|7|11|But you say, 'If a man tells his father or his mother, Whatever you would have gained from me is Corban' (that is, given to God)-
MARK|7|12|then you no longer permit him to do anything for his father or mother,
MARK|7|13|thus making void the word of God by your tradition that you have handed down. And many such things you do."
MARK|7|14|And he called the people to him again and said to them, "Hear me, all of you, and understand:
MARK|7|15|There is nothing outside a person that by going into him can defile him, but the things that come out of a person are what defile him."
MARK|7|16|***
MARK|7|17|And when he had entered the house and left the people, his disciples asked him about the parable.
MARK|7|18|And he said to them, "Then are you also without understanding? Do you not see that whatever goes into a person from outside cannot defile him,
MARK|7|19|since it enters not his heart but his stomach, and is expelled?" (Thus he declared all foods clean.)
MARK|7|20|And he said, "What comes out of a person is what defiles him.
MARK|7|21|For from within, out of the heart of man, come evil thoughts, sexual immorality, theft, murder, adultery,
MARK|7|22|coveting, wickedness, deceit, sensuality, envy, slander, pride, foolishness.
MARK|7|23|All these evil things come from within, and they defile a person."
MARK|7|24|And from there he arose and went away to the region of Tyre and Sidon. And he entered a house and did not want anyone to know, yet he could not be hidden.
MARK|7|25|But immediately a woman whose little daughter was possessed by an unclean spirit heard of him and came and fell down at his feet.
MARK|7|26|Now the woman was a Gentile, a Syrophoenician by birth. And she begged him to cast the demon out of her daughter.
MARK|7|27|And he said to her, "Let the children be fed first, for it is not right to take the children's bread and throw it to the dogs."
MARK|7|28|But she answered him, "Yes, Lord; yet even the dogs under the table eat the children's crumbs."
MARK|7|29|And he said to her, "For this statement you may go your way; the demon has left your daughter."
MARK|7|30|And she went home and found the child lying in bed and the demon gone.
MARK|7|31|Then he returned from the region of Tyre and went through Sidon to the Sea of Galilee, in the region of the Decapolis.
MARK|7|32|And they brought to him a man who was deaf and had a speech impediment, and they begged him to lay his hand on him.
MARK|7|33|And taking him aside from the crowd privately, he put his fingers into his ears, and after spitting touched his tongue.
MARK|7|34|And looking up to heaven, he sighed and said to him, "Ephphatha," that is, "Be opened."
MARK|7|35|And his ears were opened, his tongue was released, and he spoke plainly.
MARK|7|36|And Jesus charged them to tell no one. But the more he charged them, the more zealously they proclaimed it.
MARK|7|37|And they were astonished beyond measure, saying, "He has done all things well. He even makes the deaf hear and the mute speak."
MARK|8|1|In those days, when again a great crowd had gathered, and they had nothing to eat, he called his disciples to him and said to them,
MARK|8|2|"I have compassion on the crowd, because they have been with me now three days and have nothing to eat.
MARK|8|3|And if I send them away hungry to their homes, they will faint on the way. And some of them have come from far away."
MARK|8|4|And his disciples answered him, "How can one feed these people with bread here in this desolate place?"
MARK|8|5|And he asked them, "How many loaves do you have?" They said, "Seven."
MARK|8|6|And he directed the crowd to sit down on the ground. And he took the seven loaves, and having given thanks, he broke them and gave them to his disciples to set before the people; and they set them before the crowd.
MARK|8|7|And they had a few small fish. And having blessed them, he said that these also should be set before them.
MARK|8|8|And they ate and were satisfied. And they took up the broken pieces left over, seven baskets full.
MARK|8|9|And there were about four thousand people. And he sent them away.
MARK|8|10|And immediately he got into the boat with his disciples and went to the district of Dalmanutha.
MARK|8|11|The Pharisees came and began to argue with him, seeking from him a sign from heaven to test him.
MARK|8|12|And he sighed deeply in his spirit and said, "Why does this generation seek a sign? Truly, I say to you, no sign will be given to this generation."
MARK|8|13|And he left them, got into the boat again, and went to the other side.
MARK|8|14|Now they had forgotten to bring bread, and they had only one loaf with them in the boat.
MARK|8|15|And he cautioned them, saying, "Watch out; beware of the leaven of the Pharisees and the leaven of Herod."
MARK|8|16|And they began discussing with one another the fact that they had no bread.
MARK|8|17|And Jesus, aware of this, said to them, "Why are you discussing the fact that you have no bread? Do you not yet perceive or understand? Are your hearts hardened?
MARK|8|18|Having eyes do you not see, and having ears do you not hear? And do you not remember?
MARK|8|19|When I broke the five loaves for the five thousand, how many baskets full of broken pieces did you take up?" They said to him, "Twelve."
MARK|8|20|"And the seven for the four thousand, how many baskets full of broken pieces did you take up?" And they said to him, "Seven."
MARK|8|21|And he said to them, "Do you not yet understand?"
MARK|8|22|And they came to Bethsaida. And some people brought to him a blind man and begged him to touch him.
MARK|8|23|And he took the blind man by the hand and led him out of the village, and when he had spit on his eyes and laid his hands on him, he asked him, "Do you see anything?"
MARK|8|24|And he looked up and said, "I see men, but they look like trees, walking."
MARK|8|25|Then Jesus laid his hands on his eyes again; and he opened his eyes, his sight was restored, and he saw everything clearly.
MARK|8|26|And he sent him to his home, saying, "Do not even enter the village."
MARK|8|27|And Jesus went on with his disciples to the villages of Caesarea Philippi. And on the way he asked his disciples, "Who do people say that I am?"
MARK|8|28|And they told him, "John the Baptist; and others say, Elijah; and others, one of the prophets."
MARK|8|29|And he asked them, "But who do you say that I am?" Peter answered him, "You are the Christ."
MARK|8|30|And he strictly charged them to tell no one about him.
MARK|8|31|And he began to teach them that the Son of Man must suffer many things and be rejected by the elders and the chief priests and the scribes and be killed, and after three days rise again.
MARK|8|32|And he said this plainly. And Peter took him aside and began to rebuke him.
MARK|8|33|But turning and seeing his disciples, he rebuked Peter and said, "Get behind me, Satan! For you are not setting your mind on the things of God, but on the things of man."
MARK|8|34|And he called to him the crowd with his disciples and said to them, "If anyone would come after me, let him deny himself and take up his cross and follow me.
MARK|8|35|For whoever would save his life will lose it, but whoever loses his life for my sake and the gospel's will save it.
MARK|8|36|For what does it profit a man to gain the whole world and forfeit his life?
MARK|8|37|For what can a man give in return for his life?
MARK|8|38|For whoever is ashamed of me and of my words in this adulterous and sinful generation, of him will the Son of Man also be ashamed when he comes in the glory of his Father with the holy angels."
MARK|9|1|And he said to them, "Truly, I say to you, there are some standing here who will not taste death until they see the kingdom of God after it has come with power."
MARK|9|2|And after six days Jesus took with him Peter and James and John, and led them up a high mountain by themselves. And he was transfigured before them,
MARK|9|3|and his clothes became radiant, intensely white, as no one on earth could bleach them.
MARK|9|4|And there appeared to them Elijah with Moses, and they were talking with Jesus.
MARK|9|5|And Peter said to Jesus, "Rabbi, it is good that we are here. Let us make three tents, one for you and one for Moses and one for Elijah."
MARK|9|6|For he did not know what to say, for they were terrified.
MARK|9|7|And a cloud overshadowed them, and a voice came out of the cloud, "This is my beloved Son; listen to him."
MARK|9|8|And suddenly, looking around, they no longer saw anyone with them but Jesus only.
MARK|9|9|And as they were coming down the mountain, he charged them to tell no one what they had seen, until the Son of Man had risen from the dead.
MARK|9|10|So they kept the matter to themselves, questioning what this rising from the dead might mean.
MARK|9|11|And they asked him, "Why do the scribes say that first Elijah must come?"
MARK|9|12|And he said to them, "Elijah does come first to restore all things. And how is it written of the Son of Man that he should suffer many things and be treated with contempt?
MARK|9|13|But I tell you that Elijah has come, and they did to him whatever they pleased, as it is written of him."
MARK|9|14|And when they came to the disciples, they saw a great crowd around them, and scribes arguing with them.
MARK|9|15|And immediately all the crowd, when they saw him, were greatly amazed and ran up to him and greeted him.
MARK|9|16|And he asked them, "What are you arguing about with them?"
MARK|9|17|And someone from the crowd answered him, "Teacher, I brought my son to you, for he has a spirit that makes him mute.
MARK|9|18|And whenever it seizes him, it throws him down, and he foams and grinds his teeth and becomes rigid. So I asked your disciples to cast it out, and they were not able."
MARK|9|19|And he answered them, "O faithless generation, how long am I to be with you? How long am I to bear with you? Bring him to me."
MARK|9|20|And they brought the boy to him. And when the spirit saw him, immediately it convulsed the boy, and he fell on the ground and rolled about, foaming at the mouth.
MARK|9|21|And Jesus asked his father, "How long has this been happening to him?" And he said, "From childhood.
MARK|9|22|And it has often cast him into fire and into water, to destroy him. But if you can do anything, have compassion on us and help us."
MARK|9|23|And Jesus said to him, "If you can! All things are possible for one who believes."
MARK|9|24|Immediately the father of the child cried out and said, "I believe; help my unbelief!"
MARK|9|25|And when Jesus saw that a crowd came running together, he rebuked the unclean spirit, saying to it, "You mute and deaf spirit, I command you, come out of him and never enter him again."
MARK|9|26|And after crying out and convulsing him terribly, it came out, and the boy was like a corpse, so that most of them said, "He is dead."
MARK|9|27|But Jesus took him by the hand and lifted him up, and he arose.
MARK|9|28|And when he had entered the house, his disciples asked him privately, "Why could we not cast it out?"
MARK|9|29|And he said to them, "This kind cannot be driven out by anything but prayer."
MARK|9|30|They went on from there and passed through Galilee. And he did not want anyone to know,
MARK|9|31|for he was teaching his disciples, saying to them, "The Son of Man is going to be delivered into the hands of men, and they will kill him. And when he is killed, after three days he will rise."
MARK|9|32|But they did not understand the saying, and were afraid to ask him.
MARK|9|33|And they came to Capernaum. And when he was in the house he asked them, "What were you discussing on the way?"
MARK|9|34|But they kept silent, for on the way they had argued with one another about who was the greatest.
MARK|9|35|And he sat down and called the twelve. And he said to them, "If anyone would be first, he must be last of all and servant of all."
MARK|9|36|And he took a child and put him in the midst of them, and taking him in his arms, he said to them,
MARK|9|37|"Whoever receives one such child in my name receives me, and whoever receives me, receives not me but him who sent me."
MARK|9|38|John said to him, "Teacher, we saw someone casting out demons in your name, and we tried to stop him, because he was not following us."
MARK|9|39|But Jesus said, "Do not stop him, for no one who does a mighty work in my name will be able soon afterward to speak evil of me.
MARK|9|40|For the one who is not against us is for us.
MARK|9|41|For truly, I say to you, whoever gives you a cup of water to drink because you belong to Christ will by no means lose his reward.
MARK|9|42|"Whoever causes one of these little ones who believe in me to sin, it would be better for him if a great millstone were hung around his neck and he were thrown into the sea.
MARK|9|43|And if your hand causes you to sin, cut it off. It is better for you to enter life crippled than with two hands to go to hell, to the unquenchable fire.
MARK|9|44|***
MARK|9|45|And if your foot causes you to sin, cut it off. It is better for you to enter life lame than with two feet to be thrown into hell.
MARK|9|46|***
MARK|9|47|And if your eye causes you to sin, tear it out. It is better for you to enter the kingdom of God with one eye than with two eyes to be thrown into hell,
MARK|9|48|'where their worm does not die and the fire is not quenched.'
MARK|9|49|For everyone will be salted with fire.
MARK|9|50|Salt is good, but if the salt has lost its saltiness, how will you make it salty again? Have salt in yourselves, and be at peace with one another."
MARK|10|1|And he left there and went to the region of Judea and beyond the Jordan, and crowds gathered to him again. And again, as was his custom, he taught them.
MARK|10|2|And Pharisees came up and in order to test him asked, "Is it lawful for a man to divorce his wife?"
MARK|10|3|He answered them, "What did Moses command you?"
MARK|10|4|They said, "Moses allowed a man to write a certificate of divorce and to send her away."
MARK|10|5|And Jesus said to them, "Because of your hardness of heart he wrote you this commandment.
MARK|10|6|But from the beginning of creation, 'God made them male and female.'
MARK|10|7|'Therefore a man shall leave his father and mother and hold fast to his wife,
MARK|10|8|and they shall become one flesh.' So they are no longer two but one flesh.
MARK|10|9|What therefore God has joined together, let not man separate."
MARK|10|10|And in the house the disciples asked him again about this matter.
MARK|10|11|And he said to them, "Whoever divorces his wife and marries another commits adultery against her,
MARK|10|12|and if she divorces her husband and marries another, she commits adultery."
MARK|10|13|And they were bringing children to him that he might touch them, and the disciples rebuked them.
MARK|10|14|But when Jesus saw it, he was indignant and said to them, "Let the children come to me; do not hinder them, for to such belongs the kingdom of God.
MARK|10|15|Truly, I say to you, whoever does not receive the kingdom of God like a child shall not enter it."
MARK|10|16|And he took them in his arms and blessed them, laying his hands on them.
MARK|10|17|And as he was setting out on his journey, a man ran up and knelt before him and asked him, "Good Teacher, what must I do to inherit eternal life?"
MARK|10|18|And Jesus said to him, "Why do you call me good? No one is good except God alone.
MARK|10|19|You know the commandments: 'Do not murder, Do not commit adultery, Do not steal, Do not bear false witness, Do not defraud, Honor your father and mother.'"
MARK|10|20|And he said to him, "Teacher, all these I have kept from my youth."
MARK|10|21|And Jesus, looking at him, loved him, and said to him, "You lack one thing: go, sell all that you have and give to the poor, and you will have treasure in heaven; and come, follow me."
MARK|10|22|Disheartened by the saying, he went away sorrowful, for he had great possessions.
MARK|10|23|And Jesus looked around and said to his disciples, "How difficult it will be for those who have wealth to enter the kingdom of God!"
MARK|10|24|And the disciples were amazed at his words. But Jesus said to them again, "Children, how difficult it is to enter the kingdom of God!
MARK|10|25|It is easier for a camel to go through the eye of a needle than for a rich person to enter the kingdom of God."
MARK|10|26|And they were exceedingly astonished, and said to him, "Then who can be saved?"
MARK|10|27|Jesus looked at them and said, "With man it is impossible, but not with God. For all things are possible with God."
MARK|10|28|Peter began to say to him, "See, we have left everything and followed you."
MARK|10|29|Jesus said, "Truly, I say to you, there is no one who has left house or brothers or sisters or mother or father or children or lands, for my sake and for the gospel,
MARK|10|30|who will not receive a hundredfold now in this time, houses and brothers and sisters and mothers and children and lands, with persecutions, and in the age to come eternal life.
MARK|10|31|But many who are first will be last, and the last first."
MARK|10|32|And they were on the road, going up to Jerusalem, and Jesus was walking ahead of them. And they were amazed, and those who followed were afraid. And taking the twelve again, he began to tell them what was to happen to him,
MARK|10|33|saying, "See, we are going up to Jerusalem, and the Son of Man will be delivered over to the chief priests and the scribes, and they will condemn him to death and deliver him over to the Gentiles.
MARK|10|34|And they will mock him and spit on him, and flog him and kill him. And after three days he will rise."
MARK|10|35|And James and John, the sons of Zebedee, came up to him and said to him, "Teacher, we want you to do for us whatever we ask of you."
MARK|10|36|And he said to them, "What do you want me to do for you?"
MARK|10|37|And they said to him, "Grant us to sit, one at your right hand and one at your left, in your glory."
MARK|10|38|Jesus said to them, "You do not know what you are asking. Are you able to drink the cup that I drink, or to be baptized with the baptism with which I am baptized?"
MARK|10|39|And they said to him, "We are able." And Jesus said to them, "The cup that I drink you will drink, and with the baptism with which I am baptized, you will be baptized,
MARK|10|40|but to sit at my right hand or at my left is not mine to grant, but it is for those for whom it has been prepared."
MARK|10|41|And when the ten heard it, they began to be indignant at James and John.
MARK|10|42|And Jesus called them to him and said to them, "You know that those who are considered rulers of the Gentiles lord it over them, and their great ones exercise authority over them.
MARK|10|43|But it shall not be so among you. But whoever would be great among you must be your servant,
MARK|10|44|and whoever would be first among you must be slave of all.
MARK|10|45|For even the Son of Man came not to be served but to serve, and to give his life as a ransom for many."
MARK|10|46|And they came to Jericho. And as he was leaving Jericho with his disciples and a great crowd, Bartimaeus, a blind beggar, the son of Timaeus, was sitting by the roadside.
MARK|10|47|And when he heard that it was Jesus of Nazareth, he began to cry out and say, "Jesus, Son of David, have mercy on me!"
MARK|10|48|And many rebuked him, telling him to be silent. But he cried out all the more, "Son of David, have mercy on me!"
MARK|10|49|And Jesus stopped and said, "Call him." And they called the blind man, saying to him, "Take heart. Get up; he is calling you."
MARK|10|50|And throwing off his cloak, he sprang up and came to Jesus.
MARK|10|51|And Jesus said to him, "What do you want me to do for you?" And the blind man said to him, "Rabbi, let me recover my sight."
MARK|10|52|And Jesus said to him, "Go your way; your faith has made you well." And immediately he recovered his sight and followed him on the way.
MARK|11|1|Now when they drew near to Jerusalem, to Bethphage and Bethany, at the Mount of Olives, Jesus sent two of his disciples
MARK|11|2|and said to them, "Go into the village in front of you, and immediately as you enter it you will find a colt tied, on which no one has ever sat. Untie it and bring it.
MARK|11|3|If anyone says to you, 'Why are you doing this?' say, 'The Lord has need of it and will send it back here immediately.'"
MARK|11|4|And they went away and found a colt tied at a door outside in the street, and they untied it.
MARK|11|5|And some of those standing there said to them, "What are you doing, untying the colt?"
MARK|11|6|And they told them what Jesus had said, and they let them go.
MARK|11|7|And they brought the colt to Jesus and threw their cloaks on it, and he sat on it.
MARK|11|8|And many spread their cloaks on the road, and others spread leafy branches that they had cut from the fields.
MARK|11|9|And those who went before and those who followed were shouting, "Hosanna! Blessed is he who comes in the name of the Lord!
MARK|11|10|Blessed is the coming kingdom of our father David! Hosanna in the highest!"
MARK|11|11|And he entered Jerusalem and went into the temple. And when he had looked around at everything, as it was already late, he went out to Bethany with the twelve.
MARK|11|12|On the following day, when they came from Bethany, he was hungry.
MARK|11|13|And seeing in the distance a fig tree in leaf, he went to see if he could find anything on it. When he came to it, he found nothing but leaves, for it was not the season for figs.
MARK|11|14|And he said to it, "May no one ever eat fruit from you again." And his disciples heard it.
MARK|11|15|And they came to Jerusalem. And he entered the temple and began to drive out those who sold and those who bought in the temple, and he overturned the tables of the money-changers and the seats of those who sold pigeons.
MARK|11|16|And he would not allow anyone to carry anything through the temple.
MARK|11|17|And he was teaching them and saying to them, "Is it not written, 'My house shall be called a house of prayer for all the nations'? But you have made it a den of robbers."
MARK|11|18|And the chief priests and the scribes heard it and were seeking a way to destroy him, for they feared him, because all the crowd was astonished at his teaching.
MARK|11|19|And when evening came they went out of the city.
MARK|11|20|As they passed by in the morning, they saw the fig tree withered away to its roots.
MARK|11|21|And Peter remembered and said to him, "Rabbi, look! The fig tree that you cursed has withered."
MARK|11|22|And Jesus answered them, "Have faith in God.
MARK|11|23|Truly, I say to you, whoever says to this mountain, 'Be taken up and thrown into the sea,' and does not doubt in his heart, but believes that what he says will come to pass, it will be done for him.
MARK|11|24|Therefore I tell you, whatever you ask in prayer, believe that you have received it, and it will be yours.
MARK|11|25|And whenever you stand praying, forgive, if you have anything against anyone, so that your Father also who is in heaven may forgive you your trespasses."
MARK|11|26|***
MARK|11|27|And they came again to Jerusalem. And as he was walking in the temple, the chief priests and the scribes and the elders came to him,
MARK|11|28|and they said to him, "By what authority are you doing these things, or who gave you this authority to do them?"
MARK|11|29|Jesus said to them, "I will ask you one question; answer me, and I will tell you by what authority I do these things.
MARK|11|30|Was the baptism of John from heaven or from man? Answer me."
MARK|11|31|And they discussed it with one another, saying, "If we say, 'From heaven,' he will say, 'Why then did you not believe him?'
MARK|11|32|But shall we say, 'From man'?"- they were afraid of the people, for they all held that John really was a prophet.
MARK|11|33|So they answered Jesus, "We do not know." And Jesus said to them, "Neither will I tell you by what authority I do these things."
MARK|12|1|And he began to speak to them in parables. "A man planted a vineyard and put a fence around it and dug a pit for the winepress and built a tower, and leased it to tenants and went into another country.
MARK|12|2|When the season came, he sent a servant to the tenants to get from them some of the fruit of the vineyard.
MARK|12|3|And they took him and beat him and sent him away empty-handed.
MARK|12|4|Again he sent to them another servant, and they struck him on the head and treated him shamefully.
MARK|12|5|And he sent another, and him they killed. And so with many others: some they beat, and some they killed.
MARK|12|6|He had still one other, a beloved son. Finally he sent him to them, saying, 'They will respect my son.'
MARK|12|7|But those tenants said to one another, 'This is the heir. Come, let us kill him, and the inheritance will be ours.'
MARK|12|8|And they took him and killed him and threw him out of the vineyard.
MARK|12|9|What will the owner of the vineyard do? He will come and destroy the tenants and give the vineyard to others.
MARK|12|10|Have you not read this Scripture: "' The stone that the builders rejected has become the cornerstone;
MARK|12|11|this was the Lord's doing, and it is marvelous in our eyes'?"
MARK|12|12|And they were seeking to arrest him but feared the people, for they perceived that he had told the parable against them. So they left him and went away.
MARK|12|13|And they sent to him some of the Pharisees and some of the Herodians, to trap him in his talk.
MARK|12|14|And they came and said to him, "Teacher, we know that you are true and do not care about anyone's opinion. For you are not swayed by appearances, but truly teach the way of God. Is it lawful to pay taxes to Caesar, or not? Should we pay them, or should we not?"
MARK|12|15|But, knowing their hypocrisy, he said to them, "Why put me to the test? Bring me a denarius and let me look at it."
MARK|12|16|And they brought one. And he said to them, "Whose likeness and inscription is this?" They said to him, "Caesar's."
MARK|12|17|Jesus said to them, "Render to Caesar the things that are Caesar's, and to God the things that are God's." And they marveled at him.
MARK|12|18|And Sadducees came to him, who say that there is no resurrection. And they asked him a question, saying,
MARK|12|19|"Teacher, Moses wrote for us that if a man's brother dies and leaves a wife, but leaves no child, the man must take the widow and raise up offspring for his brother.
MARK|12|20|There were seven brothers; the first took a wife, and when he died left no offspring.
MARK|12|21|And the second took her, and died, leaving no offspring. And the third likewise.
MARK|12|22|And the seven left no offspring. Last of all the woman also died.
MARK|12|23|In the resurrection, when they rise again, whose wife will she be? For the seven had her as wife."
MARK|12|24|Jesus said to them, "Is this not the reason you are wrong, because you know neither the Scriptures nor the power of God?
MARK|12|25|For when they rise from the dead, they neither marry nor are given in marriage, but are like angels in heaven.
MARK|12|26|And as for the dead being raised, have you not read in the book of Moses, in the passage about the bush, how God spoke to him, saying, 'I am the God of Abraham, and the God of Isaac, and the God of Jacob'?
MARK|12|27|He is not God of the dead, but of the living. You are quite wrong."
MARK|12|28|And one of the scribes came up and heard them disputing with one another, and seeing that he answered them well, asked him, "Which commandment is the most important of all?"
MARK|12|29|Jesus answered, "The most important is, 'Hear, O Israel: The Lord our God, the Lord is one.
MARK|12|30|And you shall love the Lord your God with all your heart and with all your soul and with all your mind and with all your strength.'
MARK|12|31|The second is this: 'You shall love your neighbor as yourself.' There is no other commandment greater than these."
MARK|12|32|And the scribe said to him, "You are right, Teacher. You have truly said that he is one, and there is no other besides him.
MARK|12|33|And to love him with all the heart and with all the understanding and with all the strength, and to love one's neighbor as oneself, is much more than all whole burnt offerings and sacrifices."
MARK|12|34|And when Jesus saw that he answered wisely, he said to him, "You are not far from the kingdom of God." And after that no one dared to ask him any more questions.
MARK|12|35|And as Jesus taught in the temple, he said, "How can the scribes say that the Christ is the son of David?
MARK|12|36|David himself, in the Holy Spirit, declared, "' The Lord said to my Lord, Sit at my right hand, until I put your enemies under your feet.'
MARK|12|37|David himself calls him Lord. So how is he his son?" And the great throng heard him gladly.
MARK|12|38|And in his teaching he said, "Beware of the scribes, who like to walk around in long robes and like greetings in the marketplaces
MARK|12|39|and have the best seats in the synagogues and the places of honor at feasts,
MARK|12|40|who devour widows' houses and for a pretense make long prayers. They will receive the greater condemnation."
MARK|12|41|And he sat down opposite the treasury and watched the people putting money into the offering box. Many rich people put in large sums.
MARK|12|42|And a poor widow came and put in two small copper coins, which make a penny.
MARK|12|43|And he called his disciples to him and said to them, "Truly, I say to you, this poor widow has put in more than all those who are contributing to the offering box.
MARK|12|44|For they all contributed out of their abundance, but she out of her poverty has put in everything she had, all she had to live on."
MARK|13|1|And as he came out of the temple, one of his disciples said to him, "Look, Teacher, what wonderful stones and what wonderful buildings!"
MARK|13|2|And Jesus said to him, "Do you see these great buildings? There will not be left here one stone upon another that will not be thrown down."
MARK|13|3|And as he sat on the Mount of Olives opposite the temple, Peter and James and John and Andrew asked him privately,
MARK|13|4|"Tell us, when will these things be, and what will be the sign when all these things are about to be accomplished?"
MARK|13|5|And Jesus began to say to them, "See that no one leads you astray.
MARK|13|6|Many will come in my name, saying, 'I am he!' and they will lead many astray.
MARK|13|7|And when you hear of wars and rumors of wars, do not be alarmed. This must take place, but the end is not yet.
MARK|13|8|For nation will rise against nation, and kingdom against kingdom. There will be earthquakes in various places; there will be famines. These are but the beginning of the birth pains.
MARK|13|9|"But be on your guard. For they will deliver you over to councils, and you will be beaten in synagogues, and you will stand before governors and kings for my sake, to bear witness before them.
MARK|13|10|And the gospel must first be proclaimed to all nations.
MARK|13|11|And when they bring you to trial and deliver you over, do not be anxious beforehand what you are to say, but say whatever is given you in that hour, for it is not you who speak, but the Holy Spirit.
MARK|13|12|And brother will deliver brother over to death, and the father his child, and children will rise against parents and have them put to death.
MARK|13|13|And you will be hated by all for my name's sake. But the one who endures to the end will be saved.
MARK|13|14|"But when you see the abomination of desolation standing where it ought not to be (let the reader understand), then let those who are in Judea flee to the mountains.
MARK|13|15|Let the one who is on the housetop not go down, nor enter his house, to take anything out,
MARK|13|16|and let the one who is in the field not turn back to take his cloak.
MARK|13|17|And alas for women who are pregnant and for those who are nursing infants in those days!
MARK|13|18|Pray that it may not happen in winter.
MARK|13|19|For in those days there will be such tribulation as has not been from the beginning of the creation that God created until now, and never will be.
MARK|13|20|And if the Lord had not cut short the days, no human being would be saved. But for the sake of the elect, whom he chose, he shortened the days.
MARK|13|21|And then if anyone says to you, 'Look, here is the Christ!' or 'Look, there he is!' do not believe it.
MARK|13|22|False christs and false prophets will arise and perform signs and wonders, to lead astray, if possible, the elect.
MARK|13|23|But be on guard; I have told you all things beforehand.
MARK|13|24|"But in those days, after that tribulation, the sun will be darkened, and the moon will not give its light,
MARK|13|25|and the stars will be falling from heaven, and the powers in the heavens will be shaken.
MARK|13|26|And then they will see the Son of Man coming in clouds with great power and glory.
MARK|13|27|And then he will send out the angels and gather his elect from the four winds, from the ends of the earth to the ends of heaven.
MARK|13|28|"From the fig tree learn its lesson: as soon as its branch becomes tender and puts out its leaves, you know that summer is near.
MARK|13|29|So also, when you see these things taking place, you know that he is near, at the very gates.
MARK|13|30|Truly, I say to you, this generation will not pass away until all these things take place.
MARK|13|31|Heaven and earth will pass away, but my words will not pass away.
MARK|13|32|"But concerning that day or that hour, no one knows, not even the angels in heaven, nor the Son, but only the Father.
MARK|13|33|Be on guard, keep awake. For you do not know when the time will come.
MARK|13|34|It is like a man going on a journey, when he leaves home and puts his servants in charge, each with his work, and commands the doorkeeper to stay awake.
MARK|13|35|Therefore stay awake- for you do not know when the master of the house will come, in the evening, or at midnight, or when the cock crows, or in the morning-
MARK|13|36|lest he come suddenly and find you asleep.
MARK|13|37|And what I say to you I say to all: Stay awake."
MARK|14|1|It was now two days before the Passover and the Feast of Unleavened Bread. And the chief priests and the scribes were seeking how to arrest him by stealth and kill him,
MARK|14|2|for they said, "Not during the feast, lest there be an uproar from the people."
MARK|14|3|And while he was at Bethany in the house of Simon the leper, as he was reclining at table, a woman came with an alabaster flask of ointment of pure nard, very costly, and she broke the flask and poured it over his head.
MARK|14|4|There were some who said to themselves indignantly, "Why was the ointment wasted like that?
MARK|14|5|For this ointment could have been sold for more than three hundred denarii and given to the poor." And they scolded her.
MARK|14|6|But Jesus said, "Leave her alone. Why do you trouble her? She has done a beautiful thing to me.
MARK|14|7|For you always have the poor with you, and whenever you want, you can do good for them. But you will not always have me.
MARK|14|8|She has done what she could; she has anointed my body beforehand for burial.
MARK|14|9|And truly, I say to you, wherever the gospel is proclaimed in the whole world, what she has done will be told in memory of her."
MARK|14|10|Then Judas Iscariot, who was one of the twelve, went to the chief priests in order to betray him to them.
MARK|14|11|And when they heard it, they were glad and promised to give him money. And he sought an opportunity to betray him.
MARK|14|12|And on the first day of Unleavened Bread, when they sacrificed the Passover lamb, his disciples said to him, "Where will you have us go and prepare for you to eat the Passover?"
MARK|14|13|And he sent two of his disciples and said to them, "Go into the city, and a man carrying a jar of water will meet you. Follow him,
MARK|14|14|and wherever he enters, say to the master of the house, 'The Teacher says, Where is my guest room, where I may eat the Passover with my disciples?'
MARK|14|15|And he will show you a large upper room furnished and ready; there prepare for us."
MARK|14|16|And the disciples set out and went to the city and found it just as he had told them, and they prepared the Passover.
MARK|14|17|And when it was evening, he came with the twelve.
MARK|14|18|And as they were reclining at table and eating, Jesus said, "Truly, I say to you, one of you will betray me, one who is eating with me."
MARK|14|19|They began to be sorrowful and to say to him one after another, "Is it I?"
MARK|14|20|He said to them, "It is one of the twelve, one who is dipping bread into the dish with me.
MARK|14|21|For the Son of Man goes as it is written of him, but woe to that man by whom the Son of Man is betrayed! It would have been better for that man if he had not been born."
MARK|14|22|And as they were eating, he took bread, and after blessing it broke it and gave it to them, and said, "Take; this is my body."
MARK|14|23|And he took a cup, and when he had given thanks he gave it to them, and they all drank of it.
MARK|14|24|And he said to them, "This is my blood of the covenant, which is poured out for many.
MARK|14|25|Truly, I say to you, I will not drink again of the fruit of the vine until that day when I drink it new in the kingdom of God."
MARK|14|26|And when they had sung a hymn, they went out to the Mount of Olives.
MARK|14|27|And Jesus said to them, "You will all fall away, for it is written, 'I will strike the shepherd, and the sheep will be scattered.'
MARK|14|28|But after I am raised up, I will go before you to Galilee."
MARK|14|29|Peter said to him, "Even though they all fall away, I will not."
MARK|14|30|And Jesus said to him, "Truly, I tell you, this very night, before the rooster crows twice, you will deny me three times."
MARK|14|31|But he said emphatically, "If I must die with you, I will not deny you." And they all said the same.
MARK|14|32|And they went to a place called Gethsemane. And he said to his disciples, "Sit here while I pray."
MARK|14|33|And he took with him Peter and James and John, and began to be greatly distressed and troubled.
MARK|14|34|And he said to them, "My soul is very sorrowful, even to death. Remain here and watch."
MARK|14|35|And going a little farther, he fell on the ground and prayed that, if it were possible, the hour might pass from him.
MARK|14|36|And he said, "Abba, Father, all things are possible for you. Remove this cup from me. Yet not what I will, but what you will."
MARK|14|37|And he came and found them sleeping, and he said to Peter, "Simon, are you asleep? Could you not watch one hour?
MARK|14|38|Watch and pray that you may not enter into temptation. The spirit indeed is willing, but the flesh is weak."
MARK|14|39|And again he went away and prayed, saying the same words.
MARK|14|40|And again he came and found them sleeping, for their eyes were very heavy, and they did not know what to answer him.
MARK|14|41|And he came the third time and said to them, "Are you still sleeping and taking your rest? It is enough; the hour has come. The Son of Man is betrayed into the hands of sinners.
MARK|14|42|Rise, let us be going; see, my betrayer is at hand."
MARK|14|43|And immediately, while he was still speaking, Judas came, one of the twelve, and with him a crowd with swords and clubs, from the chief priests and the scribes and the elders.
MARK|14|44|Now the betrayer had given them a sign, saying, "The one I will kiss is the man. Seize him and lead him away under guard."
MARK|14|45|And when he came, he went up to him at once and said, "Rabbi!" And he kissed him.
MARK|14|46|And they laid hands on him and seized him.
MARK|14|47|But one of those who stood by drew his sword and struck the servant of the high priest and cut off his ear.
MARK|14|48|And Jesus said to them, "Have you come out as against a robber, with swords and clubs to capture me?
MARK|14|49|Day after day I was with you in the temple teaching, and you did not seize me. But let the Scriptures be fulfilled."
MARK|14|50|And they all left him and fled.
MARK|14|51|And a young man followed him, with nothing but a linen cloth about his body. And they seized him,
MARK|14|52|but he left the linen cloth and ran away naked.
MARK|14|53|And they led Jesus to the high priest. And all the chief priests and the elders and the scribes came together.
MARK|14|54|And Peter had followed him at a distance, right into the courtyard of the high priest. And he was sitting with the guards and warming himself at the fire.
MARK|14|55|Now the chief priests and the whole Council were seeking testimony against Jesus to put him to death, but they found none.
MARK|14|56|For many bore false witness against him, but their testimony did not agree.
MARK|14|57|And some stood up and bore false witness against him, saying,
MARK|14|58|"We heard him say, 'I will destroy this temple that is made with hands, and in three days I will build another, not made with hands.'"
MARK|14|59|Yet even about this their testimony did not agree.
MARK|14|60|And the high priest stood up in the midst and asked Jesus, "Have you no answer to make? What is it that these men testify against you?"
MARK|14|61|But he remained silent and made no answer. Again the high priest asked him, "Are you the Christ, the Son of the Blessed?"
MARK|14|62|And Jesus said, "I am, and you will see the Son of Man seated at the right hand of Power, and coming with the clouds of heaven."
MARK|14|63|And the high priest tore his garments and said, "What further witnesses do we need?
MARK|14|64|You have heard his blasphemy. What is your decision?" And they all condemned him as deserving death.
MARK|14|65|And some began to spit on him and to cover his face and to strike him, saying to him, "Prophesy!" And the guards received him with blows.
MARK|14|66|And as Peter was below in the courtyard, one of the servant girls of the high priest came,
MARK|14|67|and seeing Peter warming himself, she looked at him and said, "You also were with the Nazarene, Jesus."
MARK|14|68|But he denied it, saying, "I neither know nor understand what you mean." And he went out into the gateway and the rooster crowed.
MARK|14|69|And the servant girl saw him and began again to say to the bystanders, "This man is one of them."
MARK|14|70|But again he denied it. And after a little while the bystanders again said to Peter, "Certainly you are one of them, for you are a Galilean."
MARK|14|71|But he began to invoke a curse on himself and to swear, "I do not know this man of whom you speak."
MARK|14|72|And immediately the rooster crowed a second time. And Peter remembered how Jesus had said to him, "Before the rooster crows twice, you will deny me three times." And he broke down and wept.
MARK|15|1|And as soon as it was morning, the chief priests held a consultation with the elders and scribes and the whole Council. And they bound Jesus and led him away and delivered him over to Pilate.
MARK|15|2|And Pilate asked him, "Are you the King of the Jews?" And he answered him, "You have said so."
MARK|15|3|And the chief priests accused him of many things.
MARK|15|4|And Pilate again asked him, "Have you no answer to make? See how many charges they bring against you."
MARK|15|5|But Jesus made no further answer, so that Pilate was amazed.
MARK|15|6|Now at the feast he used to release for them one prisoner for whom they asked.
MARK|15|7|And among the rebels in prison, who had committed murder in the insurrection, there was a man called Barabbas.
MARK|15|8|And the crowd came up and began to ask Pilate to do as he usually did for them.
MARK|15|9|And he answered them, saying, "Do you want me to release for you the King of the Jews?"
MARK|15|10|For he perceived that it was out of envy that the chief priests had delivered him up.
MARK|15|11|But the chief priests stirred up the crowd to have him release for them Barabbas instead.
MARK|15|12|And Pilate again said to them, "Then what shall I do with the man you call the King of the Jews?"
MARK|15|13|And they cried out again, "Crucify him."
MARK|15|14|And Pilate said to them, "Why, what evil has he done?" But they shouted all the more, "Crucify him."
MARK|15|15|So Pilate, wishing to satisfy the crowd, released for them Barabbas, and having scourged Jesus, he delivered him to be crucified.
MARK|15|16|And the soldiers led him away inside the palace (that is, the governor's headquarters), and they called together the whole battalion.
MARK|15|17|And they clothed him in a purple cloak, and twisting together a crown of thorns, they put it on him.
MARK|15|18|And they began to salute him, "Hail, King of the Jews!"
MARK|15|19|And they were striking his head with a reed and spitting on him and kneeling down in homage to him.
MARK|15|20|And when they had mocked him, they stripped him of the purple cloak and put his own clothes on him. And they led him out to crucify him.
MARK|15|21|And they compelled a passerby, Simon of Cyrene, who was coming in from the country, the father of Alexander and Rufus, to carry his cross.
MARK|15|22|And they brought him to the place called Golgotha (which means Place of a Skull).
MARK|15|23|And they offered him wine mixed with myrrh, but he did not take it.
MARK|15|24|And they crucified him and divided his garments among them, casting lots for them, to decide what each should take.
MARK|15|25|And it was the third hour when they crucified him.
MARK|15|26|And the inscription of the charge against him read, "The King of the Jews."
MARK|15|27|And with him they crucified two robbers, one on his right and one on his left.
MARK|15|28|***
MARK|15|29|And those who passed by derided him, wagging their heads and saying, "Aha! You who would destroy the temple and rebuild it in three days,
MARK|15|30|save yourself, and come down from the cross!"
MARK|15|31|So also the chief priests with the scribes mocked him to one another, saying, "He saved others; he cannot save himself.
MARK|15|32|Let the Christ, the King of Israel, come down now from the cross that we may see and believe." Those who were crucified with him also reviled him.
MARK|15|33|And when the sixth hour had come, there was darkness over the whole land until the ninth hour.
MARK|15|34|And at the ninth hour Jesus cried with a loud voice, "Eloi, Eloi, lema sabachthani?" which means, "My God, my God, why have you forsaken me?"
MARK|15|35|And some of the bystanders hearing it said, "Behold, he is calling Elijah."
MARK|15|36|And someone ran and filled a sponge with sour wine, put it on a reed and gave it to him to drink, saying, "Wait, let us see whether Elijah will come to take him down."
MARK|15|37|And Jesus uttered a loud cry and breathed his last.
MARK|15|38|And the curtain of the temple was torn in two, from top to bottom.
MARK|15|39|And when the centurion, who stood facing him, saw that in this way he breathed his last, he said, "Truly this man was the Son of God!"
MARK|15|40|There were also women looking on from a distance, among whom were Mary Magdalene, and Mary the mother of James the younger and of Joses, and Salome.
MARK|15|41|When he was in Galilee, they followed him and ministered to him, and there were also many other women who came up with him to Jerusalem.
MARK|15|42|And when evening had come, since it was the day of Preparation, that is, the day before the Sabbath,
MARK|15|43|Joseph of Arimathea, a respected member of the Council, who was also himself looking for the kingdom of God, took courage and went to Pilate and asked for the body of Jesus.
MARK|15|44|Pilate was surprised to hear that he should have already died. And summoning the centurion, he asked him whether he was already dead.
MARK|15|45|And when he learned from the centurion that he was dead, he granted the corpse to Joseph.
MARK|15|46|And Joseph bought a linen shroud, and taking him down, wrapped him in the linen shroud and laid him in a tomb that had been cut out of the rock. And he rolled a stone against the entrance of the tomb.
MARK|15|47|Mary Magdalene and Mary the mother of Joses saw where he was laid.
MARK|16|1|When the Sabbath was past, Mary Magdalene and Mary the mother of James and Salome bought spices, so that they might go and anoint him.
MARK|16|2|And very early on the first day of the week, when the sun had risen, they went to the tomb.
MARK|16|3|And they were saying to one another, "Who will roll away the stone for us from the entrance of the tomb?"
MARK|16|4|And looking up, they saw that the stone had been rolled back- it was very large.
MARK|16|5|And entering the tomb, they saw a young man sitting on the right side, dressed in a white robe, and they were alarmed.
MARK|16|6|And he said to them, "Do not be alarmed. You seek Jesus of Nazareth, who was crucified. He has risen; he is not here. See the place where they laid him.
MARK|16|7|But go, tell his disciples and Peter that he is going before you to Galilee. There you will see him, just as he told you."
MARK|16|8|And they went out and fled from the tomb, for trembling and astonishment had seized them, and they said nothing to anyone, for they were afraid. [SOME OF THE EARLIEST MANUSCRIPTS DO NOT INCLUDE 16:9-20.]
MARK|16|9|[[Now when he rose early on the first day of the week, he appeared first to Mary Magdalene, from whom he had cast out seven demons.
MARK|16|10|She went and told those who had been with him, as they mourned and wept.
MARK|16|11|But when they heard that he was alive and had been seen by her, they would not believe it.
MARK|16|12|After these things he appeared in another form to two of them, as they were walking into the country.
MARK|16|13|And they went back and told the rest, but they did not believe them.
MARK|16|14|Afterward he appeared to the eleven themselves as they were reclining at table, and he rebuked them for their unbelief and hardness of heart, because they had not believed those who saw him after he had risen.
MARK|16|15|And he said to them, "Go into all the world and proclaim the gospel to the whole creation.
MARK|16|16|Whoever believes and is baptized will be saved, but whoever does not believe will be condemned.
MARK|16|17|And these signs will accompany those who believe: in my name they will cast out demons; they will speak in new tongues;
MARK|16|18|they will pick up serpents with their hands; and if they drink any deadly poison, it will not hurt them; they will lay their hands on the sick, and they will recover."
MARK|16|19|So then the Lord Jesus, after he had spoken to them, was taken up into heaven and sat down at the right hand of God.
MARK|16|20|And they went out and preached everywhere, while the Lord worked with them and confirmed the message by accompanying signs.]]
