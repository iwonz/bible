SONG|1|1|Да лобзает он меня лобзанием уст своих! Ибо ласки твои лучше вина.
SONG|1|2|От благовония мастей твоих имя твое – как разлитое миро; поэтому девицы любят тебя.
SONG|1|3|Влеки меня, мы побежим за тобою; – царь ввел меня в чертоги свои, – будем восхищаться и радоваться тобою, превозносить ласки твои больше, нежели вино; достойно любят тебя!
SONG|1|4|Дщери Иерусалимские! черна я, но красива, как шатры Кидарские, как завесы Соломоновы.
SONG|1|5|Не смотрите на меня, что я смугла, ибо солнце опалило меня: сыновья матери моей разгневались на меня, поставили меня стеречь виноградники, – моего собственного виноградника я не стерегла.
SONG|1|6|Скажи мне, ты, которого любит душа моя: где пасешь ты? где отдыхаешь в полдень? к чему мне быть скиталицею возле стад товарищей твоих?
SONG|1|7|Если ты не знаешь этого, прекраснейшая из женщин, то иди себе по следам овец и паси козлят твоих подле шатров пастушеских.
SONG|1|8|Кобылице моей в колеснице фараоновой я уподобил тебя, возлюбленная моя.
SONG|1|9|Прекрасны ланиты твои под подвесками, шея твоя в ожерельях;
SONG|1|10|золотые подвески мы сделаем тебе с серебряными блестками.
SONG|1|11|Доколе царь был за столом своим, нард мой издавал благовоние свое.
SONG|1|12|Мирровый пучок – возлюбленный мой у меня, у грудей моих пребывает.
SONG|1|13|Как кисть кипера, возлюбленный мой у меня в виноградниках Енгедских.
SONG|1|14|О, ты прекрасна, возлюбленная моя, ты прекрасна! глаза твои голубиные.
SONG|1|15|О, ты прекрасен, возлюбленный мой, и любезен! и ложе у нас – зелень;
SONG|1|16|кровли домов наших – кедры,
SONG|1|17|потолки наши – кипарисы.
SONG|2|1|Я нарцисс Саронский, лилия долин!
SONG|2|2|Что лилия между тернами, то возлюбленная моя между девицами.
SONG|2|3|Что яблоня между лесными деревьями, то возлюбленный мой между юношами. В тени ее люблю я сидеть, и плоды ее сладки для гортани моей.
SONG|2|4|Он ввел меня в дом пира, и знамя его надо мною – любовь.
SONG|2|5|Подкрепите меня вином, освежите меня яблоками, ибо я изнемогаю от любви.
SONG|2|6|Левая рука его у меня под головою, а правая обнимает меня.
SONG|2|7|Заклинаю вас, дщери Иерусалимские, сернами или полевыми ланями: не будите и не тревожьте возлюбленной, доколе ей угодно.
SONG|2|8|Голос возлюбленного моего! вот, он идет, скачет по горам, прыгает по холмам.
SONG|2|9|Друг мой похож на серну или на молодого оленя. Вот, он стоит у нас за стеною, заглядывает в окно, мелькает сквозь решетку.
SONG|2|10|Возлюбленный мой начал говорить мне: встань, возлюбленная моя, прекрасная моя, выйди!
SONG|2|11|Вот, зима уже прошла; дождь миновал, перестал;
SONG|2|12|цветы показались на земле; время пения настало, и голос горлицы слышен в стране нашей;
SONG|2|13|смоковницы распустили свои почки, и виноградные лозы, расцветая, издают благовоние. Встань, возлюбленная моя, прекрасная моя, выйди!
SONG|2|14|Голубица моя в ущелье скалы под кровом утеса! покажи мне лице твое, дай мне услышать голос твой, потому что голос твой сладок и лице твое приятно.
SONG|2|15|Ловите нам лисиц, лисенят, которые портят виноградники, а виноградники наши в цвете.
SONG|2|16|Возлюбленный мой принадлежит мне, а я ему; он пасет между лилиями.
SONG|2|17|Доколе день дышит [прохладою], и убегают тени, возвратись, будь подобен серне или молодому оленю на расселинах гор.
SONG|3|1|На ложе моем ночью искала я того, которого любит душа моя, искала его и не нашла его.
SONG|3|2|Встану же я, пойду по городу, по улицам и площадям, и буду искать того, которого любит душа моя; искала я его и не нашла его.
SONG|3|3|Встретили меня стражи, обходящие город: "не видали ли вы того, которого любит душа моя?"
SONG|3|4|Но едва я отошла от них, как нашла того, которого любит душа моя, ухватилась за него, и не отпустила его, доколе не привела его в дом матери моей и во внутренние комнаты родительницы моей.
SONG|3|5|Заклинаю вас, дщери Иерусалимские, сернами или полевыми ланями: не будите и не тревожьте возлюбленной, доколе ей угодно.
SONG|3|6|Кто эта, восходящая от пустыни как бы столбы дыма, окуриваемая миррою и фимиамом, всякими порошками мироварника?
SONG|3|7|Вот одр его – Соломона: шестьдесят сильных вокруг него, из сильных Израилевых.
SONG|3|8|Все они держат по мечу, опытны в бою; у каждого меч при бедре его ради страха ночного.
SONG|3|9|Носильный одр сделал себе царь Соломон из дерев Ливанских;
SONG|3|10|столпцы его сделал из серебра, локотники его из золота, седалище его из пурпуровой ткани; внутренность его убрана с любовью дщерями Иерусалимскими.
SONG|3|11|Пойдите и посмотрите, дщери Сионские, на царя Соломона в венце, которым увенчала его мать его в день бракосочетания его, в день, радостный для сердца его.
SONG|4|1|О, ты прекрасна, возлюбленная моя, ты прекрасна! глаза твои голубиные под кудрями твоими; волосы твои – как стадо коз, сходящих с горы Галаадской;
SONG|4|2|зубы твои – как стадо выстриженных овец, выходящих из купальни, из которых у каждой пара ягнят, и бесплодной нет между ними;
SONG|4|3|как лента алая губы твои, и уста твои любезны; как половинки гранатового яблока – ланиты твои под кудрями твоими;
SONG|4|4|шея твоя – как столп Давидов, сооруженный для оружий, тысяча щитов висит на нем – все щиты сильных;
SONG|4|5|два сосца твои – как двойни молодой серны, пасущиеся между лилиями.
SONG|4|6|Доколе день дышит [прохладою], и убегают тени, пойду я на гору мирровую и на холм фимиама.
SONG|4|7|Вся ты прекрасна, возлюбленная моя, и пятна нет на тебе!
SONG|4|8|Со мною с Ливана, невеста! со мною иди с Ливана! спеши с вершины Аманы, с вершины Сенира и Ермона, от логовищ львиных, от гор барсовых!
SONG|4|9|Пленила ты сердце мое, сестра моя, невеста! пленила ты сердце мое одним взглядом очей твоих, одним ожерельем на шее твоей.
SONG|4|10|О, как любезны ласки твои, сестра моя, невеста! о, как много ласки твои лучше вина, и благовоние мастей твоих лучше всех ароматов!
SONG|4|11|Сотовый мед каплет из уст твоих, невеста; мед и молоко под языком твоим, и благоухание одежды твоей подобно благоуханию Ливана!
SONG|4|12|Запертый сад – сестра моя, невеста, заключенный колодезь, запечатанный источник:
SONG|4|13|рассадники твои – сад с гранатовыми яблоками, с превосходными плодами, киперы с нардами,
SONG|4|14|нард и шафран, аир и корица со всякими благовонными деревами, мирра и алой со всякими лучшими ароматами;
SONG|4|15|садовый источник – колодезь живых вод и потоки с Ливана.
SONG|4|16|Поднимись [ветер] с севера и принесись с юга, повей на сад мой, – и польются ароматы его! – Пусть придет возлюбленный мой в сад свой и вкушает сладкие плоды его.
SONG|5|1|Пришел я в сад мой, сестра моя, невеста; набрал мирры моей с ароматами моими, поел сотов моих с медом моим, напился вина моего с молоком моим. Ешьте, друзья, пейте и насыщайтесь, возлюбленные!
SONG|5|2|Я сплю, а сердце мое бодрствует; [вот], голос моего возлюбленного, который стучится: "отвори мне, сестра моя, возлюбленная моя, голубица моя, чистая моя! потому что голова моя вся покрыта росою, кудри мои – ночною влагою".
SONG|5|3|Я скинула хитон мой; как же мне опять надевать его? Я вымыла ноги мои; как же мне марать их?
SONG|5|4|Возлюбленный мой протянул руку свою сквозь скважину, и внутренность моя взволновалась от него.
SONG|5|5|Я встала, чтобы отпереть возлюбленному моему, и с рук моих капала мирра, и с перстов моих мирра капала на ручки замка.
SONG|5|6|Отперла я возлюбленному моему, а возлюбленный мой повернулся и ушел. Души во мне не стало, когда он говорил; я искала его и не находила его; звала его, и он не отзывался мне.
SONG|5|7|Встретили меня стражи, обходящие город, избили меня, изранили меня; сняли с меня покрывало стерегущие стены.
SONG|5|8|Заклинаю вас, дщери Иерусалимские: если вы встретите возлюбленного моего, что скажете вы ему? что я изнемогаю от любви.
SONG|5|9|"Чем возлюбленный твой лучше других возлюбленных, прекраснейшая из женщин? Чем возлюбленный твой лучше других, что ты так заклинаешь нас?"
SONG|5|10|Возлюбленный мой бел и румян, лучше десяти тысяч других:
SONG|5|11|голова его – чистое золото; кудри его волнистые, черные, как ворон;
SONG|5|12|глаза его – как голуби при потоках вод, купающиеся в молоке, сидящие в довольстве;
SONG|5|13|щеки его – цветник ароматный, гряды благовонных растений; губы его – лилии, источают текучую мирру;
SONG|5|14|руки его – золотые кругляки, усаженные топазами; живот его – как изваяние из слоновой кости, обложенное сапфирами;
SONG|5|15|голени его – мраморные столбы, поставленные на золотых подножиях; вид его подобен Ливану, величествен, как кедры;
SONG|5|16|уста его – сладость, и весь он – любезность. Вот кто возлюбленный мой, и вот кто друг мой, дщери Иерусалимские!
SONG|6|1|"Куда пошел возлюбленный твой, прекраснейшая из женщин? куда обратился возлюбленный твой? мы поищем его с тобою".
SONG|6|2|Мой возлюбленный пошел в сад свой, в цветники ароматные, чтобы пасти в садах и собирать лилии.
SONG|6|3|Я принадлежу возлюбленному моему, а возлюбленный мой – мне; он пасет между лилиями.
SONG|6|4|Прекрасна ты, возлюбленная моя, как Фирца, любезна, как Иерусалим, грозна, как полки со знаменами.
SONG|6|5|Уклони очи твои от меня, потому что они волнуют меня.
SONG|6|6|Волосы твои – как стадо коз, сходящих с Галаада; зубы твои – как стадо овец, выходящих из купальни, из которых у каждой пара ягнят, и бесплодной нет между ними;
SONG|6|7|как половинки гранатового яблока – ланиты твои под кудрями твоими.
SONG|6|8|Есть шестьдесят цариц и восемьдесят наложниц и девиц без числа,
SONG|6|9|но единственная – она, голубица моя, чистая моя; единственная она у матери своей, отличенная у родительницы своей. Увидели ее девицы, и – превознесли ее, царицы и наложницы, и – восхвалили ее.
SONG|6|10|Кто эта, блистающая, как заря, прекрасная, как луна, светлая, как солнце, грозная, как полки со знаменами?
SONG|6|11|Я сошла в ореховый сад посмотреть на зелень долины, поглядеть, распустилась ли виноградная лоза, расцвели ли гранатовые яблоки?
SONG|6|12|Не знаю, как душа моя влекла меня к колесницам знатных народа моего.
SONG|7|1|"Оглянись, оглянись, Суламита! оглянись, оглянись, – и мы посмотрим на тебя". Что вам смотреть на Суламиту, как на хоровод Манаимский?
SONG|7|2|О, как прекрасны ноги твои в сандалиях, дщерь именитая! Округление бедр твоих, как ожерелье, дело рук искусного художника;
SONG|7|3|живот твой – круглая чаша, [в которой] не истощается ароматное вино; чрево твое – ворох пшеницы, обставленный лилиями;
SONG|7|4|два сосца твои – как два козленка, двойни серны;
SONG|7|5|шея твоя – как столп из слоновой кости; глаза твои – озерки Есевонские, что у ворот Батраббима; нос твой – башня Ливанская, обращенная к Дамаску;
SONG|7|6|голова твоя на тебе, как Кармил, и волосы на голове твоей, как пурпур; царь увлечен [твоими] кудрями.
SONG|7|7|Как ты прекрасна, как привлекательна, возлюбленная, твоею миловидностью!
SONG|7|8|Этот стан твой похож на пальму, и груди твои на виноградные кисти.
SONG|7|9|Подумал я: влез бы я на пальму, ухватился бы за ветви ее; и груди твои были бы вместо кистей винограда, и запах от ноздрей твоих, как от яблоков;
SONG|7|10|уста твои – как отличное вино. Оно течет прямо к другу моему, услаждает уста утомленных.
SONG|7|11|Я принадлежу другу моему, и ко мне [обращено] желание его.
SONG|7|12|Приди, возлюбленный мой, выйдем в поле, побудем в селах;
SONG|7|13|поутру пойдем в виноградники, посмотрим, распустилась ли виноградная лоза, раскрылись ли почки, расцвели ли гранатовые яблоки; там я окажу ласки мои тебе.
SONG|7|14|Мандрагоры уже пустили благовоние, и у дверей наших всякие превосходные плоды, новые и старые: [это] сберегла я для тебя, мой возлюбленный!
SONG|8|1|О, если бы ты был мне брат, сосавший груди матери моей! тогда я, встретив тебя на улице, целовала бы тебя, и меня не осуждали бы.
SONG|8|2|Повела бы я тебя, привела бы тебя в дом матери моей. Ты учил бы меня, а я поила бы тебя ароматным вином, соком гранатовых яблоков моих.
SONG|8|3|Левая рука его у меня под головою, а правая обнимает меня.
SONG|8|4|Заклинаю вас, дщери Иерусалимские, – не будите и не тревожьте возлюбленной, доколе ей угодно.
SONG|8|5|Кто это восходит от пустыни, опираясь на своего возлюбленного? Под яблоней разбудила я тебя: там родила тебя мать твоя, там родила тебя родительница твоя.
SONG|8|6|Положи меня, как печать, на сердце твое, как перстень, на руку твою: ибо крепка, как смерть, любовь; люта, как преисподняя, ревность; стрелы ее – стрелы огненные; она пламень весьма сильный.
SONG|8|7|Большие воды не могут потушить любви, и реки не зальют ее. Если бы кто давал все богатство дома своего за любовь, то он был бы отвергнут с презреньем.
SONG|8|8|Есть у нас сестра, которая еще мала, и сосцов нет у нее; что нам будет делать с сестрою нашею, когда будут свататься за нее?
SONG|8|9|Если бы она была стена, то мы построили бы на ней палаты из серебра; если бы она была дверь, то мы обложили бы ее кедровыми досками.
SONG|8|10|Я – стена, и сосцы у меня, как башни; потому я буду в глазах его, как достигшая полноты.
SONG|8|11|Виноградник был у Соломона в Ваал–Гамоне; он отдал этот виноградник сторожам; каждый должен был доставлять за плоды его тысячу сребренников.
SONG|8|12|А мой виноградник у меня при себе. Тысяча пусть тебе, Соломон, а двести – стерегущим плоды его.
SONG|8|13|Жительница садов! товарищи внимают голосу твоему, дай и мне послушать его.
SONG|8|14|Беги, возлюбленный мой; будь подобен серне или молодому оленю на горах бальзамических!
