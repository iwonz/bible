RUTH|1|1|in diebus unius iudicis quando iudices praeerant facta est fames in terra abiitque homo de Bethleem Iuda ut peregrinaretur in regione moabitide cum uxore sua ac duobus liberis
RUTH|1|2|ipse vocabatur Helimelech uxor eius Noemi e duobus filiis alter Maalon et alter Chellion Ephrathei de Bethleem Iuda ingressique regionem moabitidem morabantur ibi
RUTH|1|3|et mortuus est Helimelech maritus Noemi remansitque ipsa cum filiis
RUTH|1|4|qui acceperunt uxores moabitidas quarum una vocabatur Orpha altera Ruth manseruntque ibi decem annis
RUTH|1|5|et ambo mortui sunt Maalon videlicet et Chellion remansitque mulier orbata duobus liberis ac marito
RUTH|1|6|et surrexit ut in patriam pergeret cum utraque nuru sua de regione moabitide audierat enim quod respexisset Dominus populum suum et dedisset eis escas
RUTH|1|7|egressa est itaque de loco peregrinationis suae cum utraque nuru et iam in via posita revertendi in terram Iuda
RUTH|1|8|dixit ad eas ite in domum matris vestrae faciat Dominus vobiscum misericordiam sicut fecistis cum mortuis et mecum
RUTH|1|9|det vobis invenire requiem in domibus virorum quos sortiturae estis et osculata est eas quae elevata voce flere coeperunt
RUTH|1|10|et dicere tecum pergemus ad populum tuum
RUTH|1|11|quibus illa respondit revertimini filiae mi cur venitis mecum num ultra habeo filios in utero meo ut viros ex me sperare possitis
RUTH|1|12|revertimini filiae mi abite iam enim senectute confecta sum nec apta vinculo coniugali etiam si possem hac nocte concipere et parere filios
RUTH|1|13|si eos expectare velitis donec crescant et annos impleant pubertatis ante eritis vetulae quam nubatis nolite quaeso filiae mi quia vestra angustia me magis premit et egressa est manus Domini contra me
RUTH|1|14|elevata igitur voce rursum flere coeperunt Orpha osculata socrum est ac reversa Ruth adhesit socrui suae
RUTH|1|15|cui dixit Noemi en reversa est cognata tua ad populum suum et ad deos suos vade cum ea
RUTH|1|16|quae respondit ne adverseris mihi ut relinquam te et abeam quocumque perrexeris pergam ubi morata fueris et ego pariter morabor populus tuus populus meus et Deus tuus Deus meus
RUTH|1|17|quae te morientem terra susceperit in ea moriar ibique locum accipiam sepulturae haec mihi faciat Deus et haec addat si non sola mors me et te separaverit
RUTH|1|18|videns ergo Noemi quod obstinato Ruth animo decrevisset secum pergere adversari noluit nec ultra ad suos reditum persuadere
RUTH|1|19|profectaeque sunt simul et venerunt in Bethleem quibus urbem ingressis velox apud cunctos fama percrebuit dicebantque mulieres haec est illa Noemi
RUTH|1|20|quibus ait ne vocetis me Noemi id est pulchram sed vocate me Mara hoc est amaram quia valde me amaritudine replevit Omnipotens
RUTH|1|21|egressa sum plena et vacuam reduxit me Dominus cur igitur vocatis me Noemi quam humiliavit Dominus et adflixit Omnipotens
RUTH|1|22|venit ergo Noemi cum Ruth Moabitide nuru sua de terra peregrinationis suae ac reversa est in Bethleem quando primum hordea metebantur
RUTH|2|1|erat autem vir Helimelech consanguineus homo potens et magnarum opum nomine Booz
RUTH|2|2|dixitque Ruth Moabitis ad socrum suam si iubes vadam in agrum et colligam spicas quae metentium fugerint manus ubicumque clementis in me patris familias repperero gratiam cui illa respondit vade filia mi
RUTH|2|3|abiit itaque et colligebat spicas post terga metentium accidit autem ut ager ille haberet dominum Booz qui erat de cognatione Helimelech
RUTH|2|4|et ecce ipse veniebat de Bethleem dixitque messoribus Dominus vobiscum qui responderunt ei benedicat tibi Dominus
RUTH|2|5|dixitque Booz iuveni qui messoribus praeerat cuius est haec puella
RUTH|2|6|qui respondit haec est Moabitis quae venit cum Noemi de regione moabitide
RUTH|2|7|et rogavit ut spicas colligeret remanentes sequens messorum vestigia et de mane usque nunc stat in agro et ne ad momentum quidem domum reversa est
RUTH|2|8|et ait Booz ad Ruth audi filia ne vadas ad colligendum in alterum agrum nec recedas ab hoc loco sed iungere puellis meis
RUTH|2|9|et ubi messuerint sequere mandavi enim pueris meis ut nemo tibi molestus sit sed etiam si sitieris vade ad sarcinulas et bibe aquas de quibus et pueri bibunt
RUTH|2|10|quae cadens in faciem suam et adorans super terram dixit ad eum unde mihi hoc ut invenirem gratiam ante oculos tuos et nosse me dignareris peregrinam mulierem
RUTH|2|11|cui ille respondit nuntiata sunt mihi omnia quae feceris socrui tuae post mortem viri tui et quod dereliqueris parentes tuos et terram in qua nata es et veneris ad populum quem ante nesciebas
RUTH|2|12|reddat tibi Dominus pro opere tuo et plenam mercedem recipias a Domino Deo Israhel ad quem venisti et sub cuius confugisti alas
RUTH|2|13|quae ait inveni gratiam ante oculos tuos domine mi qui consolatus es me et locutus es ad cor ancillae tuae quae non sum similis unius puellarum tuarum
RUTH|2|14|dixitque ad eam Booz quando hora vescendi fuerit veni huc et comede panem et intingue buccellam tuam in aceto sedit itaque ad messorum latus et congessit pulentam sibi comeditque et saturata est et tulit reliquias
RUTH|2|15|atque inde surrexit ut spicas ex more colligeret praecepit autem Booz pueris suis dicens etiam si vobiscum metere voluerit ne prohibeatis eam
RUTH|2|16|et de vestris quoque manipulis proicite de industria et remanere permittite ut absque rubore colligat et colligentem nemo corripiat
RUTH|2|17|collegit ergo in agro usque ad vesperam et quae collegerat virga caedens et excutiens invenit hordei quasi oephi mensuram id est tres modios
RUTH|2|18|quos portans reversa est in civitatem et ostendit socrui suae insuper protulit et dedit ei de reliquiis cibi sui quo saturata fuerat
RUTH|2|19|dixitque ei socrus ubi hodie collegisti et ubi fecisti opus sit benedictus qui misertus est tui indicavitque ei apud quem esset operata et nomen dixit viri quod Booz vocaretur
RUTH|2|20|cui respondit Noemi benedictus sit a Domino quoniam eandem gratiam quam praebuerat vivis servavit et mortuis rursumque propinquus ait noster est homo
RUTH|2|21|et Ruth hoc quoque inquit praecepit mihi ut tamdiu messoribus eius iungerer donec omnes segetes meterentur
RUTH|2|22|cui dixit socrus melius est filia mi ut cum puellis eius exeas ad metendum ne in alieno agro quispiam resistat tibi
RUTH|2|23|iuncta est itaque puellis Booz et tamdiu cum eis messuit donec hordea et triticum in horreis conderentur
RUTH|3|1|postquam autem reversa est ad socrum suam audivit ab ea filia mi quaeram tibi requiem et providebo ut bene sit tibi
RUTH|3|2|Booz iste cuius puellis in agro iuncta es propinquus est noster et hac nocte aream hordei ventilat
RUTH|3|3|lava igitur et unguere et induere cultioribus vestimentis ac descende in aream non te videat homo donec esum potumque finierit
RUTH|3|4|quando autem ierit ad dormiendum nota locum in quo dormiat veniesque et discoperies pallium quo operitur a parte pedum et proicies te et ibi iacebis ipse autem dicet tibi quid agere debeas
RUTH|3|5|quae respondit quicquid praeceperis faciam
RUTH|3|6|descenditque in aream et fecit omnia quae sibi imperaverat socrus
RUTH|3|7|cumque comedisset Booz et bibisset et factus esset hilarior issetque ad dormiendum iuxta acervum manipulorum venit abscondite et discoperto a pedibus eius pallio se proiecit
RUTH|3|8|et ecce nocte iam media expavit homo et conturbatus est viditque mulierem iacentem ad pedes suos
RUTH|3|9|et ait illi quae es illaque respondit ego sum Ruth ancilla tua expande pallium tuum super famulam tuam quia propinquus es
RUTH|3|10|et ille benedicta inquit es Domino filia et priorem misericordiam posteriore superasti quia non es secuta iuvenes pauperes sive divites
RUTH|3|11|noli ergo metuere sed quicquid dixeris mihi faciam tibi scit enim omnis populus qui habitat intra portas urbis meae mulierem te esse virtutis
RUTH|3|12|nec abnuo me propinquum sed est alius me propinquior
RUTH|3|13|quiesce hac nocte et facto mane si te voluerit propinquitatis iure retinere bene res acta est sin autem ille noluerit ego te absque ulla dubitatione suscipiam vivit Dominus dormi usque mane
RUTH|3|14|dormivit itaque ad pedes eius usque ad noctis abscessum surrexitque antequam homines se cognoscerent mutuo et dixit Booz cave ne quis noverit quod huc veneris
RUTH|3|15|et rursum expande inquit palliolum tuum quo operiris et tene utraque manu qua extendente et tenente mensus est sex modios hordei et posuit super eam quae portans ingressa est civitatem
RUTH|3|16|et venit ad socrum suam quae dixit ei quid egisti filia narravitque ei omnia quae sibi fecisset homo
RUTH|3|17|et ait ecce sex modios hordei dedit mihi et ait nolo vacuam te reverti ad socrum tuam
RUTH|3|18|dixitque Noemi expecta filia donec videamus quem res exitum habeat neque enim cessabit homo nisi conpleverit quod locutus est
RUTH|4|1|ascendit ergo Booz ad portam et sedit ibi cumque vidisset propinquum praeterire de quo prius sermo habitus est dixit ad eum declina paulisper et sede hic vocans eum nomine suo qui devertit et sedit
RUTH|4|2|tollens autem Booz decem viros de senioribus civitatis dixit ad eos sedete hic
RUTH|4|3|quibus residentibus locutus est ad propinquum partem agri fratris nostri Helimelech vendit Noemi quae reversa est de regione moabitide
RUTH|4|4|quod audire te volui et tibi dicere coram cunctis sedentibus et maioribus natu de populo meo si vis possidere iure propinquitatis eme et posside sin autem tibi displicet hoc ipsum indica mihi ut sciam quid facere debeam nullus est enim propinquus excepto te qui prior es et me qui secundus sum at ille respondit ego agrum emam
RUTH|4|5|cui dixit Booz quando emeris agrum de manu mulieris Ruth quoque Moabitidem quae uxor defuncti fuit debes accipere ut suscites nomen propinqui tui in hereditate sua
RUTH|4|6|qui respondit cedo iure propinquitatis neque enim posteritatem familiae meae delere debeo tu meo utere privilegio quo me libenter carere profiteor
RUTH|4|7|hic autem erat mos antiquitus in Israhel inter propinquos et si quando alter alteri suo iure cedebat ut esset firma concessio solvebat homo calciamentum suum et dabat proximo suo hoc erat testimonium cessionis in Israhel
RUTH|4|8|dixit ergo propinquus Booz tolle calciamentum quod statim solvit de pede suo
RUTH|4|9|at ille maioribus natu et universo populo testes inquit vos estis hodie quod possederim omnia quae fuerunt Helimelech et Chellion et Maalon tradente Noemi
RUTH|4|10|et Ruth Moabitidem uxorem Maalon in coniugium sumpserim ut suscitem nomen defuncti in hereditate sua ne vocabulum eius de familia sua ac fratribus et populo deleatur vos inquam huius rei testes estis
RUTH|4|11|respondit omnis populus qui erat in porta et maiores natu nos testes sumus faciat Dominus hanc mulierem quae ingreditur domum tuam sicut Rachel et Liam quae aedificaverunt domum Israhel ut sit exemplum virtutis in Ephrata et habeat celebre nomen in Bethleem
RUTH|4|12|fiatque domus tua sicut domus Phares quem Thamar peperit Iudae de semine quod dederit Dominus tibi ex hac puella
RUTH|4|13|tulit itaque Booz Ruth et accepit uxorem ingressusque est ad eam et dedit illi Dominus ut conciperet et pareret filium
RUTH|4|14|dixeruntque mulieres ad Noemi benedictus Dominus qui non est passus ut deficeret successor familiae tuae et vocaretur nomen eius in Israhel
RUTH|4|15|et habeas qui consoletur animam tuam et enutriat senectutem de nuru enim tua natus est quae te diligit et multo tibi est melior quam si septem haberes filios
RUTH|4|16|susceptumque Noemi puerum posuit in sinu suo et nutricis ac gerulae officio fungebatur
RUTH|4|17|vicinae autem mulieres congratulantes ei et dicentes natus est filius Noemi vocaverunt nomen eius Obed hic est pater Isai patris David
RUTH|4|18|hae sunt generationes Phares Phares genuit Esrom
RUTH|4|19|Esrom genuit Aram Aram genuit Aminadab
RUTH|4|20|Aminadab genuit Naasson Naasson genuit Salma
RUTH|4|21|Salma genuit Booz Booz genuit Obed
