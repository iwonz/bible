LEV|1|1|І кликнув Господь до Мойсея, і промовляв до нього з скинії заповіту, говорячи:
LEV|1|2|Промовляй до Ізраїлевих синів та й скажеш до них: Коли хто з вас принесе жертву для Господа зо скотини, то з худоби великої й худоби дрібної принесете вашу жертву.
LEV|1|3|Якщо жертва його цілопалення з худоби великої, то нехай принесе його, самця безвадного; нехай приведе його до скинії заповіту, щоб він був уподобаний перед лицем Господнім.
LEV|1|4|І покладе він руку свою на голову цілопалення, і буде йому дано вподобання на очищення від гріхів його.
LEV|1|5|І заріже він ягня перед Господнім лицем. А Ааронові сини, священики, принесуть кров, і покроплять тією кров'ю на жертівника навколо, що при вході до скинії заповіту.
LEV|1|6|І здере він шкуру з жертви цілопалення, і розітне його на куски його.
LEV|1|7|І дадуть сини священика Аарона огню на жертівника, і покладуть дров на тім огні.
LEV|1|8|І порозкладають Ааронові сини, священики, ті куски, голову та товщ, на дровах, що на огні, який на жертівнику.
LEV|1|9|А його нутрощі та голінки його обмиє водою. І священик усе те спалить на жертівнику, це цілопалення, огняна жертва, пахощі любі для Господа.
LEV|1|10|А якщо його жертва з дрібної худобини, з овець або з кіз на цілопалення, то нехай приведе його, безвадного самця,
LEV|1|11|і заріже його на боці жертівника на північ, перед Господнім лицем. І покроплять сини Ааронові, священики, кров'ю його на жертівника навколо.
LEV|1|12|І розітне його на куски його, голову його, і товщ його, а священик порозкладає їх на дровах, що на огні, який на жертівнику.
LEV|1|13|А нутрощі та голінки обмиє водою. І священик принесе все це, та й спалить на жертівнику, це цілопалення, огняна жертва, пахощі любі для Господа.
LEV|1|14|А якщо цілопалення його жертва для Господа з птаства, то нехай з горлиць або з голубенят принесе жертву свою.
LEV|1|15|І принесе її священик до жертівника, і проб'є йому нігтем великим голову, та й спалить на жертівнику, а кров його буде вилита при стіні жертівника.
LEV|1|16|І здійме його воло в пір'ї його, і кине його при жертівнику на схід на місце попелу.
LEV|1|17|І роздере його між крильми його, але не відділить їх. А священик спалить його на жертівнику на дровах, що на огні, воно цілопалення, огняна жертва, пахощі любі для Господа.
LEV|2|1|А коли хто принесе жертву, жертву хлібну для Господа, то нехай пшенична мука буде жертва його, а він поллє на неї оливи, і дасть на неї ладану.
LEV|2|2|І принесе її до Ааронових синів, священиків, і візьме звідти повну свою жменю пшеничної муки її, і оливи її зо всім її ладаном, та й спалить священик на жертівнику за пригадувальну частину, це огняна жертва, пахощі любі для Господа.
LEV|2|3|А позостале з цієї хлібної жертви для Аарона та для синів його, це Найсвятіше з Господніх жертов!
LEV|2|4|А коли принесеш жертву, жертву хлібну випеченого в печі, то нехай це буде пшенична мука, прісні калачі, мішані в оливі, та прісні коржики, помазані оливою.
LEV|2|5|А якщо твоя жертва жертва хлібна на лопатці, то нехай це буде пшенична мука, мішана в оливі, прісна.
LEV|2|6|Поламати її на шматочки, і поллєш на неї оливи, це хлібна жертва.
LEV|2|7|А якщо твоя жертва жертва хлібна смаження, то нехай буде зроблена в оливі з пшеничної муки.
LEV|2|8|І принесеш хлібну жертву, що зроблена з тих речей, для Господа, і подаси її до священика, а він принесе її до жертівника.
LEV|2|9|І принесе священик із хлібної жертви за пригадувальну частину її, та й спалить на жертівнику, це огняна жертва, любі пахощі для Господа.
LEV|2|10|А позостале з цієї хлібної жертви для Аарона та для синів його: це Найсвятіше з Господніх жертов!
LEV|2|11|Кожна хлібна жертва, яку принесете Господеві, не буде зроблена квашена, бо все квашене й усякий мед не спалите з нього огняної жертви для Господа.
LEV|2|12|Як жертву первоплоду принесіть її для Господа, а на жертівника вона не приноситься на любі пахощі.
LEV|2|13|І кожну жертву, жертву хлібну, посолиш сіллю. І хлібної жертви твоєї не позбавиш соли заповіту Бога твого, на кожній жертві твоїй принесеш соли.
LEV|2|14|А якщо принесеш хлібну жертву первоплодів для Господа, то колосся, пряжене в огні, як потовчене зерно принесеш хлібну жертву своїх первоплодів.
LEV|2|15|І полий на неї оливи, і поклади на неї ладану, це жертва хлібна.
LEV|2|16|І спалить священик за пригадувальну частину її з потовченого зерна, із оливи її на всім ладані її, це огняна жертва для Господа.
LEV|3|1|А якщо його жертва мирна, якщо з великої худоби він приносить чи самця, чи самицю, він принесе її безвадну перед Господнє лице,
LEV|3|2|і покладе свою руку на голову жертви своєї, та й заріже її при вході до скинії заповіту. А Ааронові сини, священики, покроплять тією кров'ю на жертівника навколо.
LEV|3|3|І принесе він із мирної жертви огняну жертву для Господа, лій, що закриває нутрощі, та ввесь лій, що на нутрощах,
LEV|3|4|і обидві нирки, і лій, що на них, що на стегнах, а сальника на печінці здійме його з нирками.
LEV|3|5|І спалять те сини Ааронові на жертівнику на цілопалення, що на дровах, яке на огні, це огняна жертва, пахощі любі для Господа.
LEV|3|6|А якщо з дрібної худоби його жертва на мирну жертву для Господа, самець чи самиця, то безвадну принесе її.
LEV|3|7|Якщо приносить він на жертву вівцю, то принесе її перед Господнє лице,
LEV|3|8|і покладе свою руку на голову жертви своєї, та й заріже її перед скинією заповіту. А Ааронові сини покроплять кров'ю її на жертівника навколо.
LEV|3|9|І він принесе з мирної жертви огняну жертву для Господа, цілого курдюка, якого здійме при хребті, і лій, що закриває нутрощі, і ввесь лій, що на нутрощах,
LEV|3|10|і обидві нирки та лій, що на них, що на стегнах, а сальника на печінці здійме його з нирками.
LEV|3|11|І священик спалить те на жертівнику, хліб огняної жертви для Господа.
LEV|3|12|А якщо жертва його коза, то піднесе її перед лице Господнє,
LEV|3|13|і покладе свою руку на голову її, та й заріже її перед скинією заповіту. А Ааронові сини покроплять кров'ю її на жертівника навколо.
LEV|3|14|І він принесе з неї жертву свою, жертву для Господа, лій, що закриває нутрощі, та ввесь лій, що на нутрощах,
LEV|3|15|і обидві нирки, і лій, що на них, що на стегнах, а сальника на печінці здійме його з нирками.
LEV|3|16|І священик спалить їх на жертівнику, це пожива, огняна жертва на любі пахощі; увесь лій для Господа.
LEV|3|17|Оце постанова вічна для ваших родів у всіх осадах ваших: жодного лою й жодної крови не будете їсти.
LEV|4|1|І Господь промовляв до Мойсея, говорячи:
LEV|4|2|Промовляй до Ізраїлевих синів, говорячи: Коли хто невмисне згрішить проти якої зо всіх заповідей Господніх, чого не треба чинити, а він учинить проти однієї з них,
LEV|4|3|якщо помазаний священик згрішить на провину народу, то він принесе за гріх свій, що згрішив ним, бичка, молоде з худоби великої, безвадного для Господа на жертву за гріх.
LEV|4|4|І приведе він того бичка до входу скинії заповіту перед Господнє лице, і покладе свою руку на голову того бичка, та й заріже бичка перед Господнім лицем.
LEV|4|5|А помазаний священик візьме крови того бичка, та й внесе її до скинії заповіту.
LEV|4|6|І вмочить священик пальця свого в ту кров, та й покропить тією кров'ю сім раз перед Господнім лицем перед завіси святині.
LEV|4|7|І дасть священик з тієї крови на роги жертівника кадила пахощів, перед Господнім лицем, що він у скинії заповіту, а всю кров бичка виллє до підстави жертівника цілопалення, що при вході скинії заповіту.
LEV|4|8|А ввесь лій бичка жертви за гріх принесе з нього лій, що закриває нутрощі, і ввесь лій, що на нутрощах,
LEV|4|9|і обидві нирки та лій, що на них, що на стегнах, а сальника на печінці здійме його з нирками,
LEV|4|10|як приноситься з вола мирної жертви, і священик спалить те на жертівнику цілопалення.
LEV|4|11|А шкуру бичка та все м'ясо його з головою його та голінками його, і нутрощі його, і нечистість їх,
LEV|4|12|і всього бичка винесе поза табір до чистого місця, до місця висипання попелу, і спалить його на дровах в огні, на висипанні попелу буде спалений він.
LEV|4|13|А коли вся Ізраїлева громада помилково згрішить, і діло буде затаєне з очей зборів, і зроблять що проти якої зо всіх Господніх заповідей, чого не можна робити, і завинять,
LEV|4|14|а гріх буде пізнаний, що вони згрішили ним, то збори принесуть бичка, молоде з худоби великої, на жертву за гріх. І вони приведуть його перед скинію заповіту.
LEV|4|15|А старші громади покладуть свої руки на голову бичка перед Господнім лицем, та й заріже один з них бичка перед лицем Господнім.
LEV|4|16|А помазаний священик внесе крови бичка до скинії заповіту.
LEV|4|17|І вмочить священик пальця свого в ту кров, та й покропить сім раз перед Господнім лицем перед завіси.
LEV|4|18|І дасть він із тієї крови на роги жертівника, що перед Господнім лицем, що він у скинії заповіту, а всю ту кров виллє до підстави жертівника цілопалення, що при вході скинії заповіту.
LEV|4|19|А ввесь його лій принесе з нього та й спалить на жертівнику.
LEV|4|20|І зробить з тим бичком те саме, що робив бичкові жертви за гріх, так само зробить із ним. І так священик дасть очищення за них, і буде прощено їм.
LEV|4|21|І винесе бичка поза табір, та й спалить його, як палив бичка першого, він жертва за гріх зборів.
LEV|4|22|Коли згрішить начальник, і зробить що невмисне проти якої зо всіх заповідей Господа, Бога його, чого робити не можна, та й завинить,
LEV|4|23|і буде пізнаний ним гріх його, що згрішив ним, то приведе він жертву свою безвадного козла,
LEV|4|24|і покладе свою руку на голову того козла, та й заріже його в місці, де ріжеться цілопалення перед Господнім лицем, він жертва за гріх.
LEV|4|25|А священик візьме з крови жертви за гріх своїм пальцем, та й дасть на роги жертівника цілопалення, а кров його виллє до підстави жертівника цілопалення.
LEV|4|26|А ввесь лій його спалить на жертівнику, як лій мирної жертви, та й так очистить священик його з гріха його, і буде прощений йому.
LEV|4|27|А коли яка душа з народу землі невмисне згрішить, коли зробить що проти якої з заповідей Господніх, чого робити не можна, та й завинить,
LEV|4|28|і буде пізнаний ним гріх його, що згрішив, то він приведе жертву свою безвадну козу, самицю, за гріх свій, що він згрішив був,
LEV|4|29|і покладе свою руку на голову жертви за гріх, та й заріже цю жертву за гріх у місці цілопалення.
LEV|4|30|А священик візьме своїм пальцем із крови її, та й дасть на роги жертівника цілопалення, а всю її кров виллє до підстави жертівника.
LEV|4|31|А ввесь її лій він здійме, як знятий був лій із мирної жертви, і священик спалить на жертівнику на пахощі любі для Господа. І так священик очистить його, і буде прощено йому.
LEV|4|32|А якщо він приведе вівцю в жертву свою за гріх, то приведе безвадну самицю,
LEV|4|33|і покладе свою руку на голову жертви за гріх, та й заріже її на жертву за гріх у місці, де ріже він жертву цілопалення.
LEV|4|34|І візьме священик із крови жертви за гріх своїм пальцем, та й дасть на роги жертівника цілопалення, а всю кров її виллє до підстави жертівника.
LEV|4|35|А ввесь лій її здійме, як здіймається лій вівці з мирної жертви, та й спалить священик його на жертівнику на огняні жертви Господні. І так очистить його священик за гріх його, що згрішив був, і буде прощено йому.
LEV|5|1|А коли хто згрішить: почує голос прокляття, і був свідком, або бачив, або знав, але не виявив, то понесе свою провину;
LEV|5|2|або особа, що доторкнеться якої нечистої речі, або падла звірини нечистої, або падла худоби нечистої, або падла нечистого плазуючого, і буде це незнане їй, то вона нечиста й завинить;
LEV|5|3|або коли доторкнеться нечистости людини, всякої нечистости її, що нею стане нечиста, і буде це незнане їй, а вона довідається, то завинить;
LEV|5|4|або коли хто присягне, вимовляючи нерозважно устами своїми, чинити зло або чинити добро, на все, що нерозважно вимовляє людина в присязі, і буде це незнане йому, а він довідається, що завинив одним із цих,
LEV|5|5|то станеться, що завинить одним із цих, і визнає, чим він згрішив у тому.
LEV|5|6|І приведе він Господеві жертву за провину, за гріх свій, що згрішив, самицю з дрібної худоби, вівцю або козу на жертву за гріх, а священик очистить його від гріха його.
LEV|5|7|А якщо рука його не спроможна на ягня, то принесе в жертву за провину свою, що згрішив він, дві горлиці або двоє голубенят Господеві, одне на жертву за гріх, а одне на цілопалення.
LEV|5|8|І принесе їх до священика, а він перше принесе те, що на жертву за гріх, і натне великим нігтем голову його від шиї її, але не відділить.
LEV|5|9|І покропить із крови жертви за гріх на стіну жертівника, а позостала кров буде вилита до підстави жертівника, це жертва за гріх.
LEV|5|10|А другого зробить цілопаленням за уставом. І очистить його священик від гріха його, що згрішив той, і буде прощено йому.
LEV|5|11|А якщо він не спроможний на дві горлиці або на двоє голубенят, то принесе в жертву свою за те, чим згрішив, десяту частину ефи пшеничної муки на жертву за гріх, не докладе до неї оливи й не дасть на неї ладану, бо вона жертва за гріх.
LEV|5|12|І принесе її до священика, а священик візьме з неї повну свою жменю, за пригадувальну частину її, та й спалить на жертівнику на огняні жертви Господеві, вона жертва за гріх.
LEV|5|13|І очистить його священик від гріха його, що згрішив він одним із них, і буде йому прощений; і буде вона для священика, як жертва хлібна.
LEV|5|14|І Господь промовляв до Мойсея, говорячи:
LEV|5|15|Коли хто переступом спроневіриться, і невмисне згрішить проти Господніх святощів, то він приведе жертву за провину свою до Господа, безвадного барана з дрібної худоби, за твоєю оцінкою срібла шеклів, на міру шеклем святині на жертву за провину.
LEV|5|16|А те, що згрішив проти святощів, поверне, і додасть до нього п'яту частину його священикові, а священик очистить його бараном жертви за гріх, і буде прощено йому.
LEV|5|17|А якщо згрішить коли хто, і зробить що проти якої зо всіх Господніх заповідей, чого не можна робити, і не знатиме, і завинить, і понесе свій гріх,
LEV|5|18|то він приведе до священика безвадного барана з дрібної худоби в оцінці твоїй на жертву за провину. І очистить його священик за помилку його, що нею помилився, бо він не знав, і буде прощена йому.
LEV|5|19|Це жертва за провину: він справді завинив Господеві.
LEV|6|1|(5-20) І Господь промовляв до Мойсея, говорячи:
LEV|6|2|(5-21) Коли хто згрішить і переступом спроневіриться проти Господа, і скаже неправду на ближнього свого щодо даного на сховок, щодо даного в заклад, або щодо грабунку, або вимусить утиском у ближнього свого,
LEV|6|3|(5-22) або знайде якусь згубу та й скаже неправду про неї, і присягне неправдиво на одне зо всього, що робить людина, і згрішить тим,
LEV|6|4|(5-23) то станеться, коли він згрішить і завинить, нехай поверне грабунок, що заграбував, або вимушення, що був вимусив, або дане на сховок, що було зложене в нього, або згубу, що знайшов,
LEV|6|5|(5-24) або все, що присяг про нього неправдиво, і поверне його насамперед, і додасть до нього п'яту частину тому, чиє воно, дасть його в день, коли виявиться провина його.
LEV|6|6|(5-25) І він приведе Господеві до священика жертву за провину свою, безвадного барана з дрібної худоби за твоєю оцінкою на жертву за провину.
LEV|6|7|(5-26) І священик очистить його перед Господнім лицем, і буде йому прощено все до одного, що він зробив на провину.
LEV|6|8|(6-1) І Господь промовляв до Мойсея, кажучи:
LEV|6|9|(6-2) Накажи Ааронові та синам його, повідаючи: Оце закон цілопалення: Воно приноситься на огнищі своїм на жертівнику цілу ніч аж до ранку, а огонь жертівника горітиме на ньому.
LEV|6|10|(6-3) І надіне священик льняну свою шату, і льняне спіднє зодягне на тіло своє, і збере попіл, що на нього огонь спалить цілопалення на жертівнику, та й покладе його при жертівнику.
LEV|6|11|(6-4) І здійме він шати свої, і зодягне одіж іншу, та й винесе попіл поза табір до чистого місця.
LEV|6|12|(6-5) А огонь на жертівнику горітиме на ньому, не погасне, а священик палитиме на ньому дрова щоранку, і кластиме на нього цілопалення, і палитиме на ньому лій мирних жертов.
LEV|6|13|(6-6) Огонь завжди горітиме на жертівнику, не погасне.
LEV|6|14|(6-7) А оце закон про хлібну жертву: Ааронові сини принесуть її перед лице Господнє до переду жертівника.
LEV|6|15|(6-8) І візьме він із неї жменею своєю з пшеничної муки хлібної жертви, та з оливи її, та ввесь ладан, що на хлібній жертві, та й спалить на жертівнику, любі пахощі, це частина її, як пригадувальна для Господа.
LEV|6|16|(6-9) А позостале з неї їстимуть Аарон та сини його, прісне буде їджене воно в святім місці, на подвір'ї скинії заповіту будуть їсти її.
LEV|6|17|(6-10) Не буде печена вона квашеною. Їхню частину Я дав це з огняних Моїх жертов; вона Найсвятіше, як жертва за гріх та жертва за провину.
LEV|6|18|(6-11) Кожен нащадок чоловічої статі поміж Ааронових дітей буде її їсти, вічна постанова для ваших поколінь, з огняних жертов Господніх. Усе, що доторкнеться до них, освятиться.
LEV|6|19|(6-12) І Господь промовляв до Мойсея, говорячи:
LEV|6|20|(6-13) Оце жертва Аарона та синів його, що принесуть Господеві в дні помазання його: десята частина ефи пшеничної муки, це постійна хлібна жертва: половина її рано, а половина її ввечорі.
LEV|6|21|(6-14) На лопатці в оливі буде вона зроблена; принесеш її вимішану, випечену жертву хлібну в кусках принесеш, любі пахощі для Господа.
LEV|6|22|(6-15) А помазаний священик зробить її замість нього зробить її котрийсь із синів його, це вічна Господня постанова. Уся вона буде спалена.
LEV|6|23|(6-16) А кожна священикова хлібна жертва буде ціла, не буде їджена.
LEV|6|24|(6-17) І Господь промовляв до Мойсея, говорячи:
LEV|6|25|(6-18) Промовляй до Аарона та до синів його, говорячи: Оце закон про жертву за гріх: На місці, де зарізується цілопалення, буде зарізувана жертва за гріх перед лицем Господнім, Найсвятіше вона!
LEV|6|26|(6-19) Священик, що складає її як жертву за гріх, буде їсти її, на місці святому буде вона їджена, на подвір'ї скинії заповіту.
LEV|6|27|(6-20) Усе, що доторкнеться до м'яса її, стане святе; а що з її крови покропить на одежу, що покропиться нею, те випереш на місці святому.
LEV|6|28|(6-21) А глиняний посуд, що в ньому вона варена, буде розбитий. А якщо в мідянім посуді була вона варена, то буде вичищений до блиску й виполосканий водою.
LEV|6|29|(6-22) Кожен чоловічої статі із священиків буде їсти її, Найсвятіше вона.
LEV|6|30|(6-23) А кожна жертва за гріх, що з крови її буде внесено до скинії заповіту на окуплення в святині, не буде їджена, в огні буде спалена.
LEV|7|1|А оце закон жертви за провину, Найсвятіше вона.
LEV|7|2|На місці, де ріжуть цілопалення, заріжуть жертву за провину, а кров її священик покропить на жертівника навколо.
LEV|7|3|А ввесь її лій із неї він принесе, курдюка, і лій, що покриває нутрощі,
LEV|7|4|і обидві нирки, і лій, що на них, що на стегнах, а сальника на печінці здійме з нирками,
LEV|7|5|та й спалить те священик на жертівнику, це огняна жертва для Господа, жертва за провину вона.
LEV|7|6|Кожен чоловічої статі серед священиків буде їсти її, на місці святому буде вона їджена, Найсвятіше вона.
LEV|7|7|Як про жертву за гріх, так само про жертву за провини закон їм один: священикові, що очистить нею, йому вона буде.
LEV|7|8|А священик, що приносить чиєсь цілопалення, шкура цілопалення, яке приніс він, священикові, йому вона буде.
LEV|7|9|І кожна жертва хлібна, що в печі буде печена, і кожна приготовлена в горшку та на лопатці, священикові, що приносить її, йому вона буде.
LEV|7|10|А кожна хлібна жертва, мішана в оливі й суха, буде вона всім синам Аароновим, як одному, так і другому.
LEV|7|11|А оце закон про мирну жертву, що хтось принесе її Господеві.
LEV|7|12|Якщо принесе її на подяку, то він принесе на жертву подяки прісні калачі, мішані в оливі, і прісні коржі, помазані оливою, і вимішана пшенична мука, калачі, мішані в оливі.
LEV|7|13|Разом із калачами квашеного хліба принесе він жертву свою, при мирній жертві подяки його.
LEV|7|14|І принесе він щось одне з кожної жертви, приношення для Господа; це буде священикові, що кропить кров мирної жертви, буде йому.
LEV|7|15|А м'ясо мирної жертви подяки його буде їджене в дні його жертви, не позоставить із нього нічого до ранку.
LEV|7|16|А якщо жертва його приношення обітниця, або добровільний дар, то вона буде їджена в день принесення ним його жертви, а позостале з неї й назавтра буде їджене.
LEV|7|17|А позостале з м'яса кривавої жертви в третім дні буде спалене.
LEV|7|18|А якщо справді буде їджене з м'яса мирної жертви його в третім дні, то не буде вподобаний той, хто приносить її, це не буде залічене йому, буде нечисть; а хто їстиме з неї, понесе свій гріх.
LEV|7|19|А те м'ясо, що доторкнеться до чогось нечистого, не буде їджене, на огні буде спалене. А м'ясо чисте кожен чистий буде їсти м'ясо.
LEV|7|20|А душа, що буде їсти м'ясо з мирної жертви, що вона Господня, а нечисть його на ньому, то буде вона винищена з народу свого.
LEV|7|21|А коли хто доторкнеться до чогось нечистого, до нечистоти людської, або до нечистої худоби, або до всього нечистого плазуючого, та проте буде їсти з м'яса мирної жертви, що Господня вона, то буде той винищений із народу свого.
LEV|7|22|І Господь промовляв до Мойсея, говорячи:
LEV|7|23|Кажи до Ізраїлевих синів, говорячи: жодного лою волового, ані овечого, ані козиного не будете їсти.
LEV|7|24|А лій із падла й лій пошматованого буде вживаний для всякої потреби, але їсти не будете їсти його.
LEV|7|25|Бо кожен, хто їсть лій із худоби, що з неї приносить огняну жертву для Господа, то душа та, що їсть, буде винищена з народу свого.
LEV|7|26|І жодної крови птаства та худоби не будете їсти по всіх ваших оселях.
LEV|7|27|Кожна душа, що їстиме якубудь кров, то буде винищена душа та з-посеред народу свого.
LEV|7|28|І Господь промовляв до Мойсея, говорячи:
LEV|7|29|Промовляй до Ізраїлевих синів, говорячи: Хто приносить свою мирну жертву до Господа, той принесе своє приношення Господеві з своєї мирної жертви.
LEV|7|30|Руки його принесуть огняні жертви Господні, лій із грудиною, принесе грудину, щоб колихати її, як колихання перед Господнім лицем.
LEV|7|31|І священик спалить той лій на жертівнику. А та грудина буде Ааронові та синам його.
LEV|7|32|А праве стегно з мирних жертов ваших дасте священикові, як приношення.
LEV|7|33|Хто з Ааронових синів приносить кров мирних жертов та лій, йому буде на пайку праве стегно.
LEV|7|34|Бо Я взяв від Ізраїлевих синів грудину колихання й стегно приношення з мирних жертов їхніх, та й дав їх священикові Ааронові й синам його на вічну постанову від Ізраїлевих синів.
LEV|7|35|Оце частка з помазання Аарона та частка з помазання синів його з огняних жертов Господніх у день приношення їх на священнослуження Господеві,
LEV|7|36|що наказав Господь давати їм у день їхнього помазання від Ізраїлевих синів, вічна постанова на їхні покоління!
LEV|7|37|Оце закон про цілопалення, про хлібну жертву, і про жертву за гріх, і про жертву за провину, і про посвячення, та про жертву мирну,
LEV|7|38|що Господь наказав був Мойсеєві на Сінайській горі в день наказу Його Ізраїлевим синам приносити жертви свої Господеві в Сінайській пустині.
LEV|8|1|І Господь промовляв до Мойсея, говорячи:
LEV|8|2|Візьми Аарона та синів його з ним, і шати, і оливу помазання, і бичка жертви за гріх, і два барани, і коша з опрісноками.
LEV|8|3|І збери всю громаду до входу скинії заповіту.
LEV|8|4|І зробив Мойсей, як Господь наказав був йому. І зібралась громада до входу скинії заповіту.
LEV|8|5|І промовив Мойсей до громади: Оце та річ, що Господь наказав зробити.
LEV|8|6|І привів Мойсей Аарона й синів його, та й умив їх водою.
LEV|8|7|І дав він на нього хітона, й оперезав його поясом, і зодягнув його шатою, і дав на нього ефода, і оперезав його поясом ефоду, і прикріпив ним ефода на ньому.
LEV|8|8|І поклав на нього нагрудника, і дав до нагрудника урім та туммім.
LEV|8|9|І поклав завоя на голову його, і поклав на завоя спереду його золоту квітку, вінця святости, як Господь наказав був Мойсеєві.
LEV|8|10|І взяв Мойсей оливу помазання, і намастив скинію, і все, що в ній, та й освятив їх.
LEV|8|11|І покропив він із неї сім раз на жертівника, і намастив жертівника та ввесь посуд його, і вмивальницю та підставу її, щоб їх освятити.
LEV|8|12|І вилив з оливи помазання на Ааронову голову, та й помазав його, щоб його посвятити.
LEV|8|13|І привів Мойсей Ааронових синів, і зодягнув їх у хітони, й оперезав їх поясом, і поклав на них накриття голови, як Господь наказав був Мойсеєві.
LEV|8|14|І підвів він бичка жертви за гріх, і поклав Аарон та сини його свої руки на голову того бичка жертви за гріх.
LEV|8|15|І зарізав, і взяв Мойсей крови і дав своїм пальцем на роги навколо жертівника, і очистив жертівника. А кров вилив до підстави жертівника, і освятив його для очищання на ньому.
LEV|8|16|І взяв він увесь лій, що на нутрощах, і сальника на печінці, і обидві нирки та їхній лій, і Мойсей спалив на жертівнику.
LEV|8|17|А бичка, і шкуру його, і м'ясо його, і нечистість його спалив в огні поза табором, як Господь наказав був Мойсеєві.
LEV|8|18|І привів він барана цілопалення, і поклали Аарон та сини його руки свої на голову барана.
LEV|8|19|І зарізав, і покропив Мойсей кров'ю навколо жертівника.
LEV|8|20|А барана розсік на куски його, і Мойсей спалив голову, і куски, товщ.
LEV|8|21|А нутрощі та голінки пообмивав водою. І Мойсей спалив цілого барана на жертівнику, це цілопалення на пахощі любі, це огняна жертва для Господа, як Господь наказав був Мойсеєві.
LEV|8|22|І привів барана другого, барана посвячення. І поклали Аарон та сини його руки свої на голову того барана.
LEV|8|23|І зарізав, і взяв Мойсей із крови його та й дав на пипку правого вуха Ааронового й на великого пальця правої руки його, і на великого пальця правої ноги його.
LEV|8|24|І привів Ааронових синів, і дав Мойсей із крови тієї на пипку правого їхнього вуха, і на великого пальця правої руки їх, і на великого пальця правої ноги їх. І покропив Мойсей тією кров'ю жертівника навколо.
LEV|8|25|І взяв він лій, і курдюка, і ввесь лій, що на нутрощах, і сальника на печінці, і обидві нирки й їх лій, і стегно правиці.
LEV|8|26|А з коша з опрісноками, що перед лицем Господнім, узяв одного прісного калача та калача хлібного, одну оливу та одного коржика, і поклав на лої й на правім стегні.
LEV|8|27|І дав він усе на руки Аарона, і на руки синів його, і заколихав це, як колихання перед Господнім лицем.
LEV|8|28|І взяв це Мойсей із їхніх рук, та й спалив на жертівнику на цілопалення, воно жертва посвячення, на пахощі любі, воно огняна жертва для Господа.
LEV|8|29|І взяв Мойсей грудину та й заколихав її, як колихання перед Господнім лицем, із барана посвячення. Вона була для Мойсея на пайку, як Господь наказав був Мойсеєві.
LEV|8|30|І взяв Мойсей оливи помазання та крови, що на жертівнику, і покропив на Аарона, на шати його, і на синів його, і на шати синів його з ним. І посвятив Аарона, шати його, і синів його, і шати синів його з ним.
LEV|8|31|І сказав Мойсей до Аарона й до синів його: Варіть м'ясо при вході скинії заповіту, і там будете їсти його, і хліб, що в коші посвячення, як я наказав був, говорячи: Аарон та сини його будуть їсти його.
LEV|8|32|А позостале з м'яса та з хліба спалите в огні.
LEV|8|33|А із входу скинії заповіту не вийдете сім день, аж до дня виповнення днів вашого посвячення, бо Він буде сім день посвячувати вас.
LEV|8|34|Як учинив я сьогодні, так наказав Господь робити, щоб очистити вас.
LEV|8|35|А при вході скинії заповіту будете сидіти день і ніч сім день, і будете виконувати варту Господню, щоб вам не померти, бо так мені наказано.
LEV|8|36|І зробив Аарон та сини його все те, як наказав був Господь через Мойсея.
LEV|9|1|І сталося восьмого дня, закликав Мойсей Аарона та синів його, та старших Ізраїлевих,
LEV|9|2|та й сказав до Аарона: Візьми собі теля з худоби великої, на жертву за гріх, і барана на цілопалення, безвадних, і принеси перед Господнє лице.
LEV|9|3|А до синів Ізраїлевих будеш казати, говорячи: Візьміть козла на жертву за гріх, і теля й ягня однорічних, без вад, на цілопалення,
LEV|9|4|і вола, і барана на жертву мирну, на заріз перед Господнім лицем, і хлібну жертву, мішану в оливі, бо сьогодні об'явиться вам Господь.
LEV|9|5|І вони взяли, що наказав був Мойсей, перед скинію заповіту. І прийшла вся громада, та й стала перед Господнім лицем.
LEV|9|6|І сказав Мойсей: Оце та річ, що Господь наказав був, зробите, і об'явиться вам слава Господня.
LEV|9|7|І сказав Мойсей до Аарона: Підійди до жертівника, і вчини свою жертву за гріх та своє цілопалення, і очисти себе та народ, і вчини жертву за народ, і очисти їх, як наказав був Господь.
LEV|9|8|І підійшов Аарон до жертівника, та й зарізав теля жертви за свій гріх.
LEV|9|9|А сини Ааронові принесли до нього кров, і вмочив він свого пальця в кров, та й дав на роги жертівника, а кров вилив до підстави жертівника.
LEV|9|10|А лій і нирки та сальника на печінці з жертви за гріх спалив на жертівнику, як Господь наказав був Мойсеєві,
LEV|9|11|а м'ясо та шкуру спалив в огні поза табором.
LEV|9|12|І зарізав він жертву цілопалення, а Ааронові сини подали йому кров, і він покропив на жертівника навколо.
LEV|9|13|А цілопалення достачали йому його частинами, і голову, а він палив на жертівнику.
LEV|9|14|І обмив він нутрощі та голінки, і спалив на цілопаленні на жертівнику.
LEV|9|15|І приніс він жертву за народ, і взяв козла жертви за гріх народу, та й зарізав його, і склав його в жертві за гріх, як і першого.
LEV|9|16|І він приніс цілопалення, і вчинив його за постановою.
LEV|9|17|І він приніс хлібну жертву, і наповнив із неї руку свою, та й спалив на жертівнику, крім цілопалення ранкового.
LEV|9|18|І зарізав він вола й барана жертву мирну, що належить народові, а сини Ааронові принесли йому кров, і він покропив нею жертівника навколо,
LEV|9|19|і принесли лій з вола та з барана, курдюка, і лій, що покриває нутрощі, і нирки, і сальника на печінці.
LEV|9|20|І поклали вони лій на грудину, а він спалив лій на жертівнику.
LEV|9|21|А грудину та праве стегно Аарон колихав, як колихання перед Господнім лицем, як наказав був Мойсей.
LEV|9|22|І підняв Аарон свої руки до народу, та й поблагословив його, і зійшов від приношення жертви за гріх і цілопалення та мирної жертви.
LEV|9|23|І ввійшов Мойсей та Аарон до скинії заповіту; і вийшли вони, і поблагословили народ, і слава Господня показалася всьому народові.
LEV|9|24|І вийшов огонь від лиця Господнього, і спалив на жертівнику цілопалення та товщ. А ввесь народ бачив це, і закричали вони з радости, та й попадали на обличчя свої...
LEV|10|1|І взяли Ааронові сини, Надав та Авігу, кожен кадильницю свою, і дали в них огню, і поклали на ньому кадило, і принесли перед Господнє лице чужий огонь, якого Він не наказав був приносити їм.
LEV|10|2|І вийшов огонь від лиця Господнього, та й спалив їх, і вони повмирали перед Господнім лицем.
LEV|10|3|І сказав Мойсей до Аарона: Це те, про що говорив був Господь, кажучи: Серед близьких Моїх Я буду освячений, і перед усім народом буду прославлений. І замовк Аарон.
LEV|10|4|І покликав Мойсей Мисаїла та Елцафана, синів Уззіїла, Ааронового дядька, та й промовив до них: Підійдіть, винесіть братів своїх із святині поза табір.
LEV|10|5|І вони підійшли, та й винесли їх в їхніх хітонах поза табір, як наказав був Мойсей.
LEV|10|6|І сказав Мойсей до Аарона, та до Елеазара й до Ітамара, синів його: Голів ваших не відкривайте, і одеж ваших не роздирайте, щоб вам не померти, і щоб на всю громаду не розгнівався Він. А брати ваші, увесь дім Ізраїлів будуть оплакувати те спалення, що спалив Господь.
LEV|10|7|А зо входу скинії заповіту не вийдете ви, щоб не померти, бо на вас олива Господнього помазання. І зробили вони за Мойсеєвим словом.
LEV|10|8|А Господь промовляв до Аарона, говорячи:
LEV|10|9|Вина та п'янкого напою не пий ані ти, ані сини твої з тобою при вході вашім до скинії заповіту, щоб вам не померти. Це вічна постанова для ваших поколінь,
LEV|10|10|і щоб розрізняти між святістю й між несвятістю, і між нечистим та між чистим,
LEV|10|11|і щоб навчати Ізраїлевих синів усіх постанов, про що говорив до них Господь через Мойсея.
LEV|10|12|І Мойсей промовляв до Аарона та до Елеазара й до Ітамара, позосталих синів його: Візьміть хлібну жертву, полишену з огняних Господніх жертов, та й їжте її прісну при жертівнику, бо це Найсвятіше.
LEV|10|13|І будете їсти її в місці святому, бо вона уставова пайка твоя й уставова пайка синів твоїх з огняних жертов Господніх, бо так мені наказано.
LEV|10|14|А грудину колихання та стегно приношення будете їсти в місці чистому, ти й сини твої, та твої дочки з тобою, бо уставова пайка твоя й уставова пайка синів твоїх дані з мирних жертов Ізраїлевих синів.
LEV|10|15|Стегно приношення й грудину колихання на огняних жертвах лою принесуть вони, щоб колихати як колихання перед Господнім лицем. І буде це для тебе та для синів твоїх з тобою на вічну постанову, як наказав Господь.
LEV|10|16|А козла жертви за гріх пильно шукав Мойсей, і ось він був спалений. І розгнівався на Елеазара й на Ітамара, позосталих Ааронових синів, кажучи:
LEV|10|17|Чому ви не з'їли жертви за гріх у місці святому? Бо вона Найсвятіше, і її я дав вам, щоб уневажнити провину громади, щоб очистити їх перед Господнім лицем.
LEV|10|18|Тож не внесено крови її до святині всередину. Будете конче їсти її в святині, як я наказав.
LEV|10|19|І промовляв Аарон до Мойсея: От сьогодні принесли вони свою жертву за гріх і цілопалення своє перед Господнє лице, і трапилося мені оце. А буду я їсти жертву за гріх сьогодні, чи буде це добре в Господніх очах?
LEV|10|20|І почув Мойсей, і було це добре в його очах.
LEV|11|1|І Господь промовляв до Мойсея та до Аарона, говорячи їм:
LEV|11|2|Промовляйте до Ізраїлевих синів, кажучи: Оце та звірина, що будете їсти зо всієї худоби, що на землі:
LEV|11|3|Кожну з худоби, що має розділені копита, і що має копита роздвоєні розривом, що жує жуйку, її будете їсти.
LEV|11|4|Тільки цього не будете їсти з тих, що жують жуйку, і з тих, що мають розділені копита: верблюда, бо він жує жуйку, та розділених копит не має, нечистий він для вас.
LEV|11|5|І тушканчика, бо він жує жуйку, та не має розділених копит, нечистий він для вас.
LEV|11|6|І зайця, бо він жує жуйку, та не має розділених копит, нечистий він для вас.
LEV|11|7|І свині, бо вона має розділені ратиці, і має ратиці роздвоєні розривом, та жуйки не жує, нечиста вона для вас.
LEV|11|8|Їхнього м'яса не будете їсти, а до їхнього падла не будете доторкатися, нечисте воно для вас.
LEV|11|9|Оце будете їсти зо всього, що в воді: усе, що має плавці та луску в воді, у морях та в річках, їх будете їсти.
LEV|11|10|А все, що не має плавців та луски в морях і в річках, зо всього, що роїться в воді, і зо всього, що пливає в воді, гидота вони для вас!
LEV|11|11|І вони будуть гидота для вас, їхнього м'яса не будете їсти, а їхнього падла будете бридитися.
LEV|11|12|Усе, що не має плавців та луски в воді, гидота воно для вас.
LEV|11|13|А з птаства будете бридитися оцього, не будете їх їсти, гидота вони: орла, грифа й морського орла,
LEV|11|14|і коршака, і сокола за родом його,
LEV|11|15|усякого крука за родом його,
LEV|11|16|і струся, і сови, і яструба за родом його,
LEV|11|17|і пугача, і рибалки, та ібіса,
LEV|11|18|і лебедя, і пелікана, і сича,
LEV|11|19|і бусла, чаплі за родом її, і одуда, і нетопира.
LEV|11|20|Уся комашня, що ходить на чотирьох, гидота вона для вас.
LEV|11|21|Тільки те будете їсти зо всієї комашні, що ходить на чотирьох, що має голінки вище своїх ніг, щоб ними скакати на землі.
LEV|11|22|Оці серед них будете їсти: сарану за родом її, і сол'ам за родом його, і харґол за родом його, і хаґав за родом його.
LEV|11|23|А вся гадина летюча, що має чотири ноги, гидота вона для вас.
LEV|11|24|І через них ви будете ставати нечисті: кожен, хто доторкнеться до їхнього падла, буде нечистий аж до вечора.
LEV|11|25|А кожен, хто понесе що з їхнього падла, випере одежу свою, і буде нечистий аж до вечора.
LEV|11|26|Щодо всякої худоби, що має розділене копито, і що не має роздвоєного розривом копита, і жуйки не жує, нечисті вони для вас. Кожен, хто доторкнеться до них, буде нечистий.
LEV|11|27|А кожне серед усякої звірини, що ходить на лапах своїх, що ходить на чотирьох, нечисті вони для вас. Кожен, хто доторкнеться до їхнього падла, буде нечистий аж до вечора.
LEV|11|28|А хто носить їхнє падло, випере одежу свою, і буде нечистий аж до вечора. Нечисті вони для вас.
LEV|11|29|А оце вам нечисте серед плазунів, що плазують по землі: кріт, і миша, і ящірка за родом її,
LEV|11|30|і ховрах, і щур, і слимак, і їжак, і тхір.
LEV|11|31|Оці нечисті для вас серед усього плазуючого. Кожен, хто доторкнеться до них, коли вони мертві, буде нечистий аж до вечора.
LEV|11|32|І все, що впаде на нього, коли вони мертві, буде нечисте, кожна річ, з дерева, або з одежі, або зо шкури, або з грубої тканини, кожна річ, що вживається до праці, в воду треба покласти їх, і будуть нечисті аж до вечора, а потому стануть чистими.
LEV|11|33|А всякий глиняний посуд, що з них упаде що до його середини, усе, що в середині його, стане нечисте, а його розіб'єте.
LEV|11|34|Кожна їжа, що їсться, на якій була вода з такого посуду, буде нечиста; а кожен напій, що п'ється, у кожнім такім посуді стане нечистим.
LEV|11|35|І все, що на нього впаде з їхнього падла, стане нечисте: піч та огнище буде розвалене, вони нечисті, і нечисті будуть для вас.
LEV|11|36|Тільки джерело та яма, збір води, будуть чисті. А хто доторкнеться до їхнього падла, буде нечистий.
LEV|11|37|А коли що впаде з їхнього падла на всяке насіння сівби, що сіється, чисте воно.
LEV|11|38|А коли буде налита вода на насіння, і впаде на нього з їхнього падла, нечисте воно для вас.
LEV|11|39|А коли помре що з худоби, що вона на їжу для вас, то хто доторкнеться падла її, той буде нечистий аж до вечора.
LEV|11|40|А хто їсть із падла її, той випере одежу свою, і буде нечистий аж до вечора. І хто носить падло її, той випере одежу свою, і буде нечистий аж до вечора.
LEV|11|41|А все плазуюче, що плазує по землі, гидота воно, не буде їстися.
LEV|11|42|Усе, що повзає на животі, і все, що повзає на чотирьох, аж до всього, що багатоножне, усе плазуюче, що плазує по землі, не будете їх їсти, бо гидота вони.
LEV|11|43|Не занечищуйте душ своїх усім плазуючим, що плазує, і не зробитеся нечисті ними, і не станете нечисті ними.
LEV|11|44|Бо Я Господь, Бог ваш, і ви освятитеся, і будьте святі, бо святий Я, і не занечищуйте душ своїх усяким плазуючим, що плазує по землі.
LEV|11|45|Бо Я Господь, що вивів вас із єгипетського краю, щоб бути для вас Богом. І будьте святі, бо святий Я.
LEV|11|46|Оце закон про худобу, і про птаство, і про всяку живу звірину, що рухається в воді, і про всяку душу, що плазує по землі,
LEV|11|47|щоб відділювати між нечистим та між чистим, і між звіриною, що їсться, та між звіриною, що не їсться.
LEV|12|1|І Господь промовляв до Мойсея, говорячи:
LEV|12|2|Промовляй до Ізраїлевих синів, говорячи: Коли жінка зачне, і породить дитя чоловічої статі, то буде нечиста сім день; як за днів нечистоти місячного її, буде нечиста вона.
LEV|12|3|А восьмого дня буде обрізане тіло крайньої плоті його.
LEV|12|4|І буде вона сидіти в крові очищення тридцять день і три дні. До всякої святощі не буде вона доторкатися, а до святині не ввійде аж до виповнення днів очищення її.
LEV|12|5|А якщо породить дитя жіночої статі, то буде нечиста вона два тижні, як за нечистости її місячної, і буде сидіти вона на крові очищення шістдесят день і шість день.
LEV|12|6|А по виповненні днів очищення її за сина або за дочку, принесе вона однорічне ягня на цілопалення, та голубеня або горлицю на жертву за гріх, до входу скинії заповіту до священика.
LEV|12|7|І він принесе це перед Господнє лице, і очистить її, і вона очиститься від джерела своєї крови. Це закон про породіллю дитини чоловічої або жіночої статі.
LEV|12|8|А коли рука її не спроможеться на ягня, то візьме вона дві горлиці або двоє голубенят, одне на цілопалення й одне на жертву за гріх, й очистить її священик, і вона стане чиста.
LEV|13|1|І Господь промовляв до Мойсея й Аарона, говорячи:
LEV|13|2|Чоловік, коли буде на шкурі тіла його напухлина, або лишай, або біла пляма, і буде на шкурі тіла його ніби болячка прокази, то буде спроваджений він до священика Аарона або одного з синів його, священиків.
LEV|13|3|І огляне священик ту болячку на шкурі тіла, а волосся на болячці перемінилося на біле, і вигляд болячки глибший від шкури тіла його, болячка прокази воно. І огляне її священик, і визнає його за нечистого.
LEV|13|4|А якщо болячка біла вона на шкурі тіла його, а вигляд її не глибший від шкури, і волосся її не перемінилося на біле, то замкне священик хворого на сім день.
LEV|13|5|І огляне її священик сьомого дня, а ось болячка, на погляд його, спинилася, не поширилася та болячка по шкурі, то замкне його священик удруге на сім день.
LEV|13|6|І огляне його священик сьомого дня вдруге, а ось болячка поблідла, не поширилася та болячка по шкурі, то священик визнає його за чистого, лишай вона. І випере він одежу свою та й стане чистий.
LEV|13|7|А якщо справді пошириться лишай той по шкурі по явленні священику на очищення його, то явиться він удруге до священика.
LEV|13|8|І огляне священик, а ось лишай той поширився по шкурі, то священик визнає його за нечистого, проказа воно.
LEV|13|9|Коли буде на людині болячка прокази, то буде приведена до священика.
LEV|13|10|І огляне священик, а ось на шкурі біла напухлина, і вона перемінила волосся на біле, і на напухлині ріст живого м'яса,
LEV|13|11|то це стара проказа на шкурі тіла його. І священик визнає його за нечистого, але не замкне його, бо справді давно він нечистий.
LEV|13|12|А якщо справді кинеться та проказа по шкурі, і покриє та проказа всю шкуру хворого від голови його аж до ніг його, куди лиш глянуть очі священикові,
LEV|13|13|і огляне священик, а ось проказа та покрила все тіло його, то він визнає за чисту ту болячку: вся вона перемінилася на білу, чиста вона.
LEV|13|14|А того дня, коли в ній побачиться живе м'ясо, він стане нечистий.
LEV|13|15|І огляне священик живе м'ясо, і визнає його за нечистого; те живе м'ясо нечисте воно, проказа воно.
LEV|13|16|Або коли живе м'ясо знову переміниться на біле, то він прийде до священика.
LEV|13|17|І огляне його священик, а ось перемінилася болячка на білу, то священик визнає ту болячку за чисту, чиста вона.
LEV|13|18|А тіло, коли буде на ньому на шкурі його гнояк, і він вилікуваний,
LEV|13|19|а на місці гнояка буде біла напухлина, або біла, червонява пляма, то покажеться священикові.
LEV|13|20|І огляне священик, а ось вигляд її нижчий від шкури, а волосся її перемінилося на біле, то священик визнає її за нечисту, болячка прокази вона, вона кинулась на гнояку.
LEV|13|21|А якщо огляне її священик, а ось нема в ній білого волосся, і вона не нижча від шкури, і вона бліда, то замкне його священик на сім день.
LEV|13|22|А якщо справді пошириться по шкурі, то священик визнає його за нечистого, болячка прокази вона.
LEV|13|23|А якщо біла пляма спинилася на своєму місці, не поширилася, вона струп чиряка, і священик визнає його за чистого.
LEV|13|24|Або тіло, коли буде на шкурі його опалення від огню, і буде заріст того опалення плямкою білою червонявою або білою,
LEV|13|25|то огляне її священик, а ось перемінилось волосся в плямі на біле, а вид її глибший від шкури, проказа вона, в опаленні кинулась. І визнає священик його за нечистого, болячка прокази вона.
LEV|13|26|А якщо священик огляне її, а ось у плямі нема білого волосу, і вона не нижча від шкури, і вона бліда, то священик замкне його на сім день.
LEV|13|27|І огляне його священик восьмого дня. Якщо справді пошириться по шкурі, то священик визнає його за нечистого, болячка прокази вона.
LEV|13|28|А якщо пляма спиниться на своїм місці, не поширилася по шкурі, і вона бліда, вона напухлина опалення. І священик визнає його за чистого, бо струп опалення вона.
LEV|13|29|А чоловік або жінка, коли буде на кому болячка на голові або на бороді,
LEV|13|30|то священик огляне ту болячку, а ось вид її глибший від шкури, а в ній жовтий, тонкий волос, то священик визнає його за нечисту, парші вона, вона проказа голови або бороди.
LEV|13|31|А коли священик огляне болячку паршів, а ось вид її не глибший від шкури, і в ній нема чорного волосу, то священик замкне хворого на парші на сім день.
LEV|13|32|І огляне священик ту болячку сьомого дня, а ось не поширилися парші, і волосся в них не стали жовті, а вид паршів не глибший від шкури,
LEV|13|33|то він поголиться, а паршів не поголить. І замкне священик хворого на парші вдруге на сім день.
LEV|13|34|І огляне священик парші сьомого дня, а ось парші не поширилися по шкурі, і їхній вид не глибший від шкури, то священик визнає його за чистого, і він випере одежу свою, і стане чистий.
LEV|13|35|А якщо справді поширяться парші по шкурі по його очищенні,
LEV|13|36|то священик огляне його, а ось поширились парші по шкурі, то священик не буде досліджувати щодо жовтого волосся, нечистий він.
LEV|13|37|А якщо, на його погляд парші спинилися, і в них виросло чорне волосся, то парші вилікувані, він чистий. І священик визнає його за чистого.
LEV|13|38|А чоловік або жінка, коли на шкурі їхнього тіла буде багато білих плям,
LEV|13|39|то огляне священик, а ось на шкурі їхнього тіла бліді білі плями, лишай воно, кинувся на шкурі, чистий він.
LEV|13|40|А коли в кого облізе голова його, лисий він, він чистий.
LEV|13|41|А якщо голова його облізла спереду його, лисий він спереду, він чистий.
LEV|13|42|А коли на лисині ззаду або на лисині спереду буде біла червонява болячка, це проказа, кинулась вона в лисині задній його або в лисині передній його.
LEV|13|43|І огляне його священик, а ось напухлина болячки біла червонява в лисині задній його або в лисині передній його, як вигляд прокази на шкурі тіла,
LEV|13|44|то це чоловік прокажений, нечистий він. Конче визнає священик його за нечистого, на голові його болячка його.
LEV|13|45|А прокажений, що проказа на ньому, одежа його буде роздерта, а голова його буде відкрита, і по уста закриє, і буде кричати: Нечистий, нечистий!
LEV|13|46|По всі дні, коли болячка на ньому, буде нечистий, він нечистий. Самітний буде пробувати він, поза табором оселя його.
LEV|13|47|А одежа, коли буде на ній зараза прокази, на одежі вовняній або на одежі льняній,
LEV|13|48|або на нитці прямовісній, або на нитці поземій із льону та вовни, або на шкурі, або на всякім шкурянім виробі,
LEV|13|49|і буде та зараза зеленява або червонява на одежі, або на шкурі, або на нитці прямовісній, або на нитці поземій, або на всякій шкуряній речі, зараза прокази воно. І буде воно показане священикові.
LEV|13|50|І огляне священик ту заразу, та й замкне заразливе на сім день.
LEV|13|51|А дня сьомого огляне він ту заразу; коли зараза та поширилася на одежі, або на нитці прямовісній, або на нитці поземій, або на шкурі, на всьому, що зроблене зо шкури, та зараза злослива проказа, нечиста вона.
LEV|13|52|І він спалить ту одежу, або нитку прямовісну, або нитку позему в вовні або в льоні, або всяку річ шкуряну, що буде на ній зараза, бо злослива проказа це, огнем буде спалена.
LEV|13|53|А якщо священик побачить, а ось не поширилася зараза на одежі, або на нитці прямовісній, або на нитці поземій, або на всякій речі шкуряній,
LEV|13|54|то священик накаже, і виперуть те, що на ньому зараза. І він замкне те вдруге на сім день.
LEV|13|55|І огляне священик заразу по випранні, і ось, зараза не перемінила свого вигляду, і зараза не поширилася, нечиста вона, огнем її спалите; вона заглиблення на стороні його передній або на стороні його задній.
LEV|13|56|А якщо священик побачив, а ось зараза та зблідла по випранні її, то він відірве її від одежі або від шкури, або від нитки прямовісної, або від нитки поземої.
LEV|13|57|А якщо вона покажеться ще на одежі, або на нитці прямовісній, або на нитці поземій, або на якій шкуряній речі, то це шириться вона, огнем спалиш те, що на ньому та зараза.
LEV|13|58|А одежа, або нитка прямовісна, або нитка позема, або яка шкуряна річ, що випереш і зійде від них та зараза, то буде випрана вдруге, і буде чиста.
LEV|13|59|Оце закон про хворобу прокази на одежі вовняній або на льняній, або на нитці прямовісній, або на нитці поземій, або на шкурі, на очищення її або на признання її за нечисту.
LEV|14|1|І Господь промовляв до Мойсея, говорячи:
LEV|14|2|Оце буде закон про прокаженого в дні очищення його: І буде він приведений до священика.
LEV|14|3|І вийде священик поза табір, і огляне священик, а ось вилікувана хвороба прокази в прокаженого,
LEV|14|4|то священик накаже, і візьме для очищуваного двох живих чистих птахів, і кедрового дерева, і червону нитку, та ісопу.
LEV|14|5|І накаже священик, і заріже одного птаха до глиняного посуду над живою водою.
LEV|14|6|Птаха живого він візьме його, і кедрового дерева, і червону нитку, та ісопу, і вмочить їх та живого птаха в крові птаха, зарізаного над живою водою.
LEV|14|7|І покропить на очищуваного від прокази сім раз, та й очистить його, а живого птаха пустить у поле.
LEV|14|8|А очищуваний випере одежу свою й поголить усе волосся своє, і обмиється в воді, стане чистий. А потому ввійде до табору, і буде жити поза наметом своїм сім день.
LEV|14|9|І станеться сьомого дня, поголить він усе волосся своє, свою голову, і бороду свою, і брови очей своїх, і все волосся своє оголить, і випере одежу свою, і вимиє тіло своє в воді, і стане він чистий.
LEV|14|10|А восьмого дня візьме він двоє баранців безвадних, і одну однорічну безвадну вівцю і три десятих пшеничної муки, жертва хлібна, мішана в оливі, і одного лоґа оливи.
LEV|14|11|І поставить священик, що очищує, чоловіка очищуваного з ними перед Господнім лицем при вході скинії заповіту.
LEV|14|12|І візьме священик одного баранця, і принесе його на жертву за гріх, та лоґа оливи, та й буде колихати їх, як колихання перед Господнім лицем.
LEV|14|13|І він заріже того баранця в місці, де ріже жертву за гріх і цілопалення, у місці святині, бо як жертва за гріх та жертва за провину, вона для священика, найсвятіше вона.
LEV|14|14|І візьме священик крови жертви за провину, та й дасть священик на пипку правого вуха очищуваного, і на великого пальця правої руки його та на великого пальця правої ноги його.
LEV|14|15|І візьме священик з лоґу оливи, та й виллє на ліву долоню свою.
LEV|14|16|І вмочить священик правого пальця свого в оливу, що на лівій долоні його, і покропить з оливи пальцем своїм сім раз перед Господнім лицем.
LEV|14|17|А з решти оливи, що на долоні його, священик дасть на пипку правого вуха очищуваного, і на великого пальця правої руки його та на великого пальця правої ноги його на кров жертви за провину.
LEV|14|18|А позостале з оливи, що на долоні священиковій, дасть на голову очищуваного. І священик очистить його перед Господнім лицем.
LEV|14|19|І вчинить священик жертву за гріх, і очистить очищуваного з нечистоти його, а потім заріже цілопалення.
LEV|14|20|І зложить священик те цілопалення та ту хлібну жертву на жертівнику, і священик очистить його, і стане він чистий.
LEV|14|21|А якщо він бідний, і рука його неспроможна, то візьме одного баранця на жертву за провину на колихання, щоб очистити його, і одну десяту ефи пшеничної муки, мішану в оливі, і лоґа оливи,
LEV|14|22|та дві горлиці або двоє голубенят, на що спроможна рука його, і буде одне жертва за гріх, а одне цілопалення.
LEV|14|23|І він принесе їх восьмого дня на своє очищення до священика, до входу скинії заповіту перед Господнє лице.
LEV|14|24|І візьме священик ягня жертви за провину й лоґа оливи, та й буде колихати їх священик, як колихання перед Господнім лицем.
LEV|14|25|І заріже ягня жертви за провину, і візьме священик крови жертви за провину, та й дасть на пипку правого вуха очищуваного, і на великого пальця правої руки його та на великого пальця правої ноги його.
LEV|14|26|А з оливи виллє священик на ліву долоню свою.
LEV|14|27|І покропить священик своїм правим пальцем з оливи, що на лівій долоні його, сім раз перед Господнім лицем.
LEV|14|28|І дасть священик із оливи, що на долоні його, на пипку правого вуха очищуваного, і на великого пальця правої руки його та на великого пальця правої ноги його, на місце крови жертви за провину.
LEV|14|29|А позостале з оливи, що на священиковій долоні, дасть на голову очищуваного на очищення його перед Господнім лицем.
LEV|14|30|І він спорядить одну з горлиць або з голубенят із того, на що спроможна рука його,
LEV|14|31|на що спроможна рука його, одне жертва за гріх, а одне цілопалення понад жертву хлібну. І очистить священик очищуваного перед Господнім лицем.
LEV|14|32|Оце закон про того, що в ньому хвороба прокази, що рука його неспроможна при очищенні його.
LEV|14|33|І Господь промовляв до Мойсея й до Аарона, говорячи:
LEV|14|34|Коли ви ввійдете до ханаанського Краю, що Я даю вам на володіння, і наведу хворобу прокази на доми Краю вашого володіння,
LEV|14|35|то прийде той, що його той дім, та й скаже священикові, говорячи: Ніби зараза показалася мені в домі.
LEV|14|36|І накаже священик, і опорожнять той дім, поки прийде священик, щоб оглянути заразу, щоб не стало нечистим усе, що в домі. А потому ввійде священик, щоб оглянути той дім.
LEV|14|37|І він огляне заразу, і ось у стінах дому заглиблення зеленяві або червоняві, а їхній вид нижчий від стіни.
LEV|14|38|І вийде священик із того дому до виходу дому того, і замкне той дім на сім день.
LEV|14|39|І вернеться священик сьомого дня та й огляне, а ось поширилася та зараза на стінах того дому.
LEV|14|40|І накаже священик, і витягнуть каміння, що на них та зараза, та й кинуть їх поза місто, до місця нечистого.
LEV|14|41|А дім той він вишкребе зсередини кругом, а глину, що вишкребли, висиплють поза містом, до нечистого місця.
LEV|14|42|І візьмуть інше каміння, і покладуть замість того каміння, і візьме інший тинк і обтинкує той дім.
LEV|14|43|А якщо вернеться та зараза, і кинеться в домі по витягненні того каміння й по вишкребанні того дому й по обтинкуванні,
LEV|14|44|то ввійде священик і огляне, а ось поширилася та зараза в тім домі, проказа злослива вона в тім домі, нечистий він.
LEV|14|45|І розвалить той дім, і каміння його, і дерево його, і ввесь тинк дому, і винесе поза місто, до нечистого місця.
LEV|14|46|А хто входить до того дому всі дні, коли він замикав його, той буде нечистий аж до вечора.
LEV|14|47|А хто лежить у тім домі, той випере одежу свою, і хто їсть у тім домі, той випере одежу свою.
LEV|14|48|А якщо знову ввійде священик і побачить, а ось не поширилася зараза в домі по обтинкуванні дому, то священик визнає той дім за чистий, бо зараза вилікувана.
LEV|14|49|І візьме він на очищення того дому два птахи, і кедрового дерева, і червені, та ісопу.
LEV|14|50|І заріже одного птаха до глиняного посуду над живою водою.
LEV|14|51|І візьме він кедрового дерева, та ісопу, і червені, і живого птаха, та й умочить їх у крові зарізаного птаха та в живій воді, і сім раз покропить на той дім.
LEV|14|52|І очистить він той дім пташиною кров'ю, і живою водою, і птахом живим, і кедровим деревом, і ісопом, і червенню.
LEV|14|53|І пустить він живого птаха поза місто на поле, і очистить дім той, і він стане чистий.
LEV|14|54|Оце закон для всякої хвороби прокази та для паршів,
LEV|14|55|і для прокази одежі, і для дому,
LEV|14|56|і для напухлини, і для лишаю, і для білої плями,
LEV|14|57|для навчання на день занечищення й на день відчищення. Оце закон про проказу.
LEV|15|1|І Господь промовляв до Мойсея й до Аарона, говорячи:
LEV|15|2|Промовляйте до Ізраїлевих синів і скажіть їм: Кожен чоловік, коли з його тіла тектиме теча його, нечистий він.
LEV|15|3|А це буде про нечистість його в течі його: коли тіло його випускає течу свою, або коли в тілі його задержалась теча його, воно нечистість його.
LEV|15|4|Кожне ложе, що течивий ляже на ньому, буде нечисте, і кожна річ, що він сяде на ній, буде нечиста.
LEV|15|5|І кожен, хто доторкнеться ложа його, випере свою одежу й обмиється в воді, і буде нечистий аж до вечора.
LEV|15|6|А хто сяде на річ, що на ній сидів течивий, той випере одежу свою й обмиється в воді, і буде нечистий аж до вечора.
LEV|15|7|А хто доторкнеться до тіла течивого, той випере одежу свою й обмиється в воді, і буде нечистий аж до вечора.
LEV|15|8|А коли течивий плюне на чистого, то випере той одежу свою й обмиється в воді, і буде нечистий аж до вечора.
LEV|15|9|І кожен повіз, що на нім конно їде течивий, буде нечистий.
LEV|15|10|І кожен, хто доторкнеться до всього, що буде під ним, буде нечистий аж до вечора. А хто їх носить, той випере одежу свою й обмиється в воді, і буде нечистий аж до вечора.
LEV|15|11|І кожен, кого доторкнеться течивий, а рук своїх він не обілляв водою, то випере він одежу свою й обмиється в воді, і буде нечистий аж до вечора.
LEV|15|12|А глиняний посуд, що його доторкнеться течивий, буде розбитий, а кожен посуд дерев'яний буде обмитий водою.
LEV|15|13|А коли течивий стане чистий від течі своєї, то він відлічить сім день на своє очищення, і випере одежу свою, і обмиє тіло своє в живій воді, і стане чистий.
LEV|15|14|А восьмого дня він візьме собі дві горлиці або двоє голубенят, та й прийде перед лице Господнє до входу скинії заповіту, і дасть їх священикові.
LEV|15|15|І спорядить їх священик: одне жертвою за гріх, а одне цілопаленням, та й очистить священик його перед Господнім лицем від течі його.
LEV|15|16|А чоловік, коли вийде з нього насіння парування, то обмиє в воді все тіло своє, і буде нечистий аж до вечора.
LEV|15|17|А всяка одежа й всяка шкура, що на ній буде насіння парування, то вона буде випрана в воді, і буде нечиста аж до вечора.
LEV|15|18|І жінка, що чоловік лежатиме з нею на парування, то обмиються вони в воді, і будуть нечисті аж до вечора.
LEV|15|19|А жінка, коли буде течива, кров буде течею її в тілі її то сім день буде в своїй нечистості, а кожен, хто доторкнеться її, буде нечистий аж до вечора.
LEV|15|20|І все, на чому вона лежатиме в нечистості своїй, буде нечисте; і все, на чому вона сяде, буде нечисте.
LEV|15|21|А кожен, хто доторкнеться до місця лежання її, той випере одежу свою й обмиється в воді, і буде нечистий аж до вечора.
LEV|15|22|А кожен, хто доторкнеться до всякої речі, на якій вона сидить, той випере одежу свою й обмиється в воді, і буде нечистий аж до вечора.
LEV|15|23|А якщо було б щось на ложі або на тій речі, що вона сиділа на ній, і він доторкнеться того, то буде нечистий аж до вечора.
LEV|15|24|А якщо буде лежати чоловік із нею, то нечистість її буде на ньому, і буде він нечистий сім день.
LEV|15|25|А жінка, коли буде текти теча крови її багато днів не в часі нечистости її, або коли буде текти понад нечистості її, то всі дні течі нечистости її буде вона, як за днів нечистости її, нечиста вона.
LEV|15|26|Кожне ложе, на якому вона лежатиме всі дні течі її, буде для неї, як ложе її нечистости. І кожна річ, на яку вона сяде, буде нечиста, як нечистість місячного очищення її.
LEV|15|27|І кожен, хто доторкнеться до них, буде нечистий, і випере одежу свою, і обмиється в воді, і буде нечистий аж до вечора.
LEV|15|28|А якщо вона очиститься від течі своєї, то відлічить собі сім день, а потому стане чиста.
LEV|15|29|А восьмого дня візьме собі дві горлиці, або двоє голубенят, та й принесе їх до священика до входу скинії заповіту.
LEV|15|30|І спорядить священик одне жертвою за гріх, а одне цілопаленням, та й очистить священик її перед Господнім лицем від течі нечистости її.
LEV|15|31|І відділите Ізраїлевих синів від їхньої нечистости, щоб не повмирали вони в своїй нечистості через занечищення їхнє Моєї скинії, яка серед них.
LEV|15|32|Оце закон про течивого та про того, що з нього виходить насіння лежання, що ним занечищується,
LEV|15|33|і про хвору в місячнім очищенні її, і про течивого на течу свою, для чоловіка й для жінки, та для чоловіка, що буде лежати з нечистою.
LEV|16|1|І Господь промовляв до Мойсея по смерті обох Ааронових синів, коли вони були наблизилися перед Господнє лице і померли.
LEV|16|2|І сказав Господь до Мойсея: Промовляй до Аарона, брата свого, і нехай він не входить кожного часу до святині за завісу, перед віко, що на ковчезі, щоб не вмер він, бо Я в хмарі являюся над тим віком.
LEV|16|3|З оцим увійде Аарон до святині, з телям на жертву за гріх та з бараном на цілопалення.
LEV|16|4|Він зодягне священного льняного хітона, і льняна спідня одіж буде на тілі його, і підпережеться льняним поясом, і обвинеться льняним завоєм, вони священні шати. І обмиє в воді своє тіло, та й зодягне він їх.
LEV|16|5|А від громади Ізраїлевих синів візьме він два козли на жертву за гріх та одного барана на цілопалення.
LEV|16|6|І принесе Аарон теля жертви за гріх, що належить йому, та й очистить себе та свій дім.
LEV|16|7|І візьме він обох тих козлів, та й поставить їх перед Господнім лицем при вході скинії заповіту.
LEV|16|8|І кине Аарон на обох тих козлів жеребки, один жеребок для Господа, і один жеребок для Азазеля.
LEV|16|9|І принесе Аарон козла, що на нього вийшов жеребок для Господа, і вчинить його жертвою за гріх.
LEV|16|10|А козел, що на нього випав жеребок для Азазеля, буде поставлений живим перед Господнє лице, щоб очистити його, і щоб послати його до Азазеля на пустиню.
LEV|16|11|І принесе Аарон бичка жертви за гріх, що належить йому, та й очистить себе та свій дім; і заріже бичка жертви за гріх, що належить йому.
LEV|16|12|І візьме повну кадильницю горючого вугілля з-над жертівника перед Господнім лицем, і повні жмені свої тонко товченого запашного кадила, та й внесе за завісу.
LEV|16|13|І покладе він те кадило на огонь перед Господнім лицем, а хмара кадила закриє віко, що над свідоцтвом, щоб він не помер.
LEV|16|14|І візьме він крови бичка, та й покропить пальцем своїм на переді віка на схід, а перед віком покропить з крови сім раз своїм пальцем.
LEV|16|15|І заріже козла жертви за гріх, що належить народові, і внесе його кров за завісу, та й зробить із кров'ю його, як зробив був із кров'ю теляти, і покропить її на віко та перед віком.
LEV|16|16|І очистить він святиню з нечистости Ізраїлевих синів та з їхніх переступів через усі гріхи їхні. І так він зробить для скинії заповіту, що знаходиться з ними серед їхньої нечистости.
LEV|16|17|І жоден чоловік не буде в скинії заповіту, коли він входить на очищення до святині, аж до виходу його. І очистить він себе та дім свій, та всю громаду Ізраїлеву.
LEV|16|18|І вийде він до жертівника, що перед Господнім лицем, та й очистить його; і візьме крови теляти й крови козла, та й дасть на роги жертівника навколо.
LEV|16|19|І покропить на нього з крови пальцем своїм сім раз, та й очистить його, та освятить його від нечистости Ізраїлевих синів.
LEV|16|20|А коли він скінчить очищення святині й скинії заповіту та жертівника, то приведе живого козла.
LEV|16|21|І покладе Аарон обидві руки свої на голову живого козла, і визнає над ним усі гріхи Ізраїлевих синів та всі їхні провини через усі їхні гріхи, і складе їх на голову козла, та й пошле через призначеного чоловіка на пустиню.
LEV|16|22|І понесе той козел на собі всі їхні гріхи до краю неврожайного, і пустить того козла в пустиню.
LEV|16|23|І ввійде Аарон до скинії заповіту, і здійме льняні шати, що зодягнув був при вході його до святині, і покладе їх там.
LEV|16|24|І обмиє він тіло своє в воді в місці святім, і зодягне шати свої та й вийде, і вчинить цілопалення своє та цілопалення за народ, і очистить себе та народ.
LEV|16|25|А лій жертви за гріх спалить на жертівнику.
LEV|16|26|А той, хто відводив козла до Азазеля, випере одежу свою й обмиє тіло своє в воді, а потому ввійде до табору.
LEV|16|27|А теля жертви за гріх та козла жертви за гріх, що їхню кров внесено на очищення в святині, випровадять поза табір, та й спалять в огні їхні шкури, і їхнє м'ясо та їхні нечистости.
LEV|16|28|А той, хто їх палить, випере одежу свою й обмиє своє тіло в воді, а потому ввійде до табору.
LEV|16|29|І це стане для вас на вічну постанову, сьомого місяця, десятого дня місяця будете впокоряти ваші душі, і жодної праці не робитимете ви, ані тубілець, ані приходько, що мешкає серед вас,
LEV|16|30|бо того дня буде окуп ваш на очищення ваше, зо всіх гріхів ваших станете чисті перед Господом.
LEV|16|31|Субота повного відпочинку від праці вона для вас, і ви будете впокоряти душі свої, це вічна постанова.
LEV|16|32|А очистить той священик, що помазали його, і що посвятили його бути священиком замість батька свого. І зодягне він льняні шати, шати священні,
LEV|16|33|та й очистить Святеє Святих, і скинію заповіту, і жертівника очистить, і очистить священиків та ввесь народ громади.
LEV|16|34|І буде це для вас на вічну постанову на очищення Ізраїлевих синів зо всіх їхніх гріхів раз у році. І він учинив, як Господь наказав був Мойсеєві.
LEV|17|1|І Господь промовляв до Мойсея, говорячи:
LEV|17|2|Промовляй до Аарона й до синів його, та до всіх Ізраїлевих синів, та й скажеш їм: Оце та річ, що Господь наказав був, говорячи:
LEV|17|3|Кожен чоловік з Ізраїлевого дому, що заріже вола, або ягня, або козу в таборі, або щось заріже поза табором,
LEV|17|4|а до входу скинії заповіту не приведе того на принесення жертви для Господа перед скинію Господню, то кров буде полічена тому чоловікові, він пролив кров. І буде винищений чоловік той з-посеред народу свого,
LEV|17|5|щоб приводили Ізраїлеві сини свої жертви, які вони ріжуть на чистому полі, і спроваджали для Господа до входу скинії заповіту до священика, і різали їх, як мирні жертви для Господа.
LEV|17|6|І покропить священик тією кров'ю на Господнього жертівника при вході скинії заповіту, та й спалить лій на любі пахощі для Господа.
LEV|17|7|І щоб вони вже не різали своїх жертов козлам-демонам, за якими вони блудять. Це буде для них вічна постанова на їхні покоління.
LEV|17|8|А їм скажеш: Кожен чоловік із Ізраїлевого дому та з приходька, що буде мешкати серед вас, який принесе цілопалення або жертву,
LEV|17|9|а до входу скинії заповіту не принесе того, щоб учинити його для Господа, то буде знищений чоловік той з-посеред народу свого!
LEV|17|10|А кожен чоловік із Ізраїлевого дому та з приходька, що мешкає серед них, який буде їсти кров, то Я зверну лице Своє проти тієї душі, що їсть вона ту кров, і винищу її з-посеред народу її,
LEV|17|11|бо душа тіла в крові вона, а Я дав її для вас на жертівника для очищення за душі ваші, бо кров та вона очищує душу.
LEV|17|12|Тому сказав Я Ізраїлевим синам: Кожна душа з вас не буде їсти крови, і приходько, що мешкає серед вас, не буде їсти крови.
LEV|17|13|А кожен чоловік із Ізраїлевих синів та з приходька, що мешкає серед них, що вполює здобич звірини або птаства, що їджене, то він виллє кров того й закриє її піском.
LEV|17|14|Бо душа кожного тіла кров його, у душі його вона. І сказав Я Ізраїлевим синам: Крови кожного тіла ви не будете їсти, бо душа кожного тіла кров його вона. Усі, що їдять її, будуть понищені.
LEV|17|15|А всяка душа, що їстиме падло та розшарпане серед тубільця і серед приходька, нехай випере одежу свою й обмиється в воді, і буде нечистий аж до вечора, а потім стане чистий.
LEV|17|16|А якщо він не випере, а тіла свого не обмиє, то понесе свою провину.
LEV|18|1|І Господь промовляв до Мойсея, говорячи:
LEV|18|2|Промовляй до Ізраїлевих синів, і скажеш їм: Я Господь, Бог ваш!
LEV|18|3|За чином єгипетського краю, що сиділи ви в нім, не робіть, і за чином Краю ханаанського, що Я впроваджую вас туди, не зробите, і звичаями їхніми не підете.
LEV|18|4|Ви виконуватимете устави Мої, і будете додержувати постанови Мої, щоб ними ходити. Я Господь, Бог ваш!
LEV|18|5|І будете додержувати постанов Моїх та уставів Моїх, що людина їх виконує й ними живе. Я Господь!
LEV|18|6|Жоден чоловік не наблизиться до жодної однокровної своєї, щоб відкрити наготу. Я Господь!
LEV|18|7|Наготи батька свого й наготи матері своєї не відкриєш, вона мати твоя, не відкриєш наготи її!
LEV|18|8|Наготи жінки батька твого не відкриєш, вона нагота батька твого!
LEV|18|9|Наготи сестри своєї, дочки батька свого або дочки матері своєї, що народилися в домі або народилися назовні, не відкриєш їхньої наготи!
LEV|18|10|Наготу дочки сина свого або дочки дочки своєї, не відкриєш наготи їхньої, бо вони нагота твоя!
LEV|18|11|Наготи дочки жінки батька свого, народженої від батька твого, вона сестра твоя, не відкриєш наготи її!
LEV|18|12|Наготи сестри батька свого не відкриєш, вона однокровна батька твого!
LEV|18|13|Наготи сестри матері своєї не відкриєш, бо вона однокровна матері твоєї.
LEV|18|14|Наготи брата батька свого не відкриєш, до жінки його не наблизишся, вона тітка твоя!
LEV|18|15|Наготи невістки своєї не відкриєш, вона жінка сина твого, не відкриєш наготи її!
LEV|18|16|Наготи жінки брата свого не відкриєш, вона нагота брата твого!
LEV|18|17|Наготи жінки й дочки її не відкриєш; дочки сина її й дочки дочки її не візьмеш, щоб відкрити її наготу, вони однокровні її, це кровозмішання!
LEV|18|18|І жінки з сестрою її не візьмеш на суперництво, щоб відкрити наготу її при ній за життя її.
LEV|18|19|А до жінки в час відділення нечистости її не наблизишся, щоб відкрити наготу її.
LEV|18|20|А з жінкою свого ближнього не будеш лежати на насіння, щоб нею не стати нечистим.
LEV|18|21|А з насіння свого не даси на жертву Молохові, і не зневажиш Імени Бога свого. Я Господь!
LEV|18|22|А з чоловіком не будеш лежати як з жінкою, гидота воно!
LEV|18|23|І з жодною худобиною не зляжешся, щоб не стати нею нечистим. І жінка не стане перед худобиною на злягання, це паскудство!
LEV|18|24|Не занечищуйтеся тим усім, бо всім тим занечищені ті люди, яких Я виганяю перед вами.
LEV|18|25|І стала нечиста та земля, і Я полічив на ній її гріх, і та земля виригнула мешканців своїх!
LEV|18|26|І ви будете додержувати постанов Моїх та уставів Моїх, і не зробите жодної зо всіх тих гидот, як і тубілець чи приходько, що мешкає серед вас.
LEV|18|27|Бо всі ті гидоти робили люди тієї землі, які перед вами, і стала нечиста та земля.
LEV|18|28|І щоб та земля не виригнула вас через ваше занечищення її, як вона виригнула народ, який перед вами.
LEV|18|29|Бо кожен, хто зробить одну зо всіх тих гидот, то душі, що роблять, будуть винищені з-посеред їхнього народу.
LEV|18|30|І ви будете додержувати наказів Моїх, щоб не чинити чого з тих гидотних постанов, що роблені перед вами, і не споганитеся ними. Я Господь, Бог ваш!
LEV|19|1|І Господь промовляв до Мойсея, говорячи:
LEV|19|2|Промовляй до всієї громади Ізраїлевих синів, та й скажеш їм: Будьте святі, бо святий Я, Господь, Бог ваш!
LEV|19|3|Кожен буде боятися матері своєї та батька свого, а субіт Моїх будете додержувати. Я Господь, Бог ваш!
LEV|19|4|Не звертайтеся до ідолів, і не робіть собі литих божків. Я Господь Бог ваш!
LEV|19|5|А коли ви принесете мирну жертву для Господа, на вподобання вас принесете її.
LEV|19|6|Ви будете їсти її в день принесення вашого та взавтра, а позостале до дня третього огнем буде спалене.
LEV|19|7|А якщо справді буде їджене воно третього дня, нечистість воно, не буде вподобане.
LEV|19|8|А хто те їсть, понесе він свій гріх, бо споганив він святиню Господню, і буде винищена душа та з-посеред народу свого!
LEV|19|9|А коли ти будеш жати жниво своєї землі, не докінчуй жати до краю свого поля, а попадалих колосків твого жнива не будеш збирати;
LEV|19|10|а виноградника свого не вибереш дорешти, а попадалих ягід виноградника свого не будеш збирати, для вбогого та для приходька позостав їх. Я Господь, Бог ваш!
LEV|19|11|Не будете красти, і не будете неправдиво заперечувати, і не будете говорити неправди один на одного!
LEV|19|12|І не будете присягати Моїм Іменем на неправду, бо зневажиш Ім'я Бога свого. Я Господь!
LEV|19|13|Не будеш гнобити ближнього свого, і не будеш грабувати, і не задержиш в себе через ніч аж до ранку заробітку наймита.
LEV|19|14|Не будеш проклинати глухого, а перед сліпим не роби перешкоди, і будеш боятися Бога свого. Я Господь!
LEV|19|15|Не зробите кривди в суді: не будеш потурати особі вбогого, і не будеш підлещуватися до особи вельможного, за правдою суди свого ближнього!
LEV|19|16|Не будеш ходити пліткарем серед народу свого. Не будеш наставати на життя свого ближнього. Я Господь!
LEV|19|17|Не будеш ненавидіти брата свого в серці своєму. Конче вияви неправду свого ближнього, і не понесеш гріха за нього.
LEV|19|18|Не будеш мститися, і не будеш ненавидіти синів свого народу. І будеш любити ближнього свого, як самого себе! Я Господь!
LEV|19|19|Постанов Моїх будете дотримувати. Не зробиш, щоб худоба твоя злучувалася двоїсто. Поля свого не будеш обсівати двоїсто. А одежа двоїста, мішанина ниток, не ввійде на тебе.
LEV|19|20|А чоловік, коли буде злягатися з жінкою, а вона невільниця, заручена чоловікові, а справді не була вона викуплена, або визволення не було дане їй, то нехай буде кара, але не будуть вони забиті, бо не увільнена вона.
LEV|19|21|І спровадить він жертву за провину свою Господеві до входу скинії заповіту, барана жертви за провину.
LEV|19|22|І очистить його священик бараном жертви за провину перед Господнім лицем за гріх його, що він був згрішив. І проститься йому гріх його, що він був згрішив.
LEV|19|23|А коли ви ввійдете до Краю цього, і понасаджуєте всяке їстивне дерево, то плід його вважатимете за необрізаний, три роки буде воно для вас необрізане, не буде їджене.
LEV|19|24|А року четвертого ввесь плід його присвятиться для Господа.
LEV|19|25|А року п'ятого будете їсти плід його, щоб помножився для вас урожай його. Я Господь, Бог ваш.
LEV|19|26|Не будете їсти з кров'ю. Не будете ворожити, і не будете чарувати!
LEV|19|27|Не будете стригти волосся довкола голови вашої, і не будеш нищити краю бороди своєї.
LEV|19|28|І не зробите на тілі своїм нарізу за душу померлого, і не зробите на собі наколеного напису. Я Господь!
LEV|19|29|Не безчесть своєї дочки, і не роби її блудливою, щоб не стала блудливою ця земля, і не наповнилась земля розпустою.
LEV|19|30|Субіт Моїх будете додержувати, а святиню Мою будете шанувати. Я Господь!
LEV|19|31|Не звертайтесь до духів померлих та до ворожбитів, і не доводьте себе до опоганення ними. Я Господь, Бог ваш!
LEV|19|32|Перед лицем сивизни встань, і вшануй лице старого, і будеш боятися Бога свого. Я Господь!
LEV|19|33|А коли мешкатиме з тобою приходько в вашім Краї, то не будете гнобити його.
LEV|19|34|Як тубілець із вас буде для вас приходько, що мешкає з вами, і ти будеш любити його, як самого себе, бо приходьки були ви в єгипетськім краї. Я Господь, Бог ваш!
LEV|19|35|Не будете чинити кривди в суді, у мірі, у вазі та в мірі рідини.
LEV|19|36|Вага вірна, тягарці вірні, ефа вірна, гін вірний буде в вас. Я Господь, Бог ваш, що вивів вас із єгипетського краю!
LEV|19|37|І ви будете держати всі постанови Мої та всі устави Мої, і виконуватимете їх. Я Господь!
LEV|20|1|І Господь промовляв до Мойсея, говорячи:
LEV|20|2|І скажеш до Ізраїлевих синів: Кожен чоловік із Ізраїлевих синів та з приходька, що мешкає в Ізраїлі, який дасть із насіння свого Молохові, буде конче забитий, народ краю закидає його камінням.
LEV|20|3|А Я зверну лице Своє проти того чоловіка, і винищу його з-поміж народу його, бо з насіння свого дав він Молохові, щоб занечистити святиню Мою, збезчестити Моє святе Ймення.
LEV|20|4|А якщо справді люди того краю сховають свої очі від того чоловіка, коли він дасть із насіння свого Молохові, щоб не забити його,
LEV|20|5|то Я зверну Своє лице проти того чоловіка та проти родини його, і винищу його й усіх, що блудять за ним, блудячи за Молохом, з-посеред народу його.
LEV|20|6|А душа, що звертається до померлих духів та до чарівників, щоб блудити за ними, то Я зверну Своє лице проти тієї душі, і винищу того з-посеред народу його.
LEV|20|7|І ви будете освячуватися, і будьте святі, бо Я Господь, Бог ваш!
LEV|20|8|І ви будете держати постанови Мої, і будете виконувати їх. Я Господь, що освячує вас!
LEV|20|9|Бо кожен чоловік, що прокляне свого батька чи матір свою, буде конче забитий, батька свого чи матір свою він прокляв, кров його на ньому!
LEV|20|10|А кожен, хто буде чинити перелюб із чиєю жінкою, хто буде чинити перелюб із жінкою свого ближнього, буде конче забитий перелюбник та перелюбниця.
LEV|20|11|А хто буде лежати із жінкою батька свого, він відкрив наготу свого батька, будуть конче забиті обоє вони, кров їхня на них!
LEV|20|12|А хто буде лежати з невісткою своєю, будуть конче забиті обоє вони, гидоту вчинили вони, кров їхня на них!
LEV|20|13|А хто лежатиме з чоловіком як із жінкою, гидоту вчинили обоє вони, будуть конче забиті, кров їхня на них!
LEV|20|14|А хто візьме жінку й матір її, гидота це, в огні спалять його та її, і не буде кровозмішання серед вас!
LEV|20|15|А хто паруватиметься з скотиною, буде конче забитий, і скотину ту заб'єте.
LEV|20|16|А жінка, що наблизиться до якої скотини, щоб лежати з нею, то заб'єш ту жінку та скотину ту, будуть конче забиті вони, кров їхня на них!
LEV|20|17|А хто візьме сестру свою, дочку батька свого або дочку матері своєї, і побачить наготу її, а вона побачить наготу його, ганьба це! І будуть вони знищені на очах синів їхнього народу, він наготу сестри своєї відкрив, він понесе провину свою!
LEV|20|18|А хто буде лежати із жінкою, часу хвороби місячним, і відкриє її наготу, він джерело її обнажив, а вона відкрила джерело своєї крови, то будуть вони обоє знищені з-посеред народу свого!
LEV|20|19|І не відкриєш наготи сестри матері своєї й сестри батька свого, бо однокровну свою обнажив би ти, вони понесуть провину свою.
LEV|20|20|А хто буде лежати з тіткою своєю, він відкрив наготу дядька свого, гріх свій вони понесуть, бездітні помруть!
LEV|20|21|А хто візьме жінку брата свого, це нечисть, він відкрив наготу брата свого, бездітні будуть.
LEV|20|22|І ви будете додержувати всі постанови Мої й усі устави Мої, і будете виконувати їх, і не виригне вас земля та, куди Я впроваджаю вас, щоб сиділи ви в ній.
LEV|20|23|І не будете ви ходити за звичаями люду, що Я виганяю перед вами, бо все те робили вони, і Я їх обридив.
LEV|20|24|І сказав Я до вас: ви вспадкуєте їхню землю, а Я дам її вам на спадщину її, землю, що плине молоком та медом. Я Господь, Бог ваш, що відділив вас від тих народів!
LEV|20|25|І ви відділяйте між худобою чистою та нечистою, і між птаством нечистим та чистим, і не занечищуйте душ своїх худобою й птаством, і всім, що роїться на землі, що Я відділив для вас, як нечисте.
LEV|20|26|І будьте для мене святі, бо святий Я, Господь. І Я відділю вас від тих народів, щоб ви були Мої.
LEV|20|27|А чоловік або жінка, коли будуть вони викликати духа мерців або ворожити, будуть конче забиті, камінням закидають їх, кров їхня на них!
LEV|21|1|І сказав Господь до Мойсея: Говори до священиків, Ааронових синів, і скажеш їм: Ніхто з вас нехай не занечиститься через доторкнення до померлого серед свого народу.
LEV|21|2|Бо тільки через доторкнення до близьких однокровних своїх, через матір свою, і через батька свого, і через сина свого, і через дочку свою, і через брата свого,
LEV|21|3|і через сестру свою, дівчину близьку йому, що не була замужем, через тих він може занечиститися доторкненням.
LEV|21|4|Бувши одружений, нехай не занечиститься серед рідні своєї, щоб не збезчестити себе.
LEV|21|5|Не зроблять вони лисини на голові своїй, і краю бороди своєї не підстрижуть, а на тілі своїм не наріжуть надрізів.
LEV|21|6|Святі вони будуть для Бога свого, і не збезчестять вони Ймення Бога свого, бо вони приносять огняні Божі жертви, хліб свого Бога. І будуть вони святі.
LEV|21|7|Жінки блудливої та збезчещеної вони не візьмуть, і не візьмуть жінки, вигнаної від чоловіка свого, бо святий він для Бога свого.
LEV|21|8|І освятиш його, бо він приносить хліб Бога твого, святий він буде для вас, бо святий Я, Господь, що освячує вас!
LEV|21|9|А священикова дочка, коли зачне робити блуд, вона безчестить батька свого, ув огні буде спалена.
LEV|21|10|А священик, найбільший від братів своїх, що на голову його буде виллята олива помазання, і буде посвячений на одягання шат, він голови своєї не запустить і шат своїх не роздере,
LEV|21|11|і до жодного вмерлого не ввійде, навіть через батька свого та через матір свою не сміє занечиститься.
LEV|21|12|І він не відійде від святині, і не занечистить святині Бога свого, бо на ньому посвячення оливи помазання його Бога. Я Господь!
LEV|21|13|І він візьме жінку в дівоцтві її.
LEV|21|14|Удови, і розведеної, і збезчещеної, блудливої, тих він не візьме, а тільки дівицю з-поміж рідні своєї він візьме за жінку.
LEV|21|15|І не збезчестить він насіння свого в рідні своїй, бо Я Господь, що освячує його.
LEV|21|16|І Господь промовляв до Мойсея, говорячи:
LEV|21|17|Промовляй до Аарона, говорячи: Чоловік із насіння твого на їх покоління, що буде в нім вада, не приступить, щоб приносити хліб свого Бога.
LEV|21|18|Бо жоден чоловік, що в нім вада, не приступить: чоловік сліпий, або кульгавий, або кирпатий або довготелесий,
LEV|21|19|або чоловік, що матиме зламану ногу або зламану руку,
LEV|21|20|або горбатий, або висохлий, або більмо на оці його, або коростявий, або паршивий, або з розчавленими ядрами,
LEV|21|21|кожен чоловік із насіння священика Аарона, що на нім ця вада, не приступить, щоб приносити Господні огняні жертви, вада в нім, не приступить він, щоб приносити хліб свого Бога.
LEV|21|22|Він буде їсти хліб свого Бога з Найсвятішого та зо святощів.
LEV|21|23|Та до завіси не підійде він, і до жертівника не приступить, бо вада в нім, і не збезчестить святині Моєї, бо Я Господь, що освячує їх.
LEV|21|24|І Мойсей промовляв до Аарона й до синів його, та до всіх синів Ізраїлевих.
LEV|22|1|І Господь промовляв до Мойсея, говорячи:
LEV|22|2|Промовляй до Аарона й до синів його, і нехай вони обережно поводяться зо святощами Ізраїлевих синів, які вони посвячують Мені, і нехай не безчестять Мого святого Ймення. Я Господь!
LEV|22|3|Скажи їм: На ваші покоління кожен чоловік, що наблизиться зо всякого вашого насіння до святощів, які Ізраїлеві сини посвятять Господеві, а нечистість його на нім, то буде винищена душа та з-перед лиця Мого. Я Господь!
LEV|22|4|Кожен чоловік з Ааронового насіння, коли він прокажений або течивий, не буде їсти зо святощів, аж поки очиститься. А хто доторкнеться всякого нечистого від мертвого тіла, або чоловік, що з нього вийде насіння лежання,
LEV|22|5|або хто доторкнеться до всякого плазуна, через якого він стане нечистий, або до людини, через яку стане нечистий, через усяку нечистість її,
LEV|22|6|особа, що доторкнеться до того, то стане нечиста аж до вечора, і не буде їсти зо святощів, поки не обмиє свого тіла в воді.
LEV|22|7|А коли зайде сонце, то стане він чистий, а потім буде їсти зо святощів, бо це хліб його.
LEV|22|8|Падла та розшарпаного не буде він їсти, щоб не занечиститись ним. Я Господь!
LEV|22|9|І будуть вони стерегти Мої прикази, щоб не понести через те гріха на собі, і щоб не померти через нього, коли б збезчестили їх. Я Господь, що освячує їх!
LEV|22|10|А кожен чужий не буде їсти святощів; осілий у священика й наймит не будуть їсти святощів.
LEV|22|11|А коли священик купить чоловіка, купівля срібла його це, той буде їсти їх, також уроджений дому його, вони будуть їсти його хліб.
LEV|22|12|А священикова дочка, коли буде видана чужому чоловікові, вона не буде їсти принесених святощів.
LEV|22|13|А священикова дочка, коли буде вдова, або розведена, а дітей не має, і вернеться до дому свого батька, як за молодости своєї, буде їсти з хліба батька свого. А кожен чужий не буде їсти його.
LEV|22|14|А чоловік, коли з'їсть святощі через помилку, то докладе до неї п'яту частину її, і віддасть священикові ті святощі,
LEV|22|15|і священики не збезчестять святощів Ізраїлевих синів, що вони приносять Господеві,
LEV|22|16|і не стягнуть на себе вини за провину їдження своїх святощів. Бо Я Господь, що освячує їх.
LEV|22|17|І промовляв Господь до Мойсея, говорячи:
LEV|22|18|Промовляй до Аарона й до синів його, та до всіх Ізраїлевих синів, і скажеш їм: Кожен чоловік з Ізраїлевого дому та з приходька між Ізраїлем, що принесе свою жертву за всякими своїми обітницями та за всякими даруваннями своїми, що принесе Господеві на цілопалення,
LEV|22|19|то нехай принесе на вподобання ваше безвадного самця з худоби великої, з овець і з кіз.
LEV|22|20|Жодного, що в нім вада, не принесете, бо не буде воно на вподобання вас.
LEV|22|21|А чоловік, коли принесе Господеві мирну жертву на виразно висловлену обітницю або на дарунок, із худоби великої чи з худоби дрібної, безвадна буде на вподобання, жодна вада не буде в ній:
LEV|22|22|сліпа, або зламана, або скалічена, або шолудива, або коростява, або паршива, не принесете тих Господеві, і жертви огняної не дасте з них на жертівника для Господа.
LEV|22|23|А вола та вівцю з занадто довгим чи занадто коротким яким членом добровільно принесеш у жертву, а на обітницю вони не вгодні Богові.
LEV|22|24|А того, що має ядра розчавлені, чи збиті, чи відірвані, чи відрізані не піднесете Господеві, і в вашому Краї не зробите того.
LEV|22|25|І з руки чужинця не принесете хліба нашого Бога зо всіх таких, бо в них зіпсуття їх, вада в них, вони не будуть вгодні для вас.
LEV|22|26|І Господь промовляв до Мойсея, говорячи:
LEV|22|27|Віл, або вівця, або коза, коли вродиться, то буде сім день під своєю матір'ю, а від дня восьмого й далі буде вгодне на жертву огняну для Господа.
LEV|22|28|А корови та вівці, її й маля її не заріжете одного дня.
LEV|22|29|А коли будете приносити вдячну жертву для Господа, то приносьте так, щоб вона була вгодна.
LEV|22|30|Того дня буде вона з'їджена, не зоставите з неї аж до ранку. Я Господь!
LEV|22|31|І заповіді Мої будете додержувати, і будете виконувати їх. Я Господь!
LEV|22|32|І не будете безчестити Мого святого Ймення, і Я буду освячений серед Ізраїлевих синів. Я Господь, що освячує вас,
LEV|22|33|що вивів вас із єгипетського краю, щоб бути вашим Богом. Я Господь!
LEV|23|1|І Господь промовляв до Мойсея, говорячи:
LEV|23|2|Промовляй до Ізраїлевих синів і скажеш їм: Свята Господні, що в них скликатимете святі збори, оце вони, свята Мої:
LEV|23|3|Шість день буде робитись робота, а дня сьомого субота повного відпочинку, святі збори, жодної роботи не будете робити. Це субота відпочинку для Господа по всіх оселях ваших!
LEV|23|4|Оце свята Господні, святі збори, що скличете їх у їхнім означенім часі:
LEV|23|5|У місяці першім, чотирнадцятого дня місяця під вечір Пасха для Господа.
LEV|23|6|А п'ятнадцятого дня того місяця свято Опрісноків для Господа, сім день будете їсти опрісноки.
LEV|23|7|Першого дня будуть святі збори для вас, жодного робочого зайняття не будете робити.
LEV|23|8|І будете приносити для Господа жертву сім день; сьомого дня збори святі, жодного робочого зайняття не будете робити.
LEV|23|9|І Господь промовляв до Мойсея, говорячи:
LEV|23|10|Промов до Ізраїлевих синів і скажеш їм: Коли ви ввійдете до того Краю, що Я даю вам, і будете жати жниво його, то снопа первоплоду ваших жнив принесете до священика,
LEV|23|11|а він буде колихати снопа того перед лицем Господнім, щоб набути вподобання вам; першого дня по святі священик буде колихати його.
LEV|23|12|І ви прирядите в дні вашого колихання снопа однорічне безвадне ягня на цілопалення для Господа.
LEV|23|13|А хлібна його жертва дві десяті ефи пшеничної муки, мішаної в оливі, огняна жертва для Господа, пахощі любі; а жертва лита його вино, чверть гіна.
LEV|23|14|А хліба, і пряженого зерна, і свіжих зерен ви не будете їсти аж до самого того дня, аж до вашого принесення жертви для вашого Бога. Це вічна постанова для ваших поколінь по всіх ваших оселях.
LEV|23|15|І відлічите ви собі першого дня по святі, від дня вашого принесення снопа колихання, сім тижнів, повні будуть вони.
LEV|23|16|А до першого дня по сьомім тижні відлічите п'ятдесят днів, та й принесете хлібну нову жертву для Господа.
LEV|23|17|З ваших осель принесете два хліби колихання, дві десяті ефи пшеничної муки будуть вони, будуть спечені квашені, первоплоди для Господа.
LEV|23|18|І принесете понад той хліб сім ягнят безвадних у віці року, й одного бичка та два барани, вони будуть цілопалення для Господа, і жертва хлібна, і жертви литі для них, огняна жертва, пахощі любі для Господа.
LEV|23|19|І спорядите одного козла на жертву за гріх, та двоє ягнят у віці року на жертву мирну.
LEV|23|20|І священик буде колихати їх разом із хлібом первоплодів, як колихання перед Господнім лицем, над двома ягнятами. Вони будуть святощі для Господа, для священика.
LEV|23|21|І скличете того самого дня, і будуть святі збори для вас, жодного робочого зайняття не будете робити. Це вічна постанова для ваших поколінь по всіх ваших оселях!
LEV|23|22|А коли ви будете жати жниво вашої землі, не дожинай краю поля твого, а попадалих колосків жнива твого не будеш збирати, для вбогого та для приходька позоставиш їх. Я Господь, Бог ваш!
LEV|23|23|І промовив Господь до Мойсея, говорячи:
LEV|23|24|Промовляй до Ізраїлевих синів, говорячи: Сьомого місяця, першого дня місяця буде вам повний спочинок, пам'ять сурмлення, святі збори.
LEV|23|25|Жодного робочого зайняття не будете робити, і принесете огняну жертву для Господа.
LEV|23|26|І Господь промовляв до Мойсея, говорячи:
LEV|23|27|А десятого дня самого місяця день Очищення він, збори святі будуть для вас, і будете впокоряти душі ваші, і принесете огняну жертву для Господа.
LEV|23|28|І жодного зайняття не будете робити того самого дня, бо він день Очищення, щоб очистити за вас перед лицем Господа, Бога вашого.
LEV|23|29|Бо кожна душа, що не буде впокорюватись того самого дня, то буде вона винищена з своєї рідні.
LEV|23|30|А кожна душа, що буде робити яке зайняття того самого дня, то Я вигублю ту душу з-посеред народу її.
LEV|23|31|Жодного зайняття не будете робити. Це постанова вічна для ваших поколінь по всіх ваших оселях!
LEV|23|32|Він субота повного спочинку для вас, і ви будете впокоряти душі свої, ввечері дев'ятого дня місяця від вечора аж до вечора будете святкувати вашу суботу.
LEV|23|33|І Господь промовляв до Мойсея, говорячи:
LEV|23|34|Промовляй до Ізраїлевих синів, кажучи: П'ятнадцятого дня того сьомого місяця, свято Кучок, сім день для Господа.
LEV|23|35|Першого дня святі збори, жодного робочого зайняття не будете робити.
LEV|23|36|Сім день будете приносити огняну жертву для Господа; восьмого дня святі збори будуть для вас, і принесете огняну жертву для Господа; це віддання свята, жодного робочого зайняття не будете робити.
LEV|23|37|Оце свята Господні, що скликуватимете на них святі збори, щоб приносити огняну жертву для Господа, цілопалення, хлібну жертву й заколену жертву, і жертви литі, належне дневі в його дні,
LEV|23|38|окрім Господніх субіт, і окрім дарів ваших, і окрім усіх ваших обітниць, і окрім усіх ваших дарувань, що дасте Господеві.
LEV|23|39|А п'ятнадцятого дня сьомого місяця, коли ви збираєте врожай землі, будете святкувати свято Господнє сім день; першого дня повний спочинок, і восьмого повний спочинок.
LEV|23|40|І візьмете собі першого дня плоду гарного дерева, пальмові віття, і галузку многолистого дерева та припоточних тополь, і будете веселитися перед лицем Господа, Бога вашого, сім день.
LEV|23|41|І будете святкувати його, як свято для Господа, сім день у році. Постанова вічна для ваших поколінь, сьомого місяця будете святкувати його.
LEV|23|42|У кучках будете сидіти сім день, кожен тубілець в Ізраїлі сидітиме в кучках,
LEV|23|43|щоб ваші покоління пізнали що Я в кучках посадив був Ізраїлевих синів, коли виводив їх з єгипетського краю. Я Господь, Бог ваш!
LEV|23|44|І Мойсей промовляв до Ізраїлевих синів про свята Господні.
LEV|24|1|І Господь промовляв до Мойсея, говорячи:
LEV|24|2|Накажи Ізраїлевим синам, і вони принесуть тобі чистої, вичавленої оливи з оливкового дерева на освітлення, щоб запалювати вічну лямпаду.
LEV|24|3|Поза завісою свідоцтва в скинії заповіту прирядить її Аарон від вечора аж до ранку перед Господнім лицем назавжди. Це вічна постанова для ваших поколінь!
LEV|24|4|На чистім свічнику прирядить він ті лямпади перед Господнім лицем назавжди.
LEV|24|5|І візьмеш пшеничної муки, і випечеш із неї дванадцять калачів, по дві десяті ефи буде один калач.
LEV|24|6|І покладеш їх у два ряди, шість у ряд, на чистому столі перед Господнім лицем,
LEV|24|7|і поклади на ряд чистого ладану, і він стане для хліба за пригадувальну частину, огняна жертва для Господа.
LEV|24|8|Щосуботи він покладе його перед Господнім лицем завжди, від Ізраїлевих синів, вічний заповіт.
LEV|24|9|І він буде для Аарона та для синів його, і вони будуть їсти його в святому місці, бо він найсвятіше з огняних жертов Господніх. Це вічна постанова.
LEV|24|10|І вийшов син ізраїльтянки, а він був син єгиптянина, між Ізраїлевих синів. І сварився в таборі син тієї ізраїльтянки з одним ізраїльтянином.
LEV|24|11|І син тієї ізраїльтянки богозневажив Ім'я Господнє, і проклинав. І привели його до Мойсея. А ймення матері його Шеломіт, дочка Діври, з Данового племени.
LEV|24|12|І посадили його під сторожу аж до вияснення через уста Господні.
LEV|24|13|І Господь промовляв до Мойсея, говорячи:
LEV|24|14|Виведи того, що проклинав, поза табір, і покладуть усі, хто чув, свої руки на голову його, і закидає його камінням уся громада.
LEV|24|15|А до Ізраїлевих синів будеш промовляти, говорячи: Кожен чоловік, коли прокляне Бога свого, то понесе він свій гріх.
LEV|24|16|А той, хто богозневажив Господнє Ймення, буде конче забитий, конче укаменує його вся громада; чи приходько, чи тубілець, коли богозневажатиме Ймення Господнє, буде забитий.
LEV|24|17|І кожен, хто заб'є людину, буде конче забитий.
LEV|24|18|А хто заб'є яку скотину, той відшкодує її, життя за життя.
LEV|24|19|І кожен, коли зробить ваду своєму ближньому, як хто зробив, так буде зроблено йому:
LEV|24|20|зламання за зламання, око за око, зуб за зуба, яку ваду зробить хто кому, така буде зроблена йому.
LEV|24|21|А хто заб'є скотину, той відшкодує її, а хто заб'є людину, той буде забитий.
LEV|24|22|Суд один буде для вас, приходько буде як тубілець. Бо Я Господь Бог ваш!
LEV|24|23|І Мойсей промовляв до Ізраїлевих синів. І вони вивели того, хто проклинав, поза табір, та й закидали його камінням. І зробили Ізраїлеві сини, як Господь наказав був Мойсеєві.
LEV|25|1|І Господь промовляв до Мойсея на Сінайській горі, говорячи:
LEV|25|2|Промовляй до Ізраїлевих синів, та й скажеш їм: Коли ви ввійдете до землі, що Я даю вам, то святкуватиме земля та суботу для Господа.
LEV|25|3|Шість літ будеш засівати своє поле, і шість літ обтинатимеш свого виноградника, і збиратимеш урожай його,
LEV|25|4|а сьомого року субота повного відпочинку буде для землі, повний відпочинок, субота для Господа: поля свого не будеш обсіювати, а виноградника свого не будеш обтинати.
LEV|25|5|Саморослого колосу жнив твоїх не будеш жати, а ґрон з необрізаних виноградин твоїх не збиратимеш, рік повного відпочинку буде для землі.
LEV|25|6|І те, що саме вродиться в цім відпочинку землі, буде для вас на їжу, для тебе, і для раба твого, і для невільниці твоєї, і для наємника твого, і для осілого твого, що мешкають з тобою,
LEV|25|7|і для скотини твоєї, і для звірини, що в Краї твоїм, буде ввесь урожай його на їжу.
LEV|25|8|І відлічиш собі сім суботніх років, по сім років сім раз, і будуть для тебе дні семи суботніх років сорок літ і дев'ять.
LEV|25|9|І засурмите у сурми сьомого місяця, десятого дня місяця, в день Очищення засурмите в сурми по цілому Краю.
LEV|25|10|І освятите рік п'ятдесятріччя, і оголосите волю в Краю для всіх мешканців його, ювілей він буде для вас: і вернеться кожен до своєї посілости, і кожен до родини своєї вернеться.
LEV|25|11|Ювілей цей рік п'ятдесятріччя буде для вас: на будете сіяти, і не будете жати саморослі колосся її, і не будете збирати грон з необрізаних виноградин їх,
LEV|25|12|бо це ювілей, святощі будуть для вас, з поля будете їсти врожай його.
LEV|25|13|У році того ювілею вернетесь кожен до своєї посілости.
LEV|25|14|А коли продасте що своєму ближньому, або купите з руки свого ближнього, не обманюйте один одного.
LEV|25|15|За числом років по ювілеї купиш від ближнього свого, за числом років урожаю він продасть тобі.
LEV|25|16|За многістю літ побільшиш ціну тієї купівлі, а за малістю літ зменшиш ціну тієї купівлі, бо він продає тобі число літ урожаю.
LEV|25|17|І не обманите один одного, і будеш боятися Бога свого, бо Я Господь, Бог ваш!
LEV|25|18|І ви виконаєте постанови Мої, а устави Мої будете держати, і будете виконувати їх, і безпечно сидітимете на землі.
LEV|25|19|І земля дасть плід свій, а ви будете їсти досита, і безпечно сидітимете на ній.
LEV|25|20|А коли ви скажете: Що будемо їсти сьомого року, тож не будемо сіяти, не будемо збирати врожаї свої?
LEV|25|21|І зошлю Я благословення Своє на вас шостого року, і зродить врожай на три роки.
LEV|25|22|І будете сіяти восьмий той рік, і будете їсти з старих урожаїв аж до року дев'ятого, аж до виросту врожаю його будете їсти старе.
LEV|25|23|А земля не буде продаватися назавжди, бо Моя та земля, бо ви приходьки та осілі в Мене.
LEV|25|24|А ви в усій землі вашої посілости дозволяйте викуп землі.
LEV|25|25|Коли збідніє твій брат, і продасть із своєї посілости, то прийде викупник його, близький йому, і викупить продаж брата свого.
LEV|25|26|А чоловік, коли не буде йому викупника, а рука його стане спроможна, і знайде потрібне на викуп його,
LEV|25|27|то облічить він літа продажу свого, і верне позостале чоловікові, що продав йому, та й вернеться до своєї посілости.
LEV|25|28|А якщо рука його не знайде потрібного на заплату йому, то буде продаж його в руці покупця його аж до ювілейного року, і вийде він в ювілеї, та й вернеться до посілости своєї.
LEV|25|29|А коли хто продасть мешкальний дім в обмурованому місті, то викуп його буде до кінця року від часу продажу його, рік буде на викуп його.
LEV|25|30|А якщо він не буде викуплений аж до кінця року, то стане той дім, що в місті, яке має мур, назавжди для покупця його на покоління його, не вийде він в ювілеї.
LEV|25|31|А доми в оселях, що не мають муру навколо, до поля землі буде те прираховане, і буде йому викуп, і в ювілеї він вийде.
LEV|25|32|А міста Левитів, доми в містах їх посілости викуп для Левитів завжди буде можливий.
LEV|25|33|А хто викупить від Левитів, то продаж дому й міста посілости його вийде в ювілеї, бо то доми міст Левитів, їхня посілість серед Ізраїлевих синів.
LEV|25|34|А пасовисько навколо їхніх міст не буде продане, бо це вічна посілість для них.
LEV|25|35|А коли збідніє твій брат, а його рука неспроможною стане, то підтримаєш його, приходько він чи осілий, і житиме він із тобою.
LEV|25|36|Не візьмеш від нього лихви та прибутку, і будеш боятися Бога свого, і житиме брат твій з тобою.
LEV|25|37|Срібла свого не даси йому на лихву, і на прибуток не даси їжі своєї.
LEV|25|38|Я Господь, Бог ваш, що вивів вас із єгипетського краю, щоб дати вам ханаанську землю, щоб бути вашим Богом.
LEV|25|39|А коли збідніє брат твій при тобі, і буде проданий тобі, то не будеш робити ним праці раба,
LEV|25|40|як наймит, як осілий він при тобі, аж до ювілейного року буде він працювати тобі.
LEV|25|41|вийде від тебе він та сини його з ним, і вернеться він до родини своєї, і до посілости батьків своїх вернеться він:
LEV|25|42|бо вони Мої раби, що Я вивів їх з єгипетського краю, не будуть вони продані продажем раба.
LEV|25|43|Не будеш володіти ним жорстоко, і будеш боятися Бога свого.
LEV|25|44|А раб твій та невільниця твоя, що будуть твої, будуть із народів, що навколо вас, із них купите раба й невільницю.
LEV|25|45|А також із синів осілих, що мешкають з вами, з них купите та з племені їхнього, що з вами, що породили в Краї вашім, і будуть вони вам на посілість.
LEV|25|46|І передасте їх, як спадщину, вашим синам по вас на спадок посілости навіки, ними будете робити, а братами вашими, синами Ізраїлевими, один одним, не будете володіти жорстоко.
LEV|25|47|А коли рука приходька чи осілого при тобі спроможна, а брат твій збідніє при ньому, і буде проданий приходькові чи осілому в тебе, або нащадкові племени приходька,
LEV|25|48|то потім, як буде проданий, викуп буде йому, один із братів його викупить його,
LEV|25|49|або дядько його, або син дядька його викупить його, або з однокровних його, із роду його викупить його, або спроможна рука його, і буде викуплений.
LEV|25|50|І облічить він із тим, хто набув його, від року продажу його аж до ювілейного року, і буде ціна продажу його за числом літ; як за дні наймита буде полічено йому.
LEV|25|51|Якщо ще багато літ, то згідно з ними він верне свій викуп із срібла його купівлі.
LEV|25|52|А якщо позостало мало літ до ювілейного року, то облічить йому, згідно з роками його верне свого викупа.
LEV|25|53|Як щорічнии наймит він буде при ньому, він не буде жорстоко панувати над ним на твоїх очах.
LEV|25|54|А якщо він не буде викуплений у тих роках, то вийде ювілейного року він та сини його з ним,
LEV|25|55|бо Ізраїлеві сини Мої раби, Мої раби вони, що Я вивів їх із єгипетського краю. Я Господь, Бог ваш!
LEV|26|1|Не зробите собі божків та ідола, і кам'яного стовпа не поставите собі, і каменя з фіґурами не покладете в вашім Краї, щоб кланятися перед ними. Бо Я Господь, Бог ваш!
LEV|26|2|Субіт Моїх будете додержувати, а святиню Мою будете шанувати. Я Господь!
LEV|26|3|Якщо будете ходити згідно з постановами Моїми, а заповідей Моїх будете додержувати й будете виконувати їх,
LEV|26|4|то дам ваші дощі в їхнім часі, і земля дасть свій урожай, а польове дерево дасть плід свій.
LEV|26|5|І молочення досягне вам виноградобрання, а виноградобрання досягне сіяння, і ви будете їсти хліб свій досита, і будете сидіти безпечно в вашому Краї.
LEV|26|6|І дам мир у Краю, і ви будете лежати, і ніхто не вчинить, щоб ви тремтіли, бо злу звірину винищу з землі, а меч не перейде через Край ваш.
LEV|26|7|І ви будете гнати ворогів своїх, а вони попадають перед вами від меча.
LEV|26|8|І п'ятеро з вас поженуть сотню, а сотня з вас пожене десять тисяч, і попадають вороги ваші перед вами від меча.
LEV|26|9|І обернусь Я до вас, і розплоджу вас, і розмножу вас, і виконаю Свого заповіта з вами.
LEV|26|10|І ви будете їсти старе-перестаріле, і повикидаєте старе перед новим.
LEV|26|11|І поставлю місце перебування Свого серед вас, і душа Моя не обридить вами.
LEV|26|12|І Я буду ходити серед вас, і буду вам Богом, а ви будете Мені народом.
LEV|26|13|Я Господь, Бог ваш, що вивів вас з єгипетського краю, щоб ви не були їм рабами. І Я поламав занози вашого ярма, і вивів вас із піднесеною головою.
LEV|26|14|А коли ви не будете слухняні Мені, і не виконуватиме всіх тих заповідей,
LEV|26|15|і якщо постановами Моїми будете погорджувати, і якщо душа ваша бридитиметься законами Моїми, щоб не виконувати всіх заповідей Моїх, щоб ламати вам заповіта Мого,
LEV|26|16|то й Я зроблю вам оце: поставлю над вами перестрах, сухоти й пропасницю, що винищують очі й обезсилюють душу. І ви надаремно сіятимете насіння своє, бо поїдять його вороги ваші.
LEV|26|17|І зверну Я лице Своє на вас, і ви будете вдарені перед своїми ворогами. І будуть панувати над вами ненависники ваші, і ви будете втікати, хоч ніхто вас не гнатиме.
LEV|26|18|А якщо й при тому не будете слухняні Мені, то Я семикратно побільшу кару на вас за ваші гріхи.
LEV|26|19|І зломлю пиху вашої сили, і зроблю ваше небо як залізо, а землю вашу як мідь!
LEV|26|20|І надаремно буде вичерпуватися ваша сила: земля ваша не дасть свого врожаю, а дерево на землі не дасть свого плоду.
LEV|26|21|А якщо й тоді підете проти Мене, і не схочете бути слухняними Мені, то Я семикратно збільшу над вами удара Свого згідно з вашими гріхами.
LEV|26|22|І пошлю на вас пільну звірину, а вона винищить вам дітей, і вигубить вашу худобу, і зменшить кількість вашу, і попустошить ваші дороги.
LEV|26|23|А якщо цими карами не будете навчені, і будете ходити проти Мене,
LEV|26|24|то й Я піду проти вас, і вдарю вас і Я семикратно за ваші гріхи.
LEV|26|25|І приведу на вас меча, що помстить пімсту за заповіта, і ви будете зібрані до ваших міст, і Я пошлю моровицю на вас, і ви будете віддані в руку ворога.
LEV|26|26|Коли Я знищу вам хліб, підпору вашу, то десять жінок будуть пекти хліб вам в одній печі, і вернуть хліб ваш вагою, а ви будете їсти і не насититеся.
LEV|26|27|А якщо й тим не станете слухняні Мені, і будете ходити проти Мене,
LEV|26|28|то й Я з лютістю піду проти вас, і також Я семикратно покараю вас за ваші гріхи,
LEV|26|29|і ви тіло своїх синів будете їсти, і тіло дочок своїх будете поїдати...
LEV|26|30|І поруйную ваші висоти, і повитинаю ваші стовпи сонця, і поскладаю трупи ваші на трупах божків ваших, і обридить душа Моя вас!
LEV|26|31|І вчиню міста ваші руїною, і поспустошую ваші святині, і не прийму ваших пахощів любих.
LEV|26|32|І спустошу Я Край той, і будуть дивуватися з того ваші вороги, що мешкають у ньому.
LEV|26|33|А вас порозпорошую поміж народів, і вийму за вами меча, і стане Край ваш спустошенням, а міста ваші будуть руїною...
LEV|26|34|Тоді земля та надолужить собі за суботні роки по всі дні спустошення її. Коли будете в краї ваших ворогів, тоді ваша земля святкуватиме відпочинок, і надолужить собі за свої суботні роки.
LEV|26|35|По всі дні спустошення святкуватиме вона відпочинок, чого не святкувала в суботні роки, коли ви сиділи на ній.
LEV|26|36|А щодо позосталих серед вас, то впроваджу в їхні серця полохливість в краях їхніх ворогів, і буде їх гнати навіть шелест подмухненого вітром листу, і будуть вони втікати, як утікають перед мечем, та й попадають, хоч ніхто не женеться...
LEV|26|37|І будуть вони спотикатися один об одного, ніби від меча, хоч ніхто не женеться за ними. І ви не зможете стати проти ваших ворогів...
LEV|26|38|І погинете серед поганів, і пожере вас земля ваших ворогів.
LEV|26|39|А позосталі серед вас помарніють у краях ворогів ваших за гріх свій, а також за гріхи батьків своїх помарніють із ними.
LEV|26|40|І визнають вони гріх свій та гріх батьків своїх, що ними спроневірилися були Мені, а також, що ходили проти Мене.
LEV|26|41|Також і Я піду проти них, і впроваджу їх до краю їхніх ворогів. Якщо тоді впокориться їхне необрізане серце, то тоді понесуть кару за свої гріхи.
LEV|26|42|І Я згадаю заповіта Свого з Яковом, а також заповіта Свого з Ісаком, і також заповіта Свого з Авраамом згадаю, і згадаю той Край.
LEV|26|43|А Край той буде позбавлений їх, і надолужить собі свої суботні роки, опустілий від них, а вони понесуть кару за свої гріхи, а то для того, що законами Моїми погорджували, а постанови Мої огидила була їхня душа.
LEV|26|44|А проте, коли вони пробували в краю своїх ворогів, то Я не погорджував ними, і не збридив їх, щоб винищити їх, щоб зламати заповіта Свого з ними. Бо Я Господь, Бог їх!
LEV|26|45|І Я пам'ятатиму їм заповіта з предками, що Я вивів їх з єгипетського краю на очах поган, щоб бути їм Богом. Я Господь!
LEV|26|46|Оце постанови, і устави та закони, що дав Господь між Собою та між Ізраїлевими синами на Сінайскій горі через Мойсея.
LEV|27|1|І Господь промовляв до Мойсея, говорячи:
LEV|27|2|Промовляй до Ізраїлевих синів та й скажеш їм: Коли хто складає обітницю Богові за твоєю оцінкою душ для Господа,
LEV|27|3|то буде твоя оцінка: чоловіка від віку двадцяти літ і аж до віку шостидесяти літ, і буде твоя оцінка п'ятдесят шеклів срібла на міру шеклем святині;
LEV|27|4|а якщо жінка вона, то буде твоя оцінка тридцять шеклів.
LEV|27|5|А якщо від віку п'яти літ і до віку двадцяти літ, то буде твоя оцінка: чоловіка двадцять шеклів, а для жінки десять шеклів.
LEV|27|6|А якщо від віку місяця й аж до віку п'яти літ, то буде твоя оцінка: чоловіка п'ять шеклів срібла, а для жінки твоя оцінка три шеклі срібла.
LEV|27|7|А якщо від віку шостидесяти літ і вище: якщо чоловік, то буде твоя оцінка п'ятнадцять шеклів, а для жінки десять шеклів.
LEV|27|8|А якщо він обіднілий проти твоєї оцінки, то поставить його перед священиком, і священик оцінує його, за тим, що спроможна рука того, хто обіцяв, оцінує його священик.
LEV|27|9|А якщо буде худоба, що з неї приносять жертву для Господа, усе, що дається із неї для Господа, буде святощами.
LEV|27|10|Не вільно обміняти її, ані заступити її, добру злою, або злу доброю; а якщо справді заступить худобу худобою, то буде вона та заступство її буде святощами.
LEV|27|11|А якщо та всяка худоба нечиста, що з неї не приносять жертов для Господа, то він поставить ту худобу перед священиком,
LEV|27|12|і священик оцінує її чи то добре, чи недобре. Як оцінує священик, так нехай буде.
LEV|27|13|А якщо він справді викупить її, то додасть п'яту частину її над оцінку твою.
LEV|27|14|А коли хто посвятить дім свій на святість для Господа, то священик оцінує його чи то добре, чи недобре. Як оцінує його священик, так стане.
LEV|27|15|А якщо той, хто посвячує, викупить свого дома, то додасть п'яту частину срібла твоєї оцінки над нього, і буде його.
LEV|27|16|А якщо хтось посвятить Господеві з поля своєї посілости, то буде оцінка твоя посівом його, посів хомера ячменю за п'ятдесят шеклів срібла.
LEV|27|17|Якщо він посвятить своє поле від ювілейного року, то воно стане за оцінкою твоєю.
LEV|27|18|А якщо посвятить поле своє по ювілеї, то священик облічить йому те срібло за роками, позосталими до ювілейного року, і те буде відняте від оцінки твоєї.
LEV|27|19|А якщо справді викупить те поле той, хто посвячує його, то додасть п'яту частину срібла оцінки над нього, і стане воно його.
LEV|27|20|А якщо він не викупить поля того, і якщо він продасть те поле кому іншому, то вже не буде воно викуплене.
LEV|27|21|І буде те поле, коли воно вийде в ювілеї, святість для Господа, як поле закляття, для священика буде посілість ним.
LEV|27|22|А якщо він посвятить Господеві поле купівлі своєї, що не з поля посілости його,
LEV|27|23|то священик облічить йому суму твоєї оцінки аж до ювілейного року, і дасть твою оцінку того дня, як святість для Господа.
LEV|27|24|В ювілейному році вернеться те поле до того, від кого купив його, що його посілість тієї землі.
LEV|27|25|А вся оцінка твоя буде шеклем святині, двадцять ґер буде шекель.
LEV|27|26|Тільки перворідного в худобі, що визнане, як перворідне для Господа, ніхто не посвятить його, чи то віл, чи то овечка, Господеві воно!
LEV|27|27|А якщо в худобі нечистій, то викупить за твоєю оцінкою, і додасть п'яту частину над нього. А якщо не буде викуплене, то буде продане за оцінкою твоєю.
LEV|27|28|Тільки кожне закляття, що людина заклене Господеві зо всього, що його, від людини, і худоби, і від поля його посілости, не буде продане й не буде викуплене, воно найсвятіше для Господа.
LEV|27|29|Кожне закляття, що буде оголошене за закляття з-посеред людей, не буде викуплене, буде конче забите.
LEV|27|30|А всяка десятина з землі, з насіння землі, з плоду дерева, Господеві воно, святощі для Господа!
LEV|27|31|А якщо дійсно викупить хтось свою десятину, той додасть п'яту частину її над неї.
LEV|27|32|А всяка десятина худоби великої та худоби дрібної, усе, що перейде під палицею, десяте буде святість для Господа.
LEV|27|33|Не буде перебирати між добрим та злим, і не замінить його. А якщо справді заступить його, то буде воно та заступство його, буде святість, не буде викуплене.
LEV|27|34|Оце заповіді, що Господь наказав Мойсеєві для Ізраїлевих синів на Сінайській горі.
