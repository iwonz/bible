ROM|1|1|基督耶穌的僕人 保羅 ，蒙召為使徒，奉派傳上帝的福音。
ROM|1|2|這福音是上帝從前藉眾先知，在聖經上所應許的。
ROM|1|3|論到他兒子－我主耶穌基督，按肉體說，是從 大衛 後裔生的；按神聖的靈說，因從死人中復活，用大能顯明他是上帝的兒子。
ROM|1|4|
ROM|1|5|我們從他蒙恩受了使徒的職分，為他的名在萬國中使人因信而順服，
ROM|1|6|其中也有你們這蒙召屬耶穌基督的人。
ROM|1|7|我寫信給你們在 羅馬 、為上帝所愛、蒙召作聖徒的眾人。願恩惠、平安 從我們的父上帝和主耶穌基督歸給你們！
ROM|1|8|首先，我靠著耶穌基督，為你們眾人感謝我的上帝，因你們的信德傳遍了天下。
ROM|1|9|我在他兒子的福音上，用心靈所事奉的上帝可以見證，我怎樣不住地提到你們，
ROM|1|10|在我的禱告中常常懇求，或許照上帝的旨意，最終我能毫無阻礙地往你們那裏去。
ROM|1|11|因為我迫切地想見你們，要把一些屬靈的恩賜分給你們，使你們得以堅固，
ROM|1|12|也可以說，我在你們中間，因你我彼此的信心而同得安慰。
ROM|1|13|弟兄們，我不願意你們不知道，我屢次計劃往你們那裏去，要在你們中間得些果子，如同在其餘的外邦人中一樣，只是到如今仍有攔阻。
ROM|1|14|無論是 希臘 人、未開化的人、聰明人、愚拙人，我都欠他們的債，
ROM|1|15|所以願意盡我的力量把福音也傳給你們在 羅馬 的人。
ROM|1|16|我不以福音為恥；這福音本是上帝的大能，要救一切相信的，先是 猶太 人，後是 希臘 人。
ROM|1|17|因為上帝的義正在這福音上顯明出來；這義是本於信，以至於信。如經上所記：「義人必因信得生。」
ROM|1|18|原來，上帝的憤怒從天上顯明在一切不虔不義的人身上，就是那些行不義壓制真理的人。
ROM|1|19|上帝的事情，人所能知道的，原顯明在人心裏，因為上帝已經向他們顯明。
ROM|1|20|自從造天地以來，上帝的永能和神性是明明可知的，雖然眼不能見，但藉著所造之物就可以了解看見，叫人無可推諉。
ROM|1|21|因為，他們雖然知道上帝，卻不把他當作上帝榮耀他，也不感謝他。他們的思想變為虛妄，無知的心昏暗了。
ROM|1|22|他們自以為聰明，反成了愚昧，
ROM|1|23|將不能朽壞之上帝的榮耀變為偶像，仿照必朽壞的人、飛禽、走獸、爬蟲的形像。
ROM|1|24|所以，上帝任憑他們隨著心裏的情慾行污穢的事，以致彼此羞辱自己的身體。
ROM|1|25|他們將上帝的真實變為虛謊，去敬拜事奉受造之物，不敬奉那造物的主—主是可稱頌的，直到永遠。阿們！
ROM|1|26|因此，上帝任憑他們放縱可羞恥的情慾。他們的女人把自然的關係變成違反自然的；
ROM|1|27|男人也是如此，放棄了和女人自然的關係，慾火攻心，男的和男的彼此貪戀，行可恥的事，就在自己身上受這逆性行為當得的報應。
ROM|1|28|他們既然故意不認識上帝，上帝就任憑他們存扭曲的心，做那些不該做的事，
ROM|1|29|裝滿了各樣不義 、邪惡、貪婪、惡毒，滿心是嫉妒、兇殺、紛爭、詭詐、毒恨，又是毀謗的、
ROM|1|30|說人壞話的、怨恨上帝的 、侮辱人的、狂傲的、自誇的、製造是非的、忤逆父母的、
ROM|1|31|頑梗不化的、言而無信的、無情無義的、不憐憫人的。
ROM|1|32|他們雖知道上帝判定做這樣事的人是該死的，然而他們不但自己去做，還贊同別人去做。
ROM|2|1|所以，你這評斷人的人哪，無論你是誰，都無可推諉。你在甚麼事上評斷人，就在甚麼事上定自己的罪。因你這評斷人的，自己所做的卻和別人一樣。
ROM|2|2|我們知道這樣做的人，上帝必公平地審判他。
ROM|2|3|你這個人哪，你評斷做這樣事的人，自己所做的卻和別人一樣，你以為能逃脫上帝的審判嗎？
ROM|2|4|還是你藐視他豐富的恩慈、寬容、忍耐，不知道他的恩慈是領你悔改嗎？
ROM|2|5|你竟放任你剛硬不悔改的心，為自己累積憤怒！在憤怒的日子，上帝公義的審判要顯示出來。
ROM|2|6|他要照各人的行為報應各人。
ROM|2|7|凡恆心行善，尋求榮耀、尊貴和不能朽壞的，就有永生報償他們；
ROM|2|8|但是那些自私自利、不順從真理、反順從不義的人，就有惱恨、憤怒報應他們。
ROM|2|9|他要把患難、困苦加給一切作惡的人，先是 猶太 人，後是 希臘 人；
ROM|2|10|卻把榮耀、尊貴、平安加給一切行善的人，先是 猶太 人，後是 希臘 人。
ROM|2|11|因為上帝不偏待人。
ROM|2|12|凡在律法之外犯了罪的，將在律法之外滅亡；凡在律法之內犯了罪的，將按律法受審判。
ROM|2|13|原來在上帝面前，不是聽律法的為義，而是行律法的稱義。
ROM|2|14|沒有律法的外邦人若順著本性行律法上的事，他們雖然沒有律法，自己就是自己的律法。
ROM|2|15|他們顯明律法的功用刻在他們心裏，他們的良心一同作證—他們的內心掙扎，有時自責，有時為自己辯護。
ROM|2|16|在那日，上帝要藉著基督耶穌 ，按照我所傳的福音，審判人隱藏的事。
ROM|2|17|但是你，你既自稱為 猶太 人，倚靠律法，以上帝誇口，
ROM|2|18|知道上帝的旨意，從律法受了教導而能分辨是非；
ROM|2|19|你既深信自己是給盲人領路的，是在黑暗中人的光，
ROM|2|20|是無知的人的師傅，是小孩子的老師，體現了律法中的知識和真理；
ROM|2|21|那麼，你這教導別人的，還不教導自己嗎？你這宣講不可偷竊的，自己還偷竊嗎？
ROM|2|22|你這說不可姦淫的，自己還姦淫嗎？你這厭惡偶像的，自己還搶劫廟中之物嗎？
ROM|2|23|你這以律法誇口的，自己倒違犯律法，羞辱上帝！
ROM|2|24|上帝的名在外邦人中因你們受了褻瀆，正如經上所記的。
ROM|2|25|你若遵行律法，割禮固然於你有益；若違犯律法，你的割禮就算不得割禮。
ROM|2|26|所以，那未受割禮的，若遵守律法的要求，他雖然未受割禮，豈不算是受了割禮嗎？
ROM|2|27|而且那本來未受割禮的，若能全守律法，豈不是要審判你這有儀文和割禮，竟違犯律法的人嗎？
ROM|2|28|因為外表是 猶太 人的不是真 猶太 人；外表肉身的割禮也不是真割禮。
ROM|2|29|惟有內心作 猶太 人的才是真 猶太 人，真割禮也是心裏的，在乎聖靈 ，不在乎儀文。這樣的人所受的稱讚不是從人來的，而是從上帝來的。
ROM|3|1|這樣說來， 猶太 人有甚麼比別人強呢？割禮有甚麼益處呢？
ROM|3|2|很多，各方面都有。首先，上帝的聖言交託他們。
ROM|3|3|即使有不信的，這又何妨呢？難道他們的不信就廢掉上帝的信實嗎？
ROM|3|4|絕對不會！不如說，上帝是真實的，而人都是虛謊的。如經上所記： 「以致你責備的時候顯為公義； 你被指控的時候一定勝訴。」
ROM|3|5|我姑且照著人的看法來說，我們的不義若顯出上帝的義來，我們要怎麼說呢？上帝降怒是他不義嗎？
ROM|3|6|絕對不是！若是這樣，上帝怎能審判世界呢？
ROM|3|7|若上帝的真實因我的虛謊越發顯出他的榮耀，為甚麼我還像罪人一樣受審判呢？
ROM|3|8|為甚麼不說，我們可以作惡以成善呢？有人毀謗我們，說我們講過這話；這等人被定罪是應該的。
ROM|3|9|那又怎麼樣呢？我們比他們強嗎？絕不是！因我們已經指證： 猶太 人和 希臘 人都在罪惡之下。
ROM|3|10|就如經上所記： 「沒有義人，連一個也沒有。
ROM|3|11|沒有明白的， 沒有尋求上帝的。
ROM|3|12|人人偏離正路，一同走向敗壞。 沒有行善的，連一個也沒有 。
ROM|3|13|他們的喉嚨是敞開的墳墓； 他們的舌頭玩弄詭詐。 他們的嘴唇裏有毒蛇的毒液，
ROM|3|14|滿口是咒罵苦毒。
ROM|3|15|他們的腳為殺人流血飛跑；
ROM|3|16|他們的路留下毀壞和災難。
ROM|3|17|和平的路，他們不認識；
ROM|3|18|他們眼中不怕上帝。」
ROM|3|19|我們知道律法所說的話都是對律法之下的人說的，好塞住各人的口，使普世的人都伏在上帝的審判之下。
ROM|3|20|所以，凡血肉之軀沒有一個能因律法的行為而在上帝面前稱義，因為律法本是要人認識罪。
ROM|3|21|但如今，上帝的義在律法之外已經顯明出來，有律法和先知為證：
ROM|3|22|就是上帝的義，因信耶穌基督 加給一切信的人。這並沒有分別，
ROM|3|23|因為世人都犯了罪，虧缺了上帝的榮耀，
ROM|3|24|如今卻蒙上帝的恩典，藉著在基督耶穌裏的救贖，就白白地得稱為義。
ROM|3|25|上帝設立耶穌作贖罪祭，是憑耶穌的血，藉著信，要顯明上帝的義；因為他用忍耐的心寬容人先前所犯的罪，好使今時顯明他的義，讓人知道他自己為義，也稱信耶穌的人為義 。
ROM|3|26|
ROM|3|27|既是這樣，哪裏可誇口呢？沒有可誇的。是藉甚麼法呢？功德嗎？不是！是藉信主之法。
ROM|3|28|所以我們認定，人稱義是因著信，不在於律法的行為。
ROM|3|29|難道上帝只是 猶太 人的嗎？不也是外邦人的嗎？是的，他也是外邦人的上帝。
ROM|3|30|既然上帝是一位，他就要本於信稱那受割禮的為義，也要藉著信稱那未受割禮的為義。
ROM|3|31|這樣，我們藉著信廢了律法嗎？絕對不是！更是鞏固律法。
ROM|4|1|這樣，那按肉體作我們祖宗的 亞伯拉罕 ，我們要怎麼說呢？
ROM|4|2|倘若 亞伯拉罕 是因行為稱義，他就有可誇的，但是在上帝面前他一無可誇。
ROM|4|3|經上說甚麼呢？「 亞伯拉罕 信了上帝，這就算他為義。」
ROM|4|4|做工的得工資不算是恩典，而是應得的；
ROM|4|5|但那不做工的，只信那位稱不敬虔之人為義的，他的信就算為義。
ROM|4|6|正如 大衛 稱那在行為之外蒙上帝算為義的人是有福的：
ROM|4|7|「過犯得赦免，罪惡蒙遮蓋的人有福了！
ROM|4|8|主不算為有罪的，這樣的人有福了！」
ROM|4|9|如此看來，這福只加給那受割禮的人嗎？不也加給那未受割禮的人嗎？我們說，因著信，就算 亞伯拉罕 為義。
ROM|4|10|那麼，這是怎麼算的呢？是在他受割禮的時候呢？還是在他未受割禮的時候呢？不是在受割禮的時候，而是在未受割禮的時候。
ROM|4|11|並且，他受了割禮的記號，作他未受割禮的時候因信稱義的印證，為使他作一切未受割禮而信之人的父，使他們也算為義，
ROM|4|12|也使他作受割禮之人的父，就是那些不但受割禮，而且跟隨我們的祖宗 亞伯拉罕 未受割禮而信的足跡的人。
ROM|4|13|因為上帝給 亞伯拉罕 和他後裔承受世界的應許不是藉著律法，而是藉著信而得的義。
ROM|4|14|若是屬於律法的人才是後嗣，信就落空了，應許也就失效了。
ROM|4|15|因為律法是惹動憤怒的，哪裏沒有律法，哪裏就沒有過犯。
ROM|4|16|所以，人作後嗣是出於信，因此就屬乎恩，以致應許保證歸給所有的後裔，不但歸給那屬於律法的，也歸給那效法 亞伯拉罕 之信的人。 亞伯拉罕 所信的是那叫死人復活、使無變為有的上帝，在這位上帝面前 亞伯拉罕 成為我們眾人的父，如經上所記：「我已經立你作多國之父。」
ROM|4|17|
ROM|4|18|他在沒有盼望的時候，仍存著盼望來相信，就得以作多國之父，正如先前所說：「你的後裔將要如此。」
ROM|4|19|他將近百歲的時候，雖然想到 自己的身體如同已死， 撒拉 也不可能生育，他的信心還是不軟弱，
ROM|4|20|仍仰望上帝的應許，總沒有因不信而起疑惑，反倒因信而剛強，將榮耀歸給上帝，
ROM|4|21|且滿心相信上帝所應許的必能成就。
ROM|4|22|所以這也 就算他為義。
ROM|4|23|「算他為義」這句話不是單為他寫的，
ROM|4|24|也是為我們將來得算為義的人寫的，就是為我們這些信上帝使我們的主耶穌從死人中復活的人寫的。
ROM|4|25|耶穌被出賣，是為我們的過犯；他復活，是為使我們稱義。
ROM|5|1|所以，我們既因信稱義，就藉著我們的主耶穌基督得以與上帝和好。
ROM|5|2|我們又藉著他，因信 得以進入現在所站立的這恩典中，並且歡歡喜喜盼望上帝的榮耀。
ROM|5|3|不但如此，就是在患難中也是歡歡喜喜的，因為知道患難生忍耐，
ROM|5|4|忍耐生老練，老練生盼望，
ROM|5|5|盼望不至於落空，因為上帝的愛，已藉著所賜給我們的聖靈，澆灌在我們心裏。
ROM|5|6|我們還軟弱的時候，基督就在特定的時刻為不敬虔之人死。
ROM|5|7|為義人死，是少有的；為仁人死，也者有敢做的。
ROM|5|8|惟有基督在我們還作罪人的時候為我們死，上帝的愛就在此向我們顯明了。
ROM|5|9|現在我們既靠著他的血稱義，就更要藉著他得救，免受上帝的憤怒。
ROM|5|10|因為我們作仇敵的時候，尚且藉著上帝兒子的死得以與上帝和好，既已和好，就更要因他的生得救了。
ROM|5|11|不但如此，我們既藉著我們的主耶穌基督得以與上帝和好，也就藉著他以上帝為樂。
ROM|5|12|為此，正如罪是從一人進入世界，死又從罪而來，於是死就臨到所有的人，因為人人都犯了罪。
ROM|5|13|沒有律法之前，罪已經在世上，但沒有律法，罪也不算罪。
ROM|5|14|然而，從 亞當 到 摩西 ，死就掌了權，連那些不與 亞當 犯一樣罪過的，也在死的權下。 亞當 是那以後要來之人的預像。
ROM|5|15|但是過犯不如恩賜，若因一人的過犯，眾人都死了，那麼，上帝的恩典，與那因耶穌基督一人而來的恩典中的賞賜，豈不加倍地臨到眾人嗎？
ROM|5|16|因一人犯罪而來的後果，也不如賞賜，原來審判是由一人而定罪，恩賜乃是由許多過犯而稱義。
ROM|5|17|若因一人的過犯，死就因這一人掌權，那些受洪恩又蒙所賜之義的，豈不更要因耶穌基督一人在他們生命中掌權嗎？
ROM|5|18|這樣看來，因一次的過犯，所有的人都被定罪；照樣，因一次的義行，所有的人也就被稱義而得生命了。
ROM|5|19|因一人的悖逆，眾人成為罪人；照樣，因一人的順從，眾人也成為義了。
ROM|5|20|而且加添了律法，使得過犯增加，只是罪在哪裏增加，恩典就在哪裏越發豐盛了。
ROM|5|21|所以，正如罪藉著死掌權；照樣，恩典也藉著義掌權，使人因我們的主耶穌基督得永生。
ROM|6|1|這樣，我們要怎麼說呢？我們可以仍在罪中使恩典增多嗎？
ROM|6|2|絕對不可！我們向罪死了的人，豈可仍在罪中活著呢？
ROM|6|3|難道你們不知道，我們這受洗歸入基督耶穌的人，就是受洗歸入他的死嗎？
ROM|6|4|所以，我們藉著洗禮歸入死，和他一同埋葬，是要我們行事為人都有新生的樣子，像基督藉著父的榮耀從死人中復活一樣。
ROM|6|5|我們若與他合一，經歷與他一樣的死，也將經歷與他一樣的復活。
ROM|6|6|我們知道，我們的舊人和他同釘十字架，使罪身滅絕，叫我們不再作罪的奴隸，
ROM|6|7|因為已死的人是脫離了罪。
ROM|6|8|我們若與基督同死，我們信也必與他同活，
ROM|6|9|因為知道基督既從死人中復活，就不再死，死也不再作他的主了。
ROM|6|10|他死了，是對罪死，只這一次；他活，是對上帝活著。
ROM|6|11|這樣，你們也要看自己對罪是死的，在基督耶穌裏對上帝卻是活的。
ROM|6|12|所以，不要讓罪在你們必死的身上掌權，使你們順從身體的私慾。
ROM|6|13|也不要把你們的肢體獻給罪作不義的工具，倒要像從死人中活著的人，把自己獻給上帝，並把你們的肢體獻給上帝作義的工具。
ROM|6|14|罪必不能作你們的主，因你們不在律法之下，而是在恩典之下。
ROM|6|15|那又怎麼樣呢？我們在恩典之下，不在律法之下，就可以犯罪嗎？絕對不可！
ROM|6|16|難道你們不知道，你們獻自己作奴僕，順從誰就作誰的奴僕嗎？或作罪的奴隸，以至於死；或作順服的奴僕，以至於成義。
ROM|6|17|感謝上帝！因為你們從前雖然作罪的奴隸，現在卻從心裏順服了所傳給你們教導的典範。
ROM|6|18|你們既從罪裏得了釋放，就作了義的奴僕。
ROM|6|19|我因你們肉體的軟弱，就以人的觀點來說。你們從前怎樣把肢體獻給不潔不法作奴隸，以至於不法；現在也要照樣將肢體獻給義作奴僕，以至於成聖。
ROM|6|20|因為你們作罪的奴隸時，不被義所約束。
ROM|6|21|那麼，你們現在所看為羞恥的事，當時有甚麼果子呢？那些事的結局就是死。
ROM|6|22|但如今，你們既從罪裏得了釋放，作了上帝的奴僕，就結出果子，以至於成聖，那結局就是永生。
ROM|6|23|因為罪的工價乃是死；惟有上帝的恩賜，在我們的主基督耶穌裏，乃是永生。
ROM|7|1|弟兄們，我對你們這些明白律法的人說，你們豈不知道律法約束人是在他活著的時候嗎？
ROM|7|2|就如女人有了丈夫，丈夫還活著，她就被律法約束；丈夫若死了，她就從丈夫的律法中解脫了。
ROM|7|3|所以丈夫還活著，她若跟了別的男人，就叫淫婦；丈夫若死了，她就脫離了律法，雖然跟了別的男人，也不是淫婦。
ROM|7|4|我的弟兄們，這樣說來，你們藉著基督的身體對律法也是死了，使你們歸於另一位，就是歸於那從死人中復活的，為要使我們結果子給上帝。
ROM|7|5|因為我們屬肉體的時候，那因律法而生犯罪的慾望在我們肢體中發動，以致結出死亡的果子。
ROM|7|6|但如今，我們既然在捆綁我們的律法上死了，就從律法中解脫，使我們服侍主，要按著聖靈 的新樣，不按著儀文的舊樣。
ROM|7|7|這樣，我們要怎麼說呢？律法是罪嗎？絕對不是！但是，若不是藉著律法，我就不知何為罪；若不是律法說「不可貪心」，我就不知何為貪心。
ROM|7|8|然而，罪趁著機會，藉著誡命，使各樣的貪心在我裏頭發動，因為沒有律法，罪是死的。
ROM|7|9|以前沒有律法的時候，我是活的；但是誡命來到，罪活起來，
ROM|7|10|我就死了。那本該叫人活的誡命反而叫我死。
ROM|7|11|因為罪趁著機會，藉著誡命誘惑我，並且藉著誡命殺了我。
ROM|7|12|這樣看來，律法是聖的，誡命也是聖的、義的、善的。
ROM|7|13|那麼，那善的是叫我死嗎？絕對不是！叫我死的是罪。罪藉著那善的叫我死，為要顯出這真是罪，以致罪藉著誡命更顯出是惡極了。
ROM|7|14|我們原知道律法是屬靈的，我卻是屬肉體的，是已經賣給罪了。
ROM|7|15|因為我所做的，我自己不明白。我所願意的，我並不做；我所恨惡的，我反而去做。
ROM|7|16|如果我所做的是我所不願意的，我得承認律法是善的。
ROM|7|17|事實上，這不是我做的，而是住在我裏面的罪做的。
ROM|7|18|我也知道，住在我裏面的，就是我肉體之中，沒有善。因為立志為善由得我，只是行出來由不得我。
ROM|7|19|我所願意的善，我不去做；我所不願意的惡，我反而去做。
ROM|7|20|如果我去做我不願意做的，就不是我做的，而是住在我裏面的罪做的。
ROM|7|21|我覺得有個律，就是我願意行善的時候，就有惡纏著我。
ROM|7|22|因為，按著我裏面的人，我喜歡上帝的律，
ROM|7|23|但我看出肢體中另有個律和我內心的律交戰，把我擄去，使我附從那肢體中罪的律。
ROM|7|24|我真苦啊！誰能救我脫離這必死的身體呢？
ROM|7|25|感謝上帝，靠著我們的主耶穌基督就能！這樣看來，一方面，我內心順服上帝的律，另一方面，肉體卻順服罪的律了。
ROM|8|1|如今，那些在基督耶穌裏的人就不被定罪了。
ROM|8|2|因為賜生命的聖靈的律，在基督耶穌裏從罪和死的律中把你釋放出來。
ROM|8|3|律法既因肉體軟弱而無能為力，上帝就差遣自己的兒子成為罪身的樣子，為了對付罪 ，在肉體中定了罪，
ROM|8|4|為要使律法要求的義，實現在我們這不隨從肉體、只隨從聖靈去行的人身上。
ROM|8|5|因為，隨從肉體的人體貼肉體的事；隨從聖靈的人體貼聖靈的事。
ROM|8|6|體貼肉體就是死；體貼聖靈就是生命和平安 。
ROM|8|7|因為體貼肉體就是與上帝為敵，對上帝的律法不順服，事實上也無法順服。
ROM|8|8|屬肉體的人無法使上帝喜悅。
ROM|8|9|如果上帝的靈住在你們裏面，你們就不屬肉體，而是屬聖靈了。人若沒有基督的靈，就不是屬基督的。
ROM|8|10|基督若在你們裏面，身體就因罪而死，靈卻因義而活。
ROM|8|11|然而，使耶穌從死人中復活的上帝的靈若住在你們裏面，那使基督從死人中復活的，也必藉著住在你們裏面的聖靈使你們必死的身體又活過來。
ROM|8|12|弟兄們，這樣看來，我們不是欠肉體的債去順從肉體而活。
ROM|8|13|你們若順從肉體活著，必定會死；若靠著聖靈把身體的惡行處死，就必存活。
ROM|8|14|因為凡被上帝的靈引導的都是上帝的兒子。
ROM|8|15|你們所領受的不是奴僕的靈，仍舊害怕；所領受的是兒子名分的靈，因此我們呼叫：「阿爸，父！」
ROM|8|16|聖靈自己與我們的靈一同見證我們是上帝的兒女。
ROM|8|17|若是兒女，就是後嗣，是上帝的後嗣，和基督同作後嗣。如果我們和他一同受苦，是要我們和他一同得榮耀。
ROM|8|18|我認為，現在的苦楚，若比起將來要顯示給我們的榮耀，是不足介意的。
ROM|8|19|受造之物切望等候上帝的眾子顯出來。
ROM|8|20|因為受造之物屈服在虛空之下，不是自己願意，而是因那使它屈服的叫他如此。但受造之物仍然指望從敗壞的轄制下得釋放，得享上帝兒女榮耀的自由。
ROM|8|21|
ROM|8|22|我們知道，一切受造之物一同呻吟，一同忍受陣痛，直到如今。
ROM|8|23|不但如此，就是我們這有聖靈作初熟果子的，也是自己內心呻吟，等候得著兒子的名分，就是我們的身體得救贖。
ROM|8|24|我們得救是在於盼望；可是看得見的盼望就不是盼望。誰還去盼望他所看得見的呢？
ROM|8|25|但我們若盼望那看不見的，我們就耐心等候。
ROM|8|26|同樣，我們的軟弱有聖靈幫助。我們本不知道當怎樣禱告，但是聖靈親自用無可言喻的嘆息替我們祈求。
ROM|8|27|那鑒察人心的知道聖靈所體貼的，因為聖靈照著上帝的旨意替聖徒祈求。
ROM|8|28|我們知道，萬事 都互相效力，叫愛上帝的人得益處，就是按他旨意被召的人。
ROM|8|29|因為他所預知的人，他也預定他們效法他兒子的榜樣，使他兒子在許多弟兄中作長子 。
ROM|8|30|他所預定的人，他又召他們來；所召來的人，他又稱他們為義；所稱為義的人，他又叫他們得榮耀。
ROM|8|31|既是這樣，我們對這些事還要怎麼說呢？上帝若幫助我們，誰能抵擋我們呢？
ROM|8|32|上帝既不顧惜自己的兒子，為我們眾人捨了他，豈不也把萬物和他一同白白地賜給我們嗎？
ROM|8|33|誰能控告上帝所揀選的人呢？有上帝稱他們為義了。
ROM|8|34|誰能定他們的罪呢？有基督耶穌 已經死了，而且復活了，現今在上帝的右邊，也替我們祈求。
ROM|8|35|誰能使我們與基督的愛隔絕呢？難道是患難嗎？是困苦嗎？是迫害嗎？是飢餓嗎？是赤身露體嗎？是危險嗎？是刀劍嗎？
ROM|8|36|如經上所記： 「我們為你的緣故終日被殺； 人看我們如將宰的羊。」
ROM|8|37|然而，靠著愛我們的主，在這一切的事上，我們已經得勝有餘了。
ROM|8|38|因為我深信，無論是死，是活，是天使，是掌權的，是有權能的 ，是現在的事，是將來的事，
ROM|8|39|是高處的，是深處的，是別的受造之物，都不能使我們與上帝的愛隔絕，這愛是在我們的主基督耶穌裏的。
ROM|9|1|我在基督裏說真話，不說謊話；我的良心被聖靈感動為我作證。
ROM|9|2|我非常憂愁，心裏時常傷痛。
ROM|9|3|為我弟兄，我骨肉之親，就是自己被詛咒，與基督分離，我也願意。
ROM|9|4|他們是 以色列 人，那兒子的名分、榮耀、諸約、律法的頒佈、敬拜的禮儀、應許都是給他們的。
ROM|9|5|列祖是他們的，基督按肉體說也是從他們出來的。願在萬有之上的上帝被稱頌，直到永遠 。阿們！
ROM|9|6|這不是說上帝的話落了空。因為從 以色列 生的不都是 以色列 人，
ROM|9|7|也不因為是 亞伯拉罕 的後裔就都是他的兒女；惟獨「從 以撒 生的才要稱為你的後裔。」
ROM|9|8|這就是說，肉身所生的兒女不是上帝的兒女，惟獨那應許的兒女才算是後裔。
ROM|9|9|因為所應許的話是這樣：「到明年這時候我要來， 撒拉 必會生一個兒子。」
ROM|9|10|不但如此， 利百加 也是這樣。她從一個人，就是從我們的祖宗 以撒 懷了孕。
ROM|9|11|雙胞胎還沒有生下來，善惡還沒有行出來，為要貫徹上帝揀選人的旨意，
ROM|9|12|不是憑著人的行為，而是憑著那呼召人的，上帝就對 利百加 說：「將來，大的要服侍小的。」
ROM|9|13|正如經上所記：「 雅各 是我所愛的； 以掃 是我所惡的。」
ROM|9|14|這樣，我們要怎麼說呢？難道上帝有甚麼不義嗎？絕對沒有！
ROM|9|15|因他對 摩西 說： 「我要憐憫誰就憐憫誰， 要恩待誰就恩待誰。」
ROM|9|16|由此看來，這不靠人的意願，也不靠人的努力，只靠上帝的憐憫。
ROM|9|17|因為經上有話對法老說：「我將你興起來，特要在你身上彰顯我的權能，為要使我的名傳遍全地。」
ROM|9|18|由此看來，上帝要憐憫誰就憐憫誰，要使誰剛硬就使誰剛硬。
ROM|9|19|這樣，你會對我說：「那麼，他為甚麼還指責人呢？有誰能抗拒他的旨意呢？」
ROM|9|20|你這個人哪，你是誰，竟敢向上帝頂嘴呢？受造之物豈會對造他的說：「你為甚麼把我造成這樣呢？」
ROM|9|21|難道陶匠沒有權從一團泥裏拿一塊做成貴重的器皿，又拿一塊做成卑賤的器皿嗎？
ROM|9|22|倘若上帝要顯明他的憤怒，彰顯他的權能，難道不可多多忍耐寬容那應受憤怒、預備遭毀滅的器皿嗎？
ROM|9|23|這是為了要把他豐盛的榮耀彰顯在那蒙憐憫、早預備得榮耀的器皿上。
ROM|9|24|這器皿也就是我們這些蒙上帝所召的，不但是從 猶太 人中，也是從外邦人中召來的。
ROM|9|25|正如上帝在《何西阿書》上說： 「那本來不是我子民的， 我要稱為『我的子民』； 本來不是蒙愛的， 我要稱為『蒙愛的』。
ROM|9|26|從前在甚麼地方對他們說： 你們不是我的子民， 將來就在那裏稱他們為『永生上帝的兒子』。」
ROM|9|27|關於 以色列 人， 以賽亞 喊著：「雖然 以色列 人多如海沙，得救的將是剩下的餘數，
ROM|9|28|因為主要在地上施行他的話，徹底而又迅速。」
ROM|9|29|又如 以賽亞 先前說過： 「若不是萬軍之主給我們存留餘種， 我們早已變成 所多瑪 ，像 蛾摩拉 一樣了。」
ROM|9|30|這樣，我們要怎麼說呢？那不追求義的外邦人卻獲得了義，就是因信而獲得的義。
ROM|9|31|但 以色列 人追求律法的義，反而達不到律法的義。
ROM|9|32|這是甚麼緣故呢？是因為他們不憑著信心，而是憑著行為，他們正跌在那絆腳石上。
ROM|9|33|就如經上所記： 「我在 錫安 放一塊絆腳的石頭，使人跌倒的磐石； 信靠他的人必不蒙羞。」
ROM|10|1|弟兄們，我心裏所渴望的和向上帝所求的，是要 以色列 人得救。
ROM|10|2|我為他們作證，他們對上帝有熱心，但不是按著真知識。
ROM|10|3|因為不明白上帝的義，想要立自己的義，他們就不服上帝的義了。
ROM|10|4|律法的總結就是基督，使所有信他的人都得著義。
ROM|10|5|論到出於律法的義， 摩西 寫著：「行這些事的人，就必因此得生。」
ROM|10|6|但出於信的義卻如此說：「你不要心裏說：誰要升到天上去呢？（就是說，把基督領下來。）
ROM|10|7|或說：誰要下到陰間去呢？（就是說，把基督從死人中領上來。）」
ROM|10|8|他到底怎麼說呢？ 「這話語就離你近， 就在你口中，在你心裏，」 （就是說，我們傳揚所信的話語。）
ROM|10|9|你若口裏宣認耶穌為主，心裏信上帝叫他從死人中復活，就必得救。
ROM|10|10|因為，人心裏信就可以稱義，口裏宣認就可以得救。
ROM|10|11|經上說：「凡信靠他的人必不蒙羞。」
ROM|10|12|猶太 人和 希臘 人並沒有分別，因為人人都有同一位主，他也厚待求告他的每一個人。
ROM|10|13|因為「凡求告主名的就必得救」。
ROM|10|14|然而，人未曾信他，怎能求告他呢？未曾聽見他，怎能信他呢？沒有傳道的，怎能聽見呢？
ROM|10|15|若沒有奉差遣，怎能傳道呢？如經上所記：「報福音、傳喜信的人，他們的腳蹤何等佳美！」
ROM|10|16|但不是每一個人都聽從福音，因為 以賽亞 說：「主啊，我們所傳的有誰信呢？」
ROM|10|17|可見，信道是從聽道來的，聽道是從基督的話來的。
ROM|10|18|但我要問，人沒有聽見嗎？當然聽見了。 「他們的聲音傳遍全地； 他們的言語傳到地極。」
ROM|10|19|我再問， 以色列 人不知道嗎？先有 摩西 說： 「我要以不成國的激起你們嫉妒； 我要以愚頑的國惹起你們發怒。」
ROM|10|20|又有 以賽亞 放膽說： 「沒有尋找我的，我要讓他們尋見； 沒有求問我的，我要向他們顯現。」
ROM|10|21|關於 以色列 人，他說：「我整天向那悖逆頂嘴的百姓招手。」
ROM|11|1|那麼，我要問，上帝棄絕了他的百姓嗎？絕對沒有！因為我也是 以色列 人， 亞伯拉罕 的後裔，屬 便雅憫 支派的。
ROM|11|2|上帝並沒有棄絕他預先所知道的百姓。你們豈不知道經上論到 以利亞 是怎麼說的呢？他在上帝面前怎樣控告 以色列 人說：
ROM|11|3|「主啊，他們殺了你的先知，拆了你的祭壇，只剩下我一個人，他們還要我的命。」
ROM|11|4|但上帝的指示是怎麼對他說的呢？他說：「我為自己留下七千人，是未曾向 巴力 屈膝的。」
ROM|11|5|現在這時刻也是這樣，照著出於恩典的揀選，還有所留的餘數。
ROM|11|6|既是靠恩典，就不憑行為，不然，恩典就不再是恩典了。
ROM|11|7|那又怎麼說呢？ 以色列 人所尋求的，他們沒有得著。但是蒙揀選的人得著了，其餘的人卻成了頑梗不化的。
ROM|11|8|如經上所記： 「上帝給他們昏沉的靈， 眼睛看不見， 耳朵聽不到， 直到今日。」
ROM|11|9|大衛 也說： 「願他們的宴席變為羅網，變為陷阱， 變為絆腳石，作他們的報應。
ROM|11|10|願他們的眼睛昏花，看不見； 願你時常彎下他們的腰。」
ROM|11|11|那麼，我再問，他們失足是要他們跌倒嗎？絕對不是！因他們的過犯，救恩反而臨到外邦人，要激起他們嫉妒的心。
ROM|11|12|如果他們的過犯成為世界的富足，他們的缺乏成為外邦人的富足，更何況他們全數得救呢？
ROM|11|13|我對你們外邦人說，正因為我是外邦人的使徒，我敬重我的職分，
ROM|11|14|希望可以激起我骨肉之親的嫉妒，好救他們一些人。
ROM|11|15|如果他們被丟棄，世界因而得以與上帝和好；他們被收納，豈不就是從死人中復生嗎？
ROM|11|16|所獻的新麵若聖潔，整個麵團都聖潔了；樹根若聖潔，樹枝也聖潔了。
ROM|11|17|若有幾根枝子被折下來，你這野橄欖枝接上去，同享橄欖根的肥汁，
ROM|11|18|你就不可向舊枝子誇口；若是誇口，該知道不是你托著根，而是根托著你。
ROM|11|19|你會說，那些枝子被折下來是為了使我接上去。
ROM|11|20|不錯。他們因為不信，所以被折下來；你因為信，所以立得住。你不可自高，反要戰戰兢兢。
ROM|11|21|上帝既然不顧惜原來的枝子，豈會顧惜你？
ROM|11|22|可見，上帝又恩慈又嚴厲：對那跌倒的人是嚴厲的；對你是恩慈的，只要你長久在他的恩慈裏，不然，你也要被砍下來。
ROM|11|23|而且，他們若不是長久不信，仍要被接上，因為上帝能夠重新把他們接上去。
ROM|11|24|你是從那天生的野橄欖上砍下來的，尚且違反自然地接在好橄欖上，何況這些原來的枝子豈不更要接在原樹上嗎？
ROM|11|25|弟兄們，我不願意你們不知道這奧祕，恐怕你們自以為聰明。這奧祕就是有一部分 以色列 人是硬心的，等到外邦人的數目添滿了，
ROM|11|26|以色列 全家都要得救。如經上所記： 「必有一位救主從 錫安 出來， 要消除 雅各 家一切不虔不敬。」
ROM|11|27|「這就是我與他們所立的約， 那時我要除去他們的罪。」
ROM|11|28|就福音來說，他們為你們的緣故是仇敵；就揀選來說，他們因列祖的緣故是蒙愛的。
ROM|11|29|因為上帝的恩賜和選召是不會撤回的。
ROM|11|30|你們從前不順服上帝，如今因他們的不順服，你們倒蒙了憐憫。
ROM|11|31|同樣，他們現在也是不順服，叫他們因著施給你們的憐憫，現在 也就蒙憐憫。
ROM|11|32|因為上帝把眾人都圈在不順服中，為的是要憐憫眾人。
ROM|11|33|深哉，上帝的豐富、智慧和知識！ 他的判斷何其難測！ 他的蹤跡何其難尋！
ROM|11|34|誰知道主的心？ 誰作過他的謀士？
ROM|11|35|誰先給了他， 使他後來償還呢？
ROM|11|36|因為萬有都是本於他， 倚靠他，歸於他。 願榮耀歸給他，直到永遠。阿們！
ROM|12|1|所以，弟兄們，我以上帝的慈悲勸你們，將身體獻上當作活祭，是聖潔的，是上帝所喜悅的，你們如此事奉乃是理所當然的 。
ROM|12|2|不要效法這個世界，只要心意更新而變化，叫你們察驗何為上帝的善良、純全、可喜悅的旨意。
ROM|12|3|我憑著所賜我的恩對你們每一位說：不要把自己看得太高，要照著上帝所分給各人的信心來衡量，看得合乎中道。
ROM|12|4|正如我們一個身子上有好些肢體，肢體也不都有一樣的用處。
ROM|12|5|這樣，我們許多人在基督裏是一個身體，互相聯絡作肢體。
ROM|12|6|按著所得的恩典，我們各有不同的恩賜：或說預言，要按著信心的程度說預言；
ROM|12|7|或服事的，要專一服事；或教導的，要專一教導；
ROM|12|8|或勸勉的，要專一勸勉；施捨的，要誠實；治理的，要殷勤；憐憫人的，要樂意。
ROM|12|9|愛，不可虛假；惡，要厭惡；善，要親近。
ROM|12|10|愛弟兄，要相親相愛；恭敬人，要彼此推讓；
ROM|12|11|殷勤，不可懶惰。要靈裏火熱；常常服侍主。
ROM|12|12|在盼望中要喜樂；在患難中要忍耐；禱告要恆切。
ROM|12|13|聖徒有缺乏，要供給；異鄉客，要殷勤款待。
ROM|12|14|要祝福迫害你們 的，要祝福，不可詛咒。
ROM|12|15|要與喜樂的人同樂；要與哀哭的人同哭。
ROM|12|16|要彼此同心，不要心高氣傲，倒要俯就卑微的人。不要自以為聰明。
ROM|12|17|不要以惡報惡，眾人以為美的事要留心去做。
ROM|12|18|若是可行，總要盡力與眾人和睦。
ROM|12|19|各位親愛的，不要自己伸冤，寧可給主的憤怒留地步，因為經上記著：「主說：『伸冤在我，我必報應。』」
ROM|12|20|不但如此，「你的仇敵若餓了，就給他吃；若渴了，就給他喝。因為你這樣做，就是把炭火堆在他的頭上。」
ROM|12|21|不要被惡所勝，反要以善勝惡。
ROM|13|1|在上有權柄的，人人要順服，因為沒有權柄不是來自上帝的。掌權的都是上帝所立的。
ROM|13|2|所以，抗拒掌權的就是抗拒上帝所立的；抗拒的人必自招審判。
ROM|13|3|作官的原不是要使行善的懼怕，而是要使作惡的懼怕。你願意不懼怕掌權的嗎？只要行善，你就可得他的稱讚；
ROM|13|4|因為他是上帝的用人，是與你有益的。你若作惡，就該懼怕，因為他不是徒然佩劍；他是上帝的用人，為上帝的憤怒，報應作惡的。
ROM|13|5|所以，你們必須順服，不但是因上帝的憤怒，也是因著良心。
ROM|13|6|你們納糧也為這個緣故，因他們是上帝的僕役，專管這事。
ROM|13|7|凡人所當得的，就給他。當得糧的，給他納糧；當得稅的，給他上稅；當懼怕的，懼怕他；當恭敬的，恭敬他。
ROM|13|8|你們除了彼此相愛，對任何人都不可虧欠甚麼，因為那愛人的就成全了律法。
ROM|13|9|那不可姦淫，不可殺人，不可偷盜，不可貪婪，或別的誡命，都包括在「愛鄰 如己」這一句話之內了。
ROM|13|10|愛是不對鄰人作惡，所以愛就成全了律法。
ROM|13|11|還有，你們要知道，現在正是該從睡夢中醒來的時候了；因為我們得救，現在比初信的時候更近了。
ROM|13|12|黑夜已深，白晝將近。所以我們該除去暗昧的行為，帶上光明的兵器。
ROM|13|13|行事為人要端正，好像在白晝行走。不可荒宴醉酒；不可好色淫蕩；不可紛爭嫉妒。
ROM|13|14|總要披戴主耶穌基督，不要只顧滿足肉體，去放縱私慾。
ROM|14|1|信心軟弱的，你們要接納，不同的意見，不要爭論。
ROM|14|2|有人信甚麼都可吃；但那軟弱的，只吃蔬菜。
ROM|14|3|吃的人不可輕看不吃的人；不吃的人也不可評斷吃的人，因為上帝已經接納他了。
ROM|14|4|你是誰，竟評斷別人的僕人呢？他或站立或跌倒，自有他的主人在，而且他也必會站立，因為主能使他站穩。
ROM|14|5|有人看這日比那日強；有人看日日都是一樣。只是各人要在自己的心意上堅定。
ROM|14|6|守日子的人是為主守的。吃的人是為主吃的，因他感謝上帝；不吃的人是為主不吃的，他也感謝上帝。
ROM|14|7|我們沒有一個人為自己而活，也沒有一個人為自己而死。
ROM|14|8|我們若活，是為主而活；我們若死，是為主而死。所以，我們或死或活總是主的人。
ROM|14|9|為此，基督死了，又活了，為要作死人和活人的主。
ROM|14|10|可是你，你為甚麼評斷弟兄呢？你又為甚麼輕看弟兄呢？因我們都要站在上帝的審判臺前。
ROM|14|11|經上寫著： 「主說，我指著我的永生起誓： 萬膝必向我跪拜； 萬口必稱頌上帝。」
ROM|14|12|這樣看來，我們各人一定要把自己的事在上帝面前 交代。
ROM|14|13|所以，我們不可再彼此評斷，寧可決意不給弟兄放置障礙或絆腳石。
ROM|14|14|我憑著主耶穌確知深信，凡物本來沒有不潔淨的，除非人以為不潔淨的，在他就不潔淨了。
ROM|14|15|你若因食物使弟兄憂愁，就不是按著愛心行事。基督已經為他死，你不可因你的食物使他敗壞。
ROM|14|16|所以，不可讓你們的善被人毀謗。
ROM|14|17|因為上帝的國不在乎飲食，而在乎公義、和平及聖靈中的喜樂 。
ROM|14|18|凡這樣服侍基督的，就為上帝所喜悅，又為人所讚許。
ROM|14|19|所以，我們務要追求 和平與彼此造就的事。
ROM|14|20|不可因食物毀壞上帝的工作。一切都是潔淨的，但有人因食物使人跌倒，這在他就是惡了。
ROM|14|21|無論是吃肉是喝酒，是甚麼別的事，使弟兄跌倒，一概不做，才是善的。
ROM|14|22|你有信心，就要在上帝面前持守。人能在自己以為可行的事上不自責就有福了。
ROM|14|23|若有人疑惑而吃的，就被定罪，因為他吃不是出於信心。凡不出於信心的都是罪。
ROM|15|1|我們堅強的人應該分擔不堅強的人的軟弱，不求自己的喜悅。
ROM|15|2|我們各人務必要讓鄰人喜悅，使他得益處，得造就。
ROM|15|3|因為基督也不求自己的喜悅，如經上所記：「辱罵你的人的辱罵都落在我身上。」
ROM|15|4|從前所寫的聖經都是為教導我們寫的，要使我們藉著忍耐和因聖經所生的安慰，得著盼望。
ROM|15|5|但願賜忍耐和安慰的上帝使你們彼此同心，效法基督耶穌，
ROM|15|6|為使你們同心同聲榮耀我們主耶穌基督的父上帝！
ROM|15|7|所以，你們要彼此接納，如同基督接納你們一樣，歸榮耀給上帝。
ROM|15|8|我說，基督是為上帝真理作了受割禮的人的執事，要證實所應許列祖的話，
ROM|15|9|並使外邦人，因他的憐憫，榮耀上帝。如經上所記： 「因此，我要在外邦中稱頌你， 歌頌你的名。」
ROM|15|10|又說： 「外邦人哪，你們要與主的子民一同歡樂。」
ROM|15|11|又說： 「列邦啊，你們要讚美主！ 萬民哪，你們都要頌讚他！」
ROM|15|12|又有 以賽亞 說： 「將來有 耶西 的根， 就是那興起來要治理列邦的； 外邦人要仰望他。」
ROM|15|13|願賜盼望的上帝，因你們的信把各樣的喜樂、平安 充滿你們的心，使你們藉著聖靈的能力大有盼望！
ROM|15|14|我的弟兄們，我本人也深信你們自己充滿良善，有各種豐富的知識，也能彼此勸戒。
ROM|15|15|但我更大膽寫信給你們，是要在一些事上提醒你們，我因上帝所賜我的恩，
ROM|15|16|使我為外邦人作基督耶穌的僕役，作上帝福音的祭司，使所獻上的外邦人因著聖靈成為聖潔，可蒙悅納。
ROM|15|17|所以，有關上帝面前的事奉，我在基督耶穌裏是有可誇的。
ROM|15|18|除了基督藉我做的那些事，我甚麼都不敢提，只提他藉我的言語作為，用神蹟奇事的能力，並上帝的靈 的能力，使外邦人順服；甚至我從 耶路撒冷 ，直轉到 以利哩古 ，到處傳了基督的福音。
ROM|15|19|
ROM|15|20|這樣，我立了志向，不在基督的名已經傳揚過的地方傳福音，免得建造在別人的根基上；
ROM|15|21|卻如經上所記： 「未曾傳給他們的，他們必看見； 未曾聽見過的事，他們要明白。」
ROM|15|22|因此我多次被攔阻，不能到你們那裏去。
ROM|15|23|但如今，在這一帶再沒有可傳的地方，而且這許多年來，我迫切想去你們那裏，
ROM|15|24|盼望到 西班牙 去的時候經過，得見你們，先與你們彼此交往，心裏稍得滿足，然後蒙你們為我送行。
ROM|15|25|但如今我要到 耶路撒冷 去，供應聖徒的需要。
ROM|15|26|因為 馬其頓 和 亞該亞 人樂意湊出一些捐款給 耶路撒冷 聖徒中的窮人。
ROM|15|27|這固然是他們樂意的，其實也算是所欠的債；因為外邦人既然分享了他們靈性上的好處，就當把肉體上的需用供給他們。
ROM|15|28|等我辦完了這事，把這筆捐款 交付給他們，我就要路過你們那裏，到 西班牙 去。
ROM|15|29|我也知道去你們那裏的時候，我將帶著基督豐盛的恩典去。
ROM|15|30|弟兄們，我藉著我們的主耶穌基督，又藉著聖靈的愛，勸你們與我一同竭力為我祈求上帝，
ROM|15|31|使我脫離在 猶太 不順從的人，也讓我在 耶路撒冷 的事奉可蒙聖徒悅納，
ROM|15|32|並使我照著上帝的旨意歡歡喜喜地到你們那裏，與你們同得安息。
ROM|15|33|願賜平安的上帝與你們眾人同在。阿們！
ROM|16|1|我對你們推薦我們的姊妹 非比 ，她是 堅革哩 教會中的執事。
ROM|16|2|請你們在主裏用合乎聖徒的方式來接待她。她在任何事上需要你們幫助，你們就幫助她；因她素來幫助許多人，也幫助了我。
ROM|16|3|請向 百基拉 和 亞居拉 問安。他們在基督耶穌裏作我的同工，
ROM|16|4|也為我的性命把自己的生死置之度外；不但我感謝他們，就是外邦的眾教會也感謝他們。
ROM|16|5|又向在他們家中的教會問安。向我所親愛的 以拜尼土 問安，他是 亞細亞 歸於基督的初結果子。
ROM|16|6|又向 馬利亞 問安，她為你們非常辛勞。
ROM|16|7|又向與我一同坐監的親戚 安多尼古 和 猶尼亞 問安，他們在使徒中是有名望的，也是比我先在基督裏的。
ROM|16|8|又向我在主裏面所親愛的 暗伯利 問安。
ROM|16|9|又向我們在基督裏的同工 耳巴奴 和我所親愛的 士大古 問安。
ROM|16|10|又向在基督裏經過考驗的 亞比利 問安。向 亞利多布 家裏的人問安。
ROM|16|11|又向我親戚 希羅天 問安。向 拿其數 家在主裏的人問安。
ROM|16|12|又向為主辛勞的 土非拿 和 土富撒 問安。向所親愛、為主非常辛勞的 彼息 問安。
ROM|16|13|又向在主裏蒙揀選的 魯孚 和他母親問安，他的母親就是我的母親。
ROM|16|14|又向 亞遜其土 、 弗勒干 、 黑米 、 八羅巴 、 黑馬 ，和跟他們在一起的弟兄們問安。
ROM|16|15|又向 非羅羅古 和 猶利亞 ， 尼利亞 和他姊妹， 阿林巴 和跟他們在一起的眾聖徒問安。
ROM|16|16|你們要以聖潔的吻彼此問安。基督的眾教會都向你們問安！
ROM|16|17|弟兄們，那些離間你們、使你們跌倒、違背所學之道的人，我勸你們要留意躲避他們。
ROM|16|18|因為這樣的人不服侍我們的主基督，只服侍自己的肚腹，用花言巧語誘惑老實人的心。
ROM|16|19|你們的順服已經傳於眾人，所以我為你們歡喜；但我願你們在善上聰明，在惡上愚拙。
ROM|16|20|那賜平安 的上帝快要把撒但踐踏在你們腳下。願我們主耶穌基督的恩與你們同在！
ROM|16|21|我的同工 提摩太 ，和我的親戚 路求 、 耶孫 、 所西巴德 ，向你們問安。
ROM|16|22|我這代筆寫信的 德提 ，在主裏向你們問安。
ROM|16|23|那接待我，也接待全教會的 該猶 ，向你們問安。城裏的財務官 以拉都 和弟兄 括土 向你們問安。
ROM|16|24|
ROM|16|25|惟有上帝能照我所傳的福音和所講的耶穌基督，並照歷代以來隱藏的奧祕的啟示，堅固你們。
ROM|16|26|這奧祕如今顯示出來，而且按著永生上帝的命令，藉眾先知的書指示萬民，使他們因信而順服。
ROM|16|27|願榮耀，藉著耶穌基督，歸給獨一全智的上帝，直到永遠。阿們！
