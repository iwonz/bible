JOHN|1|1|太初有道，道与上帝同在，道就是上帝。
JOHN|1|2|这道太初与上帝同在。
JOHN|1|3|万物都是藉着他造的，没有一样不是藉着他造的。凡被造的，
JOHN|1|4|在他里面有生命 ，这生命就是人的光。
JOHN|1|5|光照在黑暗里，黑暗却没有胜过光 。
JOHN|1|6|有一个人，是从上帝那里差来的，名叫 约翰 。
JOHN|1|7|这人来是为了作见证，是为那光作见证，要使众人藉着他而信。
JOHN|1|8|他不是那光，而是要为那光作见证。
JOHN|1|9|那光是真光，来到世上，照亮所有的人 。
JOHN|1|10|他在世界，世界是藉着他造的，世界却不认识他。
JOHN|1|11|他来到自己的地方，自己的人并不接纳他。
JOHN|1|12|凡接纳他的，就是信他名的人，他就赐他们权柄作上帝的儿女。
JOHN|1|13|这些人不是从血生的，不是从情欲生的，也不是从人的意愿生的，而是从上帝生的。
JOHN|1|14|道成了肉身，住在我们中间，充充满满地有恩典有真理，我们也见过他的荣光，正是父独一儿子 的荣光。
JOHN|1|15|约翰 为他作见证，喊着说：“这就是我曾说：‘那在我以后来的先于我，因为在我以前，他已经存在。’”
JOHN|1|16|从他的丰富里，我们都领受了恩典，而且恩上加恩。
JOHN|1|17|律法是藉着 摩西 颁布的；恩典和真理却是由耶稣基督来的。
JOHN|1|18|从来没有人见过上帝，只有在父怀里独一的儿子将他表明出来。
JOHN|1|19|这是 约翰 的见证： 犹太 人从 耶路撒冷 差祭司和 利未 人到 约翰 那里去问他：“你是谁？”
JOHN|1|20|他就承认，并不隐瞒，承认说：“我不是基督。”
JOHN|1|21|他们又问他：“那么，你是谁？是 以利亚 吗？”他说：“我不是。”“是那位先知吗？”他回答：“不是。”
JOHN|1|22|于是他们对他说：“你到底是谁，好让我们回覆差我们来的人。你说，你自己是谁？”
JOHN|1|23|他说： “我就是那在旷野呼喊的声音： 修直主的道。” 正如 以赛亚 先知所说的。
JOHN|1|24|那些人是法利赛人差来的。
JOHN|1|25|他们就问他：“你既不是基督，不是 以利亚 ，也不是那位先知，那么，你为什么施洗呢？”
JOHN|1|26|约翰 回答：“我是用水施洗，但有一位站在你们中间，是你们不认识的，
JOHN|1|27|就是那在我以后来的，我给他解鞋带也不配。”
JOHN|1|28|这些事发生在 约旦河 东边的 伯大尼 ， 约翰 施洗的地方。
JOHN|1|29|第二天， 约翰 看见耶稣来到他那里，就说：“看哪，上帝的羔羊，除去世人的罪的！
JOHN|1|30|这就是我曾说‘那在我以后来的先于我，因为在我以前，他已经存在’的那一位。
JOHN|1|31|我先前不认识他，如今我来用水施洗，为要使他显明给 以色列 人。”
JOHN|1|32|约翰 又作见证说：“我曾看见圣灵仿佛鸽子从天降下，停留在他的身上。
JOHN|1|33|我先前不认识他，可是那差我来用水施洗的对我说：‘你看见圣灵降下来，停留在谁的身上，谁就是用圣灵施洗的。’
JOHN|1|34|我看见了，所以作证：这一位是上帝的儿子。”
JOHN|1|35|又过了一天， 约翰 同两个门徒站在那里。
JOHN|1|36|他见耶稣走过，就说：“看哪，上帝的羔羊！”
JOHN|1|37|两个门徒听见他的话，就跟从了耶稣。
JOHN|1|38|耶稣转过身来，看见他们跟着，就对他们说：“你们要什么？”他们对他说：“拉比，你在哪里住？”（“拉比”翻出来就是老师。）
JOHN|1|39|耶稣说：“你们来看。”他们就去看他在哪里住。这一天他们就跟他同住；那时大约是下午四点钟。
JOHN|1|40|听了 约翰 的话而跟从耶稣的那两个人，其中一个是 西门．彼得 的弟弟 安得烈 。
JOHN|1|41|他先找到自己的哥哥 西门 ，对他说：“我们遇见弥赛亚了。”（“弥赛亚”翻出来就是基督。）
JOHN|1|42|于是 安得烈 领 西门 去见耶稣。耶稣看着他，说：“你是 约翰 的儿子 西门 ，你要称为 矶法 。”（“矶法”翻出来就是 彼得 。）
JOHN|1|43|又过了一天，耶稣想要往 加利利 去。他找到 腓力 ，就对他说：“来跟从我！”
JOHN|1|44|这 腓力 是 伯赛大 人，是 安得烈 和 彼得 的同乡。
JOHN|1|45|腓力 找到 拿但业 ，对他说：“ 摩西 在律法书上所写的，和众先知所记的那一位，我们遇见了，就是 约瑟 的儿子 拿撒勒 人耶稣。”
JOHN|1|46|拿但业 对他说：“ 拿撒勒 还能出什么好的吗？” 腓力 说：“你来看。”
JOHN|1|47|耶稣看见 拿但业 向他走来，就论到他说：“看哪，这真是个 以色列 人！他心里是没有诡诈的。”
JOHN|1|48|拿但业 对耶稣说：“你从哪里认识我的？”耶稣回答他说：“ 腓力 还没有呼唤你，你在无花果树底下，我就看见你了。”
JOHN|1|49|拿但业 回答他说：“拉比！你是上帝的儿子，你是 以色列 的王。”
JOHN|1|50|耶稣回答他说：“因为我说在无花果树底下看见你，你就信吗？你将看见比这些更大的事呢！”
JOHN|1|51|他又说：“我实实在在地告诉你们，你们将要看见天开了，上帝的使者在人子身上，上去下来。”
JOHN|2|1|第三日，在 加利利 的 迦拿 有一个婚宴，耶稣的母亲在那里。
JOHN|2|2|耶稣和他的门徒也被请去赴宴。
JOHN|2|3|酒用完了，耶稣的母亲对他说：“他们没有酒了。”
JOHN|2|4|耶稣说：“母亲 ，我与你何干呢？我的时候还没有到。”
JOHN|2|5|他母亲对用人说：“他告诉你们什么，你们就做吧。”
JOHN|2|6|照 犹太 人洁净礼的规矩，有六口石缸摆在那里，每口可以盛两三桶 水。
JOHN|2|7|耶稣对用人说：“把缸倒满水。”他们就倒满了，直到缸口。
JOHN|2|8|耶稣又说：“现在舀出来，送给宴会总管。”他们就送了去。
JOHN|2|9|宴会总管尝了那水变的酒，并不知道是哪里来的，只有舀水的用人知道。于是宴会总管叫新郎来，
JOHN|2|10|对他说：“人家都是先摆上好酒，等客人喝够了才摆上次的，你倒把好酒留到现在！”
JOHN|2|11|这是耶稣所行的第一个神迹，是在 加利利 的 迦拿 行的，显出了他的荣耀来，他的门徒就信他了。
JOHN|2|12|这事以后，耶稣与他的母亲、兄弟 和门徒 都下 迦百农 去，在那里住了不多几天。
JOHN|2|13|犹太 人的逾越节近了，耶稣上 耶路撒冷 去。
JOHN|2|14|他看见圣殿里有卖牛羊和鸽子的，还有兑换银钱的人坐着，
JOHN|2|15|耶稣就拿绳子做成鞭子，把所有的，包括牛羊都赶出圣殿，倒出兑换银钱之人的银钱，推翻他们的桌子，
JOHN|2|16|又对卖鸽子的说：“把这些东西拿走！不要把我父的殿当作买卖的地方。”
JOHN|2|17|他的门徒就想起经上记着：“我为你的殿心里焦急，如同火烧。”
JOHN|2|18|因此 犹太 领袖问他：“你能显什么神迹给我们看，表明你可以做这些事呢？”
JOHN|2|19|耶稣回答他们说：“你们拆毁这殿，我三日内要把它重建。”
JOHN|2|20|犹太 人问：“这殿造了四十六年，你三日内就能重建吗？”
JOHN|2|21|但耶稣所说的殿是指他的身体。
JOHN|2|22|所以他从死人中复活以后，门徒想起他曾说过这事，就信了圣经和耶稣所说的话。
JOHN|2|23|耶稣在 耶路撒冷 过逾越节的时候，有许多人看见他所行的神迹，就信了他的名。
JOHN|2|24|耶稣自己却不信任他们，因为他认识所有的人，
JOHN|2|25|也用不着谁来证明人是怎样的，因为他自己认识人的内心。
JOHN|3|1|有一个法利赛人，名叫 尼哥德慕 ，是 犹太 人的官。
JOHN|3|2|这人夜里来见耶稣，对他说：“拉比，我们知道你是由上帝那里来作老师的；因为你所行的神迹，若没有上帝同在，无人能行。”
JOHN|3|3|耶稣回答他说：“我实实在在地告诉你，人若不重生 ，就不能见上帝的国。”
JOHN|3|4|尼哥德慕 对他说：“人已经老了，如何能重生呢？岂能再进母腹生出来吗？”
JOHN|3|5|耶稣回答：“我实实在在地告诉你，人若不是从水和圣灵生的，就不能进上帝的国。
JOHN|3|6|从肉身生的就是肉身；从灵生的就是灵。
JOHN|3|7|我说‘你们必须重生’，你不要惊讶。
JOHN|3|8|风 随着意思吹，你听见风的声音，却不知道是从哪里来，往哪里去；凡从圣灵生的也是如此。”
JOHN|3|9|尼哥德慕 问他：“怎么能有这些事呢？”
JOHN|3|10|耶稣回答，对他说：“你是 以色列 人的老师，还不明白这些事吗？
JOHN|3|11|我实实在在地告诉你，我们所说的是我们知道的，我们所见证的是我们见过的，你们却不领受我们的见证。
JOHN|3|12|我对你们说地上的事，你们尚且不信，若对你们说天上的事，如何能信呢？
JOHN|3|13|除了从天降下 的人子，没有人升过天。
JOHN|3|14|摩西 在旷野怎样举蛇，人子也必须照样被举起来，
JOHN|3|15|要使一切信他的人都得永生。
JOHN|3|16|“上帝爱世人，甚至将他独一的儿子 赐给他们，叫一切信他的人不致灭亡，反得永生。
JOHN|3|17|因为上帝差他的儿子到世上来，不是要定世人的罪 ，而是要使世人因他得救。
JOHN|3|18|信他的人不被定罪；不信的人已经被定罪了，因为他不信上帝独一儿子的名。
JOHN|3|19|光来到世上，世人因自己的行为是恶的，不爱光，倒爱黑暗，这就定了他们的罪。
JOHN|3|20|凡作恶的人都恨恶光，不来接近光，恐怕他的行为被暴露。
JOHN|3|21|但实行真理的人就来接近光，为要显明他的行为是靠上帝而行的。”
JOHN|3|22|这些事以后，耶稣和门徒到了 犹太 地区，在那里他和他们同住，并且施洗。
JOHN|3|23|约翰 也在靠近 撒冷 的 哀嫩 施洗，因为那里水多，众人都去受洗。
JOHN|3|24|那时 约翰 还没有下在监里。
JOHN|3|25|约翰 的门徒和一个 犹太 人辩论洁净的礼仪，
JOHN|3|26|就来见 约翰 ，对他说：“拉比，从前同你在 约旦河 的东边，你所见证的那位，你看，他在施洗，众人都到他那里去了。”
JOHN|3|27|约翰 回答说：“若不是从天上赐的，人就不能得到什么。
JOHN|3|28|你们自己可以为我作见证，我曾说，我不是基督，只是奉差遣在他前面开路的。
JOHN|3|29|娶新娘的是新郎；新郎的朋友站在一旁听，一听见新郎的声音就欢喜快乐。因此，我这喜乐得以满足了。
JOHN|3|30|他必兴旺；我必衰微。”
JOHN|3|31|“从上头来的是在万有之上；出于地的是属于地，他所说的也是属于地。从天上来的是在万有之上。
JOHN|3|32|他把所见所闻的见证出来，只是没有人领受他的见证。
JOHN|3|33|那领受他见证的，就印证上帝是真实的。
JOHN|3|34|上帝所差来的说上帝的话，因为上帝所赐给他的圣灵是没有限量的。
JOHN|3|35|父爱子，已把万有交在他手里。
JOHN|3|36|信子的人有永生；不信子的人得不到永生，而且上帝的愤怒常在他身上。”
JOHN|4|1|耶稣 知道法利赛人听见他收门徒和施洗比 约翰 还多， （
JOHN|4|2|其实不是耶稣亲自施洗，而是他的门徒施洗，）
JOHN|4|3|他就离开 犹太 ，又回 加利利 去。
JOHN|4|4|他必须经过 撒玛利亚 ，
JOHN|4|5|于是到了 撒玛利亚 的一座城，名叫 叙加 ，靠近 雅各 给他儿子 约瑟 的那块地。
JOHN|4|6|雅各井 就在那里；耶稣因旅途疲乏，坐在井旁。那时约是正午。
JOHN|4|7|有一个 撒玛利亚 妇人来打水。耶稣对她说：“请给我水喝。”
JOHN|4|8|因为那时门徒进城买食物去了。
JOHN|4|9|撒玛利亚 妇人对他说：“你是 犹太 人，怎么向我一个 撒玛利亚 女人要水喝呢？”因为 犹太 人和 撒玛利亚 人没有来往。
JOHN|4|10|耶稣回答她说：“你若知道上帝的恩赐，和对你说‘请给我水喝’的是谁，你早就会求他，他也早就会给了你活水。”
JOHN|4|11|妇人对耶稣说：“先生，你没有打水的器具，井又深，哪里去取活水呢？
JOHN|4|12|我们的祖宗 雅各 把这井留给我们，他自己和儿女以及牲畜都喝这井里的水，难道你比他还大吗？”
JOHN|4|13|耶稣回答，对她说：“凡喝这水的，还要再渴；
JOHN|4|14|谁喝我所赐的水，就永远不渴。我所赐的水要在他里面成为泉源，直涌到永生。”
JOHN|4|15|妇人对他说：“先生，请把这水赐给我，使我不渴，也不用到这里来打水。”
JOHN|4|16|耶稣对她说：“你去，叫你的丈夫，再到这里来。”
JOHN|4|17|妇人回答，对耶稣说：“我没有丈夫。”耶稣说：“你说没有丈夫是对的。
JOHN|4|18|你已经有过五个丈夫，你现在有的并不是你的丈夫。你这话是真的。”
JOHN|4|19|妇人对他说：“先生，我看你是一位先知。
JOHN|4|20|我们的祖宗在这山上敬拜上帝，你们倒说，应当敬拜的地方是在 耶路撒冷 。”
JOHN|4|21|耶稣对她说：“妇人，你要信我。时候将到，你们敬拜父，既不在这山上，也不在 耶路撒冷 。
JOHN|4|22|你们所敬拜的，你们不知道；我们所敬拜的，我们知道，因为救恩是从 犹太 人出来的。
JOHN|4|23|时候将到，现在就是了，那真正敬拜父的，要用心灵和诚实敬拜他，因为父要这样的人敬拜他。
JOHN|4|24|上帝是灵，所以敬拜他的必须用心灵和诚实敬拜他。”
JOHN|4|25|妇人对他说：“我知道弥赛亚—就是那称为基督的—要来；他来了，会把一切的事都告诉我们。”
JOHN|4|26|耶稣对她说：“我就是，正在跟你说话呢！”
JOHN|4|27|正在这时，门徒回来了。他们对耶稣正在和一个妇人说话感到惊讶，可是没有人说：“你要什么？”或说：“你为什么和她说话？”
JOHN|4|28|那妇人留下水罐，往城里去，对众人说：
JOHN|4|29|“你们来看！有一个人把我素来所做的一切事都说了出来，难道这个人就是基督吗？”
JOHN|4|30|他们就出城，来到耶稣那里。
JOHN|4|31|就在这个时候，门徒求耶稣说：“拉比，请吃吧。”
JOHN|4|32|耶稣对他们说：“我有食物吃，是你们不知道的。”
JOHN|4|33|门徒就彼此说：“难道有人拿什么给他吃了吗？”
JOHN|4|34|耶稣对他们说：“我的食物就是要遵行差我来那位的旨意，完成他的工作。
JOHN|4|35|你们不是说‘到收割的时候还有四个月’吗？我告诉你们，举目向田观看，庄稼熟了，可以收割了。
JOHN|4|36|收割的人已经得工钱 ，为永生储存五谷，使撒种的和收割的一同快乐。
JOHN|4|37|‘那人撒种，这人收割’，这话可见是真的。
JOHN|4|38|我差你们去收你们所没有辛劳的；别人辛劳，你们享受他们辛劳的成果。”
JOHN|4|39|那城里有好些 撒玛利亚 人信了耶稣，因为那妇人作见证，说：“他把我素来所做的一切事都说了出来。”
JOHN|4|40|于是 撒玛利亚 人来见耶稣，求他在他们那里住下，他就在那里住了两天。
JOHN|4|41|因为耶稣的话，信的人就更多了。
JOHN|4|42|他们对那妇人说：“现在我们信，不再是因为你的话，而是我们亲自听见了，知道这人真是世界的救主。”
JOHN|4|43|过了那两天，耶稣离开那地方，往 加利利 去。
JOHN|4|44|因为耶稣自己作过见证说：“先知在自己的家乡是没有人尊敬的。”
JOHN|4|45|到了 加利利 ， 加利利 人都欢迎他，因为他们也上 耶路撒冷 去过节，曾经看过他在节期间所做的一切事。
JOHN|4|46|耶稣又到了 加利利 的 迦拿 ，就是他从前变水为酒的地方。有一个大臣，他的儿子在 迦百农 病了。
JOHN|4|47|他听见耶稣从 犹太 到了 加利利 ，就来见他，求他下去医治他的儿子，因为他儿子快要死了。
JOHN|4|48|耶稣对他说：“若不看见神迹奇事，你们总是不信。”
JOHN|4|49|那大臣对他说：“先生，求你趁着我的孩子还没有死就下去吧。”
JOHN|4|50|耶稣对他说：“回去吧，你的儿子会活！”那人信耶稣所说的话，就回去了。
JOHN|4|51|正下去的时候，他的仆人迎面而来，说他的儿子活了。
JOHN|4|52|他就问什么时候见好的。他们对他说：“昨天下午一点钟热就退了。”
JOHN|4|53|他就知道这正是耶稣对他说“你的儿子会活”的时候；他自己和全家就都信了。
JOHN|4|54|这是耶稣从 犹太 回到 加利利 后所行的第二个神迹。
JOHN|5|1|这些事以后，到了 犹太 人的一个节期，耶稣上 耶路撒冷 去。
JOHN|5|2|在 耶路撒冷 ，靠近 羊门 有一个池子， 希伯来 话叫 毕士大 ，旁边有五个柱廊；
JOHN|5|3|里面躺着许多病人，有失明的、瘸腿的、瘫痪的 。
JOHN|5|4|
JOHN|5|5|在那里有一个人，病了三十八年。
JOHN|5|6|耶稣看见他躺着，知道他病了很久，就问他：“你要痊愈吗？”
JOHN|5|7|病人回答他：“先生，水动的时候，没有人把我放在池子里；我正要去的时候，别人比我先下去了。”
JOHN|5|8|耶稣对他说：“起来，拿起你的褥子走吧！”
JOHN|5|9|那人立刻痊愈，就拿起自己的褥子走了。 那天是安息日，
JOHN|5|10|所以 犹太 人对那被治好了的人说：“今天是安息日，你拿褥子是不合法的。”
JOHN|5|11|他却回答他们：“那使我痊愈的人对我说：‘拿起你的褥子走吧！’”
JOHN|5|12|他们问他：“对你说‘拿起褥子走’的是什么人？”
JOHN|5|13|那治好了的人不知道那人是谁，因为那里人很多，耶稣已经躲开了。
JOHN|5|14|后来耶稣在圣殿里找到他，对他说：“你已经痊愈了，不要再犯罪，免得你的遭遇更坏。”
JOHN|5|15|那人就去告诉 犹太 人，使他痊愈的是耶稣。
JOHN|5|16|所以 犹太 人迫害耶稣，因为他在安息日做了这些事。
JOHN|5|17|耶稣就回答他们：“我父做事直到如今，我也做事。”
JOHN|5|18|为了这缘故， 犹太 人越发想要杀他，因为他不但犯了安息日，而且称上帝为他的父，把自己和上帝看为同等。
JOHN|5|19|于是耶稣回答，对他们说：“我实实在在地告诉你们，子凭着自己不能做什么，惟有看见父所做的，他才做；父所做的事，子也照样做。
JOHN|5|20|父爱子，将自己所做的一切事指示给他看，还要将比这更大的事给他看，使你们惊讶。
JOHN|5|21|父怎样叫死人复活，赐他们生命，子也照样随自己的意愿赐人生命。
JOHN|5|22|父不审判任何人，而是把审判的事全交给子，
JOHN|5|23|为要使人都尊敬子，如同尊敬父一样。不尊敬子的，就是不尊敬差子来的父。
JOHN|5|24|“我实实在在地告诉你们，那听我话又信差我来那位的，就有永生，不至于被定罪，而是已经出死入生了。
JOHN|5|25|我实实在在地告诉你们，时候将到，现在就是了，死人要听见上帝儿子的声音，听见的人就要活了。
JOHN|5|26|因为父怎样自己里面有生命，也照样赐给他儿子自己里面有生命，
JOHN|5|27|并且赐给他施行审判的权柄，因为他是人子。
JOHN|5|28|你们不要对这事感到惊讶，因为时候将到，凡在坟墓里的，都要听见他的声音，
JOHN|5|29|并且要出来：行善的，复活得生命；作恶的，复活被定罪。
JOHN|5|30|“我凭着自己不能做什么。我怎么听见就怎么审判，而我的审判是公平的，因为我不寻求自己的意愿，只寻求差我来那位的旨意。”
JOHN|5|31|“我若为自己作见证，我的见证就不真。
JOHN|5|32|另有一位为我作见证，我也知道他为我作的见证是真的。
JOHN|5|33|你们曾差人到 约翰 那里，他为真理作过见证。
JOHN|5|34|其实，我所受的见证不是从人来的；然而，我说这些话是为了使你们得救。
JOHN|5|35|约翰 是点亮的明灯，你们情愿因他的光欢欣一时。
JOHN|5|36|但我有比 约翰 更大的见证：父交给我去完成的工作，就是我正在做的，为我作证是父差遣了我。
JOHN|5|37|那差我来的父也为我作了见证。你们从来没有听见他的声音，也没有看见他的形像。
JOHN|5|38|你们并没有他的道存在心里，因为你们不信他所差来的那一位。
JOHN|5|39|你们查考圣经，因你们以为其中有永生；而这经正是为我作见证的。
JOHN|5|40|然而，你们不肯到我这里来得生命。
JOHN|5|41|“我不接受从人来的荣耀，
JOHN|5|42|但我知道，你们没有爱上帝的心。
JOHN|5|43|我奉我父的名来了，你们并不接纳我；若有别人奉自己的名来，你们倒会接纳他。
JOHN|5|44|你们互相受荣耀，却不寻求从独一上帝来的荣耀，怎能信我呢？
JOHN|5|45|不要以为我会在父面前告你们；有一位告你们的，就是你们所仰望的 摩西 。
JOHN|5|46|如果你们信 摩西 ，也会信我，因为他写过关于我的事。
JOHN|5|47|你们若不信他的书，怎能信我的话呢？”
JOHN|6|1|这些事以后，耶稣渡过 加利利海 ，就是 提比哩亚海 。
JOHN|6|2|有一大群人因为看见他在病人身上所行的神迹，就跟随他。
JOHN|6|3|耶稣上了山，和门徒一同坐在那里。
JOHN|6|4|那时 犹太 人的逾越节近了。
JOHN|6|5|耶稣举目看见一大群人来，就对 腓力 说：“我们到哪里去买饼给这些人吃呢？”
JOHN|6|6|他说这话是要考验 腓力 ，他自己原知道要怎样做。
JOHN|6|7|腓力 回答他：“就是两百个银币的饼也不够给他们每人吃一点点。”
JOHN|6|8|有一个门徒，就是 西门．彼得 的弟弟 安得烈 ，对耶稣说：
JOHN|6|9|“这里有一个孩子，带着五个大麦饼和两条鱼，但是分给这么多人还算什么呢？”
JOHN|6|10|耶稣说：“你们叫大家坐下。”那地方的草多，人们就坐下，男人的数目约有五千。
JOHN|6|11|耶稣拿起饼来，祝谢了，就分给坐着的人，也同样分了鱼，都照他们所要的来分。
JOHN|6|12|他们吃饱后，耶稣对门徒说：“把剩下的碎屑收拾起来，免得糟蹋了。”
JOHN|6|13|他们就把那五个大麦饼的碎屑，就是大家吃剩的，收拾起来，装满了十二个篮子。
JOHN|6|14|人们看见耶稣所行的神迹，就说：“这真是那要到世上来的先知！”
JOHN|6|15|耶稣知道他们要来强迫他作王，就独自又退到山上去了。
JOHN|6|16|到了晚上，他的门徒下到海边，
JOHN|6|17|上了船，要过海往 迦百农 去。天已经黑了，耶稣还没有来到他们那里。
JOHN|6|18|忽然狂风大作，海浪翻腾。
JOHN|6|19|门徒摇橹，约行了十里多 ，看见耶稣在海面上走，渐渐靠近了船，他们就害怕。
JOHN|6|20|耶稣对他们说：“是我，不要怕！”
JOHN|6|21|门徒就欣然接他上船，船立刻到了他们所要去的地方。
JOHN|6|22|第二天，留在海的对岸的众人发觉那里原来只有一条小船，而且耶稣没有同他的门徒上船，是门徒自己去的。
JOHN|6|23|另外有几条从 提比哩亚 来的小船，却停靠在主祝谢后给他们吃饼的地方附近。
JOHN|6|24|这时众人见耶稣和门徒都不在那里，就上了船，往 迦百农 去找耶稣。
JOHN|6|25|他们在海的对岸找到他后，对他说：“拉比，你几时到这里来的？”
JOHN|6|26|耶稣回答他们说：“我实实在在地告诉你们，你们找我，并不是因见了神迹，而是因吃饼吃饱了。
JOHN|6|27|不要为那会坏的食物操劳，而要为那存到永生的食物操劳。这食物是人子要赐给你们的，因为父上帝已印证了。”
JOHN|6|28|于是他们问他：“我们该做什么才算是做上帝的工作呢？”
JOHN|6|29|耶稣回答，对他们说：“信上帝所差来的，这就是上帝的工作。”
JOHN|6|30|于是他们对他说：“你行什么神迹，好让我们看见而信你呢？你到底要做什么呢？
JOHN|6|31|我们的祖宗在旷野吃过吗哪，如经上写着：‘他从天上赐下粮食来给他们吃。’”
JOHN|6|32|于是耶稣对他们说：“我实实在在地告诉你们，那从天上来的粮不是 摩西 赐给你们的，那从天上来的真粮是我父赐给你们的。
JOHN|6|33|因为上帝的粮就是那位从天上降下来，并且赐生命给世界的。”
JOHN|6|34|于是他们对他说：“主啊，请常常把这粮赐给我们！”
JOHN|6|35|耶稣对他们说：“我就是生命的粮。到我这里来的，绝不饥饿；信我的，永不干渴。
JOHN|6|36|可是，我告诉过你们，你们已经看见我 ，还是不信。
JOHN|6|37|凡父所赐给我的人，必到我这里来；到我这里来的，我总不丢弃他。
JOHN|6|38|因为我从天上降下来，不是要按自己的意愿行，而是要遵行差我来那位的旨意。
JOHN|6|39|差我来那位的旨意就是：他所赐给我的，要我一个也不失落，并且在末日使他复活。
JOHN|6|40|因为我父的旨意是要使每一个见了子而信的人得永生，并且在末日我要使他复活。”
JOHN|6|41|犹太 人因为耶稣说“我是从天上降下来的粮”，就私下议论他，
JOHN|6|42|说：“这不是 约瑟 的儿子耶稣吗？我们岂不认得他的父母吗？现在他怎么说‘我是从天上降下来的’呢？”
JOHN|6|43|耶稣回答，对他们说：“你们不要彼此私下议论。
JOHN|6|44|若不是差我来的父吸引人，就没有人能到我这里来；到我这里来的，在末日我要使他复活。
JOHN|6|45|在先知书上写着：‘他们都要蒙上帝教导。’凡听了父的教导而学习的，都到我这里来。
JOHN|6|46|这不是说有人看见过父，惟独从上帝来的，他才看见过父。
JOHN|6|47|我实实在在地告诉你们，信的人有永生。
JOHN|6|48|我就是生命的粮。
JOHN|6|49|你们的祖宗在旷野吃过吗哪，还是死了。
JOHN|6|50|这是从天上降下来的粮，使人吃了就不死。
JOHN|6|51|我就是从天上降下来生命的粮；人若吃这粮，必永远活着。我为世人的生命所赐下的粮就是我的肉。”
JOHN|6|52|因此， 犹太 人彼此争论说：“这个人怎能把他的肉给我们吃呢？”
JOHN|6|53|耶稣对他们说：“我实实在在地告诉你们，你们若不吃人子的肉，不喝人子的血，在你们里面就没有生命。
JOHN|6|54|吃我肉、喝我血的人就有永生，并且在末日我要使他复活。
JOHN|6|55|我的肉是真正可吃的；我的血是真正可喝的。
JOHN|6|56|吃我肉、喝我血的人常在我里面，我也常在他里面。
JOHN|6|57|永生的父怎样差我来，我又怎样因父活着，照样，吃我肉的人也要因我活着。
JOHN|6|58|这是从天上降下来的粮，不像你们的祖宗吃过吗哪还是死了；吃这粮的人将永远活着。”
JOHN|6|59|这些话是耶稣在 迦百农 会堂里教导人的时候说的。
JOHN|6|60|他的门徒中有好些人听见了，就说：“这话很难，谁听得进呢？”
JOHN|6|61|耶稣心里知道门徒为这话私下议论，就对他们说：“这话成了你们的绊脚石吗？
JOHN|6|62|如果你们看见人子升到他原来所在之处，会怎么样呢？
JOHN|6|63|圣灵赐人生命，肉体毫无用处。我对你们所说的话就是灵，就是生命。
JOHN|6|64|可是你们中间有些人不信。”耶稣起初就知道哪些人不信他，哪一个要出卖他。
JOHN|6|65|于是耶稣说：“所以，我对你们说过，若不是蒙我父的恩赐，没有人能到我这里来。”
JOHN|6|66|从此，他门徒中有很多退却了，不再和他同行。
JOHN|6|67|耶稣就对那十二使徒说：“你们也要离开吗？”
JOHN|6|68|西门．彼得 回答他：“主啊，你有永生之道，我们还跟从谁呢？
JOHN|6|69|我们已经信了，又知道你是上帝的圣者。”
JOHN|6|70|耶稣回答他们：“我不是拣选了你们十二个吗？但你们中间有一个是魔鬼。”
JOHN|6|71|耶稣这话是指着要出卖他的 加略 人 西门 的儿子 犹大 说的；他本是十二使徒里的一个。
JOHN|7|1|这些事以后，耶稣周游 加利利 ，不愿在 犹太 往来，因为 犹太 人想要杀他。
JOHN|7|2|这时 犹太 人的住棚节近了。
JOHN|7|3|耶稣的兄弟们对他说：“你离开这里上 犹太 去吧，好让你的门徒也看见你所做的事。
JOHN|7|4|因为人要扬名，没有在隐秘的地方行事的，如果你要做这些事，该把自己显明给世人看。”
JOHN|7|5|原来连他的兄弟们也不信他。
JOHN|7|6|于是耶稣对他们说：“我的时机还没有到，你们的时机却随时都有。
JOHN|7|7|世人不会恨你们，却是恨我，因为我指证他们的行为是恶的。
JOHN|7|8|你们上去过节吧！我现在不上去过这节 ，因为我的时机还没有成熟。”
JOHN|7|9|耶稣说了这些话，仍然留在 加利利 。
JOHN|7|10|但他的兄弟们上去过节以后，他也上去，不是公开去，却似乎 是秘密地去的。
JOHN|7|11|节期间， 犹太 人寻找耶稣，说：“他在哪里？”
JOHN|7|12|人群中有许多人对他议论纷纷，另有的说：“他是好人。”有的说：“不，他是迷惑群众的。”
JOHN|7|13|可是没有人公开谈论他，因为他们怕 犹太 人。
JOHN|7|14|节期已过了一半，耶稣上圣殿去教导人。
JOHN|7|15|犹太 人惊讶地说：“这个人没有学过，怎么那样熟悉经典呢？”
JOHN|7|16|于是耶稣回答他们，说：“我的教导不是我自己的，而是差我来那位的。
JOHN|7|17|人若立志要遵行上帝的旨意，就会知道这教导究竟是出于上帝，还是我凭着自己说的。
JOHN|7|18|凭着自己说的人是寻求自己的荣耀；但那寻求差他来那位的荣耀的人，他是真诚的，在他心里没有不义。
JOHN|7|19|摩西 不是传了律法给你们吗？你们却没有一个人守律法。为什么想要杀我呢？”
JOHN|7|20|众人回答：“你是被鬼附了！谁想要杀你呢？”
JOHN|7|21|耶稣回答，对他们说：“我做了一件事，你们都惊讶。
JOHN|7|22|摩西 传割礼给你们（其实割礼不是从 摩西 开始，而是从列祖开始的），你们就在安息日给人行割礼。
JOHN|7|23|人若在安息日受割礼，是为了不违背 摩西 的律法，我在安息日使一个人痊愈了，你们就向我发怒吗？
JOHN|7|24|不要凭外表断定是非，总要按公平断定是非。”
JOHN|7|25|于是 耶路撒冷 人中有的说：“这个人不是他们想要杀的吗？
JOHN|7|26|你看，他还公开讲道，他们也不对他说什么。难道官长真的认为这是基督吗？
JOHN|7|27|然而，我们知道这个人从哪里来；可是基督来的时候，没有人知道他从哪里来。”
JOHN|7|28|那时，耶稣在圣殿里教导人，喊着说：“你们认识我，也知道我从哪里来；我并不是凭着自己来的。但差我来的那位是真实的，你们不认识他。
JOHN|7|29|我却认识他，因为我从他那里来，是他差遣了我。”
JOHN|7|30|于是他们想要捉拿耶稣，只是没有人下手，因为他的时候还没有到。
JOHN|7|31|但人群中有好些人信他，他们说：“基督来的时候，他所行的神迹难道会比这人行的更多吗？”
JOHN|7|32|法利赛人听见群众对耶稣这样议论纷纷，祭司长和法利赛人就打发圣殿警卫去捉拿他。
JOHN|7|33|于是耶稣说：“我跟你们在一起的时候不会太久了，我要回到那差我来的那里去。
JOHN|7|34|你们要找我，却找不到；我所在的地方，你们不能去。”
JOHN|7|35|于是 犹太 人彼此问：“这人要往哪里去，使我们找不到他呢？难道他要往散居在 希腊 的 犹太 人那里去教导 希腊 人吗？
JOHN|7|36|他说‘你们要找我，却找不到；我所在的地方，你们不能去’这话是什么意思呢？”
JOHN|7|37|节期的最后一天，就是最隆重的一天，耶稣站着，喊着说：“人若渴了，到我这里来喝！
JOHN|7|38|信我的人，就如经上所说：‘从他腹中将流出活水的江河来。’”
JOHN|7|39|耶稣这话是指信他的人要受圣灵说的；那时还没有赐下圣灵，因为耶稣还没有得到荣耀。
JOHN|7|40|众人听见这些话，有的说：“这真是那先知。”
JOHN|7|41|另有的说：“这是基督。”但也有的说：“难道基督是出自 加利利 吗？
JOHN|7|42|经上不是说‘基督是 大卫 的后裔，出自 大卫 的本乡 伯利恒 ’吗？”
JOHN|7|43|于是众人因耶稣而分裂了。
JOHN|7|44|其中有人要捉拿他，只是没有人下手。
JOHN|7|45|警卫们回到祭司长和法利赛人那里。他们对警卫说：“你们为什么没有带他来呢？”
JOHN|7|46|警卫回答：“从来没有像他这样说话的！”
JOHN|7|47|于是法利赛人说：“你们也受了迷惑吗？
JOHN|7|48|难道官长或法利赛人中有信他的吗？
JOHN|7|49|但这些不明白律法的众人是被诅咒的！”
JOHN|7|50|其中有 尼哥德慕 ，就是从前去见过耶稣的，对他们说：
JOHN|7|51|“不先听本人的口供，查明他所做的事，难道我们的律法还定他的罪吗？”
JOHN|7|52|他们回答他说：“你也是出自 加利利 吗？你去查考就知道， 加利利 是不出先知的。” 〔
JOHN|7|53|于是各人都回家去了，
JOHN|8|1|耶稣却到 橄榄山 去。
JOHN|8|2|清早，他又回到圣殿里。众百姓都到他那里去，他就坐下，教导他们。
JOHN|8|3|文士和法利赛人带着一个犯奸淫时被捉的女人来，叫她站在当中，
JOHN|8|4|然后对耶稣说：“老师，这女人是正在犯奸淫的时候被捉到的。
JOHN|8|5|摩西 在律法书上命令我们把这样的女人用石头打死。那么，你怎么说呢？”
JOHN|8|6|他们说这话是要试探耶稣，要抓到控告他的把柄。耶稣却弯下腰，用指头在地上写字。
JOHN|8|7|他们还是不住地问他，耶稣就直起腰来，对他们说：“你们中间谁没有罪，谁就先拿石头打她！”
JOHN|8|8|于是他又弯着腰，用指头在地上写字。
JOHN|8|9|他们听见这话，从老的开始，一个一个都走开了，只剩下耶稣一人和那仍然站在中间的女人。
JOHN|8|10|耶稣就直起腰来，对她说：“妇人，那些人在哪里呢？没有任何人定你的罪吗？”
JOHN|8|11|她说：“主啊，没有。”耶稣说：“我也不定你的罪。去吧！从今以后不要再犯罪了。”〕
JOHN|8|12|耶稣又对众人说：“我就是世界的光。跟从我的，必不在黑暗里走，却要得着生命的光。”
JOHN|8|13|法利赛人对他说：“你是为自己作见证，你的见证不真。”
JOHN|8|14|耶稣回答他们，对他们说：“即使我为自己作见证，我的见证还是真的，因为我知道我从哪里来，到哪里去。你们却不知道我从哪里来，到哪里去。
JOHN|8|15|你们是以人的标准来判断人，我不判断任何人。
JOHN|8|16|即使我判断人，我的判断也是真确的，因为不是我独自在判断，而是差我来的父与我一同判断。
JOHN|8|17|你们的律法也记着说：‘两个人的见证才算为真’。
JOHN|8|18|我是为自己作见证，还有差我来的父也为我作见证。”
JOHN|8|19|于是他们问他：“你的父在哪里？”耶稣回答：“你们不认识我，也不认识我的父；若是认识我，也会认识我的父。”
JOHN|8|20|这些话是耶稣在圣殿的银库房里教导人的时候说的。当时没有人捉拿他，因为他的时候还没有到。
JOHN|8|21|于是耶稣又对他们说：“我去了，你们会找我，而你们会死在自己的罪中；我所去的地方，你们不能去。”
JOHN|8|22|犹太 人说：“他说‘我所去的地方，你们不能去’，难道他要自杀吗？”
JOHN|8|23|耶稣对他们说：“你们是从下面来的，我是从上面来的；你们是属这世界的，我不是属这世界的。
JOHN|8|24|所以我对你们说，你们会死在自己的罪中，你们若不信我就是那位，就会死在自己的罪中。”
JOHN|8|25|他们就问他：“你到底是谁？”耶稣对他们说：“我从起初就告诉你们了。
JOHN|8|26|我有许多事要讲论你们，判断你们；但差我来的那位是真实的，我从他那里所听见的，就告诉世人。”
JOHN|8|27|他们不明白耶稣是对他们讲父的事。
JOHN|8|28|所以耶稣说：“你们举起人子以后就会知道我就是那位了，并且知道我没有一件事是凭着自己做的。我说这些话是照着父所教导我的。
JOHN|8|29|差我来的那位与我同在；他没有撇下我独自一人，因为我一直行他所喜悦的事。”
JOHN|8|30|耶稣说这些话的时候，有许多人信了他。
JOHN|8|31|耶稣对信他的 犹太 人说：“你们若继续遵守我的道，就真是我的门徒了。
JOHN|8|32|你们将认识真理，真理会使你们自由。”
JOHN|8|33|他们回答他：“我们是 亚伯拉罕 的后裔，从来没有作过谁的奴隶，你怎么说‘会使你们自由’呢？”
JOHN|8|34|耶稣回答他们：“我实实在在地告诉你们，所有犯罪的人就是罪的奴隶。
JOHN|8|35|奴隶不能永远住在家里；儿子才永远住在家里。
JOHN|8|36|所以，上帝的儿子若使你们自由，你们就真正自由了。”
JOHN|8|37|“我知道，你们是 亚伯拉罕 的后裔，你们却想要杀我，因为你们心里容不下我的道。
JOHN|8|38|我所说的是在我父那里看见的；你们所做的是在你们的父那里听到的。”
JOHN|8|39|他们回答耶稣：“我们的父是 亚伯拉罕 。”耶稣对他们说：“你们若是 亚伯拉罕 的儿女，就会做 亚伯拉罕 所做的事。
JOHN|8|40|我把在上帝那里所听见的真理告诉了你们，现在你们却想要杀我； 亚伯拉罕 没有做过这样的事。
JOHN|8|41|你们是做你们父的工作。”他们就对他说：“我们不是从淫乱生的，我们只有一位父，就是上帝。”
JOHN|8|42|耶稣对他们说：“假如上帝是你们的父，你们会爱我，因为我本是出于上帝，也是从上帝而来，我不是凭着自己来，而是他差我来的。
JOHN|8|43|你们为什么不明白我的话呢？无非是你们听不进我的道。
JOHN|8|44|你们是出于你们的父魔鬼，你们宁愿随着你们父的欲念而行。他从起初就是杀人的，不守真理，因他心里没有真理。他说谎是出于自己的本性，因他本来是说谎的，也是说谎者之父。
JOHN|8|45|但是，因为我讲真理，你们就不信我。
JOHN|8|46|你们中间谁能指证我有罪呢？既然我讲真理，你们为什么不信我呢？
JOHN|8|47|出于上帝的，必听上帝的话；你们不听，因为你们不是出于上帝。”
JOHN|8|48|犹太 人回答他：“我们说你是 撒玛利亚 人，并且是被鬼附的，这话不是很对吗？”
JOHN|8|49|耶稣回答：“我没有被鬼附的；我尊敬我的父，你们却不尊敬我。
JOHN|8|50|我不寻求自己的荣耀，但有一位为我寻求荣耀，判断是非。
JOHN|8|51|我实实在在地告诉你们，人若遵守我的道，就永远不经历死亡。”
JOHN|8|52|于是 犹太 人对他说：“现在我们知道你是被鬼附了。 亚伯拉罕 死了，众先知也死了，你还说：‘人若遵守我的道，就永远不经历死亡。’
JOHN|8|53|难道你比我们的祖宗 亚伯拉罕 还大吗？他死了，众先知也死了，你把自己当作什么人呢？”
JOHN|8|54|耶稣回答：“我若荣耀自己，我的荣耀就算不了什么；荣耀我的是我的父，就是你们所说的你们的上帝。
JOHN|8|55|你们不认识他，我却认识他。我若说不认识他，我就是说谎的，像你们一样；但我认识他，也遵守他的道。
JOHN|8|56|你们的祖宗 亚伯拉罕 欢欢喜喜地仰望我的日子，他看见了，就快乐。”
JOHN|8|57|犹太 人就对他说：“你还没有五十岁，难道见过 亚伯拉罕 吗？”
JOHN|8|58|耶稣对他们说：“我实实在在地告诉你们，还没有 亚伯拉罕 我就存在了。”
JOHN|8|59|于是他们拿石头要打他，耶稣却躲开，走出了圣殿。
JOHN|9|1|耶稣往前走的时候，看见一个生来就失明的人。
JOHN|9|2|门徒问耶稣：“拉比，这人生来失明，是谁犯了罪？是这人还是他的父母呢？”
JOHN|9|3|耶稣回答：“既不是这人犯了罪，也不是他的父母，而是要在他身上显出上帝的作为来。
JOHN|9|4|趁着白日，我们 必须做差我 来的那位的工；黑夜来到，就没有人能做工了。
JOHN|9|5|我在世上的时候，是世上的光。”
JOHN|9|6|耶稣说了这些话，就吐唾沫在地上，用唾沫和了泥抹在盲人的眼睛上，
JOHN|9|7|对他说：“你到 西罗亚 池子里去洗。”（ 西罗亚 翻出来就是“奉差遣”。）于是他去，洗了，回来就看见了。
JOHN|9|8|他的邻舍和素常见他讨饭的人，就说：“这不是那从前坐着讨饭的人吗？”
JOHN|9|9|有的说：“是他”；又有的说：“不是，却是像他。”他自己说：“是我。”
JOHN|9|10|于是他们对他说：“你的眼睛是怎么开的呢？”
JOHN|9|11|那人回答：“有一个名叫耶稣的，他和了泥抹我的眼睛，对我说：‘你到 西罗亚 池子去洗。’我去一洗，就看见了。”
JOHN|9|12|他们对他说：“那个人在哪里？”他说：“我不知道。”
JOHN|9|13|他们把以前失明的那个人带到法利赛人那里。
JOHN|9|14|耶稣和泥开他眼睛的那一天是安息日。
JOHN|9|15|法利赛人又问他是怎么得看见的。他对他们说：“他把泥抹在我的眼睛上，我一洗，就看见了。”
JOHN|9|16|于是法利赛人中有的说：“这个人不是从上帝来的，因为他不守安息日。”另有的说：“一个罪人怎能行这样的神迹呢？”他们之间就产生了分裂。
JOHN|9|17|于是他们又对那盲人说：“他开了你的眼睛，你说他是怎样的人呢？”他说：“他是个先知。”
JOHN|9|18|犹太 人不信他以前是失明，后来能看见的，等到叫了他的父母来，
JOHN|9|19|问他们说：“这是你们的儿子吗？你们说他生来是失明的，现在怎么看见了呢？”
JOHN|9|20|他的父母就回答说：“他是我们的儿子，生来就失明，这是我们知道的。
JOHN|9|21|至于他现在怎么能看见，我们却不知道；是谁开了他的眼睛，我们也不知道。他已经是成人，你们问他吧，他自己会说。”
JOHN|9|22|他父母说这些话，是怕 犹太 人，因为 犹太 人已经商定，若有宣认耶稣是基督的，要把他赶出会堂。
JOHN|9|23|因此他父母说“他已经是成人，你们问他吧”。
JOHN|9|24|于是法利赛人第二次叫了那以前失明的人来，对他说：“你要将荣耀归给上帝，我们知道这人是个罪人。”
JOHN|9|25|那人就回答：“他是不是个罪人，我不知道；有一件事我知道，我本来是失明的，现在我看见了。”
JOHN|9|26|他们就问他：“他给你做了什么？是怎么开了你的眼睛？”
JOHN|9|27|他回答他们：“我已经告诉你们了，你们不听，为什么又要听呢？难道你们也要作他的门徒吗？”
JOHN|9|28|他们就骂他：“你是他的门徒，而我们是 摩西 的门徒。
JOHN|9|29|上帝对 摩西 说话是我们知道的，可是这个人，我们不知道他从哪里来。”
JOHN|9|30|那人回答，对他们说：“他开了我的眼睛，你们竟不知道他从哪里来，这真是奇怪！
JOHN|9|31|我们知道上帝不听罪人，惟有敬奉上帝、遵行他旨意的，上帝才听他。
JOHN|9|32|从创世以来，未曾听见有人开了生来就失明的人的眼睛。
JOHN|9|33|这人若不是从上帝来的，什么也不能做。”
JOHN|9|34|他们回答他说：“你完全是生在罪中的，还要来教训我们吗？”于是他们把他赶出去了。
JOHN|9|35|耶稣听说他们把他赶出去，就找到他，说：“你信人子 吗？”
JOHN|9|36|那人回答说：“主啊，人子是谁？告诉我，好让我信他。”
JOHN|9|37|耶稣对他说：“你已经看见他，现在和你说话的就是他。”
JOHN|9|38|他说：“主啊，我信！”他就拜耶稣。
JOHN|9|39|耶稣说：“我为审判到这世上来，使不能看见的看见，能看见的反而失明。”
JOHN|9|40|同他在那里的法利赛人听见这些话，就对他说：“难道我们也失明了吗？”
JOHN|9|41|耶稣对他们说：“你们若是失明的，就没有罪了；但现在你们说‘我们能看见’，你们的罪还在。”
JOHN|10|1|“我实实在在地告诉你们，那不从门进羊圈，倒从别处爬进去的，就是贼，就是强盗。
JOHN|10|2|那从门进去的才是羊的牧人。
JOHN|10|3|看门的给他开门，羊也听他的声音。他按著名叫自己的羊，把羊领出来。
JOHN|10|4|当他把自己的羊都放出来，就走在前面，羊也跟着他，因为它们认得他的声音。
JOHN|10|5|羊绝不跟陌生人，反而会逃走，因为不认得陌生人的声音。”
JOHN|10|6|耶稣把这比方告诉他们，但他们不明白他所说的是什么。
JOHN|10|7|所以，耶稣又对他们说：“我实实在在地告诉你们，我就是羊的门。
JOHN|10|8|凡在我以前 来的都是贼，是强盗；羊没有听从他们。
JOHN|10|9|我就是门，凡从我进来的，必得安全 ，并且可进出，找到草吃。
JOHN|10|10|盗贼来，无非要偷窃，杀害，毁坏；我来了，是要羊得生命，并且得的更丰盛。
JOHN|10|11|“我是好牧人，好牧人为羊舍命。
JOHN|10|12|雇工不是牧人，羊不是他自己的，他一看见狼来，就撇下羊群逃跑；狼抓住羊，把它们赶散。
JOHN|10|13|雇工逃走，因为他是雇工，对羊毫不关心。
JOHN|10|14|我是好牧人；我认识我的羊，我的羊也认识我，
JOHN|10|15|正如父认识我，我也认识父一样；并且我为羊舍命。
JOHN|10|16|我另外有羊，不属这圈里的，我必须领它们来，它们也要听我的声音，并且要合成一群，归一个牧人。
JOHN|10|17|为此，我父爱我，因为我把命舍去，好再取回来。
JOHN|10|18|没有人夺去我的命，是我自己舍的；我有权舍弃，也有权再取回。这是我从我父所受的命令。”
JOHN|10|19|犹太 人为这些话又起了分裂。
JOHN|10|20|其中有好些人说：“他是被鬼附了，而且疯了，为什么听他的呢？”
JOHN|10|21|另有的说：“这不是被鬼附的人所说的话。鬼岂能开盲人的眼睛呢？”
JOHN|10|22|那时正是冬天，在 耶路撒冷 有献殿节。
JOHN|10|23|耶稣在圣殿里的 所罗门 廊下行走。
JOHN|10|24|犹太 人围着他，对他说：“你让我们犹豫不定到几时呢？你若是基督，就明白地告诉我们。”
JOHN|10|25|耶稣回答他们：“我已经告诉你们，你们却不信。我奉我父的名所行的事可以为我作见证。
JOHN|10|26|但是你们不信，因为你们不是我的羊。
JOHN|10|27|我的羊听我的声音，我认识它们，它们也跟从我。
JOHN|10|28|并且，我赐给他们永生；他们永不灭亡，谁也不能从我手里把他们夺去。
JOHN|10|29|我父所赐给我的比万有都大 ，谁也不能从我父手里把他们夺去。
JOHN|10|30|我与父原为一。”
JOHN|10|31|犹太 人又拿起石头来要打他。
JOHN|10|32|耶稣回应他们：“我做了许多从父那里来的善事给你们看，你们是为哪一件拿石头打我呢？”
JOHN|10|33|犹太 人回答他：“我们不是为了善事拿石头打你，而是为了你说亵渎的话；因为你是个人，却把自己当作上帝。”
JOHN|10|34|耶稣回答他们：“你们的律法书上不是写着‘我曾说你们是诸神’吗？
JOHN|10|35|经上的话是不能废的；如果那些领受上帝的道的人，上帝尚且称他们为诸神，
JOHN|10|36|那么父所分别为圣又差到世上来的那位说‘我是上帝的儿子’，你们还对他说‘你说亵渎的话’吗？
JOHN|10|37|我若不做我父的工作，你们就不必信我；
JOHN|10|38|我若做了，你们即使不信我，也当信这些工作，好让你们知道并且明白父在我里面，我也在父里面。”
JOHN|10|39|于是，他们又要捉拿他，他却从他们手中逃脱了。
JOHN|10|40|耶稣又往 约旦河 的东边去，到了 约翰 起初施洗的地方，就住在那里。
JOHN|10|41|有许多人来到他那里，说：“ 约翰 没有行过一件神迹，但 约翰 所说有关这人的一切话都是真的。”
JOHN|10|42|在那里，许多人信了耶稣。
JOHN|11|1|有一个患病的人，名叫 拉撒路 ，住在 伯大尼 ，就是 马利亚 和她姐姐 马大 的村庄。
JOHN|11|2|这 马利亚 就是那用香膏抹主，又用头发擦他脚的；患病的 拉撒路 是她的弟弟。
JOHN|11|3|姊妹两个就打发人去见耶稣，说：“主啊，你所爱的人病了。”
JOHN|11|4|耶稣听见后却说：“这病不至于死，而是为了上帝的荣耀，为要使上帝的儿子藉此得荣耀。”
JOHN|11|5|耶稣素来爱 马大 和她妹妹，以及 拉撒路 。
JOHN|11|6|他听见 拉撒路 病了，仍在原地住了两天，
JOHN|11|7|然后对门徒说：“我们再到 犹太 去吧！”
JOHN|11|8|门徒对他说：“拉比， 犹太 人近来要拿石头打你，你还再到那里去吗？”
JOHN|11|9|耶稣回答：“白天不是有十二小时吗？人若在白天行走，就不致跌倒，因为他看见这世上的光。
JOHN|11|10|人若在黑夜行走，就会跌倒，因为他没有光。”
JOHN|11|11|耶稣说了这些话，随后对他们说：“我们的朋友 拉撒路 睡了，我去叫醒他。”
JOHN|11|12|门徒就说：“主啊，他若睡了，就会好的。”
JOHN|11|13|耶稣说这话是指 拉撒路 死了，他们却以为他是指通常的睡眠。
JOHN|11|14|于是耶稣就明白地告诉他们：“ 拉撒路 死了。
JOHN|11|15|为了你们的缘故，我不在那里反而欢喜，为要使你们信。现在我们到他那里去吧。”
JOHN|11|16|于是那称为 低土马 的 多马 对其他的门徒说：“我们也去和他同死吧！”
JOHN|11|17|耶稣到了，知道 拉撒路 在坟墓里已经四天了。
JOHN|11|18|伯大尼 离 耶路撒冷 不远，约有六里 路。
JOHN|11|19|有好些 犹太 人来看 马大 和 马利亚 ，要为她们弟弟的缘故安慰她们。
JOHN|11|20|马大 听见耶稣来了，就出去迎接他； 马利亚 却仍然坐在家里。
JOHN|11|21|马大 对耶稣说：“主啊，你若早在这里，我弟弟就不会死了。
JOHN|11|22|我也知道，即使现在，你无论向上帝求什么，上帝也必赐给你。”
JOHN|11|23|耶稣对她说：“你弟弟会复活的。”
JOHN|11|24|马大 对他说：“我知道在末日复活的时候，他会复活。”
JOHN|11|25|耶稣对她说：“复活...也在我 。信我的人虽然死了，也必复活；
JOHN|11|26|凡活着信我的人必永远不死。你信这话吗？”
JOHN|11|27|马大 对他说：“主啊，是的。我信你是基督，是上帝的儿子，就是那要临到世界的。”
JOHN|11|28|马大 说了这话就回去，叫她妹妹 马利亚 ，私下说：“老师来了，他在叫你。”
JOHN|11|29|马利亚 听见了，急忙起来，到耶稣那里去。
JOHN|11|30|那时，耶稣还没有进村子，仍在 马大 迎接他的地方。
JOHN|11|31|那些同 马利亚 在家里安慰她的 犹太 人，见她急忙起来，出去，就跟着她，以为她要往坟墓那里去哭。
JOHN|11|32|马利亚 到了耶稣那里，看见他，就俯伏在他脚前，对他说：“主啊，你若早在这里，我弟弟就不会死了。”
JOHN|11|33|耶稣看见她哭，并看见与她同来的 犹太 人也哭，就心里悲叹，又甚忧愁，
JOHN|11|34|就说：“你们把他安放在哪里？”他们对他说：“主啊，请你来看。”
JOHN|11|35|耶稣哭了。
JOHN|11|36|犹太 人就说：“你看，他多么爱他！”
JOHN|11|37|其中有人说：“他既然开了盲人的眼睛，难道不能叫这人不死吗？”
JOHN|11|38|耶稣又心里悲叹，来到坟墓前。那坟墓是个穴，有一块石头挡着。
JOHN|11|39|耶稣说：“把石头挪开！”那死者的姐姐 马大 对他说：“主啊，他现在必定臭了，因为他已经死了四天了。”
JOHN|11|40|耶稣对她说：“我不是对你说过，你若信就必看见上帝的荣耀吗？”
JOHN|11|41|于是他们把石头挪开。耶稣举目望天，说：“父啊，我感谢你，因为你已经听了我。
JOHN|11|42|我知道你常常听我，但我说这话是为了周围站着的众人，要使他们信是你差了我来的。”
JOHN|11|43|说了这些话，他大声呼叫说：“ 拉撒路 ，出来！”
JOHN|11|44|那死了的人就出来了，手脚都裹着布，脸上包着头巾。耶稣对他们说：“解开他，让他走！”
JOHN|11|45|于是来看 马利亚 的 犹太 人中，有很多人见了耶稣所做的事，就信了他。
JOHN|11|46|但其中也有人去见法利赛人，把耶稣所做的事告诉他们。
JOHN|11|47|祭司长和法利赛人召开议会，说：“这人行好些神迹，我们怎么办呢？
JOHN|11|48|若让他这样做，人人都要信他； 罗马 人也要来毁灭我们的圣殿 和我们的民族。”
JOHN|11|49|其中有一个人，名叫 该亚法 ，那年当大祭司，对他们说：“你们什么都不知道，
JOHN|11|50|也不想想，一个人替百姓死，免得整个民族灭亡，这对你们是有利的。”
JOHN|11|51|他这话不是出于自己的意思，而是因他那年当大祭司，所以预言耶稣将为这民族而死。
JOHN|11|52|他不但替这民族死，还要把上帝四散的儿女都聚集起来，合成一群。
JOHN|11|53|从那日起，他们就商议要杀耶稣。
JOHN|11|54|所以，耶稣不再公开在 犹太 人中走动，却离开那里，往靠近旷野的乡间去，到了一座城，名叫 以法莲 ，就在那里和门徒住下来。
JOHN|11|55|犹太 人的逾越节近了，有许多人从乡下上 耶路撒冷 去，要在过节前洁净自己。
JOHN|11|56|于是他们寻找耶稣，站在圣殿里彼此说：“你们认为怎样，他不会来过节吧？”
JOHN|11|57|那时，祭司长和法利赛人早已下令，若有人知道耶稣的下落，就要报告，他们好去捉拿他。
JOHN|12|1|逾越节前六天，耶稣来到 伯大尼 ，就是他使 拉撒路 从死人中复活的地方。
JOHN|12|2|有人在那里为耶稣预备宴席； 马大 伺候， 拉撒路 也在同耶稣坐席的人中间。
JOHN|12|3|马利亚 拿着一斤极贵的纯哪哒 香膏，抹耶稣的脚，又用自己头发去擦，屋里充满了膏的香气。
JOHN|12|4|有一个门徒，就是那将要出卖耶稣的 加略 人 犹大 ，说：
JOHN|12|5|“为什么不把这香膏卖三百个银币去周济穷人呢？”
JOHN|12|6|他说这话，并不是关心穷人，而是因为他是个贼，又管钱囊，常偷取钱囊中所存的。
JOHN|12|7|耶稣说：“由她吧！她这香膏本是为我的安葬之日留着的。
JOHN|12|8|因为常有穷人和你们在一起，但是你们不常有我。”
JOHN|12|9|有一大群 犹太 人知道耶稣在那里，就来了，不但是为耶稣的缘故，也是要看耶稣使他从死人中复活的 拉撒路 。
JOHN|12|10|于是众祭司长商议连 拉撒路 也要杀了，
JOHN|12|11|因为有许多 犹太 人为了 拉撒路 的缘故，开始背离他们，信了耶稣。
JOHN|12|12|第二天，有一大群上来过节的人听见耶稣要来 耶路撒冷 ，
JOHN|12|13|就拿着棕树枝出去迎接他，喊着： “和散那 ， 以色列 的王！ 奉主名来的是应当称颂的！”
JOHN|12|14|耶稣找到了一匹驴驹，就骑上，如经上所记：
JOHN|12|15|“ 锡安 的儿女 啊，不要惧怕！ 看哪，你的王来了； 他骑在驴驹上。”
JOHN|12|16|门徒当初不明白这些事，等到耶稣得了荣耀后才想起这些话是指他写的，并且人们果然对他做了这些事。
JOHN|12|17|当耶稣呼唤 拉撒路 ，使他从死人中复活出坟墓的时候，同耶稣在那里的众人就作见证。
JOHN|12|18|众人因听见耶稣行了这神迹，就去迎接他。
JOHN|12|19|法利赛人彼此说：“你们看，你们一事无成，世人都随着他去了。”
JOHN|12|20|那时，上来过节礼拜的人中，有几个 希腊 人。
JOHN|12|21|他们来见 加利利 的 伯赛大 人 腓力 ，请求他说：“先生，我们想见耶稣。”
JOHN|12|22|腓力 去告诉 安得烈 ，然后 安得烈 同 腓力 去告诉耶稣。
JOHN|12|23|耶稣回答他们说：“人子得荣耀的时候到了。
JOHN|12|24|我实实在在地告诉你们，一粒麦子不落在地里死了，仍旧是一粒；若是死了，就结出许多子粒来。
JOHN|12|25|爱惜自己性命的，就丧失性命；那恨恶自己在这世上的性命的，要保全性命到永生。
JOHN|12|26|若有人服事我，就当跟从我；我在哪里，服事我的人也要在哪里；若有人服事我，我父必尊重他。”
JOHN|12|27|“我现在心里忧愁，我说什么才好呢？说‘父啊，救我脱离这时候’吗？但我正是为这时候来的。
JOHN|12|28|父啊，愿你荣耀你的名！”于是有声音从天上来，说：“我已经荣耀了我的名，还要再荣耀。”
JOHN|12|29|站在旁边的众人听见，就说：“打雷了。”另有的说：“有天使对他说话。”
JOHN|12|30|耶稣回答说：“这声音不是为我，而是为你们来的。
JOHN|12|31|现在正是这世界受审判的时候；现在这世界的统治者要被赶出去。
JOHN|12|32|我从地上被举起来的时候，我要吸引万人来归我。”
JOHN|12|33|耶稣这话是指自己将要怎样死说的。
JOHN|12|34|众人就回答他：“我们听见律法书上说，基督是永存的；你怎么说，人子必须被举起来呢？这人子是谁呢？”
JOHN|12|35|耶稣对他们说：“光在你们中间为时不多了，应该趁着有光的时候行走，免得黑暗临到你们；那在黑暗里行走的，不知道往何处去。
JOHN|12|36|你们趁着有光，要信从这光，使你们成为光明之子。” 耶稣说了这些话，就离开他们隐藏了。
JOHN|12|37|他虽然在他们面前行了许多神迹，他们还是不信他。
JOHN|12|38|这是要应验 以赛亚 先知所说的话： “主啊，我们所传的有谁信呢？ 主的膀臂向谁显露呢？”
JOHN|12|39|他们所以不能信，因为 以赛亚 又说：
JOHN|12|40|“主使他们瞎了眼， 使他们硬了心， 免得他们眼睛看见， 他们心里明白，回转过来， 我会医治他们。”
JOHN|12|41|以赛亚 因看见了他的荣耀，就说了关于他的这话。
JOHN|12|42|虽然如此，官长中却有好些信他的，只因法利赛人的缘故不敢承认，恐怕被赶出会堂。
JOHN|12|43|这是因他们爱人给的尊荣过于爱上帝给的尊荣。
JOHN|12|44|耶稣喊着说：“信我的人不是信我，而是信差我来的那位。
JOHN|12|45|看见我的，就是看见差我来的那位。
JOHN|12|46|我就是来到世上的光，使凡信我的不住在黑暗里。
JOHN|12|47|若有人听见我的话而不遵守，我不审判他，因为我来不是要审判世人，而是要拯救世人。
JOHN|12|48|弃绝我、不领受我话的人自有审判他的；我所讲的道在末日要审判他。
JOHN|12|49|因为我没有凭着自己讲，而是差我来的父已经给我命令，叫我说什么，讲什么。
JOHN|12|50|我也知道他的命令就是永生。所以，我讲的正是照着父所告诉我的，我就这么讲了。”
JOHN|13|1|逾越节以前，耶稣知道自己离世归父的时候到了。他一向爱世间属自己的人，就爱他们到底。
JOHN|13|2|晚餐的时候，魔鬼已把出卖耶稣的意思放在 加略 人 西门 的儿子 犹大 心里。
JOHN|13|3|耶稣知道父已把万有交在他手里，且知道自己是从上帝出来的，又要回到上帝那里去，
JOHN|13|4|就离席站起来，脱了衣服，拿一条手巾束腰，
JOHN|13|5|随后把水倒在盆里，开始洗门徒的脚，并用束腰的手巾擦干。
JOHN|13|6|到了 西门．彼得 跟前， 彼得 对他说：“主啊，你洗我的脚吗？”
JOHN|13|7|耶稣回答他说：“我所做的，你现在不知道，但以后会明白。”
JOHN|13|8|彼得 对他说：“你绝对不可以洗我的脚！”耶稣回答他：“我若不洗你，你就与我无份了。”
JOHN|13|9|西门．彼得 对他说：“主啊，不仅是我的脚，连手和头也要洗！”
JOHN|13|10|耶稣对他说：“凡洗过澡的人不需要再洗，只要把脚一洗，全身就干净了。你们是干净的，然而不都是干净的。”
JOHN|13|11|耶稣已知道要出卖他的是谁，因此说“你们不都是干净的”。
JOHN|13|12|耶稣洗完了他们的脚，就穿上衣服，又坐下，对他们说：“我为你们所做的，你们明白吗？
JOHN|13|13|你们称呼我老师，称呼我主，你们说的不错，我本来就是。
JOHN|13|14|我是你们的主，你们的老师，尚且洗你们的脚，你们也应当彼此洗脚。
JOHN|13|15|我给你们作了榜样，为要你们照着我为你们所做的去做。
JOHN|13|16|我实实在在地告诉你们，仆人不大于主人；奉差的人也不大于差他的人。
JOHN|13|17|你们既知道这些事，若是去实行就有福了。
JOHN|13|18|我不是指着你们众人说的，我知道我所拣选的是谁；但是要应验经上的话：‘吃我饭的人 用脚踢我。’
JOHN|13|19|事情还没有发生，我现在先告诉你们，让你们到事情发生的时候好信我就是那位。
JOHN|13|20|我实实在在地告诉你们，接纳我所差遣的就是接纳我；接纳我的就是接纳差遣我的那位。”
JOHN|13|21|耶稣说了这些话，心里忧愁，于是明确地说：“我实实在在地告诉你们，你们中间有一个人要出卖我。”
JOHN|13|22|门徒彼此相看，猜不出他说的是谁。
JOHN|13|23|门徒中有一个人，是耶稣所爱的，侧身挨近耶稣的胸怀。
JOHN|13|24|西门．彼得 就对这个人示意，要问耶稣是指着谁说的。
JOHN|13|25|于是那人紧靠着耶稣的胸膛，问他：“主啊，是谁呢？”
JOHN|13|26|耶稣回答：“我蘸一点饼给谁，就是谁。”耶稣就蘸了一点饼，递给 加略 人 西门 的儿子 犹大 。
JOHN|13|27|他接 了那饼以后，撒但就进入他的心。于是耶稣对他说：“你要做的，快做吧！”
JOHN|13|28|同席的人没有一个知道耶稣为什么对他说这话。
JOHN|13|29|有人因 犹大 管钱囊，以为耶稣是对他说“你去买我们过节所需要的东西”，或是叫他拿些什么给穷人。
JOHN|13|30|犹大 受 了那点饼以后立刻出去。那时候是夜间了。
JOHN|13|31|犹大 出去后，耶稣说：“如今人子得了荣耀，上帝在人子身上也得了荣耀。
JOHN|13|32|如果上帝因人子得了荣耀 ，上帝也要因自己荣耀人子，并且要立刻荣耀他。
JOHN|13|33|孩子们！我与你们同在的时候不多了；你们会找我，但我所去的地方，你们不能去。这话我曾对 犹太 人说过，现在也照样对你们说。
JOHN|13|34|我赐给你们一条新命令，乃是叫你们彼此相爱；我怎样爱你们，你们也要怎样彼此相爱。
JOHN|13|35|你们若彼此相爱，众人因此就认出你们是我的门徒了。”
JOHN|13|36|西门．彼得 问耶稣：“主啊，你去哪里？”耶稣回答：“我所去的地方，你现在不能跟我去，以后却要跟我去。”
JOHN|13|37|彼得 对他说：“主啊，为什么我现在不能跟你去？我愿意为你舍命。”
JOHN|13|38|耶稣回答：“你愿意为我舍命吗？我实实在在地告诉你，鸡叫以前，你要三次不认我。”
JOHN|14|1|“你们心里不要忧愁；你们信上帝，也当信我。
JOHN|14|2|在我父的家里有许多住处；若是没有，我就早已告诉你们了。我去原是为你们预备地去方。
JOHN|14|3|我若去为你们预备了地方，就必再来接你们到我那里去，我在哪里，叫你们也在哪里。
JOHN|14|4|我往哪里去，你们知道那条路。”
JOHN|14|5|多马 对他说：“主啊，我们不知道你去哪里，怎么能知道那条路呢？”
JOHN|14|6|耶稣对他说：“我就是道路、真理、生命；若不藉着我，没有人能到父那里去。
JOHN|14|7|既然你们认识了我，也会认识我的父。从今以后，你们就认识他，并且已经看见他了。”
JOHN|14|8|腓力 对他说：“主啊，将父显给我们看，我们就知足了。”
JOHN|14|9|耶稣对他说：“ 腓力 ，我与你们在一起这么久了，你还不认识我吗？看见我的就是看见了父，你怎么还说‘将父显给我们看’呢？
JOHN|14|10|我在父里面，父在我里面，你不信吗？我对你们所说的话不是凭着自己说的，而是住在我里面的父在做他的工作。
JOHN|14|11|你们要信我，我在父里面，父在我里面；即使不信，也要因我所做的工作信我。
JOHN|14|12|我实实在在地告诉你们，我所做的工作，信我的人也要做，并且要做得比这些更大，因为我到父那里去。
JOHN|14|13|你们奉我的名无论求什么，我必成全，为了使父因儿子得荣耀。
JOHN|14|14|你们若奉我的名向我求什么，我必成全。”
JOHN|14|15|“你们若爱我，就会遵守我的命令。
JOHN|14|16|我要求父，父就赐给你们另外一位保惠师 ，使他永远与你们同在。
JOHN|14|17|他就是真理的灵，是世人不能接受的。因为他们既看不见他，也不认识他；你们却认识他，因他常与你们同在，也要在你们里面。
JOHN|14|18|我不会撇下你们为孤儿，我必到你们这里来。
JOHN|14|19|再过不久，世人不再看见我，你们却会看见我，因为我活着，你们也要活着。
JOHN|14|20|到那日，你们就会知道我在父里面，你们在我里面，我也在你们里面。
JOHN|14|21|有了我的命令而又遵守的人，就是爱我的；爱我的人，我父要爱他，我也要爱他，并且要亲自向他显现。”
JOHN|14|22|犹大 （不是 加略 人 犹大 ）问耶稣：“主啊，为什么亲自向我们显现，而不向世人显现呢？”
JOHN|14|23|耶稣回答他说：“凡爱我的人就会遵守我的道，我父也会爱他，并且我们要到他那里去，与他同住。
JOHN|14|24|不爱我的人就不遵守我的道。你们所听见的道不是我的，而是差我来之父的。
JOHN|14|25|“我还与你们在一起的时候，已对你们说了这些事。
JOHN|14|26|但保惠师，就是父因我的名所要差来的圣灵，他要把一切的事教导你们，并且要使你们想起我对你们所说的一切话。
JOHN|14|27|我留下平安给你们，我把我的平安赐给你们。我所赐给你们的，不像世人所赐的。你们心里不要忧愁，也不要胆怯。
JOHN|14|28|你们听见我对你们说过，我去了还要回到你们这里来。你们若爱我，就会因我到父那里去而喜乐，因为父比我大。
JOHN|14|29|现在事情还没有发生，我预先告诉你们，使你们在事情发生的时候会信。
JOHN|14|30|我不再和你们多说了，因为这世界的统治者将到，他在我身上一无所能。
JOHN|14|31|我这么做是照着父命令我的，为了让世人知道我爱父。起来，我们走吧！”
JOHN|15|1|“我就是真葡萄树，我父是栽培的人。
JOHN|15|2|凡属我不结果子的枝子，他就剪掉；凡结果子的，他就修剪干净，使枝子结果子更多。
JOHN|15|3|现在你们因我讲给你们的道已经洁净了。
JOHN|15|4|你们要常在我里面，我也常在你们里面。枝子若不常在葡萄树上，自己就不能结果子；你们若不常在我里面，也是这样。
JOHN|15|5|我就是葡萄树，你们是枝子。常在我里面的，我也常在他里面，这人就多结果子，因为离了我，你们就不能做什么。
JOHN|15|6|人若不常在我里面，就像枝子被丢在外面，枯干了，人捡起来，扔进火里烧了。
JOHN|15|7|你们若常在我里面，我的话也常在你们里面，凡你们想要的，祈求，就给你们成全。
JOHN|15|8|你们多结果子，我父就因此得荣耀，你们也就是 我的门徒了。
JOHN|15|9|我爱你们，正如父爱我一样；你们要常在我的爱里。
JOHN|15|10|你们若遵守我的命令，就会常在我的爱里，正如我遵守了我父的命令，常在他的爱里。
JOHN|15|11|“我已对你们说了这些事，是要让我的喜乐存在你们心里，并让你们的喜乐得以满足。
JOHN|15|12|你们要彼此相爱，像我爱你们一样，这是我的命令。
JOHN|15|13|人为朋友舍命，人的爱心没有比这个更大的了。
JOHN|15|14|你们若遵行我所命令的，就是我的朋友。
JOHN|15|15|以后我不再称你们为仆人，因为仆人不知道主人所做的事；但我称你们为朋友，因为我从我父所听见的一切都已经让你们知道了。
JOHN|15|16|不是你们拣选了我，而是我拣选了你们，并且派你们去结果子，让你们的果子得以长存，好使你们奉我的名，无论向父求什么，他会赐给你们。
JOHN|15|17|我这样命令你们，是要你们彼此相爱。”
JOHN|15|18|“世人若恨你们，你们要知道，他们在恨你们以前已经恨我了。
JOHN|15|19|你们若属世界，世界会爱属自己的；只因你们不属世界，而是我从世界中拣选了你们，所以世界就恨你们。
JOHN|15|20|你们要记得我对你们说过的话：‘仆人不大于主人。’他们若迫害了我，也会迫害你们，他们若遵守了我的话，也会遵守你们的话。
JOHN|15|21|但他们要因我的名向你们做这一切的事，因为他们不认识差我来的那位。
JOHN|15|22|我若没有来教导他们，他们就没有罪；但如今他们的罪无可推诿了。
JOHN|15|23|恨我的也恨我的父。
JOHN|15|24|我若没有在他们中间做过别人未曾做的事，他们就没有罪；但如今连我与我的父，他们也看见了，也恨恶了。
JOHN|15|25|这是要应验他们律法上所写的话：‘他们无故地恨我。’
JOHN|15|26|“但我要从父那里差保惠师来，就是从父出来的那真理的灵，他来的时候要为我作见证。
JOHN|15|27|你们也要作见证，因为你们从起初就与我同在。”
JOHN|16|1|“我对你们说了这些事，是要使你们不至于跌倒。
JOHN|16|2|人要把你们赶出会堂，而且时候将到，凡杀你们的还以为是在事奉上帝。
JOHN|16|3|他们这样做，是因为没有认识父，也没有认识我。
JOHN|16|4|我对你们说了这些事，是要在他们做这些事的时候，你们会想起我对你们说过的话。” “我起先没有对你们说这些事，因为我一直与你们同在。
JOHN|16|5|现在我要到差我来的父那里去，你们中间却没有人问我‘你去哪里？’
JOHN|16|6|只因我对你们说了这些事，你们就满心忧愁。
JOHN|16|7|然而，我把真情告诉你们，我去对你们是有益的。我若不去，保惠师就不会到你们这里来；我若去，就差他到你们这里来。
JOHN|16|8|他来的时候，要为罪、为义，为审判，指证世人；
JOHN|16|9|为罪，是因他们不信我；
JOHN|16|10|为义，是因我到父那里去，你们将不再见到我；
JOHN|16|11|为审判，是因这世界的统治者已受了审判。
JOHN|16|12|“我还有好些事要告诉你们，但你们现在担当不了 。
JOHN|16|13|但真理的灵来的时候，他要引导你们进入一切真理。因为他不是凭着自己说的，而是把他所听见的都说出来，并且要把将要来的事向你们传达。
JOHN|16|14|他要荣耀我，因为他要把从我领受的向你们传达。
JOHN|16|15|凡父所有的都是我的，所以我说，他要把从我领受的向你们传达。”
JOHN|16|16|“不久，你们将不再见到我；再过不久，你们还要见到我。”
JOHN|16|17|有几个门徒彼此说：“他对我们说‘不久，你们将不再见到我；再过不久，你们还要见到我’；又说‘因我到父那里去’。这是什么意思呢？”
JOHN|16|18|于是门徒说：“他说 ‘不久’到底是什么意思呢？我们不明白他说什么。”
JOHN|16|19|耶稣看出他们要问他，就对他们说：“我说‘不久，你们将不再见到我；再过不久，你们还要见到我’，你们为这话彼此询问吗？
JOHN|16|20|我实实在在地告诉你们，你们将要痛哭，哀号，世人反要欢喜。你们将要忧愁，然而你们的忧愁要变成喜乐。
JOHN|16|21|妇人生产的时候会忧愁，因为她的时候到了；但孩子一生出来，就不再记得那痛苦了，因为欢喜有一个人生在世上了。
JOHN|16|22|你们现在也是忧愁，但我要再见到你们，你们的心就会有喜乐了；这喜乐没有人能夺去。
JOHN|16|23|到那日，你们什么也不会问我了。我实实在在地告诉你们，你们奉我的名无论向父求什么，他会赐给你们 。
JOHN|16|24|直到现在，你们没有奉我的名求什么，如今你们求就必得着，使你们的喜乐得以满足。”
JOHN|16|25|“这些事，我是用比方对你们说的；时候将到，我不再用比方对你们说，而是要把父的事明白地告诉你们。
JOHN|16|26|到那日，你们要奉我的名祈求；我并不对你们说，我要为你们向父祈求。
JOHN|16|27|父自己爱你们，因为你们已经爱我，又信我是从上帝 而来的。
JOHN|16|28|我从父而来，到了世界 ，又离开世界，到父那里去。”
JOHN|16|29|门徒说：“你看，如今你是明说，不用比方了。
JOHN|16|30|现在我们晓得你凡事都知道，也不需要有人问你；从此我们信你是从上帝而来的。”
JOHN|16|31|耶稣回答他们：“现在你们信了吗？
JOHN|16|32|看哪，时候将到，其实已经到了，你们要分散，各归自己的地方，留下我独自一人；然而我不是独自一人，因为有父与我同在。
JOHN|16|33|我对你们说了这些事，是要使你们在我里面有平安。在世上你们有苦难，但你们要有勇气 ，我已经胜过世界。”
JOHN|17|1|耶稣说了这些话，就举目望天，说：“父啊，时候到了，愿你荣耀你的儿子，使儿子也荣耀你；
JOHN|17|2|因为你曾赐给他权柄掌管凡血肉之躯的，使他把永生赐给你所赐给他的人。
JOHN|17|3|认识你—独一的真神，并且认识你所差来的耶稣基督，这就是永生。
JOHN|17|4|我在地上已经荣耀你，你交给我做的工作，我已完成了。
JOHN|17|5|父啊，现在求你使我在你面前得荣耀，就是在未有世界以前，我同你享有的荣耀。
JOHN|17|6|“你从世上赐给我的人，我已把你的名显明给他们。他们本是你的，你把他们赐给我，他们也遵守了你的道。
JOHN|17|7|现在他们知道，你所赐给我的一切都是从你那里来的；
JOHN|17|8|因为你所赐给我的话，我已经赐给他们，他们也领受了，又确实知道，我是从你出来的，并且信你差了我来。
JOHN|17|9|我为他们祈求，不为世人祈求，却为你所赐给我的人祈求，因他们本是你的。
JOHN|17|10|凡是我的都是你的，你的也是我的，并且我因他们得了荣耀。
JOHN|17|11|我到你那里去；我不再留在世上，他们却在世上。圣父啊，求你因你的名，就是你所赐给我的名，保守他们，使他们像我们一样合而为一。
JOHN|17|12|我与他们同在的时候，我奉你的名，就是你所赐给我的名，保守了他们，我也护卫了他们；其中除了那灭亡之子，没有一个灭亡的，好使经上的话得以应验。
JOHN|17|13|现在我到你那里去，我在世上说这些话，是要他们心里充满了我的喜乐。
JOHN|17|14|我已把你的道赐给他们；世界恨他们，因为他们不属世界，正如我不属世界一样。
JOHN|17|15|我不求你把他们从世上接走，只求你保全他们，使他们脱离那恶者。
JOHN|17|16|他们不属世界，正如我不属世界一样。
JOHN|17|17|求你用真理使他们成圣；你的道就是真理。
JOHN|17|18|你怎样差我到世上，我也照样差他们到世上。
JOHN|17|19|我为他们的缘故使自己分别为圣，为要使他们也因真理成圣。
JOHN|17|20|“我不但为这些人祈求，也为那些藉着他们的话信我的人祈求，
JOHN|17|21|使他们都合而为一。正如父你在我里面，我在你里面，使他们也在我们里面，好让世人信是你差我来的。
JOHN|17|22|你所赐给我的荣耀，我已赐给他们，使他们合而为一，像我们合而为一。
JOHN|17|23|我在他们里面，你在我里面，使他们完完全全合而为一，让世人知道是你差我来的，也知道你爱他们，如同爱我一样。
JOHN|17|24|父啊，我在哪里，愿你所赐给我的人也同我在哪里，使他们看见你所赐给我的荣耀，因为创世以前，你已经爱我了。
JOHN|17|25|公义的父啊，世人未曾认识你，我却认识你，这些人也知道是你差我来的。
JOHN|17|26|我已让他们认识你的名，还要让他们认识，好让你爱我的爱在他们里面，我也在他们里面。”
JOHN|18|1|耶稣说了这些话，就同门徒出去，过了 汲沦溪 。在那里有一个园子，他和门徒进去了。
JOHN|18|2|出卖耶稣的 犹大 也知道那地方，因为耶稣和门徒屡次在那里聚集。
JOHN|18|3|犹大 领了一队兵，以及祭司长和法利赛人的圣殿警卫，拿着灯笼、火把和兵器来到园里。
JOHN|18|4|耶稣知道将要临到自己的一切事，就出来对他们说：“你们找谁？”
JOHN|18|5|他们回答他：“ 拿撒勒 人耶稣。”耶稣对他们说：“我就是。”出卖他的 犹大 也同他们站在一起。
JOHN|18|6|耶稣一对他们说“我就是”，他们就退后，倒在地上。
JOHN|18|7|他又问他们：“你们找谁？”他们说：“ 拿撒勒 人耶稣。”
JOHN|18|8|耶稣回答：“我已经告诉你们，我就是。你们若找的是我，就让这些人走吧。”
JOHN|18|9|这要应验耶稣说过的话：“你所赐给我的人，我一个也不失落。”
JOHN|18|10|西门．彼得 带着一把刀，就拔出来，把大祭司的仆人砍了一刀，削掉了他的右耳，那仆人名叫 马勒古 。
JOHN|18|11|于是耶稣对 彼得 说：“收刀入鞘吧！我父给我的杯，我岂可不喝呢？”
JOHN|18|12|那队兵、千夫长和 犹太 人的警卫拿住耶稣，把他捆绑了，
JOHN|18|13|先带到 亚那 面前，因为他是那年的大祭司 该亚法 的岳父。
JOHN|18|14|这 该亚法 就是从前向 犹太 人忠告说“一个人替百姓死是有利的”那个人。
JOHN|18|15|西门．彼得 跟着耶稣，另一个门徒也跟着；那门徒是大祭司所认识的，他就同耶稣进了大祭司的院子。
JOHN|18|16|彼得 却站在门外。大祭司所认识的那个门徒出来，对看门的使女说了一声，就领 彼得 进去。
JOHN|18|17|那看门的使女对 彼得 说：“你不也是这人的门徒吗？”他说：“我不是。”
JOHN|18|18|仆人和警卫因为天冷生了炭火，站在那里取暖； 彼得 也同他们站着取暖。
JOHN|18|19|于是，大祭司盘问耶稣有关他的门徒和他教导的事。
JOHN|18|20|耶稣回答他：“我一向都是公开地对世人讲话，我常在会堂和圣殿里，就是 犹太 人聚集的地方教导人，我私下并没有讲什么。
JOHN|18|21|你为什么问我呢？去问那些听过我讲话的人，我所说的，他们都知道。”
JOHN|18|22|耶稣说了这些话，旁边站着的一个警卫打了他一耳光，说：“你这样回答大祭司吗？”
JOHN|18|23|耶稣回答他：“假如我说的不对，你指证不对的地方；假如我说的对，你为什么打我呢？”
JOHN|18|24|于是 亚那 把耶稣绑着押解到大祭司 该亚法 那里。
JOHN|18|25|西门．彼得 正站着取暖，有人对他说：“你不也是他的门徒吗？” 彼得 不承认，说：“我不是。”
JOHN|18|26|大祭司的一个仆人，是被 彼得 削掉耳朵那人的亲属，说：“我不是看见你同他在园子里吗？”
JOHN|18|27|彼得 又不承认，立刻鸡就叫了。
JOHN|18|28|他们把耶稣从 该亚法 那里押解到总督府。那时是清早。他们自己却不进总督府，恐怕染了污秽，不能吃逾越节的宴席。
JOHN|18|29|于是 彼拉多 出来，到他们那里，说：“你们告这人是为什么事呢？”
JOHN|18|30|他们回答他说：“这人若不作恶，我们就不会把他交给你了。”
JOHN|18|31|彼拉多 对他们说：“你们自己带他去，按着你们的律法问他吧！” 犹太 人说：“我们没有杀人的权柄。”
JOHN|18|32|这是要应验耶稣所说，指自己将要怎样死的话。
JOHN|18|33|于是 彼拉多 又进了总督府，叫耶稣来，对他说：“你是 犹太 人的王吗？”
JOHN|18|34|耶稣回答：“这话是你说的，还是别人论到我时对你说的呢？”
JOHN|18|35|彼拉多 回答：“难道我是 犹太 人吗？你的同胞和祭司长把你交给我。你做了什么事呢？”
JOHN|18|36|耶稣回答：“我的国不属于这世界；我的国若属于这世界，我的部下就会为我战斗，使我不至于被交给 犹太 人。只是我的国不属于这世界。”
JOHN|18|37|于是 彼拉多 对他说：“那么，你是王了？”耶稣回答：“是你说我是王。我为此而生，也为此来到世界，为了给真理作见证。凡属真理的人都听我的话。”
JOHN|18|38|彼拉多 对他说：“真理是什么呢？” 说了这话， 彼拉多 又出来到 犹太 人那里，对他们说：“我查不出他有什么罪状。
JOHN|18|39|但你们有个规矩，在逾越节要我给你们释放一个人，你们要我给你们释放这 犹太 人的王吗？”
JOHN|18|40|他们又再喊着说：“不要这人！要 巴拉巴 ！”这 巴拉巴 是个强盗。
JOHN|19|1|于是， 彼拉多 命令把耶稣带去鞭打了。
JOHN|19|2|士兵用荆棘编了冠冕，戴在他头上，给他穿上紫袍，
JOHN|19|3|又走到他面前，说：“万岁， 犹太 人的王！”他们就打他耳光。
JOHN|19|4|彼拉多 又出来对众人说：“看，我带他出来见你们，让你们知道我查不出他有什么罪状。”
JOHN|19|5|耶稣出来，戴着荆棘冠冕，穿着紫袍。 彼拉多 对他们说：“看哪，这个人！”
JOHN|19|6|祭司长和圣殿警卫看见他，就喊着说：“钉十字架！钉十字架！” 彼拉多 对他们说：“你们自己把他带去钉十字架吧！我查不出他有什么罪状。”
JOHN|19|7|犹太 人回答他：“我们有律法，按照律法，他是该死的，因为他自以为是上帝的儿子。”
JOHN|19|8|彼拉多 听见这话，越发害怕，
JOHN|19|9|又进了总督府，对耶稣说：“你是哪里来的？”耶稣却不回答。
JOHN|19|10|于是 彼拉多 对他说：“你不对我说话吗？难道你不知道我有权柄释放你，也有权柄把你钉十字架吗？”
JOHN|19|11|耶稣回答他：“若不是从上头赐给你的，你就毫无权柄办我，所以，把我交给你的那人罪更重了。”
JOHN|19|12|从此， 彼拉多 想要释放耶稣，无奈 犹太 人喊着说：“你若释放这个人，你就不是凯撒的忠臣 。凡自立为王的就是背叛凯撒。”
JOHN|19|13|彼拉多 听见这些话，就带耶稣出来，到了一个地方，叫“铺华石处”， 希伯来 话叫 厄巴大 ，就在那里坐堂。
JOHN|19|14|那日是逾越节的预备日，约在正午。 彼拉多 对 犹太 人说：“看哪，你们的王！”
JOHN|19|15|他们就喊着：“除掉他！除掉他！把他钉十字架！” 彼拉多 对他们说：“要我把你们的王钉十字架吗？”祭司长回答：“除了凯撒，我们没有王。”
JOHN|19|16|于是 彼拉多 把耶稣交给他们去钉十字架。 他们就把耶稣带了去。
JOHN|19|17|耶稣背着自己的十字架出来，到了一个地方，名叫“髑髅地”， 希伯来 话叫 各各他 。
JOHN|19|18|他们就在那里把他钉在十字架上，还有两个人和他一同被钉，一边一个，耶稣在中间。
JOHN|19|19|彼拉多 又写了一个牌子，钉在十字架上，写的是：“ 犹太 人的王， 拿撒勒 人耶稣。”
JOHN|19|20|有许多 犹太 人念这牌子，因为耶稣被钉十字架的地方靠近城，而且牌子是用 希伯来 、 罗马 、 希腊 三种文字写的。
JOHN|19|21|犹太 人的祭司长就对 彼拉多 说：“不要写‘ 犹太 人的王’，要写‘那人说：我是 犹太 人的王’。”
JOHN|19|22|彼拉多 回答：“我写了就写了。”
JOHN|19|23|士兵把耶稣钉在十字架上以后，把他的衣服拿来分为四份，每人一份。他们又拿他的内衣，这件内衣没有缝，是上下一片织成的。
JOHN|19|24|他们就彼此说：“我们不要撕开，我们抽签，看是谁的。”这要应验经上的话说： “他们分了我的外衣， 为我的内衣抽签。” 士兵果然做了这些事。
JOHN|19|25|站在耶稣十字架旁边的，有他的母亲、姨母、 革罗罢 的妻子 马利亚 ，和 抹大拉 的 马利亚 。
JOHN|19|26|耶稣见母亲和他所爱的那门徒站在旁边，就对母亲说：“母亲 ，看，你的儿子！”
JOHN|19|27|又对那门徒说：“看，你的母亲！”从那刻起，那门徒就接她到自己家里去了。
JOHN|19|28|这事以后，耶稣知道各样的事已经成了，为使经上的话应验，就说：“我渴了。”
JOHN|19|29|有一个盛满了醋的罐子放在那里，他们就拿海绵蘸满了醋，绑在牛膝草上，送到他嘴边。
JOHN|19|30|耶稣尝了那醋，说：“成了！”就低下头，断了气 。
JOHN|19|31|因为这日是预备日，又因为那安息日是个大日子， 犹太 人就来求 彼拉多 叫人打断他们的腿，把他们搬走，免得尸首在安息日留在十字架上。
JOHN|19|32|于是士兵来，把第一个人的腿，和与耶稣同钉的另一个人的腿，都打断了。
JOHN|19|33|当他们来到耶稣那里，见他已经死了，就没有打断他的腿。
JOHN|19|34|然而有一个士兵拿枪扎他的肋旁，立刻有血和水流出来。
JOHN|19|35|看见这事的人作了见证—他的见证是真的，他知道自己所说的是真的—好让你们也信。
JOHN|19|36|这些事发生，为要应验经上的话：“他的骨头一根也不可折断。”
JOHN|19|37|另有经文也说：“他们要仰望自己所扎的人。”
JOHN|19|38|这些事以后， 亚利马太 的 约瑟 来求 彼拉多 ，要把耶稣的身体领去。他是耶稣的门徒，只因怕 犹太 人，就暗地里作门徒。 彼拉多 准许了，他就把耶稣的身体领走。
JOHN|19|39|尼哥德慕 也来了，就是先前夜里去见耶稣的那位，他带着约一百斤的没药和沉香。
JOHN|19|40|他们照 犹太 人丧葬的规矩，用细麻布加上香料，把耶稣的身体裹好了。
JOHN|19|41|在耶稣钉十字架的地方有一个园子，园子里有一座新墓穴，是从来没有葬过人的。
JOHN|19|42|因为那天是 犹太 人的预备日，而那坟墓又在附近，他们就把耶稣安放在那里。
JOHN|20|1|七日的第一日清早，天还黑的时候， 抹大拉 的 马利亚 来到坟墓，看见石头已从坟墓挪开了，
JOHN|20|2|就跑来见 西门．彼得 和耶稣所爱的那个门徒，对他们说：“有人从坟墓里把主移走了，我们不知道他们把他放在哪里。”
JOHN|20|3|彼得 和那门徒就出来，往坟墓去。
JOHN|20|4|两个人同跑，那门徒比 彼得 跑得快，先到了坟墓，
JOHN|20|5|低头往里看，看见细麻布还放在那里，只是没有进去。
JOHN|20|6|西门．彼得 随后也到了，进了坟墓，看见细麻布放在那里，
JOHN|20|7|又看见耶稣的裹头巾没有和细麻布放在一起，是另在一处卷着。
JOHN|20|8|然后先到坟墓的那门徒也进去，他看见就信了。
JOHN|20|9|他们还不明白圣经所说耶稣必须从死人中复活的意思。
JOHN|20|10|于是两个门徒回自己的住处去了。
JOHN|20|11|马利亚 却站在坟墓外面哭。她哭的时候，低头往坟墓里看，
JOHN|20|12|看见两个天使穿着白衣，在安放耶稣身体的地方坐着，一个在头，一个在脚。
JOHN|20|13|天使对她说：“妇人，你为什么哭？”她对他们说：“因为有人把我主移走了，我不知道他们把他放在哪里。”
JOHN|20|14|说了这些话，她转过身来，看见耶稣站在那里，却不知道他是耶稣。
JOHN|20|15|耶稣问她：“妇人，你为什么哭？你找谁？” 马利亚 以为他是看园子的，就对他说：“先生，若是你把他移了去，请告诉我，你把他放在哪里，我去把他移回来。”
JOHN|20|16|耶稣对她说：“ 马利亚 。” 马利亚 转过身来，用 希伯来 话对他说：“拉波尼！”（“拉波尼”就是老师的意思。）
JOHN|20|17|耶稣对她说：“不要拉住我，因为我还没有升上去见我的父。你到我弟兄那里去告诉他们，我要升上去见我的父，也是你们的父，见我的上帝，也是你们的上帝。”
JOHN|20|18|抹大拉 的 马利亚 就向门徒报信：“我已经看见了主。”她又把主对她说的话告诉他们。
JOHN|20|19|那日（就是七日的第一日）晚上，门徒因怕 犹太 人，所在的地方门都关了。耶稣来，站在当中，对他们说：“愿你们平安！”
JOHN|20|20|说了这话，他把手和肋旁给他们看。门徒一看见主就喜乐了。
JOHN|20|21|于是耶稣又对他们说：“愿你们平安！父怎样差遣了我，我也照样差遣你们。”
JOHN|20|22|说了这话，他向他们吹一口气，说：“领受圣灵吧！
JOHN|20|23|你们赦免谁的罪，谁的罪就得赦免；你们不赦免谁的罪，谁的罪就不得赦免。”
JOHN|20|24|那十二使徒中，有个叫 低土马 的 多马 ，耶稣来的时候，他没有和他们在一起。
JOHN|20|25|其他的门徒就对他说：“我们已经看见主了。” 多马 却对他们说：“除非我看见他手上的钉痕，用我的指头探入那钉痕，用我的手探入他的肋旁，我绝不信。”
JOHN|20|26|过了八日，门徒又在屋里， 多马 也和他们在一起。门都关了，耶稣来，站在当中，说：“愿你们平安！”
JOHN|20|27|然后他对 多马 说：“把你的指头伸到这里来，看看我的手；把你的手伸过来，探入我的肋旁。不要疑惑，总要信！”
JOHN|20|28|多马 回答，对他说：“我的主！我的上帝！”
JOHN|20|29|耶稣对他说：“你因为看见了我才信吗？那没有看见却信的有福了。”
JOHN|20|30|耶稣在他门徒面前另外行了许多神迹，没有记录在这书上。
JOHN|20|31|但记载这些事是要使你们信 耶稣是基督，是上帝的儿子，并且使你们信他，好因着他的名得生命。
JOHN|21|1|这些事以后，耶稣在 提比哩亚 海边又向门徒显现。他怎样显现记在下面。
JOHN|21|2|西门．彼得 、叫 低土马 的 多马 、 加利利 的 迦拿 人 拿但业 、 西庇太 的两个儿子，和另外两个门徒，都在一起。
JOHN|21|3|西门．彼得 对他们说：“我打鱼去。”他们对他说：“我们也和你一起去。”他们就出去，上了船；那一夜并没有打着什么。
JOHN|21|4|天刚亮的时候，耶稣站在岸上，门徒却不知道他是耶稣。
JOHN|21|5|耶稣就对他们说：“孩子们！你们有吃的没有？”他们回答他：“没有。”
JOHN|21|6|耶稣对他们说：“你们把网撒在船的右边，就会得到。”于是他们撒下网去，竟拉不上来了，因为鱼很多。
JOHN|21|7|耶稣所爱的那门徒对 彼得 说：“是主！”那时 西门．彼得 赤着身子，一听见是主，就束上外衣，跳进海里。
JOHN|21|8|其余的门徒因离岸不远，约有二百肘，就坐着小船把那网鱼拉过来。
JOHN|21|9|他们上了岸，看见那里有炭火，上面有鱼和饼。
JOHN|21|10|耶稣对他们说：“把刚才打的鱼拿几条来。”
JOHN|21|11|西门．彼得 就上船，把网拉到岸上，网里满了大鱼，共一百五十三条；虽然鱼这样多，网却没有破。
JOHN|21|12|耶稣对他们说：“你们来吃早饭。”门徒中没有一个敢问他：“你是谁？”因为他们知道他是主。
JOHN|21|13|耶稣走过来，拿饼给他们，也照样拿鱼给他们。
JOHN|21|14|耶稣从死人中复活后向门徒显现，这是第三次。
JOHN|21|15|他们吃完了早饭，耶稣对 西门．彼得 说：“ 约翰 的儿子 西门 ，你爱我比这些更深吗？” 彼得 对他说：“主啊，是的，你知道我爱你。”耶稣对他说：“你喂养我的小羊。”
JOHN|21|16|耶稣第二次又对他说：“ 约翰 的儿子 西门 ，你爱我吗？” 彼得 对他说：“主啊，是的，你知道我爱你。”耶稣说：“你牧养我的羊。”
JOHN|21|17|耶稣第三次对他说：“ 约翰 的儿子 西门 ，你爱我吗？” 彼得 因为耶稣第三次对他说“你爱我吗”，就忧愁，对耶稣说：“主啊，你无所不知，你知道我爱你。”耶稣说：“你喂养我的羊。
JOHN|21|18|我实实在在地告诉你，你年轻的时候，自己束上带子，随意往来；但年老的时候，你要伸出手来，别人要把你束上，带你到不愿意去的地方。”
JOHN|21|19|耶稣说这话，是指 彼得 会怎样死来荣耀上帝。说了这话，耶稣对他说：“你跟从我吧！”
JOHN|21|20|彼得 转过身来，看见耶稣所爱的那门徒跟着，就是在晚餐时靠着耶稣胸膛说“主啊，出卖你的是谁”的那门徒。
JOHN|21|21|彼得 看见他，就问耶稣：“主啊，这个人怎样呢？”
JOHN|21|22|耶稣对他说：“假如我要他等到我来的时候还在，跟你有什么关系呢？你跟从我吧！”
JOHN|21|23|于是这话在弟兄中间流传，说那门徒不死。其实，耶稣不是说他不死，而是对 彼得 说：“假如我要他等到我来的时候还在，跟你有什么关系呢？ ”
JOHN|21|24|这门徒就是为这些事作见证、并且记载这些事的，我们知道他的见证是真的。
JOHN|21|25|耶稣所行的事还有许多，若是一一都写出来，我想，就是全世界也容不下所要写的书。
