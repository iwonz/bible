MATT|1|1|liber generationis Iesu Christi filii David filii Abraham
MATT|1|2|Abraham genuit Isaac Isaac autem genuit Iacob Iacob autem genuit Iudam et fratres eius
MATT|1|3|Iudas autem genuit Phares et Zara de Thamar Phares autem genuit Esrom Esrom autem genuit Aram
MATT|1|4|Aram autem genuit Aminadab Aminadab autem genuit Naasson Naasson autem genuit Salmon
MATT|1|5|Salmon autem genuit Booz de Rachab Booz autem genuit Obed ex Ruth Obed autem genuit Iesse Iesse autem genuit David regem
MATT|1|6|David autem rex genuit Salomonem ex ea quae fuit Uriae
MATT|1|7|Salomon autem genuit Roboam Roboam autem genuit Abiam Abia autem genuit Asa
MATT|1|8|Asa autem genuit Iosaphat Iosaphat autem genuit Ioram Ioram autem genuit Oziam
MATT|1|9|Ozias autem genuit Ioatham Ioatham autem genuit Achaz Achaz autem genuit Ezechiam
MATT|1|10|Ezechias autem genuit Manassen Manasses autem genuit Amon Amon autem genuit Iosiam
MATT|1|11|Iosias autem genuit Iechoniam et fratres eius in transmigratione Babylonis
MATT|1|12|et post transmigrationem Babylonis Iechonias genuit Salathihel Salathihel autem genuit Zorobabel
MATT|1|13|Zorobabel autem genuit Abiud Abiud autem genuit Eliachim Eliachim autem genuit Azor
MATT|1|14|Azor autem genuit Saddoc Saddoc autem genuit Achim Achim autem genuit Eliud
MATT|1|15|Eliud autem genuit Eleazar Eleazar autem genuit Matthan Matthan autem genuit Iacob
MATT|1|16|Iacob autem genuit Ioseph virum Mariae de qua natus est Iesus qui vocatur Christus
MATT|1|17|omnes ergo generationes ab Abraham usque ad David generationes quattuordecim et a David usque ad transmigrationem Babylonis generationes quattuordecim et a transmigratione Babylonis usque ad Christum generationes quattuordecim
MATT|1|18|Christi autem generatio sic erat cum esset desponsata mater eius Maria Ioseph antequam convenirent inventa est in utero habens de Spiritu Sancto
MATT|1|19|Ioseph autem vir eius cum esset iustus et nollet eam traducere voluit occulte dimittere eam
MATT|1|20|haec autem eo cogitante ecce angelus Domini in somnis apparuit ei dicens Ioseph fili David noli timere accipere Mariam coniugem tuam quod enim in ea natum est de Spiritu Sancto est
MATT|1|21|pariet autem filium et vocabis nomen eius Iesum ipse enim salvum faciet populum suum a peccatis eorum
MATT|1|22|hoc autem totum factum est ut adimpleretur id quod dictum est a Domino per prophetam dicentem
MATT|1|23|ecce virgo in utero habebit et pariet filium et vocabunt nomen eius Emmanuhel quod est interpretatum Nobiscum Deus
MATT|1|24|exsurgens autem Ioseph a somno fecit sicut praecepit ei angelus Domini et accepit coniugem suam
MATT|1|25|et non cognoscebat eam donec peperit filium suum primogenitum et vocavit nomen eius Iesum
MATT|2|1|cum ergo natus esset Iesus in Bethleem Iudaeae in diebus Herodis regis ecce magi ab oriente venerunt Hierosolymam
MATT|2|2|dicentes ubi est qui natus est rex Iudaeorum vidimus enim stellam eius in oriente et venimus adorare eum
MATT|2|3|audiens autem Herodes rex turbatus est et omnis Hierosolyma cum illo
MATT|2|4|et congregans omnes principes sacerdotum et scribas populi sciscitabatur ab eis ubi Christus nasceretur
MATT|2|5|at illi dixerunt ei in Bethleem Iudaeae sic enim scriptum est per prophetam
MATT|2|6|et tu Bethleem terra Iuda nequaquam minima es in principibus Iuda ex te enim exiet dux qui reget populum meum Israhel
MATT|2|7|tunc Herodes clam vocatis magis diligenter didicit ab eis tempus stellae quae apparuit eis
MATT|2|8|et mittens illos in Bethleem dixit ite et interrogate diligenter de puero et cum inveneritis renuntiate mihi ut et ego veniens adorem eum
MATT|2|9|qui cum audissent regem abierunt et ecce stella quam viderant in oriente antecedebat eos usque dum veniens staret supra ubi erat puer
MATT|2|10|videntes autem stellam gavisi sunt gaudio magno valde
MATT|2|11|et intrantes domum invenerunt puerum cum Maria matre eius et procidentes adoraverunt eum et apertis thesauris suis obtulerunt ei munera aurum tus et murram
MATT|2|12|et responso accepto in somnis ne redirent ad Herodem per aliam viam reversi sunt in regionem suam
MATT|2|13|qui cum recessissent ecce angelus Domini apparuit in somnis Ioseph dicens surge et accipe puerum et matrem eius et fuge in Aegyptum et esto ibi usque dum dicam tibi futurum est enim ut Herodes quaerat puerum ad perdendum eum
MATT|2|14|qui consurgens accepit puerum et matrem eius nocte et recessit in Aegyptum
MATT|2|15|et erat ibi usque ad obitum Herodis ut adimpleretur quod dictum est a Domino per prophetam dicentem ex Aegypto vocavi filium meum
MATT|2|16|tunc Herodes videns quoniam inlusus esset a magis iratus est valde et mittens occidit omnes pueros qui erant in Bethleem et in omnibus finibus eius a bimatu et infra secundum tempus quod exquisierat a magis
MATT|2|17|tunc adimpletum est quod dictum est per Hieremiam prophetam dicentem
MATT|2|18|vox in Rama audita est ploratus et ululatus multus Rachel plorans filios suos et noluit consolari quia non sunt
MATT|2|19|defuncto autem Herode ecce apparuit angelus Domini in somnis Ioseph in Aegypto
MATT|2|20|dicens surge et accipe puerum et matrem eius et vade in terram Israhel defuncti sunt enim qui quaerebant animam pueri
MATT|2|21|qui surgens accepit puerum et matrem eius et venit in terram Israhel
MATT|2|22|audiens autem quod Archelaus regnaret in Iudaea pro Herode patre suo timuit illo ire et admonitus in somnis secessit in partes Galilaeae
MATT|2|23|et veniens habitavit in civitate quae vocatur Nazareth ut adimpleretur quod dictum est per prophetas quoniam Nazareus vocabitur
MATT|3|1|in diebus autem illis venit Iohannes Baptista praedicans in deserto Iudaeae
MATT|3|2|et dicens paenitentiam agite adpropinquavit enim regnum caelorum
MATT|3|3|hic est enim qui dictus est per Esaiam prophetam dicentem vox clamantis in deserto parate viam Domini rectas facite semitas eius
MATT|3|4|ipse autem Iohannes habebat vestimentum de pilis camelorum et zonam pelliciam circa lumbos suos esca autem eius erat lucustae et mel silvestre
MATT|3|5|tunc exiebat ad eum Hierosolyma et omnis Iudaea et omnis regio circa Iordanen
MATT|3|6|et baptizabantur in Iordane ab eo confitentes peccata sua
MATT|3|7|videns autem multos Pharisaeorum et Sadducaeorum venientes ad baptismum suum dixit eis progenies viperarum quis demonstravit vobis fugere a futura ira
MATT|3|8|facite ergo fructum dignum paenitentiae
MATT|3|9|et ne velitis dicere intra vos patrem habemus Abraham dico enim vobis quoniam potest Deus de lapidibus istis suscitare filios Abrahae
MATT|3|10|iam enim securis ad radicem arborum posita est omnis ergo arbor quae non facit fructum bonum exciditur et in ignem mittitur
MATT|3|11|ego quidem vos baptizo in aqua in paenitentiam qui autem post me venturus est fortior me est cuius non sum dignus calciamenta portare ipse vos baptizabit in Spiritu Sancto et igni
MATT|3|12|cuius ventilabrum in manu sua et permundabit aream suam et congregabit triticum suum in horreum paleas autem conburet igni inextinguibili
MATT|3|13|tunc venit Iesus a Galilaea in Iordanen ad Iohannem ut baptizaretur ab eo
MATT|3|14|Iohannes autem prohibebat eum dicens ego a te debeo baptizari et tu venis ad me
MATT|3|15|respondens autem Iesus dixit ei sine modo sic enim decet nos implere omnem iustitiam tunc dimisit eum
MATT|3|16|baptizatus autem confestim ascendit de aqua et ecce aperti sunt ei caeli et vidit Spiritum Dei descendentem sicut columbam venientem super se
MATT|3|17|et ecce vox de caelis dicens hic est Filius meus dilectus in quo mihi conplacui
MATT|4|1|tunc Iesus ductus est in desertum ab Spiritu ut temptaretur a diabolo
MATT|4|2|et cum ieiunasset quadraginta diebus et quadraginta noctibus postea esuriit
MATT|4|3|et accedens temptator dixit ei si Filius Dei es dic ut lapides isti panes fiant
MATT|4|4|qui respondens dixit scriptum est non in pane solo vivet homo sed in omni verbo quod procedit de ore Dei
MATT|4|5|tunc adsumit eum diabolus in sanctam civitatem et statuit eum supra pinnaculum templi
MATT|4|6|et dixit ei si Filius Dei es mitte te deorsum scriptum est enim quia angelis suis mandabit de te et in manibus tollent te ne forte offendas ad lapidem pedem tuum
MATT|4|7|ait illi Iesus rursum scriptum est non temptabis Dominum Deum tuum
MATT|4|8|iterum adsumit eum diabolus in montem excelsum valde et ostendit ei omnia regna mundi et gloriam eorum
MATT|4|9|et dixit illi haec tibi omnia dabo si cadens adoraveris me
MATT|4|10|tunc dicit ei Iesus vade Satanas scriptum est Dominum Deum tuum adorabis et illi soli servies
MATT|4|11|tunc reliquit eum diabolus et ecce angeli accesserunt et ministrabant ei
MATT|4|12|cum autem audisset quod Iohannes traditus esset secessit in Galilaeam
MATT|4|13|et relicta civitate Nazareth venit et habitavit in Capharnaum maritimam in finibus Zabulon et Nepthalim
MATT|4|14|ut adimpleretur quod dictum est per Esaiam prophetam
MATT|4|15|terra Zabulon et terra Nepthalim via maris trans Iordanen Galilaeae gentium
MATT|4|16|populus qui sedebat in tenebris lucem vidit magnam et sedentibus in regione et umbra mortis lux orta est eis
MATT|4|17|exinde coepit Iesus praedicare et dicere paenitentiam agite adpropinquavit enim regnum caelorum
MATT|4|18|ambulans autem iuxta mare Galilaeae vidit duos fratres Simonem qui vocatur Petrus et Andream fratrem eius mittentes rete in mare erant enim piscatores
MATT|4|19|et ait illis venite post me et faciam vos fieri piscatores hominum
MATT|4|20|at illi continuo relictis retibus secuti sunt eum
MATT|4|21|et procedens inde vidit alios duos fratres Iacobum Zebedaei et Iohannem fratrem eius in navi cum Zebedaeo patre eorum reficientes retia sua et vocavit eos
MATT|4|22|illi autem statim relictis retibus et patre secuti sunt eum
MATT|4|23|et circumibat Iesus totam Galilaeam docens in synagogis eorum et praedicans evangelium regni et sanans omnem languorem et omnem infirmitatem in populo
MATT|4|24|et abiit opinio eius in totam Syriam et obtulerunt ei omnes male habentes variis languoribus et tormentis conprehensos et qui daemonia habebant et lunaticos et paralyticos et curavit eos
MATT|4|25|et secutae sunt eum turbae multae de Galilaea et Decapoli et Hierosolymis et Iudaea et de trans Iordanen
MATT|5|1|videns autem turbas ascendit in montem et cum sedisset accesserunt ad eum discipuli eius
MATT|5|2|et aperiens os suum docebat eos dicens
MATT|5|3|beati pauperes spiritu quoniam ipsorum est regnum caelorum
MATT|5|4|beati mites quoniam ipsi possidebunt terram
MATT|5|5|beati qui lugent quoniam ipsi consolabuntur
MATT|5|6|beati qui esuriunt et sitiunt iustitiam quoniam ipsi saturabuntur
MATT|5|7|beati misericordes quia ipsi misericordiam consequentur
MATT|5|8|beati mundo corde quoniam ipsi Deum videbunt
MATT|5|9|beati pacifici quoniam filii Dei vocabuntur
MATT|5|10|beati qui persecutionem patiuntur propter iustitiam quoniam ipsorum est regnum caelorum
MATT|5|11|beati estis cum maledixerint vobis et persecuti vos fuerint et dixerint omne malum adversum vos mentientes propter me
MATT|5|12|gaudete et exultate quoniam merces vestra copiosa est in caelis sic enim persecuti sunt prophetas qui fuerunt ante vos
MATT|5|13|vos estis sal terrae quod si sal evanuerit in quo sallietur ad nihilum valet ultra nisi ut mittatur foras et conculcetur ab hominibus
MATT|5|14|vos estis lux mundi non potest civitas abscondi supra montem posita
MATT|5|15|neque accendunt lucernam et ponunt eam sub modio sed super candelabrum ut luceat omnibus qui in domo sunt
MATT|5|16|sic luceat lux vestra coram hominibus ut videant vestra bona opera et glorificent Patrem vestrum qui in caelis est
MATT|5|17|nolite putare quoniam veni solvere legem aut prophetas non veni solvere sed adimplere
MATT|5|18|amen quippe dico vobis donec transeat caelum et terra iota unum aut unus apex non praeteribit a lege donec omnia fiant
MATT|5|19|qui ergo solverit unum de mandatis istis minimis et docuerit sic homines minimus vocabitur in regno caelorum qui autem fecerit et docuerit hic magnus vocabitur in regno caelorum
MATT|5|20|dico enim vobis quia nisi abundaverit iustitia vestra plus quam scribarum et Pharisaeorum non intrabitis in regnum caelorum
MATT|5|21|audistis quia dictum est antiquis non occides qui autem occiderit reus erit iudicio
MATT|5|22|ego autem dico vobis quia omnis qui irascitur fratri suo reus erit iudicio qui autem dixerit fratri suo racha reus erit concilio qui autem dixerit fatue reus erit gehennae ignis
MATT|5|23|si ergo offeres munus tuum ad altare et ibi recordatus fueris quia frater tuus habet aliquid adversum te
MATT|5|24|relinque ibi munus tuum ante altare et vade prius reconciliare fratri tuo et tunc veniens offers munus tuum
MATT|5|25|esto consentiens adversario tuo cito dum es in via cum eo ne forte tradat te adversarius iudici et iudex tradat te ministro et in carcerem mittaris
MATT|5|26|amen dico tibi non exies inde donec reddas novissimum quadrantem
MATT|5|27|audistis quia dictum est antiquis non moechaberis
MATT|5|28|ego autem dico vobis quoniam omnis qui viderit mulierem ad concupiscendum eam iam moechatus est eam in corde suo
MATT|5|29|quod si oculus tuus dexter scandalizat te erue eum et proice abs te expedit enim tibi ut pereat unum membrorum tuorum quam totum corpus tuum mittatur in gehennam
MATT|5|30|et si dextera manus tua scandalizat te abscide eam et proice abs te expedit tibi ut pereat unum membrorum tuorum quam totum corpus tuum eat in gehennam
MATT|5|31|dictum est autem quicumque dimiserit uxorem suam det illi libellum repudii
MATT|5|32|ego autem dico vobis quia omnis qui dimiserit uxorem suam excepta fornicationis causa facit eam moechari et qui dimissam duxerit adulterat
MATT|5|33|iterum audistis quia dictum est antiquis non peierabis reddes autem Domino iuramenta tua
MATT|5|34|ego autem dico vobis non iurare omnino neque per caelum quia thronus Dei est
MATT|5|35|neque per terram quia scabillum est pedum eius neque per Hierosolymam quia civitas est magni Regis
MATT|5|36|neque per caput tuum iuraveris quia non potes unum capillum album facere aut nigrum
MATT|5|37|sit autem sermo vester est est non non quod autem his abundantius est a malo est
MATT|5|38|audistis quia dictum est oculum pro oculo et dentem pro dente
MATT|5|39|ego autem dico vobis non resistere malo sed si quis te percusserit in dextera maxilla tua praebe illi et alteram
MATT|5|40|et ei qui vult tecum iudicio contendere et tunicam tuam tollere remitte ei et pallium
MATT|5|41|et quicumque te angariaverit mille passus vade cum illo alia duo
MATT|5|42|qui petit a te da ei et volenti mutuari a te ne avertaris
MATT|5|43|audistis quia dictum est diliges proximum tuum et odio habebis inimicum tuum
MATT|5|44|ego autem dico vobis diligite inimicos vestros benefacite his qui oderunt vos et orate pro persequentibus et calumniantibus vos
MATT|5|45|ut sitis filii Patris vestri qui in caelis est qui solem suum oriri facit super bonos et malos et pluit super iustos et iniustos
MATT|5|46|si enim diligatis eos qui vos diligunt quam mercedem habebitis nonne et publicani hoc faciunt
MATT|5|47|et si salutaveritis fratres vestros tantum quid amplius facitis nonne et ethnici hoc faciunt
MATT|5|48|estote ergo vos perfecti sicut et Pater vester caelestis perfectus est
MATT|6|1|adtendite ne iustitiam vestram faciatis coram hominibus ut videamini ab eis alioquin mercedem non habebitis apud Patrem vestrum qui in caelis est
MATT|6|2|cum ergo facies elemosynam noli tuba canere ante te sicut hypocritae faciunt in synagogis et in vicis ut honorificentur ab hominibus amen dico vobis receperunt mercedem suam
MATT|6|3|te autem faciente elemosynam nesciat sinistra tua quid faciat dextera tua
MATT|6|4|ut sit elemosyna tua in abscondito et Pater tuus qui videt in abscondito reddet tibi
MATT|6|5|et cum oratis non eritis sicut hypocritae qui amant in synagogis et in angulis platearum stantes orare ut videantur ab hominibus amen dico vobis receperunt mercedem suam
MATT|6|6|tu autem cum orabis intra in cubiculum tuum et cluso ostio tuo ora Patrem tuum in abscondito et Pater tuus qui videt in abscondito reddet tibi
MATT|6|7|orantes autem nolite multum loqui sicut ethnici putant enim quia in multiloquio suo exaudiantur
MATT|6|8|nolite ergo adsimilari eis scit enim Pater vester quibus opus sit vobis antequam petatis eum
MATT|6|9|sic ergo vos orabitis Pater noster qui in caelis es sanctificetur nomen tuum
MATT|6|10|veniat regnum tuum fiat voluntas tua sicut in caelo et in terra
MATT|6|11|panem nostrum supersubstantialem da nobis hodie
MATT|6|12|et dimitte nobis debita nostra sicut et nos dimisimus debitoribus nostris
MATT|6|13|et ne inducas nos in temptationem sed libera nos a malo
MATT|6|14|si enim dimiseritis hominibus peccata eorum dimittet et vobis Pater vester caelestis delicta vestra
MATT|6|15|si autem non dimiseritis hominibus nec Pater vester dimittet peccata vestra
MATT|6|16|cum autem ieiunatis nolite fieri sicut hypocritae tristes demoliuntur enim facies suas ut pareant hominibus ieiunantes amen dico vobis quia receperunt mercedem suam
MATT|6|17|tu autem cum ieiunas ungue caput tuum et faciem tuam lava
MATT|6|18|ne videaris hominibus ieiunans sed Patri tuo qui est in abscondito et Pater tuus qui videt in abscondito reddet tibi
MATT|6|19|nolite thesaurizare vobis thesauros in terra ubi erugo et tinea demolitur ubi fures effodiunt et furantur
MATT|6|20|thesaurizate autem vobis thesauros in caelo ubi neque erugo neque tinea demolitur et ubi fures non effodiunt nec furantur
MATT|6|21|ubi enim est thesaurus tuus ibi est et cor tuum
MATT|6|22|lucerna corporis est oculus si fuerit oculus tuus simplex totum corpus tuum lucidum erit
MATT|6|23|si autem oculus tuus nequam fuerit totum corpus tuum tenebrosum erit si ergo lumen quod in te est tenebrae sunt tenebrae quantae erunt
MATT|6|24|nemo potest duobus dominis servire aut enim unum odio habebit et alterum diliget aut unum sustinebit et alterum contemnet non potestis Deo servire et mamonae
MATT|6|25|ideo dico vobis ne solliciti sitis animae vestrae quid manducetis neque corpori vestro quid induamini nonne anima plus est quam esca et corpus plus est quam vestimentum
MATT|6|26|respicite volatilia caeli quoniam non serunt neque metunt neque congregant in horrea et Pater vester caelestis pascit illa nonne vos magis pluris estis illis
MATT|6|27|quis autem vestrum cogitans potest adicere ad staturam suam cubitum unum
MATT|6|28|et de vestimento quid solliciti estis considerate lilia agri quomodo crescunt non laborant nec nent
MATT|6|29|dico autem vobis quoniam nec Salomon in omni gloria sua coopertus est sicut unum ex istis
MATT|6|30|si autem faenum agri quod hodie est et cras in clibanum mittitur Deus sic vestit quanto magis vos minimae fidei
MATT|6|31|nolite ergo solliciti esse dicentes quid manducabimus aut quid bibemus aut quo operiemur
MATT|6|32|haec enim omnia gentes inquirunt scit enim Pater vester quia his omnibus indigetis
MATT|6|33|quaerite autem primum regnum et iustitiam eius et omnia haec adicientur vobis
MATT|6|34|nolite ergo esse solliciti in crastinum crastinus enim dies sollicitus erit sibi ipse sufficit diei malitia sua
MATT|7|1|nolite iudicare ut non iudicemini
MATT|7|2|in quo enim iudicio iudicaveritis iudicabimini et in qua mensura mensi fueritis metietur vobis
MATT|7|3|quid autem vides festucam in oculo fratris tui et trabem in oculo tuo non vides
MATT|7|4|aut quomodo dicis fratri tuo sine eiciam festucam de oculo tuo et ecce trabis est in oculo tuo
MATT|7|5|hypocrita eice primum trabem de oculo tuo et tunc videbis eicere festucam de oculo fratris tui
MATT|7|6|nolite dare sanctum canibus neque mittatis margaritas vestras ante porcos ne forte conculcent eas pedibus suis et conversi disrumpant vos
MATT|7|7|petite et dabitur vobis quaerite et invenietis pulsate et aperietur vobis
MATT|7|8|omnis enim qui petit accipit et qui quaerit invenit et pulsanti aperietur
MATT|7|9|aut quis est ex vobis homo quem si petierit filius suus panem numquid lapidem porriget ei
MATT|7|10|aut si piscem petet numquid serpentem porriget ei
MATT|7|11|si ergo vos cum sitis mali nostis bona dare filiis vestris quanto magis Pater vester qui in caelis est dabit bona petentibus se
MATT|7|12|omnia ergo quaecumque vultis ut faciant vobis homines et vos facite eis haec est enim lex et prophetae
MATT|7|13|intrate per angustam portam quia lata porta et spatiosa via quae ducit ad perditionem et multi sunt qui intrant per eam
MATT|7|14|quam angusta porta et arta via quae ducit ad vitam et pauci sunt qui inveniunt eam
MATT|7|15|adtendite a falsis prophetis qui veniunt ad vos in vestimentis ovium intrinsecus autem sunt lupi rapaces
MATT|7|16|a fructibus eorum cognoscetis eos numquid colligunt de spinis uvas aut de tribulis ficus
MATT|7|17|sic omnis arbor bona fructus bonos facit mala autem arbor fructus malos facit
MATT|7|18|non potest arbor bona fructus malos facere neque arbor mala fructus bonos facere
MATT|7|19|omnis arbor quae non facit fructum bonum exciditur et in ignem mittitur
MATT|7|20|igitur ex fructibus eorum cognoscetis eos
MATT|7|21|non omnis qui dicit mihi Domine Domine intrabit in regnum caelorum sed qui facit voluntatem Patris mei qui in caelis est ipse intrabit in regnum caelorum
MATT|7|22|multi dicent mihi in illa die Domine Domine nonne in nomine tuo prophetavimus et in tuo nomine daemonia eiecimus et in tuo nomine virtutes multas fecimus
MATT|7|23|et tunc confitebor illis quia numquam novi vos discedite a me qui operamini iniquitatem
MATT|7|24|omnis ergo qui audit verba mea haec et facit ea adsimilabitur viro sapienti qui aedificavit domum suam supra petram
MATT|7|25|et descendit pluvia et venerunt flumina et flaverunt venti et inruerunt in domum illam et non cecidit fundata enim erat super petram
MATT|7|26|et omnis qui audit verba mea haec et non facit ea similis erit viro stulto qui aedificavit domum suam supra harenam
MATT|7|27|et descendit pluvia et venerunt flumina et flaverunt venti et inruerunt in domum illam et cecidit et fuit ruina eius magna
MATT|7|28|et factum est cum consummasset Iesus verba haec admirabantur turbae super doctrinam eius
MATT|7|29|erat enim docens eos sicut potestatem habens non sicut scribae eorum et Pharisaei
MATT|8|1|cum autem descendisset de monte secutae sunt eum turbae multae
MATT|8|2|et ecce leprosus veniens adorabat eum dicens Domine si vis potes me mundare
MATT|8|3|et extendens manum tetigit eum Iesus dicens volo mundare et confestim mundata est lepra eius
MATT|8|4|et ait illi Iesus vide nemini dixeris sed vade ostende te sacerdoti et offer munus quod praecepit Moses in testimonium illis
MATT|8|5|cum autem introisset Capharnaum accessit ad eum centurio rogans eum
MATT|8|6|et dicens Domine puer meus iacet in domo paralyticus et male torquetur
MATT|8|7|et ait illi Iesus ego veniam et curabo eum
MATT|8|8|et respondens centurio ait Domine non sum dignus ut intres sub tectum meum sed tantum dic verbo et sanabitur puer meus
MATT|8|9|nam et ego homo sum sub potestate habens sub me milites et dico huic vade et vadit et alio veni et venit et servo meo fac hoc et facit
MATT|8|10|audiens autem Iesus miratus est et sequentibus se dixit amen dico vobis non inveni tantam fidem in Israhel
MATT|8|11|dico autem vobis quod multi ab oriente et occidente venient et recumbent cum Abraham et Isaac et Iacob in regno caelorum
MATT|8|12|filii autem regni eicientur in tenebras exteriores ibi erit fletus et stridor dentium
MATT|8|13|et dixit Iesus centurioni vade et sicut credidisti fiat tibi et sanatus est puer in hora illa
MATT|8|14|et cum venisset Iesus in domum Petri vidit socrum eius iacentem et febricitantem
MATT|8|15|et tetigit manum eius et dimisit eam febris et surrexit et ministrabat eis
MATT|8|16|vespere autem facto obtulerunt ei multos daemonia habentes et eiciebat spiritus verbo et omnes male habentes curavit
MATT|8|17|ut adimpleretur quod dictum est per Esaiam prophetam dicentem ipse infirmitates nostras accepit et aegrotationes portavit
MATT|8|18|videns autem Iesus turbas multas circum se iussit ire trans fretum
MATT|8|19|et accedens unus scriba ait illi magister sequar te quocumque ieris
MATT|8|20|et dicit ei Iesus vulpes foveas habent et volucres caeli tabernacula Filius autem hominis non habet ubi caput reclinet
MATT|8|21|alius autem de discipulis eius ait illi Domine permitte me primum ire et sepelire patrem meum
MATT|8|22|Iesus autem ait illi sequere me et dimitte mortuos sepelire mortuos suos
MATT|8|23|et ascendente eo in navicula secuti sunt eum discipuli eius
MATT|8|24|et ecce motus magnus factus est in mari ita ut navicula operiretur fluctibus ipse vero dormiebat
MATT|8|25|et accesserunt et suscitaverunt eum dicentes Domine salva nos perimus
MATT|8|26|et dicit eis quid timidi estis modicae fidei tunc surgens imperavit ventis et mari et facta est tranquillitas magna
MATT|8|27|porro homines mirati sunt dicentes qualis est hic quia et venti et mare oboediunt ei
MATT|8|28|et cum venisset trans fretum in regionem Gerasenorum occurrerunt ei duo habentes daemonia de monumentis exeuntes saevi nimis ita ut nemo posset transire per viam illam
MATT|8|29|et ecce clamaverunt dicentes quid nobis et tibi Fili Dei venisti huc ante tempus torquere nos
MATT|8|30|erat autem non longe ab illis grex porcorum multorum pascens
MATT|8|31|daemones autem rogabant eum dicentes si eicis nos mitte nos in gregem porcorum
MATT|8|32|et ait illis ite at illi exeuntes abierunt in porcos et ecce impetu abiit totus grex per praeceps in mare et mortui sunt in aquis
MATT|8|33|pastores autem fugerunt et venientes in civitatem nuntiaverunt omnia et de his qui daemonia habuerant
MATT|8|34|et ecce tota civitas exiit obviam Iesu et viso eo rogabant ut transiret a finibus eorum
MATT|9|1|et ascendens in naviculam transfretavit et venit in civitatem suam
MATT|9|2|et ecce offerebant ei paralyticum iacentem in lecto et videns Iesus fidem illorum dixit paralytico confide fili remittuntur tibi peccata tua
MATT|9|3|et ecce quidam de scribis dixerunt intra se hic blasphemat
MATT|9|4|et cum vidisset Iesus cogitationes eorum dixit ut quid cogitatis mala in cordibus vestris
MATT|9|5|quid est facilius dicere dimittuntur tibi peccata aut dicere surge et ambula
MATT|9|6|ut sciatis autem quoniam Filius hominis habet potestatem in terra dimittendi peccata tunc ait paralytico surge tolle lectum tuum et vade in domum tuam
MATT|9|7|et surrexit et abiit in domum suam
MATT|9|8|videntes autem turbae timuerunt et glorificaverunt Deum qui dedit potestatem talem hominibus
MATT|9|9|et cum transiret inde Iesus vidit hominem sedentem in teloneo Mattheum nomine et ait illi sequere me et surgens secutus est eum
MATT|9|10|et factum est discumbente eo in domo ecce multi publicani et peccatores venientes discumbebant cum Iesu et discipulis eius
MATT|9|11|et videntes Pharisaei dicebant discipulis eius quare cum publicanis et peccatoribus manducat magister vester
MATT|9|12|at Iesus audiens ait non est opus valentibus medico sed male habentibus
MATT|9|13|euntes autem discite quid est misericordiam volo et non sacrificium non enim veni vocare iustos sed peccatores
MATT|9|14|tunc accesserunt ad eum discipuli Iohannis dicentes quare nos et Pharisaei ieiunamus frequenter discipuli autem tui non ieiunant
MATT|9|15|et ait illis Iesus numquid possunt filii sponsi lugere quamdiu cum illis est sponsus venient autem dies cum auferetur ab eis sponsus et tunc ieiunabunt
MATT|9|16|nemo autem inmittit commissuram panni rudis in vestimentum vetus tollit enim plenitudinem eius a vestimento et peior scissura fit
MATT|9|17|neque mittunt vinum novum in utres veteres alioquin rumpuntur utres et vinum effunditur et utres pereunt sed vinum novum in utres novos mittunt et ambo conservantur
MATT|9|18|haec illo loquente ad eos ecce princeps unus accessit et adorabat eum dicens filia mea modo defuncta est sed veni inpone manum super eam et vivet
MATT|9|19|et surgens Iesus sequebatur eum et discipuli eius
MATT|9|20|et ecce mulier quae sanguinis fluxum patiebatur duodecim annis accessit retro et tetigit fimbriam vestimenti eius
MATT|9|21|dicebat enim intra se si tetigero tantum vestimentum eius salva ero
MATT|9|22|at Iesus conversus et videns eam dixit confide filia fides tua te salvam fecit et salva facta est mulier ex illa hora
MATT|9|23|et cum venisset Iesus in domum principis et vidisset tibicines et turbam tumultuantem
MATT|9|24|dicebat recedite non est enim mortua puella sed dormit et deridebant eum
MATT|9|25|et cum eiecta esset turba intravit et tenuit manum eius et surrexit puella
MATT|9|26|et exiit fama haec in universam terram illam
MATT|9|27|et transeunte inde Iesu secuti sunt eum duo caeci clamantes et dicentes miserere nostri Fili David
MATT|9|28|cum autem venisset domum accesserunt ad eum caeci et dicit eis Iesus creditis quia possum hoc facere vobis dicunt ei utique Domine
MATT|9|29|tunc tetigit oculos eorum dicens secundum fidem vestram fiat vobis
MATT|9|30|et aperti sunt oculi illorum et comminatus est illis Iesus dicens videte ne quis sciat
MATT|9|31|illi autem exeuntes diffamaverunt eum in tota terra illa
MATT|9|32|egressis autem illis ecce obtulerunt ei hominem mutum daemonium habentem
MATT|9|33|et eiecto daemone locutus est mutus et miratae sunt turbae dicentes numquam paruit sic in Israhel
MATT|9|34|Pharisaei autem dicebant in principe daemoniorum eicit daemones
MATT|9|35|et circumibat Iesus civitates omnes et castella docens in synagogis eorum et praedicans evangelium regni et curans omnem languorem et omnem infirmitatem
MATT|9|36|videns autem turbas misertus est eis quia erant vexati et iacentes sicut oves non habentes pastorem
MATT|9|37|tunc dicit discipulis suis messis quidem multa operarii autem pauci
MATT|9|38|rogate ergo dominum messis ut eiciat operarios in messem suam
MATT|10|1|et convocatis duodecim discipulis suis dedit illis potestatem spirituum inmundorum ut eicerent eos et curarent omnem languorem et omnem infirmitatem
MATT|10|2|duodecim autem apostolorum nomina sunt haec primus Simon qui dicitur Petrus et Andreas frater eius
MATT|10|3|Iacobus Zebedaei et Iohannes frater eius Philippus et Bartholomeus Thomas et Mattheus publicanus et Iacobus Alphei et Thaddeus
MATT|10|4|Simon Cananeus et Iudas Scariotes qui et tradidit eum
MATT|10|5|hos duodecim misit Iesus praecipiens eis et dicens in viam gentium ne abieritis et in civitates Samaritanorum ne intraveritis
MATT|10|6|sed potius ite ad oves quae perierunt domus Israhel
MATT|10|7|euntes autem praedicate dicentes quia adpropinquavit regnum caelorum
MATT|10|8|infirmos curate mortuos suscitate leprosos mundate daemones eicite gratis accepistis gratis date
MATT|10|9|nolite possidere aurum neque argentum neque pecuniam in zonis vestris
MATT|10|10|non peram in via neque duas tunicas neque calciamenta neque virgam dignus enim est operarius cibo suo
MATT|10|11|in quamcumque civitatem aut castellum intraveritis interrogate quis in ea dignus sit et ibi manete donec exeatis
MATT|10|12|intrantes autem in domum salutate eam
MATT|10|13|et siquidem fuerit domus digna veniat pax vestra super eam si autem non fuerit digna pax vestra ad vos revertatur
MATT|10|14|et quicumque non receperit vos neque audierit sermones vestros exeuntes foras de domo vel de civitate excutite pulverem de pedibus vestris
MATT|10|15|amen dico vobis tolerabilius erit terrae Sodomorum et Gomorraeorum in die iudicii quam illi civitati
MATT|10|16|ecce ego mitto vos sicut oves in medio luporum estote ergo prudentes sicut serpentes et simplices sicut columbae
MATT|10|17|cavete autem ab hominibus tradent enim vos in conciliis et in synagogis suis flagellabunt vos
MATT|10|18|et ad praesides et ad reges ducemini propter me in testimonium illis et gentibus
MATT|10|19|cum autem tradent vos nolite cogitare quomodo aut quid loquamini dabitur enim vobis in illa hora quid loquamini
MATT|10|20|non enim vos estis qui loquimini sed Spiritus Patris vestri qui loquitur in vobis
MATT|10|21|tradet autem frater fratrem in mortem et pater filium et insurgent filii in parentes et morte eos adficient
MATT|10|22|et eritis odio omnibus propter nomen meum qui autem perseveraverit in finem hic salvus erit
MATT|10|23|cum autem persequentur vos in civitate ista fugite in aliam amen enim dico vobis non consummabitis civitates Israhel donec veniat Filius hominis
MATT|10|24|non est discipulus super magistrum nec servus super dominum suum
MATT|10|25|sufficit discipulo ut sit sicut magister eius et servus sicut dominus eius si patrem familias Beelzebub vocaverunt quanto magis domesticos eius
MATT|10|26|ne ergo timueritis eos nihil enim opertum quod non revelabitur et occultum quod non scietur
MATT|10|27|quod dico vobis in tenebris dicite in lumine et quod in aure auditis praedicate super tecta
MATT|10|28|et nolite timere eos qui occidunt corpus animam autem non possunt occidere sed potius eum timete qui potest et animam et corpus perdere in gehennam
MATT|10|29|nonne duo passeres asse veneunt et unus ex illis non cadet super terram sine Patre vestro
MATT|10|30|vestri autem et capilli capitis omnes numerati sunt
MATT|10|31|nolite ergo timere multis passeribus meliores estis vos
MATT|10|32|omnis ergo qui confitebitur me coram hominibus confitebor et ego eum coram Patre meo qui est in caelis
MATT|10|33|qui autem negaverit me coram hominibus negabo et ego eum coram Patre meo qui est in caelis
MATT|10|34|nolite arbitrari quia venerim mittere pacem in terram non veni pacem mittere sed gladium
MATT|10|35|veni enim separare hominem adversus patrem suum et filiam adversus matrem suam et nurum adversus socrum suam
MATT|10|36|et inimici hominis domestici eius
MATT|10|37|qui amat patrem aut matrem plus quam me non est me dignus et qui amat filium aut filiam super me non est me dignus
MATT|10|38|et qui non accipit crucem suam et sequitur me non est me dignus
MATT|10|39|qui invenit animam suam perdet illam et qui perdiderit animam suam propter me inveniet eam
MATT|10|40|qui recipit vos me recipit et qui me recipit recipit eum qui me misit
MATT|10|41|qui recipit prophetam in nomine prophetae mercedem prophetae accipiet et qui recipit iustum in nomine iusti mercedem iusti accipiet
MATT|10|42|et quicumque potum dederit uni ex minimis istis calicem aquae frigidae tantum in nomine discipuli amen dico vobis non perdet mercedem suam
MATT|11|1|et factum est cum consummasset Iesus praecipiens duodecim discipulis suis transiit inde ut doceret et praedicaret in civitatibus eorum
MATT|11|2|Iohannes autem cum audisset in vinculis opera Christi mittens duos de discipulis suis
MATT|11|3|ait illi tu es qui venturus es an alium expectamus
MATT|11|4|et respondens Iesus ait illis euntes renuntiate Iohanni quae auditis et videtis
MATT|11|5|caeci vident claudi ambulant leprosi mundantur surdi audiunt mortui resurgunt pauperes evangelizantur
MATT|11|6|et beatus est qui non fuerit scandalizatus in me
MATT|11|7|illis autem abeuntibus coepit Iesus dicere ad turbas de Iohanne quid existis in desertum videre harundinem vento agitatam
MATT|11|8|sed quid existis videre hominem mollibus vestitum ecce qui mollibus vestiuntur in domibus regum sunt
MATT|11|9|sed quid existis videre prophetam etiam dico vobis et plus quam prophetam
MATT|11|10|hic enim est de quo scriptum est ecce ego mitto angelum meum ante faciem tuam qui praeparabit viam tuam ante te
MATT|11|11|amen dico vobis non surrexit inter natos mulierum maior Iohanne Baptista qui autem minor est in regno caelorum maior est illo
MATT|11|12|a diebus autem Iohannis Baptistae usque nunc regnum caelorum vim patitur et violenti rapiunt illud
MATT|11|13|omnes enim prophetae et lex usque ad Iohannem prophetaverunt
MATT|11|14|et si vultis recipere ipse est Helias qui venturus est
MATT|11|15|qui habet aures audiendi audiat
MATT|11|16|cui autem similem aestimabo generationem istam similis est pueris sedentibus in foro qui clamantes coaequalibus
MATT|11|17|dicunt cecinimus vobis et non saltastis lamentavimus et non planxistis
MATT|11|18|venit enim Iohannes neque manducans neque bibens et dicunt daemonium habet
MATT|11|19|venit Filius hominis manducans et bibens et dicunt ecce homo vorax et potator vini publicanorum et peccatorum amicus et iustificata est sapientia a filiis suis
MATT|11|20|tunc coepit exprobrare civitatibus in quibus factae sunt plurimae virtutes eius quia non egissent paenitentiam
MATT|11|21|vae tibi Corazain vae tibi Bethsaida quia si in Tyro et Sidone factae essent virtutes quae factae sunt in vobis olim in cilicio et cinere paenitentiam egissent
MATT|11|22|verumtamen dico vobis Tyro et Sidoni remissius erit in die iudicii quam vobis
MATT|11|23|et tu Capharnaum numquid usque in caelum exaltaberis usque in infernum descendes quia si in Sodomis factae fuissent virtutes quae factae sunt in te forte mansissent usque in hunc diem
MATT|11|24|verumtamen dico vobis quia terrae Sodomorum remissius erit in die iudicii quam tibi
MATT|11|25|in illo tempore respondens Iesus dixit confiteor tibi Pater Domine caeli et terrae quia abscondisti haec a sapientibus et prudentibus et revelasti ea parvulis
MATT|11|26|ita Pater quoniam sic fuit placitum ante te
MATT|11|27|omnia mihi tradita sunt a Patre meo et nemo novit Filium nisi Pater neque Patrem quis novit nisi Filius et cui voluerit Filius revelare
MATT|11|28|venite ad me omnes qui laboratis et onerati estis et ego reficiam vos
MATT|11|29|tollite iugum meum super vos et discite a me quia mitis sum et humilis corde et invenietis requiem animabus vestris
MATT|11|30|iugum enim meum suave est et onus meum leve est
MATT|12|1|in illo tempore abiit Iesus sabbato per sata discipuli autem eius esurientes coeperunt vellere spicas et manducare
MATT|12|2|Pharisaei autem videntes dixerunt ei ecce discipuli tui faciunt quod non licet eis facere sabbatis
MATT|12|3|at ille dixit eis non legistis quid fecerit David quando esuriit et qui cum eo erant
MATT|12|4|quomodo intravit in domum Dei et panes propositionis comedit quos non licebat ei edere neque his qui cum eo erant nisi solis sacerdotibus
MATT|12|5|aut non legistis in lege quia sabbatis sacerdotes in templo sabbatum violant et sine crimine sunt
MATT|12|6|dico autem vobis quia templo maior est hic
MATT|12|7|si autem sciretis quid est misericordiam volo et non sacrificium numquam condemnassetis innocentes
MATT|12|8|dominus est enim Filius hominis etiam sabbati
MATT|12|9|et cum inde transisset venit in synagogam eorum
MATT|12|10|et ecce homo manum habens aridam et interrogabant eum dicentes si licet sabbatis curare ut accusarent eum
MATT|12|11|ipse autem dixit illis quis erit ex vobis homo qui habeat ovem unam et si ceciderit haec sabbatis in foveam nonne tenebit et levabit eam
MATT|12|12|quanto magis melior est homo ove itaque licet sabbatis benefacere
MATT|12|13|tunc ait homini extende manum tuam et extendit et restituta est sanitati sicut altera
MATT|12|14|exeuntes autem Pharisaei consilium faciebant adversus eum quomodo eum perderent
MATT|12|15|Iesus autem sciens recessit inde et secuti sunt eum multi et curavit eos omnes
MATT|12|16|et praecepit eis ne manifestum eum facerent
MATT|12|17|ut adimpleretur quod dictum est per Esaiam prophetam dicentem
MATT|12|18|ecce puer meus quem elegi dilectus meus in quo bene placuit animae meae ponam spiritum meum super eum et iudicium gentibus nuntiabit
MATT|12|19|non contendet neque clamabit neque audiet aliquis in plateis vocem eius
MATT|12|20|harundinem quassatam non confringet et linum fumigans non extinguet donec eiciat ad victoriam iudicium
MATT|12|21|et in nomine eius gentes sperabunt
MATT|12|22|tunc oblatus est ei daemonium habens caecus et mutus et curavit eum ita ut loqueretur et videret
MATT|12|23|et stupebant omnes turbae et dicebant numquid hic est Filius David
MATT|12|24|Pharisaei autem audientes dixerunt hic non eicit daemones nisi in Beelzebub principe daemoniorum
MATT|12|25|Iesus autem sciens cogitationes eorum dixit eis omne regnum divisum contra se desolatur et omnis civitas vel domus divisa contra se non stabit
MATT|12|26|et si Satanas Satanan eicit adversus se divisus est quomodo ergo stabit regnum eius
MATT|12|27|et si ego in Beelzebub eicio daemones filii vestri in quo eiciunt ideo ipsi iudices erunt vestri
MATT|12|28|si autem ego in Spiritu Dei eicio daemones igitur pervenit in vos regnum Dei
MATT|12|29|aut quomodo potest quisquam intrare in domum fortis et vasa eius diripere nisi prius alligaverit fortem et tunc domum illius diripiat
MATT|12|30|qui non est mecum contra me est et qui non congregat mecum spargit
MATT|12|31|ideo dico vobis omne peccatum et blasphemia remittetur hominibus Spiritus autem blasphemia non remittetur
MATT|12|32|et quicumque dixerit verbum contra Filium hominis remittetur ei qui autem dixerit contra Spiritum Sanctum non remittetur ei neque in hoc saeculo neque in futuro
MATT|12|33|aut facite arborem bonam et fructum eius bonum aut facite arborem malam et fructum eius malum siquidem ex fructu arbor agnoscitur
MATT|12|34|progenies viperarum quomodo potestis bona loqui cum sitis mali ex abundantia enim cordis os loquitur
MATT|12|35|bonus homo de bono thesauro profert bona et malus homo de malo thesauro profert mala
MATT|12|36|dico autem vobis quoniam omne verbum otiosum quod locuti fuerint homines reddent rationem de eo in die iudicii
MATT|12|37|ex verbis enim tuis iustificaberis et ex verbis tuis condemnaberis
MATT|12|38|tunc responderunt ei quidam de scribis et Pharisaeis dicentes magister volumus a te signum videre
MATT|12|39|qui respondens ait illis generatio mala et adultera signum quaerit et signum non dabitur ei nisi signum Ionae prophetae
MATT|12|40|sicut enim fuit Ionas in ventre ceti tribus diebus et tribus noctibus sic erit Filius hominis in corde terrae tribus diebus et tribus noctibus
MATT|12|41|viri ninevitae surgent in iudicio cum generatione ista et condemnabunt eam quia paenitentiam egerunt in praedicatione Ionae et ecce plus quam Iona hic
MATT|12|42|regina austri surget in iudicio cum generatione ista et condemnabit eam quia venit a finibus terrae audire sapientiam Salomonis et ecce plus quam Salomon hic
MATT|12|43|cum autem inmundus spiritus exierit ab homine ambulat per loca arida quaerens requiem et non invenit
MATT|12|44|tunc dicit revertar in domum meam unde exivi et veniens invenit vacantem scopis mundatam et ornatam
MATT|12|45|tunc vadit et adsumit septem alios spiritus secum nequiores se et intrantes habitant ibi et fiunt novissima hominis illius peiora prioribus sic erit et generationi huic pessimae
MATT|12|46|adhuc eo loquente ad turbas ecce mater eius et fratres stabant foris quaerentes loqui ei
MATT|12|47|dixit autem ei quidam ecce mater tua et fratres tui foris stant quaerentes te
MATT|12|48|at ipse respondens dicenti sibi ait quae est mater mea et qui sunt fratres mei
MATT|12|49|et extendens manum in discipulos suos dixit ecce mater mea et fratres mei
MATT|12|50|quicumque enim fecerit voluntatem Patris mei qui in caelis est ipse meus et frater et soror et mater est
MATT|13|1|in illo die exiens Iesus de domo sedebat secus mare
MATT|13|2|et congregatae sunt ad eum turbae multae ita ut in naviculam ascendens sederet et omnis turba stabat in litore
MATT|13|3|et locutus est eis multa in parabolis dicens ecce exiit qui seminat seminare
MATT|13|4|et dum seminat quaedam ceciderunt secus viam et venerunt volucres et comederunt ea
MATT|13|5|alia autem ceciderunt in petrosa ubi non habebat terram multam et continuo exorta sunt quia non habebant altitudinem terrae
MATT|13|6|sole autem orto aestuaverunt et quia non habebant radicem aruerunt
MATT|13|7|alia autem ceciderunt in spinas et creverunt spinae et suffocaverunt ea
MATT|13|8|alia vero ceciderunt in terram bonam et dabant fructum aliud centesimum aliud sexagesimum aliud tricesimum
MATT|13|9|qui habet aures audiendi audiat
MATT|13|10|et accedentes discipuli dixerunt ei quare in parabolis loqueris eis
MATT|13|11|qui respondens ait illis quia vobis datum est nosse mysteria regni caelorum illis autem non est datum
MATT|13|12|qui enim habet dabitur ei et abundabit qui autem non habet et quod habet auferetur ab eo
MATT|13|13|ideo in parabolis loquor eis quia videntes non vident et audientes non audiunt neque intellegunt
MATT|13|14|et adimpletur eis prophetia Esaiae dicens auditu audietis et non intellegetis et videntes videbitis et non videbitis
MATT|13|15|incrassatum est enim cor populi huius et auribus graviter audierunt et oculos suos cluserunt nequando oculis videant et auribus audiant et corde intellegant et convertantur et sanem eos
MATT|13|16|vestri autem beati oculi quia vident et aures vestrae quia audiunt
MATT|13|17|amen quippe dico vobis quia multi prophetae et iusti cupierunt videre quae videtis et non viderunt et audire quae auditis et non audierunt
MATT|13|18|vos ergo audite parabolam seminantis
MATT|13|19|omnis qui audit verbum regni et non intellegit venit malus et rapit quod seminatum est in corde eius hic est qui secus viam seminatus est
MATT|13|20|qui autem supra petrosa seminatus est hic est qui verbum audit et continuo cum gaudio accipit illud
MATT|13|21|non habet autem in se radicem sed est temporalis facta autem tribulatione et persecutione propter verbum continuo scandalizatur
MATT|13|22|qui autem est seminatus in spinis hic est qui verbum audit et sollicitudo saeculi istius et fallacia divitiarum suffocat verbum et sine fructu efficitur
MATT|13|23|qui vero in terra bona seminatus est hic est qui audit verbum et intellegit et fructum adfert et facit aliud quidem centum aliud autem sexaginta porro aliud triginta
MATT|13|24|aliam parabolam proposuit illis dicens simile factum est regnum caelorum homini qui seminavit bonum semen in agro suo
MATT|13|25|cum autem dormirent homines venit inimicus eius et superseminavit zizania in medio tritici et abiit
MATT|13|26|cum autem crevisset herba et fructum fecisset tunc apparuerunt et zizania
MATT|13|27|accedentes autem servi patris familias dixerunt ei domine nonne bonum semen seminasti in agro tuo unde ergo habet zizania
MATT|13|28|et ait illis inimicus homo hoc fecit servi autem dixerunt ei vis imus et colligimus ea
MATT|13|29|et ait non ne forte colligentes zizania eradicetis simul cum eis et triticum
MATT|13|30|sinite utraque crescere usque ad messem et in tempore messis dicam messoribus colligite primum zizania et alligate ea fasciculos ad conburendum triticum autem congregate in horreum meum
MATT|13|31|aliam parabolam proposuit eis dicens simile est regnum caelorum grano sinapis quod accipiens homo seminavit in agro suo
MATT|13|32|quod minimum quidem est omnibus seminibus cum autem creverit maius est omnibus holeribus et fit arbor ita ut volucres caeli veniant et habitent in ramis eius
MATT|13|33|aliam parabolam locutus est eis simile est regnum caelorum fermento quod acceptum mulier abscondit in farinae satis tribus donec fermentatum est totum
MATT|13|34|haec omnia locutus est Iesus in parabolis ad turbas et sine parabolis non loquebatur eis
MATT|13|35|ut impleretur quod dictum erat per prophetam dicentem aperiam in parabolis os meum eructabo abscondita a constitutione mundi
MATT|13|36|tunc dimissis turbis venit in domum et accesserunt ad eum discipuli eius dicentes dissere nobis parabolam zizaniorum agri
MATT|13|37|qui respondens ait qui seminat bonum semen est Filius hominis
MATT|13|38|ager autem est mundus bonum vero semen hii sunt filii regni zizania autem filii sunt nequam
MATT|13|39|inimicus autem qui seminavit ea est diabolus messis vero consummatio saeculi est messores autem angeli sunt
MATT|13|40|sicut ergo colliguntur zizania et igni conburuntur sic erit in consummatione saeculi
MATT|13|41|mittet Filius hominis angelos suos et colligent de regno eius omnia scandala et eos qui faciunt iniquitatem
MATT|13|42|et mittent eos in caminum ignis ibi erit fletus et stridor dentium
MATT|13|43|tunc iusti fulgebunt sicut sol in regno Patris eorum qui habet aures audiat
MATT|13|44|simile est regnum caelorum thesauro abscondito in agro quem qui invenit homo abscondit et prae gaudio illius vadit et vendit universa quae habet et emit agrum illum
MATT|13|45|iterum simile est regnum caelorum homini negotiatori quaerenti bonas margaritas
MATT|13|46|inventa autem una pretiosa margarita abiit et vendidit omnia quae habuit et emit eam
MATT|13|47|iterum simile est regnum caelorum sagenae missae in mare et ex omni genere congreganti
MATT|13|48|quam cum impleta esset educentes et secus litus sedentes elegerunt bonos in vasa malos autem foras miserunt
MATT|13|49|sic erit in consummatione saeculi exibunt angeli et separabunt malos de medio iustorum
MATT|13|50|et mittent eos in caminum ignis ibi erit fletus et stridor dentium
MATT|13|51|intellexistis haec omnia dicunt ei etiam
MATT|13|52|ait illis ideo omnis scriba doctus in regno caelorum similis est homini patri familias qui profert de thesauro suo nova et vetera
MATT|13|53|et factum est cum consummasset Iesus parabolas istas transiit inde
MATT|13|54|et veniens in patriam suam docebat eos in synagogis eorum ita ut mirarentur et dicerent unde huic sapientia haec et virtutes
MATT|13|55|nonne hic est fabri filius nonne mater eius dicitur Maria et fratres eius Iacobus et Ioseph et Simon et Iudas
MATT|13|56|et sorores eius nonne omnes apud nos sunt unde ergo huic omnia ista
MATT|13|57|et scandalizabantur in eo Iesus autem dixit eis non est propheta sine honore nisi in patria sua et in domo sua
MATT|13|58|et non fecit ibi virtutes multas propter incredulitatem illorum
MATT|14|1|in illo tempore audiit Herodes tetrarcha famam Iesu
MATT|14|2|et ait pueris suis hic est Iohannes Baptista ipse surrexit a mortuis et ideo virtutes inoperantur in eo
MATT|14|3|Herodes enim tenuit Iohannem et alligavit eum et posuit in carcere propter Herodiadem uxorem fratris sui
MATT|14|4|dicebat enim illi Iohannes non licet tibi habere eam
MATT|14|5|et volens illum occidere timuit populum quia sicut prophetam eum habebant
MATT|14|6|die autem natalis Herodis saltavit filia Herodiadis in medio et placuit Herodi
MATT|14|7|unde cum iuramento pollicitus est ei dare quodcumque postulasset ab eo
MATT|14|8|at illa praemonita a matre sua da mihi inquit hic in disco caput Iohannis Baptistae
MATT|14|9|et contristatus est rex propter iuramentum autem et eos qui pariter recumbebant iussit dari
MATT|14|10|misitque et decollavit Iohannem in carcere
MATT|14|11|et adlatum est caput eius in disco et datum est puellae et tulit matri suae
MATT|14|12|et accedentes discipuli eius tulerunt corpus et sepelierunt illud et venientes nuntiaverunt Iesu
MATT|14|13|quod cum audisset Iesus secessit inde in navicula in locum desertum seorsum et cum audissent turbae secutae sunt eum pedestres de civitatibus
MATT|14|14|et exiens vidit turbam multam et misertus est eius et curavit languidos eorum
MATT|14|15|vespere autem facto accesserunt ad eum discipuli eius dicentes desertus est locus et hora iam praeteriit dimitte turbas ut euntes in castella emant sibi escas
MATT|14|16|Iesus autem dixit eis non habent necesse ire date illis vos manducare
MATT|14|17|responderunt ei non habemus hic nisi quinque panes et duos pisces
MATT|14|18|qui ait eis adferte illos mihi huc
MATT|14|19|et cum iussisset turbam discumbere supra faenum acceptis quinque panibus et duobus piscibus aspiciens in caelum benedixit et fregit et dedit discipulis panes discipuli autem turbis
MATT|14|20|et manducaverunt omnes et saturati sunt et tulerunt reliquias duodecim cofinos fragmentorum plenos
MATT|14|21|manducantium autem fuit numerus quinque milia virorum exceptis mulieribus et parvulis
MATT|14|22|et statim iussit discipulos ascendere in navicula et praecedere eum trans fretum donec dimitteret turbas
MATT|14|23|et dimissa turba ascendit in montem solus orare vespere autem facto solus erat ibi
MATT|14|24|navicula autem in medio mari iactabatur fluctibus erat enim contrarius ventus
MATT|14|25|quarta autem vigilia noctis venit ad eos ambulans supra mare
MATT|14|26|et videntes eum supra mare ambulantem turbati sunt dicentes quia fantasma est et prae timore clamaverunt
MATT|14|27|statimque Iesus locutus est eis dicens habete fiduciam ego sum nolite timere
MATT|14|28|respondens autem Petrus dixit Domine si tu es iube me venire ad te super aquas
MATT|14|29|at ipse ait veni et descendens Petrus de navicula ambulabat super aquam ut veniret ad Iesum
MATT|14|30|videns vero ventum validum timuit et cum coepisset mergi clamavit dicens Domine salvum me fac
MATT|14|31|et continuo Iesus extendens manum adprehendit eum et ait illi modicae fidei quare dubitasti
MATT|14|32|et cum ascendissent in naviculam cessavit ventus
MATT|14|33|qui autem in navicula erant venerunt et adoraverunt eum dicentes vere Filius Dei es
MATT|14|34|et cum transfretassent venerunt in terram Gennesar
MATT|14|35|et cum cognovissent eum viri loci illius miserunt in universam regionem illam et obtulerunt ei omnes male habentes
MATT|14|36|et rogabant eum ut vel fimbriam vestimenti eius tangerent et quicumque tetigerunt salvi facti sunt
MATT|15|1|tunc accesserunt ad eum ab Hierosolymis scribae et Pharisaei dicentes
MATT|15|2|quare discipuli tui transgrediuntur traditionem seniorum non enim lavant manus suas cum panem manducant
MATT|15|3|ipse autem respondens ait illis quare et vos transgredimini mandatum Dei propter traditionem vestram
MATT|15|4|nam Deus dixit honora patrem et matrem et qui maledixerit patri vel matri morte moriatur
MATT|15|5|vos autem dicitis quicumque dixerit patri vel matri munus quodcumque est ex me tibi proderit
MATT|15|6|et non honorificabit patrem suum aut matrem et irritum fecistis mandatum Dei propter traditionem vestram
MATT|15|7|hypocritae bene prophetavit de vobis Esaias dicens
MATT|15|8|populus hic labiis me honorat cor autem eorum longe est a me
MATT|15|9|sine causa autem colunt me docentes doctrinas mandata hominum
MATT|15|10|et convocatis ad se turbis dixit eis audite et intellegite
MATT|15|11|non quod intrat in os coinquinat hominem sed quod procedit ex ore hoc coinquinat hominem
MATT|15|12|tunc accedentes discipuli eius dixerunt ei scis quia Pharisaei audito verbo scandalizati sunt
MATT|15|13|at ille respondens ait omnis plantatio quam non plantavit Pater meus caelestis eradicabitur
MATT|15|14|sinite illos caeci sunt duces caecorum caecus autem si caeco ducatum praestet ambo in foveam cadunt
MATT|15|15|respondens autem Petrus dixit ei edissere nobis parabolam istam
MATT|15|16|at ille dixit adhuc et vos sine intellectu estis
MATT|15|17|non intellegitis quia omne quod in os intrat in ventrem vadit et in secessum emittitur
MATT|15|18|quae autem procedunt de ore de corde exeunt et ea coinquinant hominem
MATT|15|19|de corde enim exeunt cogitationes malae homicidia adulteria fornicationes furta falsa testimonia blasphemiae
MATT|15|20|haec sunt quae coinquinant hominem non lotis autem manibus manducare non coinquinat hominem
MATT|15|21|et egressus inde Iesus secessit in partes Tyri et Sidonis
MATT|15|22|et ecce mulier chananea a finibus illis egressa clamavit dicens ei miserere mei Domine Fili David filia mea male a daemonio vexatur
MATT|15|23|qui non respondit ei verbum et accedentes discipuli eius rogabant eum dicentes dimitte eam quia clamat post nos
MATT|15|24|ipse autem respondens ait non sum missus nisi ad oves quae perierunt domus Israhel
MATT|15|25|at illa venit et adoravit eum dicens Domine adiuva me
MATT|15|26|qui respondens ait non est bonum sumere panem filiorum et mittere canibus
MATT|15|27|at illa dixit etiam Domine nam et catelli edunt de micis quae cadunt de mensa dominorum suorum
MATT|15|28|tunc respondens Iesus ait illi o mulier magna est fides tua fiat tibi sicut vis et sanata est filia illius ex illa hora
MATT|15|29|et cum transisset inde Iesus venit secus mare Galilaeae et ascendens in montem sedebat ibi
MATT|15|30|et accesserunt ad eum turbae multae habentes secum mutos clodos caecos debiles et alios multos et proiecerunt eos ad pedes eius et curavit eos
MATT|15|31|ita ut turbae mirarentur videntes mutos loquentes clodos ambulantes caecos videntes et magnificabant Deum Israhel
MATT|15|32|Iesus autem convocatis discipulis suis dixit misereor turbae quia triduo iam perseverant mecum et non habent quod manducent et dimittere eos ieiunos nolo ne deficiant in via
MATT|15|33|et dicunt ei discipuli unde ergo nobis in deserto panes tantos ut saturemus turbam tantam
MATT|15|34|et ait illis Iesus quot panes habetis at illi dixerunt septem et paucos pisciculos
MATT|15|35|et praecepit turbae ut discumberet super terram
MATT|15|36|et accipiens septem panes et pisces et gratias agens fregit et dedit discipulis suis et discipuli dederunt populo
MATT|15|37|et comederunt omnes et saturati sunt et quod superfuit de fragmentis tulerunt septem sportas plenas
MATT|15|38|erant autem qui manducaverant quattuor milia hominum extra parvulos et mulieres
MATT|15|39|et dimissa turba ascendit in naviculam et venit in fines Magedan
MATT|16|1|et accesserunt ad eum Pharisaei et Sadducaei temptantes et rogaverunt eum ut signum de caelo ostenderet eis
MATT|16|2|at ille respondens ait eis facto vespere dicitis serenum erit rubicundum est enim caelum
MATT|16|3|et mane hodie tempestas rutilat enim triste caelum
MATT|16|4|faciem ergo caeli diiudicare nostis signa autem temporum non potestis generatio mala et adultera signum quaerit et signum non dabitur ei nisi signum Ionae et relictis illis abiit
MATT|16|5|et cum venissent discipuli eius trans fretum obliti sunt panes accipere
MATT|16|6|qui dixit illis intuemini et cavete a fermento Pharisaeorum et Sadducaeorum
MATT|16|7|at illi cogitabant inter se dicentes quia panes non accepimus
MATT|16|8|sciens autem Iesus dixit quid cogitatis inter vos modicae fidei quia panes non habetis
MATT|16|9|nondum intellegitis neque recordamini quinque panum quinque milium hominum et quot cofinos sumpsistis
MATT|16|10|neque septem panum quattuor milium hominum et quot sportas sumpsistis
MATT|16|11|quare non intellegitis quia non de pane dixi vobis cavete a fermento Pharisaeorum et Sadducaeorum
MATT|16|12|tunc intellexerunt quia non dixerit cavendum a fermento panum sed a doctrina Pharisaeorum et Sadducaeorum
MATT|16|13|venit autem Iesus in partes Caesareae Philippi et interrogabat discipulos suos dicens quem dicunt homines esse Filium hominis
MATT|16|14|at illi dixerunt alii Iohannem Baptistam alii autem Heliam alii vero Hieremiam aut unum ex prophetis
MATT|16|15|dicit illis vos autem quem me esse dicitis
MATT|16|16|respondens Simon Petrus dixit tu es Christus Filius Dei vivi
MATT|16|17|respondens autem Iesus dixit ei beatus es Simon Bar Iona quia caro et sanguis non revelavit tibi sed Pater meus qui in caelis est
MATT|16|18|et ego dico tibi quia tu es Petrus et super hanc petram aedificabo ecclesiam meam et portae inferi non praevalebunt adversum eam
MATT|16|19|et tibi dabo claves regni caelorum et quodcumque ligaveris super terram erit ligatum in caelis et quodcumque solveris super terram erit solutum in caelis
MATT|16|20|tunc praecepit discipulis suis ut nemini dicerent quia ipse esset Iesus Christus
MATT|16|21|exinde coepit Iesus ostendere discipulis suis quia oporteret eum ire Hierosolymam et multa pati a senioribus et scribis et principibus sacerdotum et occidi et tertia die resurgere
MATT|16|22|et adsumens eum Petrus coepit increpare illum dicens absit a te Domine non erit tibi hoc
MATT|16|23|qui conversus dixit Petro vade post me Satana scandalum es mihi quia non sapis ea quae Dei sunt sed ea quae hominum
MATT|16|24|tunc Iesus dixit discipulis suis si quis vult post me venire abneget semet ipsum et tollat crucem suam et sequatur me
MATT|16|25|qui enim voluerit animam suam salvam facere perdet eam qui autem perdiderit animam suam propter me inveniet eam
MATT|16|26|quid enim prodest homini si mundum universum lucretur animae vero suae detrimentum patiatur aut quam dabit homo commutationem pro anima sua
MATT|16|27|Filius enim hominis venturus est in gloria Patris sui cum angelis suis et tunc reddet unicuique secundum opus eius
MATT|16|28|amen dico vobis sunt quidam de hic stantibus qui non gustabunt mortem donec videant Filium hominis venientem in regno suo
MATT|17|1|et post dies sex adsumpsit Iesus Petrum et Iacobum et Iohannem fratrem eius et ducit illos in montem excelsum seorsum
MATT|17|2|et transfiguratus est ante eos et resplenduit facies eius sicut sol vestimenta autem eius facta sunt alba sicut nix
MATT|17|3|et ecce apparuit illis Moses et Helias cum eo loquentes
MATT|17|4|respondens autem Petrus dixit ad Iesum Domine bonum est nos hic esse si vis faciamus hic tria tabernacula tibi unum et Mosi unum et Heliae unum
MATT|17|5|adhuc eo loquente ecce nubes lucida obumbravit eos et ecce vox de nube dicens hic est Filius meus dilectus in quo mihi bene conplacuit ipsum audite
MATT|17|6|et audientes discipuli ceciderunt in faciem suam et timuerunt valde
MATT|17|7|et accessit Iesus et tetigit eos dixitque eis surgite et nolite timere
MATT|17|8|levantes autem oculos suos neminem viderunt nisi solum Iesum
MATT|17|9|et descendentibus illis de monte praecepit Iesus dicens nemini dixeritis visionem donec Filius hominis a mortuis resurgat
MATT|17|10|et interrogaverunt eum discipuli dicentes quid ergo scribae dicunt quod Heliam oporteat primum venire
MATT|17|11|at ille respondens ait eis Helias quidem venturus est et restituet omnia
MATT|17|12|dico autem vobis quia Helias iam venit et non cognoverunt eum sed fecerunt in eo quaecumque voluerunt sic et Filius hominis passurus est ab eis
MATT|17|13|tunc intellexerunt discipuli quia de Iohanne Baptista dixisset eis
MATT|17|14|et cum venisset ad turbam accessit ad eum homo genibus provolutus ante eum dicens Domine miserere filii mei quia lunaticus est et male patitur nam saepe cadit in ignem et crebro in aquam
MATT|17|15|et obtuli eum discipulis tuis et non potuerunt curare eum
MATT|17|16|respondens Iesus ait o generatio incredula et perversa quousque ero vobiscum usquequo patiar vos adferte huc illum ad me
MATT|17|17|et increpavit ei Iesus et exiit ab eo daemonium et curatus est puer ex illa hora
MATT|17|18|tunc accesserunt discipuli ad Iesum secreto et dixerunt quare nos non potuimus eicere illum
MATT|17|19|dicit illis propter incredulitatem vestram amen quippe dico vobis si habueritis fidem sicut granum sinapis dicetis monti huic transi hinc et transibit et nihil inpossibile erit vobis
MATT|17|20|hoc autem genus non eicitur nisi per orationem et ieiunium
MATT|17|21|conversantibus autem eis in Galilaea dixit illis Iesus Filius hominis tradendus est in manus hominum
MATT|17|22|et occident eum et tertio die resurget et contristati sunt vehementer
MATT|17|23|et cum venissent Capharnaum accesserunt qui didragma accipiebant ad Petrum et dixerunt magister vester non solvit didragma
MATT|17|24|ait etiam et cum intrasset domum praevenit eum Iesus dicens quid tibi videtur Simon reges terrae a quibus accipiunt tributum vel censum a filiis suis an ab alienis
MATT|17|25|et ille dixit ab alienis dixit illi Iesus ergo liberi sunt filii
MATT|17|26|ut autem non scandalizemus eos vade ad mare et mitte hamum et eum piscem qui primus ascenderit tolle et aperto ore eius invenies staterem illum sumens da eis pro me et te
MATT|17|27|
MATT|18|1|in illa hora accesserunt discipuli ad Iesum dicentes quis putas maior est in regno caelorum
MATT|18|2|et advocans Iesus parvulum statuit eum in medio eorum
MATT|18|3|et dixit amen dico vobis nisi conversi fueritis et efficiamini sicut parvuli non intrabitis in regnum caelorum
MATT|18|4|quicumque ergo humiliaverit se sicut parvulus iste hic est maior in regno caelorum
MATT|18|5|et qui susceperit unum parvulum talem in nomine meo me suscipit
MATT|18|6|qui autem scandalizaverit unum de pusillis istis qui in me credunt expedit ei ut suspendatur mola asinaria in collo eius et demergatur in profundum maris
MATT|18|7|vae mundo ab scandalis necesse est enim ut veniant scandala verumtamen vae homini per quem scandalum venit
MATT|18|8|si autem manus tua vel pes tuus scandalizat te abscide eum et proice abs te bonum tibi est ad vitam ingredi debilem vel clodum quam duas manus vel duos pedes habentem mitti in ignem aeternum
MATT|18|9|et si oculus tuus scandalizat te erue eum et proice abs te bonum tibi est unoculum in vitam intrare quam duos oculos habentem mitti in gehennam ignis
MATT|18|10|videte ne contemnatis unum ex his pusillis dico enim vobis quia angeli eorum in caelis semper vident faciem Patris mei qui in caelis est
MATT|18|11|venit enim Filius hominis salvare quod perierat
MATT|18|12|quid vobis videtur si fuerint alicui centum oves et erraverit una ex eis nonne relinquet nonaginta novem in montibus et vadit quaerere eam quae erravit
MATT|18|13|et si contigerit ut inveniat eam amen dico vobis quia gaudebit super eam magis quam super nonaginta novem quae non erraverunt
MATT|18|14|sic non est voluntas ante Patrem vestrum qui in caelis est ut pereat unus de pusillis istis
MATT|18|15|si autem peccaverit in te frater tuus vade et corripe eum inter te et ipsum solum si te audierit lucratus es fratrem tuum
MATT|18|16|si autem non te audierit adhibe tecum adhuc unum vel duos ut in ore duorum testium vel trium stet omne verbum
MATT|18|17|quod si non audierit eos dic ecclesiae si autem et ecclesiam non audierit sit tibi sicut ethnicus et publicanus
MATT|18|18|amen dico vobis quaecumque alligaveritis super terram erunt ligata et in caelo et quaecumque solveritis super terram erunt soluta et in caelo
MATT|18|19|iterum dico vobis quia si duo ex vobis consenserint super terram de omni re quacumque petierint fiet illis a Patre meo qui in caelis est
MATT|18|20|ubi enim sunt duo vel tres congregati in nomine meo ibi sum in medio eorum
MATT|18|21|tunc accedens Petrus ad eum dixit Domine quotiens peccabit in me frater meus et dimittam ei usque septies
MATT|18|22|dicit illi Iesus non dico tibi usque septies sed usque septuagies septies
MATT|18|23|ideo adsimilatum est regnum caelorum homini regi qui voluit rationem ponere cum servis suis
MATT|18|24|et cum coepisset rationem ponere oblatus est ei unus qui debebat decem milia talenta
MATT|18|25|cum autem non haberet unde redderet iussit eum dominus venundari et uxorem eius et filios et omnia quae habebat et reddi
MATT|18|26|procidens autem servus ille orabat eum dicens patientiam habe in me et omnia reddam tibi
MATT|18|27|misertus autem dominus servi illius dimisit eum et debitum dimisit ei
MATT|18|28|egressus autem servus ille invenit unum de conservis suis qui debebat ei centum denarios et tenens suffocabat eum dicens redde quod debes
MATT|18|29|et procidens conservus eius rogabat eum dicens patientiam habe in me et omnia reddam tibi
MATT|18|30|ille autem noluit sed abiit et misit eum in carcerem donec redderet debitum
MATT|18|31|videntes autem conservi eius quae fiebant contristati sunt valde et venerunt et narraverunt domino suo omnia quae facta erant
MATT|18|32|tunc vocavit illum dominus suus et ait illi serve nequam omne debitum dimisi tibi quoniam rogasti me
MATT|18|33|non ergo oportuit et te misereri conservi tui sicut et ego tui misertus sum
MATT|18|34|et iratus dominus eius tradidit eum tortoribus quoadusque redderet universum debitum
MATT|18|35|sic et Pater meus caelestis faciet vobis si non remiseritis unusquisque fratri suo de cordibus vestris
MATT|19|1|et factum est cum consummasset Iesus sermones istos migravit a Galilaea et venit in fines Iudaeae trans Iordanen
MATT|19|2|et secutae sunt eum turbae multae et curavit eos ibi
MATT|19|3|et accesserunt ad eum Pharisaei temptantes eum et dicentes si licet homini dimittere uxorem suam quacumque ex causa
MATT|19|4|qui respondens ait eis non legistis quia qui fecit ab initio masculum et feminam fecit eos
MATT|19|5|et dixit propter hoc dimittet homo patrem et matrem et adherebit uxori suae et erunt duo in carne una
MATT|19|6|itaque iam non sunt duo sed una caro quod ergo Deus coniunxit homo non separet
MATT|19|7|dicunt illi quid ergo Moses mandavit dari libellum repudii et dimittere
MATT|19|8|ait illis quoniam Moses ad duritiam cordis vestri permisit vobis dimittere uxores vestras ab initio autem non sic fuit
MATT|19|9|dico autem vobis quia quicumque dimiserit uxorem suam nisi ob fornicationem et aliam duxerit moechatur et qui dimissam duxerit moechatur
MATT|19|10|dicunt ei discipuli eius si ita est causa homini cum uxore non expedit nubere
MATT|19|11|qui dixit non omnes capiunt verbum istud sed quibus datum est
MATT|19|12|sunt enim eunuchi qui de matris utero sic nati sunt et sunt eunuchi qui facti sunt ab hominibus et sunt eunuchi qui se ipsos castraverunt propter regnum caelorum qui potest capere capiat
MATT|19|13|tunc oblati sunt ei parvuli ut manus eis inponeret et oraret discipuli autem increpabant eis
MATT|19|14|Iesus vero ait eis sinite parvulos et nolite eos prohibere ad me venire talium est enim regnum caelorum
MATT|19|15|et cum inposuisset eis manus abiit inde
MATT|19|16|et ecce unus accedens ait illi magister bone quid boni faciam ut habeam vitam aeternam
MATT|19|17|qui dixit ei quid me interrogas de bono unus est bonus Deus si autem vis ad vitam ingredi serva mandata
MATT|19|18|dicit illi quae Iesus autem dixit non homicidium facies non adulterabis non facies furtum non falsum testimonium dices
MATT|19|19|honora patrem et matrem et diliges proximum tuum sicut te ipsum
MATT|19|20|dicit illi adulescens omnia haec custodivi quid adhuc mihi deest
MATT|19|21|ait illi Iesus si vis perfectus esse vade vende quae habes et da pauperibus et habebis thesaurum in caelo et veni sequere me
MATT|19|22|cum audisset autem adulescens verbum abiit tristis erat enim habens multas possessiones
MATT|19|23|Iesus autem dixit discipulis suis amen dico vobis quia dives difficile intrabit in regnum caelorum
MATT|19|24|et iterum dico vobis facilius est camelum per foramen acus transire quam divitem intrare in regnum caelorum
MATT|19|25|auditis autem his discipuli mirabantur valde dicentes quis ergo poterit salvus esse
MATT|19|26|aspiciens autem Iesus dixit illis apud homines hoc inpossibile est apud Deum autem omnia possibilia sunt
MATT|19|27|tunc respondens Petrus dixit ei ecce nos reliquimus omnia et secuti sumus te quid ergo erit nobis
MATT|19|28|Iesus autem dixit illis amen dico vobis quod vos qui secuti estis me in regeneratione cum sederit Filius hominis in sede maiestatis suae sedebitis et vos super sedes duodecim iudicantes duodecim tribus Israhel
MATT|19|29|et omnis qui reliquit domum vel fratres aut sorores aut patrem aut matrem aut uxorem aut filios aut agros propter nomen meum centuplum accipiet et vitam aeternam possidebit
MATT|19|30|multi autem erunt primi novissimi et novissimi primi
MATT|20|1|simile est enim regnum caelorum homini patri familias qui exiit primo mane conducere operarios in vineam suam
MATT|20|2|conventione autem facta cum operariis ex denario diurno misit eos in vineam suam
MATT|20|3|et egressus circa horam tertiam vidit alios stantes in foro otiosos
MATT|20|4|et illis dixit ite et vos in vineam et quod iustum fuerit dabo vobis
MATT|20|5|illi autem abierunt iterum autem exiit circa sextam et nonam horam et fecit similiter
MATT|20|6|circa undecimam vero exiit et invenit alios stantes et dicit illis quid hic statis tota die otiosi
MATT|20|7|dicunt ei quia nemo nos conduxit dicit illis ite et vos in vineam
MATT|20|8|cum sero autem factum esset dicit dominus vineae procuratori suo voca operarios et redde illis mercedem incipiens a novissimis usque ad primos
MATT|20|9|cum venissent ergo qui circa undecimam horam venerant acceperunt singulos denarios
MATT|20|10|venientes autem et primi arbitrati sunt quod plus essent accepturi acceperunt autem et ipsi singulos denarios
MATT|20|11|et accipientes murmurabant adversus patrem familias
MATT|20|12|dicentes hii novissimi una hora fecerunt et pares illos nobis fecisti qui portavimus pondus diei et aestus
MATT|20|13|at ille respondens uni eorum dixit amice non facio tibi iniuriam nonne ex denario convenisti mecum
MATT|20|14|tolle quod tuum est et vade volo autem et huic novissimo dare sicut et tibi
MATT|20|15|aut non licet mihi quod volo facere an oculus tuus nequam est quia ego bonus sum
MATT|20|16|sic erunt novissimi primi et primi novissimi multi sunt enim vocati pauci autem electi
MATT|20|17|et ascendens Iesus Hierosolymam adsumpsit duodecim discipulos secreto et ait illis
MATT|20|18|ecce ascendimus Hierosolymam et Filius hominis tradetur principibus sacerdotum et scribis et condemnabunt eum morte
MATT|20|19|et tradent eum gentibus ad deludendum et flagellandum et crucifigendum et tertia die resurget
MATT|20|20|tunc accessit ad eum mater filiorum Zebedaei cum filiis suis adorans et petens aliquid ab eo
MATT|20|21|qui dixit ei quid vis ait illi dic ut sedeant hii duo filii mei unus ad dexteram tuam et unus ad sinistram in regno tuo
MATT|20|22|respondens autem Iesus dixit nescitis quid petatis potestis bibere calicem quem ego bibiturus sum dicunt ei possumus
MATT|20|23|ait illis calicem quidem meum bibetis sedere autem ad dexteram meam et sinistram non est meum dare vobis sed quibus paratum est a Patre meo
MATT|20|24|et audientes decem indignati sunt de duobus fratribus
MATT|20|25|Iesus autem vocavit eos ad se et ait scitis quia principes gentium dominantur eorum et qui maiores sunt potestatem exercent in eos
MATT|20|26|non ita erit inter vos sed quicumque voluerit inter vos maior fieri sit vester minister
MATT|20|27|et qui voluerit inter vos primus esse erit vester servus
MATT|20|28|sicut Filius hominis non venit ministrari sed ministrare et dare animam suam redemptionem pro multis
MATT|20|29|et egredientibus eis ab Hiericho secuta est eum turba multa
MATT|20|30|et ecce duo caeci sedentes secus viam audierunt quia Iesus transiret et clamaverunt dicentes Domine miserere nostri Fili David
MATT|20|31|turba autem increpabat eos ut tacerent at illi magis clamabant dicentes Domine miserere nostri Fili David
MATT|20|32|et stetit Iesus et vocavit eos et ait quid vultis ut faciam vobis
MATT|20|33|dicunt illi Domine ut aperiantur oculi nostri
MATT|20|34|misertus autem eorum Iesus tetigit oculos eorum et confestim viderunt et secuti sunt eum
MATT|21|1|et cum adpropinquassent Hierosolymis et venissent Bethfage ad montem Oliveti tunc Iesus misit duos discipulos
MATT|21|2|dicens eis ite in castellum quod contra vos est et statim invenietis asinam alligatam et pullum cum ea solvite et adducite mihi
MATT|21|3|et si quis vobis aliquid dixerit dicite quia Dominus his opus habet et confestim dimittet eos
MATT|21|4|hoc autem factum est ut impleretur quod dictum est per prophetam dicentem
MATT|21|5|dicite filiae Sion ecce rex tuus venit tibi mansuetus et sedens super asinam et pullum filium subiugalis
MATT|21|6|euntes autem discipuli fecerunt sicut praecepit illis Iesus
MATT|21|7|et adduxerunt asinam et pullum et inposuerunt super eis vestimenta sua et eum desuper sedere fecerunt
MATT|21|8|plurima autem turba straverunt vestimenta sua in via alii autem caedebant ramos de arboribus et sternebant in via
MATT|21|9|turbae autem quae praecedebant et quae sequebantur clamabant dicentes osanna Filio David benedictus qui venturus est in nomine Domini osanna in altissimis
MATT|21|10|et cum intrasset Hierosolymam commota est universa civitas dicens quis est hic
MATT|21|11|populi autem dicebant hic est Iesus propheta a Nazareth Galilaeae
MATT|21|12|et intravit Iesus in templum Dei et eiciebat omnes vendentes et ementes in templo et mensas nummulariorum et cathedras vendentium columbas evertit
MATT|21|13|et dicit eis scriptum est domus mea domus orationis vocabitur vos autem fecistis eam speluncam latronum
MATT|21|14|et accesserunt ad eum caeci et claudi in templo et sanavit eos
MATT|21|15|videntes autem principes sacerdotum et scribae mirabilia quae fecit et pueros clamantes in templo et dicentes osanna Filio David indignati sunt
MATT|21|16|et dixerunt ei audis quid isti dicant Iesus autem dicit eis utique numquam legistis quia ex ore infantium et lactantium perfecisti laudem
MATT|21|17|et relictis illis abiit foras extra civitatem in Bethaniam ibique mansit
MATT|21|18|mane autem revertens in civitatem esuriit
MATT|21|19|et videns fici arborem unam secus viam venit ad eam et nihil invenit in ea nisi folia tantum et ait illi numquam ex te fructus nascatur in sempiternum et arefacta est continuo ficulnea
MATT|21|20|et videntes discipuli mirati sunt dicentes quomodo continuo aruit
MATT|21|21|respondens autem Iesus ait eis amen dico vobis si habueritis fidem et non haesitaveritis non solum de ficulnea facietis sed et si monti huic dixeritis tolle et iacta te in mare fiet
MATT|21|22|et omnia quaecumque petieritis in oratione credentes accipietis
MATT|21|23|et cum venisset in templum accesserunt ad eum docentem principes sacerdotum et seniores populi dicentes in qua potestate haec facis et quis tibi dedit hanc potestatem
MATT|21|24|respondens Iesus dixit illis interrogabo vos et ego unum sermonem quem si dixeritis mihi et ego vobis dicam in qua potestate haec facio
MATT|21|25|baptismum Iohannis unde erat e caelo an ex hominibus at illi cogitabant inter se dicentes si dixerimus e caelo dicet nobis quare ergo non credidistis illi
MATT|21|26|si autem dixerimus ex hominibus timemus turbam omnes enim habent Iohannem sicut prophetam
MATT|21|27|et respondentes Iesu dixerunt nescimus ait illis et ipse nec ego dico vobis in qua potestate haec facio
MATT|21|28|quid autem vobis videtur homo habebat duos filios et accedens ad primum dixit fili vade hodie operare in vinea mea
MATT|21|29|ille autem respondens ait nolo postea autem paenitentia motus abiit
MATT|21|30|accedens autem ad alterum dixit similiter at ille respondens ait eo domine et non ivit
MATT|21|31|quis ex duobus fecit voluntatem patris dicunt novissimus dicit illis Iesus amen dico vobis quia publicani et meretrices praecedunt vos in regno Dei
MATT|21|32|venit enim ad vos Iohannes in via iustitiae et non credidistis ei publicani autem et meretrices crediderunt ei vos autem videntes nec paenitentiam habuistis postea ut crederetis ei
MATT|21|33|aliam parabolam audite homo erat pater familias qui plantavit vineam et sepem circumdedit ei et fodit in ea torcular et aedificavit turrem et locavit eam agricolis et peregre profectus est
MATT|21|34|cum autem tempus fructuum adpropinquasset misit servos suos ad agricolas ut acciperent fructus eius
MATT|21|35|et agricolae adprehensis servis eius alium ceciderunt alium occiderunt alium vero lapidaverunt
MATT|21|36|iterum misit alios servos plures prioribus et fecerunt illis similiter
MATT|21|37|novissime autem misit ad eos filium suum dicens verebuntur filium meum
MATT|21|38|agricolae autem videntes filium dixerunt intra se hic est heres venite occidamus eum et habebimus hereditatem eius
MATT|21|39|et adprehensum eum eiecerunt extra vineam et occiderunt
MATT|21|40|cum ergo venerit dominus vineae quid faciet agricolis illis
MATT|21|41|aiunt illi malos male perdet et vineam locabit aliis agricolis qui reddant ei fructum temporibus suis
MATT|21|42|dicit illis Iesus numquam legistis in scripturis lapidem quem reprobaverunt aedificantes hic factus est in caput anguli a Domino factum est istud et est mirabile in oculis nostris
MATT|21|43|ideo dico vobis quia auferetur a vobis regnum Dei et dabitur genti facienti fructus eius
MATT|21|44|et qui ceciderit super lapidem istum confringetur super quem vero ceciderit conteret eum
MATT|21|45|et cum audissent principes sacerdotum et Pharisaei parabolas eius cognoverunt quod de ipsis diceret
MATT|21|46|et quaerentes eum tenere timuerunt turbas quoniam sicut prophetam eum habebant
MATT|22|1|et respondens Iesus dixit iterum in parabolis eis dicens
MATT|22|2|simile factum est regnum caelorum homini regi qui fecit nuptias filio suo
MATT|22|3|et misit servos suos vocare invitatos ad nuptias et nolebant venire
MATT|22|4|iterum misit alios servos dicens dicite invitatis ecce prandium meum paravi tauri mei et altilia occisa et omnia parata venite ad nuptias
MATT|22|5|illi autem neglexerunt et abierunt alius in villam suam alius vero ad negotiationem suam
MATT|22|6|reliqui vero tenuerunt servos eius et contumelia adfectos occiderunt
MATT|22|7|rex autem cum audisset iratus est et missis exercitibus suis perdidit homicidas illos et civitatem illorum succendit
MATT|22|8|tunc ait servis suis nuptiae quidem paratae sunt sed qui invitati erant non fuerunt digni
MATT|22|9|ite ergo ad exitus viarum et quoscumque inveneritis vocate ad nuptias
MATT|22|10|et egressi servi eius in vias congregaverunt omnes quos invenerunt malos et bonos et impletae sunt nuptiae discumbentium
MATT|22|11|intravit autem rex ut videret discumbentes et vidit ibi hominem non vestitum veste nuptiali
MATT|22|12|et ait illi amice quomodo huc intrasti non habens vestem nuptialem at ille obmutuit
MATT|22|13|tunc dixit rex ministris ligatis pedibus eius et manibus mittite eum in tenebras exteriores ibi erit fletus et stridor dentium
MATT|22|14|multi autem sunt vocati pauci vero electi
MATT|22|15|tunc abeuntes Pharisaei consilium inierunt ut caperent eum in sermone
MATT|22|16|et mittunt ei discipulos suos cum Herodianis dicentes magister scimus quia verax es et viam Dei in veritate doces et non est tibi cura de aliquo non enim respicis personam hominum
MATT|22|17|dic ergo nobis quid tibi videatur licet censum dare Caesari an non
MATT|22|18|cognita autem Iesus nequitia eorum ait quid me temptatis hypocritae
MATT|22|19|ostendite mihi nomisma census at illi obtulerunt ei denarium
MATT|22|20|et ait illis Iesus cuius est imago haec et suprascriptio
MATT|22|21|dicunt ei Caesaris tunc ait illis reddite ergo quae sunt Caesaris Caesari et quae sunt Dei Deo
MATT|22|22|et audientes mirati sunt et relicto eo abierunt
MATT|22|23|in illo die accesserunt ad eum Sadducaei qui dicunt non esse resurrectionem et interrogaverunt eum
MATT|22|24|dicentes magister Moses dixit si quis mortuus fuerit non habens filium ut ducat frater eius uxorem illius et suscitet semen fratri suo
MATT|22|25|erant autem apud nos septem fratres et primus uxore ducta defunctus est et non habens semen reliquit uxorem suam fratri suo
MATT|22|26|similiter secundus et tertius usque ad septimum
MATT|22|27|novissime autem omnium et mulier defuncta est
MATT|22|28|in resurrectione ergo cuius erit de septem uxor omnes enim habuerunt eam
MATT|22|29|respondens autem Iesus ait illis erratis nescientes scripturas neque virtutem Dei
MATT|22|30|in resurrectione enim neque nubent neque nubentur sed sunt sicut angeli Dei in caelo
MATT|22|31|de resurrectione autem mortuorum non legistis quod dictum est a Deo dicente vobis
MATT|22|32|ego sum Deus Abraham et Deus Isaac et Deus Iacob non est Deus mortuorum sed viventium
MATT|22|33|et audientes turbae mirabantur in doctrina eius
MATT|22|34|Pharisaei autem audientes quod silentium inposuisset Sadducaeis convenerunt in unum
MATT|22|35|et interrogavit eum unus ex eis legis doctor temptans eum
MATT|22|36|magister quod est mandatum magnum in lege
MATT|22|37|ait illi Iesus diliges Dominum Deum tuum ex toto corde tuo et in tota anima tua et in tota mente tua
MATT|22|38|hoc est maximum et primum mandatum
MATT|22|39|secundum autem simile est huic diliges proximum tuum sicut te ipsum
MATT|22|40|in his duobus mandatis universa lex pendet et prophetae
MATT|22|41|congregatis autem Pharisaeis interrogavit eos Iesus
MATT|22|42|dicens quid vobis videtur de Christo cuius filius est dicunt ei David
MATT|22|43|ait illis quomodo ergo David in spiritu vocat eum Dominum dicens
MATT|22|44|dixit Dominus Domino meo sede a dextris meis donec ponam inimicos tuos scabillum pedum tuorum
MATT|22|45|si ergo David vocat eum Dominum quomodo filius eius est
MATT|22|46|et nemo poterat respondere ei verbum neque ausus fuit quisquam ex illa die eum amplius interrogare
MATT|23|1|tunc Iesus locutus est ad turbas et discipulos suos
MATT|23|2|dicens super cathedram Mosi sederunt scribae et Pharisaei
MATT|23|3|omnia ergo quaecumque dixerint vobis servate et facite secundum opera vero eorum nolite facere dicunt enim et non faciunt
MATT|23|4|alligant autem onera gravia et inportabilia et inponunt in umeros hominum digito autem suo nolunt ea movere
MATT|23|5|omnia vero opera sua faciunt ut videantur ab hominibus dilatant enim phylacteria sua et magnificant fimbrias
MATT|23|6|amant autem primos recubitus in cenis et primas cathedras in synagogis
MATT|23|7|et salutationes in foro et vocari ab hominibus rabbi
MATT|23|8|vos autem nolite vocari rabbi unus enim est magister vester omnes autem vos fratres estis
MATT|23|9|et patrem nolite vocare vobis super terram unus enim est Pater vester qui in caelis est
MATT|23|10|nec vocemini magistri quia magister vester unus est Christus
MATT|23|11|qui maior est vestrum erit minister vester
MATT|23|12|qui autem se exaltaverit humiliabitur et qui se humiliaverit exaltabitur
MATT|23|13|vae autem vobis scribae et Pharisaei hypocritae quia clauditis regnum caelorum ante homines vos enim non intratis nec introeuntes sinitis intrare
MATT|23|14|
MATT|23|15|vae vobis scribae et Pharisaei hypocritae quia circuitis mare et aridam ut faciatis unum proselytum et cum fuerit factus facitis eum filium gehennae duplo quam vos
MATT|23|16|vae vobis duces caeci qui dicitis quicumque iuraverit per templum nihil est qui autem iuraverit in aurum templi debet
MATT|23|17|stulti et caeci quid enim maius est aurum an templum quod sanctificat aurum
MATT|23|18|et quicumque iuraverit in altari nihil est quicumque autem iuraverit in dono quod est super illud debet
MATT|23|19|caeci quid enim maius est donum an altare quod sanctificat donum
MATT|23|20|qui ergo iurat in altare iurat in eo et in omnibus quae super illud sunt
MATT|23|21|et qui iuraverit in templo iurat in illo et in eo qui inhabitat in ipso
MATT|23|22|et qui iurat in caelo iurat in throno Dei et in eo qui sedet super eum
MATT|23|23|vae vobis scribae et Pharisaei hypocritae quia decimatis mentam et anethum et cyminum et reliquistis quae graviora sunt legis iudicium et misericordiam et fidem haec oportuit facere et illa non omittere
MATT|23|24|duces caeci excolantes culicem camelum autem gluttientes
MATT|23|25|vae vobis scribae et Pharisaei hypocritae quia mundatis quod de foris est calicis et parapsidis intus autem pleni sunt rapina et inmunditia
MATT|23|26|Pharisaee caece munda prius quod intus est calicis et parapsidis ut fiat et id quod de foris est mundum
MATT|23|27|vae vobis scribae et Pharisaei hypocritae quia similes estis sepulchris dealbatis quae a foris parent hominibus speciosa intus vero plena sunt ossibus mortuorum et omni spurcitia
MATT|23|28|sic et vos a foris quidem paretis hominibus iusti intus autem pleni estis hypocrisi et iniquitate
MATT|23|29|vae vobis scribae et Pharisaei hypocritae quia aedificatis sepulchra prophetarum et ornatis monumenta iustorum
MATT|23|30|et dicitis si fuissemus in diebus patrum nostrorum non essemus socii eorum in sanguine prophetarum
MATT|23|31|itaque testimonio estis vobismet ipsis quia filii estis eorum qui prophetas occiderunt
MATT|23|32|et vos implete mensuram patrum vestrorum
MATT|23|33|serpentes genimina viperarum quomodo fugietis a iudicio gehennae
MATT|23|34|ideo ecce ego mitto ad vos prophetas et sapientes et scribas ex illis occidetis et crucifigetis et ex eis flagellabitis in synagogis vestris et persequemini de civitate in civitatem
MATT|23|35|ut veniat super vos omnis sanguis iustus qui effusus est super terram a sanguine Abel iusti usque ad sanguinem Zacchariae filii Barachiae quem occidistis inter templum et altare
MATT|23|36|amen dico vobis venient haec omnia super generationem istam
MATT|23|37|Hierusalem Hierusalem quae occidis prophetas et lapidas eos qui ad te missi sunt quotiens volui congregare filios tuos quemadmodum gallina congregat pullos suos sub alas et noluisti
MATT|23|38|ecce relinquitur vobis domus vestra deserta
MATT|23|39|dico enim vobis non me videbitis amodo donec dicatis benedictus qui venit in nomine Domini
MATT|24|1|et egressus Iesus de templo ibat et accesserunt discipuli eius ut ostenderent ei aedificationes templi
MATT|24|2|ipse autem respondens dixit eis videtis haec omnia amen dico vobis non relinquetur hic lapis super lapidem qui non destruatur
MATT|24|3|sedente autem eo super montem Oliveti accesserunt ad eum discipuli secreto dicentes dic nobis quando haec erunt et quod signum adventus tui et consummationis saeculi
MATT|24|4|et respondens Iesus dixit eis videte ne quis vos seducat
MATT|24|5|multi enim venient in nomine meo dicentes ego sum Christus et multos seducent
MATT|24|6|audituri autem estis proelia et opiniones proeliorum videte ne turbemini oportet enim haec fieri sed nondum est finis
MATT|24|7|consurget enim gens in gentem et regnum in regnum et erunt pestilentiae et fames et terraemotus per loca
MATT|24|8|haec autem omnia initia sunt dolorum
MATT|24|9|tunc tradent vos in tribulationem et occident vos et eritis odio omnibus gentibus propter nomen meum
MATT|24|10|et tunc scandalizabuntur multi et invicem tradent et odio habebunt invicem
MATT|24|11|et multi pseudoprophetae surgent et seducent multos
MATT|24|12|et quoniam abundabit iniquitas refrigescet caritas multorum
MATT|24|13|qui autem permanserit usque in finem hic salvus erit
MATT|24|14|et praedicabitur hoc evangelium regni in universo orbe in testimonium omnibus gentibus et tunc veniet consummatio
MATT|24|15|cum ergo videritis abominationem desolationis quae dicta est a Danihelo propheta stantem in loco sancto qui legit intellegat
MATT|24|16|tunc qui in Iudaea sunt fugiant ad montes
MATT|24|17|et qui in tecto non descendat tollere aliquid de domo sua
MATT|24|18|et qui in agro non revertatur tollere tunicam suam
MATT|24|19|vae autem praegnatibus et nutrientibus in illis diebus
MATT|24|20|orate autem ut non fiat fuga vestra hieme vel sabbato
MATT|24|21|erit enim tunc tribulatio magna qualis non fuit ab initio mundi usque modo neque fiet
MATT|24|22|et nisi breviati fuissent dies illi non fieret salva omnis caro sed propter electos breviabuntur dies illi
MATT|24|23|tunc si quis vobis dixerit ecce hic Christus aut illic nolite credere
MATT|24|24|surgent enim pseudochristi et pseudoprophetae et dabunt signa magna et prodigia ita ut in errorem inducantur si fieri potest etiam electi
MATT|24|25|ecce praedixi vobis
MATT|24|26|si ergo dixerint vobis ecce in deserto est nolite exire ecce in penetrabilibus nolite credere
MATT|24|27|sicut enim fulgur exit ab oriente et paret usque in occidente ita erit et adventus Filii hominis
MATT|24|28|ubicumque fuerit corpus illuc congregabuntur aquilae
MATT|24|29|statim autem post tribulationem dierum illorum sol obscurabitur et luna non dabit lumen suum et stellae cadent de caelo et virtutes caelorum commovebuntur
MATT|24|30|et tunc parebit signum Filii hominis in caelo et tunc plangent omnes tribus terrae et videbunt Filium hominis venientem in nubibus caeli cum virtute multa et maiestate
MATT|24|31|et mittet angelos suos cum tuba et voce magna et congregabunt electos eius a quattuor ventis a summis caelorum usque ad terminos eorum
MATT|24|32|ab arbore autem fici discite parabolam cum iam ramus eius tener fuerit et folia nata scitis quia prope est aestas
MATT|24|33|ita et vos cum videritis haec omnia scitote quia prope est in ianuis
MATT|24|34|amen dico vobis quia non praeteribit haec generatio donec omnia haec fiant
MATT|24|35|caelum et terra transibunt verba vero mea non praeteribunt
MATT|24|36|de die autem illa et hora nemo scit neque angeli caelorum nisi Pater solus
MATT|24|37|sicut autem in diebus Noe ita erit et adventus Filii hominis
MATT|24|38|sicut enim erant in diebus ante diluvium comedentes et bibentes nubentes et nuptum tradentes usque ad eum diem quo introivit in arcam Noe
MATT|24|39|et non cognoverunt donec venit diluvium et tulit omnes ita erit et adventus Filii hominis
MATT|24|40|tunc duo erunt in agro unus adsumetur et unus relinquetur
MATT|24|41|duae molentes in mola una adsumetur et una relinquetur
MATT|24|42|vigilate ergo quia nescitis qua hora Dominus vester venturus sit
MATT|24|43|illud autem scitote quoniam si sciret pater familias qua hora fur venturus esset vigilaret utique et non sineret perfodiri domum suam
MATT|24|44|ideoque et vos estote parati quia qua nescitis hora Filius hominis venturus est
MATT|24|45|quis putas est fidelis servus et prudens quem constituit dominus suus supra familiam suam ut det illis cibum in tempore
MATT|24|46|beatus ille servus quem cum venerit dominus eius invenerit sic facientem
MATT|24|47|amen dico vobis quoniam super omnia bona sua constituet eum
MATT|24|48|si autem dixerit malus servus ille in corde suo moram facit dominus meus venire
MATT|24|49|et coeperit percutere conservos suos manducet autem et bibat cum ebriis
MATT|24|50|veniet dominus servi illius in die qua non sperat et hora qua ignorat
MATT|24|51|et dividet eum partemque eius ponet cum hypocritis illic erit fletus et stridor dentium
MATT|25|1|tunc simile erit regnum caelorum decem virginibus quae accipientes lampadas suas exierunt obviam sponso et sponsae
MATT|25|2|quinque autem ex eis erant fatuae et quinque prudentes
MATT|25|3|sed quinque fatuae acceptis lampadibus non sumpserunt oleum secum
MATT|25|4|prudentes vero acceperunt oleum in vasis suis cum lampadibus
MATT|25|5|moram autem faciente sponso dormitaverunt omnes et dormierunt
MATT|25|6|media autem nocte clamor factus est ecce sponsus venit exite obviam ei
MATT|25|7|tunc surrexerunt omnes virgines illae et ornaverunt lampades suas
MATT|25|8|fatuae autem sapientibus dixerunt date nobis de oleo vestro quia lampades nostrae extinguntur
MATT|25|9|responderunt prudentes dicentes ne forte non sufficiat nobis et vobis ite potius ad vendentes et emite vobis
MATT|25|10|dum autem irent emere venit sponsus et quae paratae erant intraverunt cum eo ad nuptias et clausa est ianua
MATT|25|11|novissime veniunt et reliquae virgines dicentes domine domine aperi nobis
MATT|25|12|at ille respondens ait amen dico vobis nescio vos
MATT|25|13|vigilate itaque quia nescitis diem neque horam
MATT|25|14|sicut enim homo proficiscens vocavit servos suos et tradidit illis bona sua
MATT|25|15|et uni dedit quinque talenta alii autem duo alii vero unum unicuique secundum propriam virtutem et profectus est statim
MATT|25|16|abiit autem qui quinque talenta acceperat et operatus est in eis et lucratus est alia quinque
MATT|25|17|similiter qui duo acceperat lucratus est alia duo
MATT|25|18|qui autem unum acceperat abiens fodit in terra et abscondit pecuniam domini sui
MATT|25|19|post multum vero temporis venit dominus servorum illorum et posuit rationem cum eis
MATT|25|20|et accedens qui quinque talenta acceperat obtulit alia quinque talenta dicens domine quinque talenta mihi tradidisti ecce alia quinque superlucratus sum
MATT|25|21|ait illi dominus eius euge bone serve et fidelis quia super pauca fuisti fidelis super multa te constituam intra in gaudium domini tui
MATT|25|22|accessit autem et qui duo talenta acceperat et ait domine duo talenta tradidisti mihi ecce alia duo lucratus sum
MATT|25|23|ait illi dominus eius euge serve bone et fidelis quia super pauca fuisti fidelis supra multa te constituam intra in gaudium domini tui
MATT|25|24|accedens autem et qui unum talentum acceperat ait domine scio quia homo durus es metis ubi non seminasti et congregas ubi non sparsisti
MATT|25|25|et timens abii et abscondi talentum tuum in terra ecce habes quod tuum est
MATT|25|26|respondens autem dominus eius dixit ei serve male et piger sciebas quia meto ubi non semino et congrego ubi non sparsi
MATT|25|27|oportuit ergo te mittere pecuniam meam nummulariis et veniens ego recepissem utique quod meum est cum usura
MATT|25|28|tollite itaque ab eo talentum et date ei qui habet decem talenta
MATT|25|29|omni enim habenti dabitur et abundabit ei autem qui non habet et quod videtur habere auferetur ab eo
MATT|25|30|et inutilem servum eicite in tenebras exteriores illic erit fletus et stridor dentium
MATT|25|31|cum autem venerit Filius hominis in maiestate sua et omnes angeli cum eo tunc sedebit super sedem maiestatis suae
MATT|25|32|et congregabuntur ante eum omnes gentes et separabit eos ab invicem sicut pastor segregat oves ab hedis
MATT|25|33|et statuet oves quidem a dextris suis hedos autem a sinistris
MATT|25|34|tunc dicet rex his qui a dextris eius erunt venite benedicti Patris mei possidete paratum vobis regnum a constitutione mundi
MATT|25|35|esurivi enim et dedistis mihi manducare sitivi et dedistis mihi bibere hospes eram et collexistis me
MATT|25|36|nudus et operuistis me infirmus et visitastis me in carcere eram et venistis ad me
MATT|25|37|tunc respondebunt ei iusti dicentes Domine quando te vidimus esurientem et pavimus sitientem et dedimus tibi potum
MATT|25|38|quando autem te vidimus hospitem et colleximus te aut nudum et cooperuimus
MATT|25|39|aut quando te vidimus infirmum aut in carcere et venimus ad te
MATT|25|40|et respondens rex dicet illis amen dico vobis quamdiu fecistis uni de his fratribus meis minimis mihi fecistis
MATT|25|41|tunc dicet et his qui a sinistris erunt discedite a me maledicti in ignem aeternum qui paratus est diabolo et angelis eius
MATT|25|42|esurivi enim et non dedistis mihi manducare sitivi et non dedistis mihi potum
MATT|25|43|hospes eram et non collexistis me nudus et non operuistis me infirmus et in carcere et non visitastis me
MATT|25|44|tunc respondebunt et ipsi dicentes Domine quando te vidimus esurientem aut sitientem aut hospitem aut nudum aut infirmum vel in carcere et non ministravimus tibi
MATT|25|45|tunc respondebit illis dicens amen dico vobis quamdiu non fecistis uni de minoribus his nec mihi fecistis
MATT|25|46|et ibunt hii in supplicium aeternum iusti autem in vitam aeternam
MATT|26|1|et factum est cum consummasset Iesus sermones hos omnes dixit discipulis suis
MATT|26|2|scitis quia post biduum pascha fiet et Filius hominis tradetur ut crucifigatur
MATT|26|3|tunc congregati sunt principes sacerdotum et seniores populi in atrium principis sacerdotum qui dicebatur Caiaphas
MATT|26|4|et consilium fecerunt ut Iesum dolo tenerent et occiderent
MATT|26|5|dicebant autem non in die festo ne forte tumultus fieret in populo
MATT|26|6|cum autem esset Iesus in Bethania in domo Simonis leprosi
MATT|26|7|accessit ad eum mulier habens alabastrum unguenti pretiosi et effudit super caput ipsius recumbentis
MATT|26|8|videntes autem discipuli indignati sunt dicentes ut quid perditio haec
MATT|26|9|potuit enim istud venundari multo et dari pauperibus
MATT|26|10|sciens autem Iesus ait illis quid molesti estis mulieri opus bonum operata est in me
MATT|26|11|nam semper pauperes habetis vobiscum me autem non semper habetis
MATT|26|12|mittens enim haec unguentum hoc in corpus meum ad sepeliendum me fecit
MATT|26|13|amen dico vobis ubicumque praedicatum fuerit hoc evangelium in toto mundo dicetur et quod haec fecit in memoriam eius
MATT|26|14|tunc abiit unus de duodecim qui dicitur Iudas Scarioth ad principes sacerdotum
MATT|26|15|et ait illis quid vultis mihi dare et ego vobis eum tradam at illi constituerunt ei triginta argenteos
MATT|26|16|et exinde quaerebat oportunitatem ut eum traderet
MATT|26|17|prima autem azymorum accesserunt discipuli ad Iesum dicentes ubi vis paremus tibi comedere pascha
MATT|26|18|at Iesus dixit ite in civitatem ad quendam et dicite ei magister dicit tempus meum prope est apud te facio pascha cum discipulis meis
MATT|26|19|et fecerunt discipuli sicut constituit illis Iesus et paraverunt pascha
MATT|26|20|vespere autem facto discumbebat cum duodecim discipulis
MATT|26|21|et edentibus illis dixit amen dico vobis quia unus vestrum me traditurus est
MATT|26|22|et contristati valde coeperunt singuli dicere numquid ego sum Domine
MATT|26|23|at ipse respondens ait qui intinguit mecum manum in parapside hic me tradet
MATT|26|24|Filius quidem hominis vadit sicut scriptum est de illo vae autem homini illi per quem Filius hominis traditur bonum erat ei si natus non fuisset homo ille
MATT|26|25|respondens autem Iudas qui tradidit eum dixit numquid ego sum rabbi ait illi tu dixisti
MATT|26|26|cenantibus autem eis accepit Iesus panem et benedixit ac fregit deditque discipulis suis et ait accipite et comedite hoc est corpus meum
MATT|26|27|et accipiens calicem gratias egit et dedit illis dicens bibite ex hoc omnes
MATT|26|28|hic est enim sanguis meus novi testamenti qui pro multis effunditur in remissionem peccatorum
MATT|26|29|dico autem vobis non bibam amodo de hoc genimine vitis usque in diem illum cum illud bibam vobiscum novum in regno Patris mei
MATT|26|30|et hymno dicto exierunt in montem Oliveti
MATT|26|31|tunc dicit illis Iesus omnes vos scandalum patiemini in me in ista nocte scriptum est enim percutiam pastorem et dispergentur oves gregis
MATT|26|32|postquam autem resurrexero praecedam vos in Galilaeam
MATT|26|33|respondens autem Petrus ait illi et si omnes scandalizati fuerint in te ego numquam scandalizabor
MATT|26|34|ait illi Iesus amen dico tibi quia in hac nocte antequam gallus cantet ter me negabis
MATT|26|35|ait illi Petrus etiam si oportuerit me mori tecum non te negabo similiter et omnes discipuli dixerunt
MATT|26|36|tunc venit Iesus cum illis in villam quae dicitur Gethsemani et dixit discipulis suis sedete hic donec vadam illuc et orem
MATT|26|37|et adsumpto Petro et duobus filiis Zebedaei coepit contristari et maestus esse
MATT|26|38|tunc ait illis tristis est anima mea usque ad mortem sustinete hic et vigilate mecum
MATT|26|39|et progressus pusillum procidit in faciem suam orans et dicens mi Pater si possibile est transeat a me calix iste verumtamen non sicut ego volo sed sicut tu
MATT|26|40|et venit ad discipulos et invenit eos dormientes et dicit Petro sic non potuistis una hora vigilare mecum
MATT|26|41|vigilate et orate ut non intretis in temptationem spiritus quidem promptus est caro autem infirma
MATT|26|42|iterum secundo abiit et oravit dicens Pater mi si non potest hic calix transire nisi bibam illum fiat voluntas tua
MATT|26|43|et venit iterum et invenit eos dormientes erant enim oculi eorum gravati
MATT|26|44|et relictis illis iterum abiit et oravit tertio eundem sermonem dicens
MATT|26|45|tunc venit ad discipulos suos et dicit illis dormite iam et requiescite ecce adpropinquavit hora et Filius hominis traditur in manus peccatorum
MATT|26|46|surgite eamus ecce adpropinquavit qui me tradit
MATT|26|47|adhuc ipso loquente ecce Iudas unus de duodecim venit et cum eo turba multa cum gladiis et fustibus a principibus sacerdotum et senioribus populi
MATT|26|48|qui autem tradidit eum dedit illis signum dicens quemcumque osculatus fuero ipse est tenete eum
MATT|26|49|et confestim accedens ad Iesum dixit have rabbi et osculatus est eum
MATT|26|50|dixitque illi Iesus amice ad quod venisti tunc accesserunt et manus iniecerunt in Iesum et tenuerunt eum
MATT|26|51|et ecce unus ex his qui erant cum Iesu extendens manum exemit gladium suum et percutiens servum principis sacerdotum amputavit auriculam eius
MATT|26|52|tunc ait illi Iesus converte gladium tuum in locum suum omnes enim qui acceperint gladium gladio peribunt
MATT|26|53|an putas quia non possum rogare Patrem meum et exhibebit mihi modo plus quam duodecim legiones angelorum
MATT|26|54|quomodo ergo implebuntur scripturae quia sic oportet fieri
MATT|26|55|in illa hora dixit Iesus turbis tamquam ad latronem existis cum gladiis et fustibus conprehendere me cotidie apud vos sedebam docens in templo et non me tenuistis
MATT|26|56|hoc autem totum factum est ut implerentur scripturae prophetarum tunc discipuli omnes relicto eo fugerunt
MATT|26|57|at illi tenentes Iesum duxerunt ad Caiaphan principem sacerdotum ubi scribae et seniores convenerant
MATT|26|58|Petrus autem sequebatur eum a longe usque in atrium principis sacerdotum et ingressus intro sedebat cum ministris ut videret finem
MATT|26|59|principes autem sacerdotum et omne concilium quaerebant falsum testimonium contra Iesum ut eum morti traderent
MATT|26|60|et non invenerunt cum multi falsi testes accessissent novissime autem venerunt duo falsi testes
MATT|26|61|et dixerunt hic dixit possum destruere templum Dei et post triduum aedificare illud
MATT|26|62|et surgens princeps sacerdotum ait illi nihil respondes ad ea quae isti adversum te testificantur
MATT|26|63|Iesus autem tacebat et princeps sacerdotum ait illi adiuro te per Deum vivum ut dicas nobis si tu es Christus Filius Dei
MATT|26|64|dicit illi Iesus tu dixisti verumtamen dico vobis amodo videbitis Filium hominis sedentem a dextris virtutis et venientem in nubibus caeli
MATT|26|65|tunc princeps sacerdotum scidit vestimenta sua dicens blasphemavit quid adhuc egemus testibus ecce nunc audistis blasphemiam
MATT|26|66|quid vobis videtur at illi respondentes dixerunt reus est mortis
MATT|26|67|tunc expuerunt in faciem eius et colaphis eum ceciderunt alii autem palmas in faciem ei dederunt
MATT|26|68|dicentes prophetiza nobis Christe quis est qui te percussit
MATT|26|69|Petrus vero sedebat foris in atrio et accessit ad eum una ancilla dicens et tu cum Iesu Galilaeo eras
MATT|26|70|at ille negavit coram omnibus dicens nescio quid dicis
MATT|26|71|exeunte autem illo ianuam vidit eum alia et ait his qui erant ibi et hic erat cum Iesu Nazareno
MATT|26|72|et iterum negavit cum iuramento quia non novi hominem
MATT|26|73|et post pusillum accesserunt qui stabant et dixerunt Petro vere et tu ex illis es nam et loquella tua manifestum te facit
MATT|26|74|tunc coepit detestari et iurare quia non novisset hominem et continuo gallus cantavit
MATT|26|75|et recordatus est Petrus verbi Iesu quod dixerat priusquam gallus cantet ter me negabis et egressus foras ploravit amare
MATT|27|1|mane autem facto consilium inierunt omnes principes sacerdotum et seniores populi adversus Iesum ut eum morti traderent
MATT|27|2|et vinctum adduxerunt eum et tradiderunt Pontio Pilato praesidi
MATT|27|3|tunc videns Iudas qui eum tradidit quod damnatus esset paenitentia ductus rettulit triginta argenteos principibus sacerdotum et senioribus
MATT|27|4|dicens peccavi tradens sanguinem iustum at illi dixerunt quid ad nos tu videris
MATT|27|5|et proiectis argenteis in templo recessit et abiens laqueo se suspendit
MATT|27|6|principes autem sacerdotum acceptis argenteis dixerunt non licet mittere eos in corbanan quia pretium sanguinis est
MATT|27|7|consilio autem inito emerunt ex illis agrum figuli in sepulturam peregrinorum
MATT|27|8|propter hoc vocatus est ager ille Acheldemach ager sanguinis usque in hodiernum diem
MATT|27|9|tunc impletum est quod dictum est per Hieremiam prophetam dicentem et acceperunt triginta argenteos pretium adpretiati quem adpretiaverunt a filiis Israhel
MATT|27|10|et dederunt eos in agrum figuli sicut constituit mihi Dominus
MATT|27|11|Iesus autem stetit ante praesidem et interrogavit eum praeses dicens tu es rex Iudaeorum dicit ei Iesus tu dicis
MATT|27|12|et cum accusaretur a principibus sacerdotum et senioribus nihil respondit
MATT|27|13|tunc dicit illi Pilatus non audis quanta adversum te dicant testimonia
MATT|27|14|et non respondit ei ad ullum verbum ita ut miraretur praeses vehementer
MATT|27|15|per diem autem sollemnem consueverat praeses dimittere populo unum vinctum quem voluissent
MATT|27|16|habebat autem tunc vinctum insignem qui dicebatur Barabbas
MATT|27|17|congregatis ergo illis dixit Pilatus quem vultis dimittam vobis Barabban an Iesum qui dicitur Christus
MATT|27|18|sciebat enim quod per invidiam tradidissent eum
MATT|27|19|sedente autem illo pro tribunali misit ad illum uxor eius dicens nihil tibi et iusto illi multa enim passa sum hodie per visum propter eum
MATT|27|20|princeps autem sacerdotum et seniores persuaserunt populis ut peterent Barabban Iesum vero perderent
MATT|27|21|respondens autem praeses ait illis quem vultis vobis de duobus dimitti at illi dixerunt Barabban
MATT|27|22|dicit illis Pilatus quid igitur faciam de Iesu qui dicitur Christus
MATT|27|23|dicunt omnes crucifigatur ait illis praeses quid enim mali fecit at illi magis clamabant dicentes crucifigatur
MATT|27|24|videns autem Pilatus quia nihil proficeret sed magis tumultus fieret accepta aqua lavit manus coram populo dicens innocens ego sum a sanguine iusti huius vos videritis
MATT|27|25|et respondens universus populus dixit sanguis eius super nos et super filios nostros
MATT|27|26|tunc dimisit illis Barabban Iesum autem flagellatum tradidit eis ut crucifigeretur
MATT|27|27|tunc milites praesidis suscipientes Iesum in praetorio congregaverunt ad eum universam cohortem
MATT|27|28|et exuentes eum clamydem coccineam circumdederunt ei
MATT|27|29|et plectentes coronam de spinis posuerunt super caput eius et harundinem in dextera eius et genu flexo ante eum inludebant dicentes have rex Iudaeorum
MATT|27|30|et expuentes in eum acceperunt harundinem et percutiebant caput eius
MATT|27|31|et postquam inluserunt ei exuerunt eum clamydem et induerunt eum vestimentis eius et duxerunt eum ut crucifigerent
MATT|27|32|exeuntes autem invenerunt hominem cyreneum nomine Simonem hunc angariaverunt ut tolleret crucem eius
MATT|27|33|et venerunt in locum qui dicitur Golgotha quod est Calvariae locus
MATT|27|34|et dederunt ei vinum bibere cum felle mixtum et cum gustasset noluit bibere
MATT|27|35|postquam autem crucifixerunt eum diviserunt vestimenta eius sortem mittentes
MATT|27|36|et sedentes servabant eum
MATT|27|37|et inposuerunt super caput eius causam ipsius scriptam hic est Iesus rex Iudaeorum
MATT|27|38|tunc crucifixi sunt cum eo duo latrones unus a dextris et unus a sinistris
MATT|27|39|praetereuntes autem blasphemabant eum moventes capita sua
MATT|27|40|et dicentes qui destruit templum et in triduo illud reaedificat salva temet ipsum si Filius Dei es descende de cruce
MATT|27|41|similiter et principes sacerdotum inludentes cum scribis et senioribus dicentes
MATT|27|42|alios salvos fecit se ipsum non potest salvum facere si rex Israhel est descendat nunc de cruce et credemus ei
MATT|27|43|confidet in Deo liberet nunc eum si vult dixit enim quia Dei Filius sum
MATT|27|44|id ipsum autem et latrones qui fixi erant cum eo inproperabant ei
MATT|27|45|a sexta autem hora tenebrae factae sunt super universam terram usque ad horam nonam
MATT|27|46|et circa horam nonam clamavit Iesus voce magna dicens Heli Heli lema sabacthani hoc est Deus meus Deus meus ut quid dereliquisti me
MATT|27|47|quidam autem illic stantes et audientes dicebant Heliam vocat iste
MATT|27|48|et continuo currens unus ex eis acceptam spongiam implevit aceto et inposuit harundini et dabat ei bibere
MATT|27|49|ceteri vero dicebant sine videamus an veniat Helias liberans eum
MATT|27|50|Iesus autem iterum clamans voce magna emisit spiritum
MATT|27|51|et ecce velum templi scissum est in duas partes a summo usque deorsum et terra mota est et petrae scissae sunt
MATT|27|52|et monumenta aperta sunt et multa corpora sanctorum qui dormierant surrexerunt
MATT|27|53|et exeuntes de monumentis post resurrectionem eius venerunt in sanctam civitatem et apparuerunt multis
MATT|27|54|centurio autem et qui cum eo erant custodientes Iesum viso terraemotu et his quae fiebant timuerunt valde dicentes vere Dei Filius erat iste
MATT|27|55|erant autem ibi mulieres multae a longe quae secutae erant Iesum a Galilaea ministrantes ei
MATT|27|56|inter quas erat Maria Magdalene et Maria Iacobi et Ioseph mater et mater filiorum Zebedaei
MATT|27|57|cum sero autem factum esset venit quidam homo dives ab Arimathia nomine Ioseph qui et ipse discipulus erat Iesu
MATT|27|58|hic accessit ad Pilatum et petiit corpus Iesu tunc Pilatus iussit reddi corpus
MATT|27|59|et accepto corpore Ioseph involvit illud sindone munda
MATT|27|60|et posuit illud in monumento suo novo quod exciderat in petra et advolvit saxum magnum ad ostium monumenti et abiit
MATT|27|61|erat autem ibi Maria Magdalene et altera Maria sedentes contra sepulchrum
MATT|27|62|altera autem die quae est post parasceven convenerunt principes sacerdotum et Pharisaei ad Pilatum
MATT|27|63|dicentes domine recordati sumus quia seductor ille dixit adhuc vivens post tres dies resurgam
MATT|27|64|iube ergo custodiri sepulchrum usque in diem tertium ne forte veniant discipuli eius et furentur eum et dicant plebi surrexit a mortuis et erit novissimus error peior priore
MATT|27|65|ait illis Pilatus habetis custodiam ite custodite sicut scitis
MATT|27|66|illi autem abeuntes munierunt sepulchrum signantes lapidem cum custodibus
MATT|28|1|vespere autem sabbati quae lucescit in primam sabbati venit Maria Magdalene et altera Maria videre sepulchrum
MATT|28|2|et ecce terraemotus factus est magnus angelus enim Domini descendit de caelo et accedens revolvit lapidem et sedebat super eum
MATT|28|3|erat autem aspectus eius sicut fulgur et vestimentum eius sicut nix
MATT|28|4|prae timore autem eius exterriti sunt custodes et facti sunt velut mortui
MATT|28|5|respondens autem angelus dixit mulieribus nolite timere vos scio enim quod Iesum qui crucifixus est quaeritis
MATT|28|6|non est hic surrexit enim sicut dixit venite videte locum ubi positus erat Dominus
MATT|28|7|et cito euntes dicite discipulis eius quia surrexit et ecce praecedit vos in Galilaeam ibi eum videbitis ecce praedixi vobis
MATT|28|8|et exierunt cito de monumento cum timore et magno gaudio currentes nuntiare discipulis eius
MATT|28|9|et ecce Iesus occurrit illis dicens havete illae autem accesserunt et tenuerunt pedes eius et adoraverunt eum
MATT|28|10|tunc ait illis Iesus nolite timere ite nuntiate fratribus meis ut eant in Galilaeam ibi me videbunt
MATT|28|11|quae cum abissent ecce quidam de custodibus venerunt in civitatem et nuntiaverunt principibus sacerdotum omnia quae facta fuerant
MATT|28|12|et congregati cum senioribus consilio accepto pecuniam copiosam dederunt militibus
MATT|28|13|dicentes dicite quia discipuli eius nocte venerunt et furati sunt eum nobis dormientibus
MATT|28|14|et si hoc auditum fuerit a praeside nos suadebimus ei et securos vos faciemus
MATT|28|15|at illi accepta pecunia fecerunt sicut erant docti et divulgatum est verbum istud apud Iudaeos usque in hodiernum diem
MATT|28|16|undecim autem discipuli abierunt in Galilaeam in montem ubi constituerat illis Iesus
MATT|28|17|et videntes eum adoraverunt quidam autem dubitaverunt
MATT|28|18|et accedens Iesus locutus est eis dicens data est mihi omnis potestas in caelo et in terra
MATT|28|19|euntes ergo docete omnes gentes baptizantes eos in nomine Patris et Filii et Spiritus Sancti
MATT|28|20|docentes eos servare omnia quaecumque mandavi vobis et ecce ego vobiscum sum omnibus diebus usque ad consummationem saeculi
