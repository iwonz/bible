OBAD|1|1|俄巴底亚 所见的异象。 我们从耶和华那里得到消息， 有使者被差往列国去： “起来吧， 我们要起来与 以东 争战！” 主耶和华论 以东 如此说：
OBAD|1|2|看哪，我要使你在列国中为最小， 被人大大藐视。
OBAD|1|3|你狂傲的心欺骗了你， 你住在岩穴， 居所在高处， 心里说： “谁能把我拉下来到地上呢？”
OBAD|1|4|你虽如鹰高飞， 在星宿之间搭窝， 我必从那里拉你下来。 这是耶和华说的。
OBAD|1|5|盗贼若来到你那里， 小偷夜间来到， 岂不是只偷他们所需要的吗？ 摘葡萄的若来到你那里， 岂不留下几串吗？ 你竟全然灭绝！
OBAD|1|6|以扫 遭到搜查， 他隐藏的宝物竟被寻出！
OBAD|1|7|与你结盟的都驱赶你，直到边界， 与你和好的欺骗你，胜过你， 吃你饭的人设下圈套陷害你─ 他却毫无聪明 。
OBAD|1|8|到那日， 我岂不从 以东 除灭智慧人？ 从 以扫山 除灭聪明人？ 这是耶和华说的。
OBAD|1|9|提幔 哪， 你的勇士必惊惶， 以致 以扫山 的人都被杀戮剪除。
OBAD|1|10|因你向兄弟 雅各 施暴， 你必蒙羞， 永被剪除。
OBAD|1|11|当陌生人掳掠 雅各 的财物， 当外邦人进入他的城门， 为 耶路撒冷 抽签分取财物的日子， 你竟站在一旁，像与他们同伙。
OBAD|1|12|你兄弟遭难的日子， 你不该瞪着眼看； 犹大 人被灭的日子， 你不该幸灾乐祸； 他们遭难的日子， 你不该说狂傲的话。
OBAD|1|13|我子民遭灾的日子， 你不该进他们的城门； 他们遭灾的日子， 你不该瞪着眼看他们受苦； 他们遭灾的日子， 你不该伸手抢他们的财物。
OBAD|1|14|他们遭难的日子， 你不该站在岔路口 剪除他们逃脱的人， 你不该交出他们的幸存者。
OBAD|1|15|耶和华的日子临近万国； 你所做的，人也必向你照样做， 你的报应必归到自己头上。
OBAD|1|16|你们在我圣山怎样喝了苦杯， 万国必照样不停地喝， 且喝且吞， 他们就必归于无有。
OBAD|1|17|但在 锡安山 必有逃脱的人， 那山必成为圣； 雅各 家必得原有的产业 。
OBAD|1|18|雅各 家必成为大火， 约瑟 家成为火焰； 以扫 家必如碎秸， 遭燃烧，被吞灭， 以扫 家必无幸存者。 这是耶和华说的。
OBAD|1|19|他们必得 尼革夫 和 以扫山 ， 得 谢非拉 ， 非利士 人之地， 他们必得 以法莲 地和 撒玛利亚 地， 得 便雅悯 和 基列 ；
OBAD|1|20|被掳的 以色列 大军 必得 迦南 人的地，直到 撒勒法 ， 在 西法拉 被掳的 耶路撒冷 人 必得 尼革夫 的城镇。
OBAD|1|21|必有一些解救者 上到 锡安山 ，审判 以扫山 ， 国度就归耶和华了。
