2KGS|1|1|After the death of Ahab, Moab rebelled against Israel.
2KGS|1|2|Now Ahaziah fell through the lattice in his upper chamber in Samaria, and lay sick; so he sent messengers, telling them, "Go, inquire of Baal-zebub, the god of Ekron, whether I shall recover from this sickness."
2KGS|1|3|But the angel of the LORD said to Elijah the Tishbite, "Arise, go up to meet the messengers of the king of Samaria, and say to them, 'Is it because there is no God in Israel that you are going to inquire of Baal-zebub, the god of Ekron?
2KGS|1|4|Now therefore thus says the LORD, You shall not come down from the bed to which you have gone up, but you shall surely die.'"So Elijah went.
2KGS|1|5|The messengers returned to the king, and he said to them, "Why have you returned?"
2KGS|1|6|And they said to him, "There came a man to meet us, and said to us, 'Go back to the king who sent you, and say to him, Thus says the LORD, Is it because there is no God in Israel that you are sending to inquire of Baal-zebub, the god of Ekron? Therefore you shall not come down from the bed to which you have gone up, but you shall surely die.'"
2KGS|1|7|He said to them, "What kind of man was he who came to meet you and told you these things?"
2KGS|1|8|They answered him, "He wore a garment of hair, with a belt of leather about his waist." And he said, "It is Elijah the Tishbite."
2KGS|1|9|Then the king sent to him a captain of fifty men with his fifty. He went up to Elijah, who was sitting on the top of a hill, and said to him, "O man of God, the king says, 'Come down.'"
2KGS|1|10|But Elijah answered the captain of fifty, "If I am a man of God, let fire come down from heaven and consume you and your fifty." Then fire came down from heaven and consumed him and his fifty.
2KGS|1|11|Again the king sent to him another captain of fifty men with his fifty. And he answered and said to him, "O man of God, this is the king's order, 'Come down quickly!'"
2KGS|1|12|But Elijah answered them, "If I am a man of God, let fire come down from heaven and consume you and your fifty." Then the fire of God came down from heaven and consumed him and his fifty.
2KGS|1|13|Again the king sent the captain of a third fifty with his fifty. And the third captain of fifty went up and came and fell on his knees before Elijah and entreated him, "O man of God, please let my life, and the life of these fifty servants of yours, be precious in your sight.
2KGS|1|14|Behold, fire came down from heaven and consumed the two former captains of fifty men with their fifties, but now let my life be precious in your sight."
2KGS|1|15|Then the angel of the LORD said to Elijah, "Go down with him; do not be afraid of him." So he arose and went down with him to the king
2KGS|1|16|and said to him, "Thus says the LORD, 'Because you have sent messengers to inquire of Baal-zebub, the god of Ekron- is it because there is no God in Israel to inquire of his word?- therefore you shall not come down from the bed to which you have gone up, but you shall surely die.'"
2KGS|1|17|So he died according to the word of the LORD that Elijah had spoken. Jehoram became king in his place in the second year of Jehoram the son of Jehoshaphat, king of Judah, because Ahaziah had no son.
2KGS|1|18|Now the rest of the acts of Ahaziah that he did, are they not written in the Book of the Chronicles of the Kings of Israel?
2KGS|2|1|Now when the LORD was about to take Elijah up to heaven by a whirlwind, Elijah and Elisha were on their way from Gilgal.
2KGS|2|2|And Elijah said to Elisha, "Please stay here, for the LORD has sent me as far as Bethel." But Elisha said, "As the LORD lives, and as you yourself live, I will not leave you." So they went down to Bethel.
2KGS|2|3|And the sons of the prophets who were in Bethel came out to Elisha and said to him, "Do you know that today the LORD will take away your master from over you?" And he said, "Yes, I know it; keep quiet."
2KGS|2|4|Elijah said to him, "Elisha, please stay here, for the LORD has sent me to Jericho." But he said, "As the LORD lives, and as you yourself live, I will not leave you." So they came to Jericho.
2KGS|2|5|The sons of the prophets who were at Jericho drew near to Elisha and said to him, "Do you know that today the LORD will take away your master from over you?" And he answered, "Yes, I know it; keep quiet."
2KGS|2|6|Then Elijah said to him, "Please stay here, for the LORD has sent me to the Jordan." But he said, "As the LORD lives, and as you yourself live, I will not leave you." So the two of them went on.
2KGS|2|7|Fifty men of the sons of the prophets also went and stood at some distance from them, as they both were standing by the Jordan.
2KGS|2|8|Then Elijah took his cloak and rolled it up and struck the water, and the water was parted to the one side and to the other, till the two of them could go over on dry ground.
2KGS|2|9|When they had crossed, Elijah said to Elisha, "Ask what I shall do for you, before I am taken from you." And Elisha said, "Please let there be a double portion of your spirit on me."
2KGS|2|10|And he said, "You have asked a hard thing; yet, if you see me as I am being taken from you, it shall be so for you, but if you do not see me, it shall not be so."
2KGS|2|11|And as they still went on and talked, behold, chariots of fire and horses of fire separated the two of them. And Elijah went up by a whirlwind into heaven.
2KGS|2|12|And Elisha saw it and he cried, "My father, my father! The chariots of Israel and its horsemen!" And he saw him no more. Then he took hold of his own clothes and tore them in two pieces.
2KGS|2|13|And he took up the cloak of Elijah that had fallen from him and went back and stood on the bank of the Jordan.
2KGS|2|14|Then he took the cloak of Elijah that had fallen from him and struck the water, saying, "Where is the LORD, the God of Elijah?" And when he had struck the water, the water was parted to the one side and to the other, and Elisha went over.
2KGS|2|15|Now when the sons of the prophets who were at Jericho saw him opposite them, they said, "The spirit of Elijah rests on Elisha." And they came to meet him and bowed to the ground before him.
2KGS|2|16|And they said to him, "Behold now, there are with your servants fifty strong men. Please let them go and seek your master. It may be that the Spirit of the LORD has caught him up and cast him upon some mountain or into some valley." And he said, "You shall not send."
2KGS|2|17|But when they urged him till he was ashamed, he said, "Send." They sent therefore fifty men. And for three days they sought him but did not find him.
2KGS|2|18|And they came back to him while he was staying at Jericho, and he said to them, "Did I not say to you, 'Do not go'?"
2KGS|2|19|Now the men of the city said to Elisha, "Behold, the situation of this city is pleasant, as my lord sees, but the water is bad, and the land is unfruitful."
2KGS|2|20|He said, "Bring me a new bowl, and put salt in it." So they brought it to him.
2KGS|2|21|Then he went to the spring of water and threw salt in it and said, "Thus says the LORD, I have healed this water; from now on neither death nor miscarriage shall come from it."
2KGS|2|22|So the water has been healed to this day, according to the word that Elisha spoke.
2KGS|2|23|He went up from there to Bethel, and while he was going up on the way, some small boys came out of the city and jeered at him, saying, "Go up, you baldhead! Go up, you baldhead!"
2KGS|2|24|And he turned around, and when he saw them, he cursed them in the name of the LORD. And two she-bears came out of the woods and tore forty-two of the boys.
2KGS|2|25|From there he went on to Mount Carmel, and from there he returned to Samaria.
2KGS|3|1|In the eighteenth year of Jehoshaphat king of Judah, Jehoram the son of Ahab became king over Israel in Samaria, and he reigned twelve years.
2KGS|3|2|He did what was evil in the sight of the LORD, though not like his father and mother, for he put away the pillar of Baal that his father had made.
2KGS|3|3|Nevertheless, he clung to the sin of Jeroboam the son of Nebat, which he made Israel to sin; he did not depart from it.
2KGS|3|4|Now Mesha king of Moab was a sheep breeder, and he had to deliver to the king of Israel 100,000 lambs and the wool of 100,000 rams.
2KGS|3|5|But when Ahab died, the king of Moab rebelled against the king of Israel.
2KGS|3|6|So King Jehoram marched out of Samaria at that time and mustered all Israel.
2KGS|3|7|And he went and sent word to Jehoshaphat king of Judah, "The king of Moab has rebelled against me. Will you go with me to battle against Moab?" And he said, "I will go. I am as you are, my people as your people, my horses as your horses."
2KGS|3|8|Then he said, "By which way shall we march?" Jehoram answered, "By the way of the wilderness of Edom."
2KGS|3|9|So the king of Israel went with the king of Judah and the king of Edom. And when they had made a circuitous march of seven days, there was no water for the army or for the animals that followed them.
2KGS|3|10|Then the king of Israel said, "Alas! The LORD has called these three kings to give them into the hand of Moab."
2KGS|3|11|And Jehoshaphat said, "Is there no prophet of the LORD here, through whom we may inquire of the LORD?" Then one of the king of Israel's servants answered, "Elisha the son of Shaphat is here, who poured water on the hands of Elijah."
2KGS|3|12|And Jehoshaphat said, "The word of the LORD is with him." So the king of Israel and Jehoshaphat and the king of Edom went down to him.
2KGS|3|13|And Elisha said to the king of Israel, "What have I to do with you? Go to the prophets of your father and to the prophets of your mother." But the king of Israel said to him, "No; it is the LORD who has called these three kings to give them into the hand of Moab."
2KGS|3|14|And Elisha said, "As the LORD of hosts lives, before whom I stand, were it not that I have regard for Jehoshaphat the king of Judah, I would neither look at you nor see you.
2KGS|3|15|But now bring me a musician." And when the musician played, the hand of the LORD came upon him.
2KGS|3|16|And he said, "Thus says the LORD, 'I will make this dry streambed full of pools.'
2KGS|3|17|For thus says the LORD, 'You shall not see wind or rain, but that streambed shall be filled with water, so that you shall drink, you, your livestock, and your animals.'
2KGS|3|18|This is a light thing in the sight of the LORD. He will also give the Moabites into your hand,
2KGS|3|19|and you shall attack every fortified city and every choice city, and shall fell every good tree and stop up all springs of water and ruin every good piece of land with stones."
2KGS|3|20|The next morning, about the time of offering the sacrifice, behold, water came from the direction of Edom, till the country was filled with water.
2KGS|3|21|When all the Moabites heard that the kings had come up to fight against them, all who were able to put on armor, from the youngest to the oldest, were called out and were drawn up at the border.
2KGS|3|22|And when they rose early in phe morning and the sun shone on the water, the Moabites saw the water opposite them as red as blood.
2KGS|3|23|And they said, "This is blood; the kings have surely fought together and struck one another down. Now then, Moab, to the spoil!"
2KGS|3|24|But when they came to the camp of Israel, the Israelites rose and struck the Moabites, till they fled before them. And they went forward, striking the Moabites as they went.
2KGS|3|25|And they overthrew the cities, and on every good piece of land every man threw a stone until it was covered. They stopped every spring of water and felled all the good trees, till only its stones were left in Kir-hareseth, and the slingers surrounded and attacked it.
2KGS|3|26|When the king of Moab saw that the battle was going against him, he took with him 700 swordsmen to break through, opposite the king of Edom, but they could not.
2KGS|3|27|Then he took his oldest son who was to reign in his place and offered him for a burnt offering on the wall. And there came great wrath against Israel. And they withdrew from him and returned to their own land.
2KGS|4|1|Now the wife of one of the sons of the prophets cried to Elisha, "Your servant my husband is dead, and you know that your servant feared the LORD, but the creditor has come to take my two children to be his slaves."
2KGS|4|2|And Elisha said to her, "What shall I do for you? Tell me; what have you in the house?" And she said, "Your servant has nothing in the house except a jar of oil."
2KGS|4|3|Then he said, "Go outside, borrow vessels from all your neighbors, empty vessels and not too few.
2KGS|4|4|Then go in and shut the door behind yourself and your sons and pour into all these vessels. And when one is full, set it aside."
2KGS|4|5|So she went from him and shut the door behind herself and her sons. And as she poured they brought the vessels to her.
2KGS|4|6|When the vessels were full, she said to her son, "Bring me another vessel." And he said to her, "There is not another." Then the oil stopped flowing.
2KGS|4|7|She came and told the man of God, and he said, "Go, sell the oil and pay your debts, and you and your sons can live on the rest."
2KGS|4|8|One day Elisha went on to Shunem, where a wealthy woman lived, who urged him to eat some food. So whenever he passed that way, he would turn in there to eat food.
2KGS|4|9|And she said to her husband, "Behold now, I know that this is a holy man of God who is continually passing our way.
2KGS|4|10|Let us make a small room on the roof with walls and put there for him a bed, a table, a chair, and a lamp, so that whenever he comes to us, he can go in there."
2KGS|4|11|One day he came there, and he turned into the chamber and rested there.
2KGS|4|12|And he said to Gehazi his servant, "Call this Shunammite." When he had called her, she stood before him.
2KGS|4|13|And he said to him, "Say now to her, 'See, you have taken all this trouble for us; what is to be done for you? Would you have a word spoken on your behalf to the king or to the commander of the army?'"She answered, "I dwell among my own people."
2KGS|4|14|And he said, "What then is to be done for her?" Gehazi answered, "Well, she has no son, and her husband is old."
2KGS|4|15|He said, "Call her." And when he had called her, she stood in the doorway.
2KGS|4|16|And he said, "At this season, about this time next year, you shall embrace a son." And she said, "No, my lord, O man of God; do not lie to your servant."
2KGS|4|17|But the woman conceived, and she bore a son about that time the following spring, as Elisha had said to her.
2KGS|4|18|When the child had grown, he went out one day to his father among the reapers.
2KGS|4|19|And he said to his father, "Oh, my head, my head!" The father said to his servant, "Carry him to his mother."
2KGS|4|20|And when he had lifted him and brought him to his mother, the child sat on her lap till noon, and then he died.
2KGS|4|21|And she went up and laid him on the bed of the man of God and shut the door behind him and went out.
2KGS|4|22|Then she called to her husband and said, "Send me one of the servants and one of the donkeys, that I may quickly go to the man of God and come back again."
2KGS|4|23|And he said, "Why will you go to him today? It is neither new moon nor Sabbath." She said, "All is well."
2KGS|4|24|Then she saddled the donkey, and she said to her servant, "Urge the animal on; do not slacken the pace for me unless I tell you."
2KGS|4|25|So she set out and came to the man of God at Mount Carmel. When the man of God saw her coming, he said to Gehazi his servant, "Look, there is the Shunammite.
2KGS|4|26|Run at once to meet her and say to her, 'Is all well with you? Is all well with your husband? Is all well with the child?'"And she answered, "All is well."
2KGS|4|27|And when she came to the mountain to the man of God, she caught hold of his feet. And Gehazi came to push her away. But the man of God said, "Leave her alone, for she is in bitter distress, and the LORD has hidden it from me and has not told me."
2KGS|4|28|Then she said, "Did I ask my lord for a son? Did I not say, 'Do not deceive me?'"
2KGS|4|29|He said to Gehazi, "Tie up your garment and take my staff in your hand and go. If you meet anyone, do not greet him, and if anyone greets you, do not reply. And lay my staff on the face of the child."
2KGS|4|30|Then the mother of the child said, "As the LORD lives and as you yourself live, I will not leave you." So he arose and followed her.
2KGS|4|31|Gehazi went on ahead and laid the staff on the face of the child, but there was no sound or sign of life. Therefore he returned to meet him and told him, "The child has not awakened."
2KGS|4|32|When Elisha came into the house, he saw the child lying dead on his bed.
2KGS|4|33|So he went in and shut the door behind the two of them and prayed to the LORD.
2KGS|4|34|Then he went up and lay on the child, putting his mouth on his mouth, his eyes on his eyes, and his hands on his hands. And as he stretched himself upon him, the flesh of the child became warm.
2KGS|4|35|Then he got up again and walked once back and forth in the house, and went up and stretched himself upon him. The child sneezed seven times, and the child opened his eyes.
2KGS|4|36|Then he summoned Gehazi and said, "Call this Shunammite." So he called her. And when she came to him, he said, "Pick up your son."
2KGS|4|37|She came and fell at his feet, bowing to the ground. Then she picked up her son and went out.
2KGS|4|38|And Elisha came again to Gilgal when there was a famine in the land. And as the sons of the prophets were sitting before him, he said to his servant, "Set on the large pot, and boil stew for the sons of the prophets."
2KGS|4|39|One of them went out into the field to gather herbs, and found a wild vine and gathered from it his lap full of wild gourds, and came and cut them up into the pot of stew, not knowing what they were.
2KGS|4|40|And they poured out some for the men to eat. But while they were eating of the stew, they cried out, "O man of God, there is death in the pot!" And they could not eat it.
2KGS|4|41|He said, "Then bring flour." And he threw it into the pot and said, "Pour some out for the men, that they may eat." And there was no harm in the pot.
2KGS|4|42|A man came from Baal-shalishah, bringing the man of God bread of the firstfruits, twenty loaves of barley and fresh ears of grain in his sack. And Elisha said, "Give to the men, that they may eat."
2KGS|4|43|But his servant said, "How can I set this before a hundred men?" So he repeated, "Give them to the men, that they may eat, for thus says the LORD, 'They shall eat and have some left.'"
2KGS|4|44|So he set it before them. And they ate and had some left, according to the word of the LORD.
2KGS|5|1|Naaman, commander of the army of the king of Syria, was a great man with his master and in high favor, because by him the LORD had given victory to Syria. He was a mighty man of valor, but he was a leper.
2KGS|5|2|Now the Syrians on one of their raids had carried off a little girl from the land of Israel, and she worked in the service of Naaman's wife.
2KGS|5|3|She said to her mistress, "Would that my lord were with the prophet who is in Samaria! He would cure him of his leprosy."
2KGS|5|4|So Naaman went in and told his lord, "Thus and so spoke the girl from the land of Israel."
2KGS|5|5|And the king of Syria said, "Go now, and I will send a letter to the king of Israel." So he went, taking with him ten talents of silver, six thousand shekels of gold, and ten changes of clothes.
2KGS|5|6|And he brought the letter to the king of Israel, which read, "When this letter reaches you, know that I have sent to you Naaman my servant, that you may cure him of his leprosy."
2KGS|5|7|And when the king of Israel read the letter, he tore his clothes and said, "Am I God, to kill and to make alive, that this man sends word to me to cure a man of his leprosy? Only consider, and see how he is seeking a quarrel with me."
2KGS|5|8|But when Elisha the man of God heard that the king of Israel had torn his clothes, he sent to the king, saying, "Why have you torn your clothes? Let him come now to me, that he may know that there is a prophet in Israel."
2KGS|5|9|So Naaman came with his horses and chariots and stood at the door of Elisha's house.
2KGS|5|10|And Elisha sent a messenger to him, saying, "Go and wash in the Jordan seven times, and your flesh shall be restored, and you shall be clean."
2KGS|5|11|But Naaman was angry and went away, saying, "Behold, I thought that he would surely come out to me and stand and call upon the name of the LORD his God, and wave his hand over the place and cure the leper.
2KGS|5|12|Are not Abana and Pharpar, the rivers of Damascus, better than all the waters of Israel? Could I not wash in them and be clean?" So he turned and went away in a rage.
2KGS|5|13|But his servants came near and said to him, "My father, it is a great word the prophet has spoken to you; will you not do it? Has he actually said to you, 'Wash, and be clean'?"
2KGS|5|14|So he went down and dipped himself seven times in the Jordan, according to the word of the man of God, and his flesh was restored like the flesh of a little child, and he was clean.
2KGS|5|15|Then he returned to the man of God, he and all his company, and he came and stood before him. And he said, "Behold, I know that there is no God in all the earth but in Israel; so accept now a present from your servant."
2KGS|5|16|But he said, "As the LORD lives, before whom I stand, I will receive none." And he urged him to take it, but he refused.
2KGS|5|17|Then Naaman said, "If not, please let there be given to your servant two mules' load of earth, for from now on your servant will not offer burnt offering or sacrifice to any god but the LORD.
2KGS|5|18|In this matter may the LORD pardon your servant: when my master goes into the house of Rimmon to worship there, leaning on my arm, and I bow myself in the house of Rimmon, when I bow myself in the house of Rimmon, the LORD pardon your servant in this matter."
2KGS|5|19|He said to him, "Go in peace." But when Naaman had gone from him a short distance,
2KGS|5|20|Gehazi, the servant of Elisha the man of God, said, "See, my master has spared this Naaman the Syrian, in not accepting from his hand what he brought. As the LORD lives, I will run after him and get something from him."
2KGS|5|21|So Gehazi followed Naaman. And when Naaman saw someone running after him, he got down from the chariot to meet him and said, "Is all well?"
2KGS|5|22|And he said, "All is well. My master has sent me to say, 'There have just now come to me from the hill country of Ephraim two young men of the sons of the prophets. Please give them a talent of silver and two festal garments.'"
2KGS|5|23|And Naaman said, "Be pleased to accept two talents." And he urged him and tied up two talents of silver in two bags, with two festal garments, and laid them on two of his servants. And they carried them before Gehazi.
2KGS|5|24|And when he came to the hill, he took them from their hand and put them in the house, and he sent the men away, and they departed.
2KGS|5|25|He went in and stood before his master, and Elisha said to him, "Where have you been, Gehazi?" And he said, "Your servant went nowhere."
2KGS|5|26|But he said to him, "Did not my heart go when the man turned from his chariot to meet you? Was it a time to accept money and garments, olive orchards and vineyards, sheep and oxen, male servants and female servants?
2KGS|5|27|Therefore the leprosy of Naaman shall cling to you and to your descendants forever." So he went out from his presence a leper, like snow.
2KGS|6|1|Now the sons of the prophets said to Elisha, "See, the place where we dwell under your charge is too small for us.
2KGS|6|2|Let us go to the Jordan and each of us get there a log, and let us make a place for us to dwell there." And he answered, "Go."
2KGS|6|3|Then one of them said, "Be pleased to go with your servants." And he answered, "I will go."
2KGS|6|4|So he went with them. And when they came to the Jordan, they cut down trees.
2KGS|6|5|But as one was felling a log, his axe head fell into the water, and he cried out, "Alas, my master! It was borrowed."
2KGS|6|6|Then the man of God said, "Where did it fall?" When he showed him the place, he cut off a stick and threw it in there and made the iron float.
2KGS|6|7|And he said, "Take it up." So he reached out his hand and took it.
2KGS|6|8|Once when the king of Syria was warring against Israel, he took counsel with his servants, saying, "At such and such a place shall be my camp."
2KGS|6|9|But the man of God sent word to the king of Israel, "Beware that you do not pass this place, for the Syrians are going down there."
2KGS|6|10|And the king of Israel sent to the place about which the man of God told him. Thus he used to warn him, so that he saved himself there more than once or twice.
2KGS|6|11|And the mind of the king of Syria was greatly troubled because of this thing, and he called his servants and said to them, "Will you not show me who of us is for the king of Israel?"
2KGS|6|12|And one of his servants said, "None, my lord, O king; but Elisha, the prophet who is in Israel, tells the king of Israel the words that you speak in your bedroom."
2KGS|6|13|And he said, "Go and see where he is, that I may send and seize him." It was told him, "Behold, he is in Dothan."
2KGS|6|14|So he sent there horses and chariots and a great army, and they came by night and surrounded the city.
2KGS|6|15|When the servant of the man of God rose early in the morning and went out, behold, an army with horses and chariots was all around the city. And the servant said, "Alas, my master! What shall we do?"
2KGS|6|16|He said, "Do not be afraid, for those who are with us are more than those who are with them."
2KGS|6|17|Then Elisha prayed and said, "O LORD, please open his eyes that he may see." So the LORD opened the eyes of the young man, and he saw, and behold, the mountain was full of horses and chariots of fire all around Elisha.
2KGS|6|18|And when the Syrians came down against him, Elisha prayed to the LORD and said, "Please strike this people with blindness." So he struck them with blindness in accordance with the prayer of Elisha.
2KGS|6|19|And Elisha said to them, "This is not the way, and this is not the city. Follow me, and I will bring you to the man whom you seek." And he led them to Samaria.
2KGS|6|20|As soon as they entered Samaria, Elisha said, "O LORD, open the eyes of these men, that they may see." So the LORD opened their eyes and they saw, and behold, they were in the midst of Samaria.
2KGS|6|21|As soon as the king of Israel saw them, he said to Elisha, "My father, shall I strike them down? Shall I strike them down?"
2KGS|6|22|He answered, "You shall not strike them down. Would you strike down those whom you have taken captive with your sword and with your bow? Set bread and water before them, that they may eat and drink and go to their master."
2KGS|6|23|So he prepared for them a great feast, and when they had eaten and drunk, he sent them away, and they went to their master. And the Syrians did not come again on raids into the land of Israel.
2KGS|6|24|Afterward Ben-hadad king of Syria mustered his entire army and went up and besieged Samaria.
2KGS|6|25|And there was a great famine in Samaria, as they besieged it, until a donkey's head was sold for eighty shekels of silver, and the fourth part of a kab of dove's dung for five shekels of silver.
2KGS|6|26|Now as the king of Israel was passing by on the wall, a woman cried out to him, saying, "Help, my lord, O king!"
2KGS|6|27|And he said, "If the LORD will not help you, how shall I help you? From the threshing floor, or from the winepress?"
2KGS|6|28|And the king asked her, "What is your trouble?" She answered, "This woman said to me, 'Give your son, that we may eat him today, and we will eat my son tomorrow.'
2KGS|6|29|So we boiled my son and ate him. And on the next day I said to her, 'Give your son, that we may eat him.' But she has hidden her son."
2KGS|6|30|When the king heard the words of the woman, he tore his clothes- now he was passing by on the wall- and the people looked, and behold, he had sackcloth beneath on his body-
2KGS|6|31|and he said, "May God do so to me and more also, if the head of Elisha the son of Shaphat remains on his shoulders today."
2KGS|6|32|Elisha was sitting in his house, and the elders were sitting with him. Now the king had dispatched a man from his presence, but before the messenger arrived Elisha said to the elders, "Do you see how this murderer has sent to take off my head? Look, when the messenger comes, shut the door and hold the door fast against him. Is not the sound of his master's feet behind him?"
2KGS|6|33|And while he was still speaking with them, the messenger came down to him and said, "This trouble is from the LORD! Why should I wait for the LORD any longer?"
2KGS|7|1|But Elisha said, "Hear the word of the LORD: thus says the LORD, Tomorrow about this time a seah of fine flour shall be sold for a shekel, and two seahs of barley for a shekel, at the gate of Samaria."
2KGS|7|2|Then the captain on whose hand the king leaned said to the man of God, "If the LORD himself should make windows in heaven, could this thing be?" But he said, "You shall see it with your own eyes, but you shall not eat of it."
2KGS|7|3|Now there were four men who were lepers at the entrance to the gate. And they said to one another, "Why are we sitting here until we die?
2KGS|7|4|If we say, 'Let us enter the city,' the famine is in the city, and we shall die there. And if we sit here, we die also. So now come, let us go over to the camp of the Syrians. If they spare our lives we shall live, and if they kill us we shall but die."
2KGS|7|5|So they arose at twilight to go to the camp of the Syrians. But when they came to the edge of the camp of the Syrians, behold, there was no one there.
2KGS|7|6|For the Lord had made the army of the Syrians hear the sound of chariots and of horses, the sound of a great army, so that they said to one another, "Behold, the king of Israel has hired against us the kings of the Hittites and the kings of Egypt to come against us."
2KGS|7|7|So they fled away in the twilight and abandoned their tents, their horses, and their donkeys, leaving the camp as it was, and fled for their lives.
2KGS|7|8|And when these lepers came to the edge of the camp, they went into a tent and ate and drank, and they carried off silver and gold and clothing and went and hid them. Then they came back and entered another tent and carried off things from it and went and hid them.
2KGS|7|9|Then they said to one another, "We are not doing right. This day is a day of good news. If we are silent and wait until the morning light, punishment will overtake us. Now therefore come; let us go and tell the king's household."
2KGS|7|10|So they came and called to the gatekeepers of the city and told them, "We came to the camp of the Syrians, and behold, there was no one to be seen or heard there, nothing but the horses tied and the donkeys tied and the tents as they were."
2KGS|7|11|Then the gatekeepers called out, and it was told within the king's household.
2KGS|7|12|And the king rose in the night and said to his servants, "I will tell you what the Syrians have done to us. They know that we are hungry. Therefore they have gone out of the camp to hide themselves in the open country, thinking, 'When they come out of the city, we shall take them alive and get into the city.'"
2KGS|7|13|And one of his servants said, "Let some men take five of the remaining horses, seeing that those who are left here will fare like the whole multitude of Israel who have already perished. Let us send and see."
2KGS|7|14|So they took two horsemen, and the king sent them after the army of the Syrians, saying, "Go and see."
2KGS|7|15|So they went after them as far as the Jordan, and behold, all the way was littered with garments and equipment that the Syrians had thrown away in their haste. And the messengers returned and told the king.
2KGS|7|16|Then the people went out and plundered the camp of the Syrians. So a seah of fine flour was sold for a shekel, and two seahs of barley for a shekel, according to the word of the LORD.
2KGS|7|17|Now the king had appointed the captain on whose hand he leaned to have charge of the gate. And the people trampled him in the gate, so that he died, as the man of God had said when the king came down to him.
2KGS|7|18|For when the man of God had said to the king, "Two seahs of barley shall be sold for a shekel, and a seah of fine flour for a shekel, about this time tomorrow in the gate of Samaria,"
2KGS|7|19|the captain had answered the man of God, "If the LORD himself should make windows in heaven, could such a thing be?" And he had said, "You shall see it with your own eyes, but you shall not eat of it."
2KGS|7|20|And so it happened to him, for the people trampled him in the gate and he died.
2KGS|8|1|Now Elisha had said to the woman whose son he had restored to life, "Arise, and depart with your household, and sojourn wherever you can, for the LORD has called for a famine, and it will come upon the land for seven years."
2KGS|8|2|So the woman arose and did according to the word of the man of God. She went with her household and sojourned in the land of the Philistines seven years.
2KGS|8|3|And at the end of the seven years, when the woman returned from the land of the Philistines, she went to appeal to the king for her house and her land.
2KGS|8|4|Now the king was talking with Gehazi the servant of the man of God, saying, "Tell me all the great things that Elisha has done."
2KGS|8|5|And while he was telling the king how Elisha had restored the dead to life, behold, the woman whose son he had restored to life appealed to the king for her house and her land. And Gehazi said, "My lord, O king, here is the woman, and here is her son whom Elisha restored to life."
2KGS|8|6|And when the king asked the woman, she told him. So the king appointed an official for her, saying, "Restore all that was hers, together with all the produce of the fields from the day that she left the land until now."
2KGS|8|7|Now Elisha came to Damascus. Ben-hadad the king of Syria was sick. And when it was told him, "The man of God has come here,"
2KGS|8|8|the king said to Hazael, "Take a present with you and go to meet the man of God, and inquire of the LORD through him, saying, 'Shall I recover from this sickness?'"
2KGS|8|9|So Hazael went to meet him, and took a present with him, all kinds of goods of Damascus, forty camel loads. When he came and stood before him, he said, "Your son Ben-hadad king of Syria has sent me to you, saying, 'Shall I recover from this sickness?'"
2KGS|8|10|And Elisha said to him, "Go, say to him, 'You shall certainly recover,' but the LORD has shown me that he shall certainly die."
2KGS|8|11|And he fixed his gaze and stared at him, until he was embarrassed. And the man of God wept.
2KGS|8|12|And Hazael said, "Why does my lord weep?" He answered, "Because I know the evil that you will do to the people of Israel. You will set on fire their fortresses, and you will kill their young men with the sword and dash in pieces their little ones and rip open their pregnant women."
2KGS|8|13|And Hazael said, "What is your servant, who is but a dog, that he should do this great thing?" Elisha answered, "The LORD has shown me that you are to be king over Syria."
2KGS|8|14|Then he departed from Elisha and came to his master, who said to him, "What did Elisha say to you?" And he answered, "He told me that you would certainly recover."
2KGS|8|15|But the next day he took the bed cloth and dipped it in water and spread it over his face, till he died. And Hazael became king in his place.
2KGS|8|16|In the fifth year of Joram the son of Ahab, king of Israel, when Jehoshaphat was king of Judah, Jehoram the son of Jehoshaphat, king of Judah, began to reign.
2KGS|8|17|He was thirty-two years old when he became king, and he reigned eight years in Jerusalem.
2KGS|8|18|And he walked in the way of the kings of Israel, as the house of Ahab had done, for the daughter of Ahab was his wife. And he did what was evil in the sight of the LORD.
2KGS|8|19|Yet the LORD was not willing to destroy Judah, for the sake of David his servant, since he promised to give a lamp to him and to his sons forever.
2KGS|8|20|In his days Edom revolted from the rule of Judah and set up a king of their own.
2KGS|8|21|Then Joram passed over to Zair with all his chariots and rose by night, and he and his chariot commanders struck the Edomites who had surrounded him, but his army fled home.
2KGS|8|22|So Edom revolted from the rule of Judah to this day. Then Libnah revolted at the same time.
2KGS|8|23|Now the rest of the acts of Joram, and all that he did, are they not written in the Book of the Chronicles of the Kings of Judah?
2KGS|8|24|So Joram slept with his fathers and was buried with his fathers in the city of David, and Ahaziah his son reigned in his place.
2KGS|8|25|In the twelfth year of Joram the son of Ahab, king of Israel, Ahaziah the son of Jehoram, king of Judah, began to reign.
2KGS|8|26|Ahaziah was twenty-two years old when he began to reign, and he reigned one year in Jerusalem. His mother's name was Athaliah; she was a granddaughter of Omri king of Israel.
2KGS|8|27|He also walked in the way of the house of Ahab and did what was evil in the sight of the LORD, as the house of Ahab had done, for he was son-in-law to the house of Ahab.
2KGS|8|28|He went with Joram the son of Ahab to make war against Hazael king of Syria at Ramoth-gilead, and the Syrians wounded Joram.
2KGS|8|29|And King Joram returned to be healed in Jezreel of the wounds that the Syrians had given him at Ramah, when he fought against Hazael king of Syria. And Ahaziah the son of Jehoram king of Judah went down to see Joram the son of Ahab in Jezreel, because he was sick.
2KGS|9|1|Then Elisha the prophet called one of the sons of the prophets and said to him, "Tie up your garments, and take this flask of oil in your hand, and go to Ramoth-gilead.
2KGS|9|2|And when you arrive, look there for Jehu the son of Jehoshaphat, son of Nimshi. And go in and have him rise from among his fellows, and lead him to an inner chamber.
2KGS|9|3|Then take the flask of oil and pour it on his head and say, 'Thus says the LORD, I anoint you king over Israel.' Then open the door and flee; do not linger."
2KGS|9|4|So the young man, the servant of the prophet, went to Ramoth-gilead.
2KGS|9|5|And when he came, behold, the commanders of the army were in council. And he said, "I have a word for you, O commander." And Jehu said, "To which of us all?" And he said, "To you, O commander."
2KGS|9|6|So he arose and went into the house. And the young man poured the oil on his head, saying to him, "Thus says the LORD the God of Israel, I anoint you king over the people of the LORD, over Israel.
2KGS|9|7|And you shall strike down the house of Ahab your master, so that I may avenge on Jezebel the blood of my servants the prophets, and the blood of all the servants of the LORD.
2KGS|9|8|For the whole house of Ahab shall perish, and I will cut off from Ahab every male, bond or free, in Israel.
2KGS|9|9|And I will make the house of Ahab like the house of Jeroboam the son of Nebat, and like the house of Baasha the son of Ahijah.
2KGS|9|10|And the dogs shall eat Jezebel in the territory of Jezreel, and none shall bury her." Then he opened the door and fled.
2KGS|9|11|When Jehu came out to the servants of his master, they said to him, "Is all well? Why did this mad fellow come to you?" And he said to them, "You know the fellow and his talk."
2KGS|9|12|And they said, "That is not true; tell us now." And he said, "Thus and so he spoke to me, saying, 'Thus says the LORD, I anoint you king over Israel.'"
2KGS|9|13|Then in haste every man of them took his garment and put it under him on the bare steps, and they blew the trumpet and proclaimed, "Jehu is king."
2KGS|9|14|Thus Jehu the son of Jehoshaphat the son of Nimshi conspired against Joram. (Now Joram with all Israel had been on guard at Ramoth-gilead against Hazael king of Syria,
2KGS|9|15|but King Joram had returned to be healed in Jezreel of the wounds that the Syrians had given him, when he fought with Hazael king of Syria.) So Jehu said, "If this is your decision, then let no one slip out of the city to go and tell the news in Jezreel."
2KGS|9|16|Then Jehu mounted his chariot and went to Jezreel, for Joram lay there. And Ahaziah king of Judah had come down to visit Joram.
2KGS|9|17|Now the watchman was standing on the tower in Jezreel, and he saw the company of Jehu as he came and said, "I see a company." And Joram said, "Take a horseman and send to meet them, and let him say, 'Is it peace?'"
2KGS|9|18|So a man on horseback went to meet him and said, "Thus says the king, 'Is it peace?'"And Jehu said, "What do you have to do with peace? Turn around and ride behind me." And the watchman reported, saying, "The messenger reached them, but he is not coming back."
2KGS|9|19|Then he sent out a second horseman, who came to them and said, "Thus the king has said, 'Is it peace?'"And Jehu answered, "What do you have to do with peace? Turn around and ride behind me."
2KGS|9|20|Again the watchman reported, "He reached them, but he is not coming back. And the driving is like the driving of Jehu the son of Nimshi, for he drives furiously."
2KGS|9|21|Joram said, "Make ready." And they made ready his chariot. Then Joram king of Israel and Ahaziah king of Judah set out, each in his chariot, and went to meet Jehu, and met him at the property of Naboth the Jezreelite.
2KGS|9|22|And when Joram saw Jehu, he said, "Is it peace, Jehu?" He answered, "What peace can there be, so long as the whorings and the sorceries of your mother Jezebel are so many?"
2KGS|9|23|Then Joram reined about and fled, saying to Ahaziah, "Treachery, O Ahaziah!"
2KGS|9|24|And Jehu drew his bow with his full strength, and shot Joram between the shoulders, so that the arrow pierced his heart, and he sank in his chariot.
2KGS|9|25|Jehu said to Bidkar his aide, "Take him up and throw him on the plot of ground belonging to Naboth the Jezreelite. For remember, when you and I rode side by side behind Ahab his father, how the LORD made this pronouncement against him:
2KGS|9|26|'As surely as I saw yesterday the blood of Naboth and the blood of his sons- declares the LORD- I will repay you on this plot of ground.' Now therefore take him up and throw him on the plot of ground, in accordance with the word of the LORD."
2KGS|9|27|When Ahaziah the king of Judah saw this, he fled in the direction of Beth-haggan. And Jehu pursued him and said, "Shoot him also." And they shot him in the chariot at the ascent of Gur, which is by Ibleam. And he fled to Megiddo and died there.
2KGS|9|28|His servants carried him in a chariot to Jerusalem, and buried him in his tomb with his fathers in the city of David.
2KGS|9|29|In the eleventh year of Joram the son of Ahab, Ahaziah began to reign over Judah.
2KGS|9|30|When Jehu came to Jezreel, Jezebel heard of it. And she painted her eyes and adorned her head and looked out of the window.
2KGS|9|31|And as Jehu entered the gate, she said, "Is it peace, you Zimri, murderer of your master?"
2KGS|9|32|And he lifted up his face to the window and said, "Who is on my side? Who?" Two or three eunuchs looked out at him.
2KGS|9|33|He said, "Throw her down." So they threw her down. And some of her blood spattered on the wall and on the horses, and they trampled on her.
2KGS|9|34|Then he went in and ate and drank. And he said, "See now to this cursed woman and bury her, for she is a king's daughter."
2KGS|9|35|But when they went to bury her, they found no more of her than the skull and the feet and the palms of her hands.
2KGS|9|36|When they came back and told him, he said, "This is the word of the LORD, which he spoke by his servant Elijah the Tishbite, 'In the territory of Jezreel the dogs shall eat the flesh of Jezebel,
2KGS|9|37|and the corpse of Jezebel shall be as dung on the face of the field in the territory of Jezreel, so that no one can say, This is Jezebel.'"
2KGS|10|1|Now Ahab had seventy sons in Samaria. So Jehu wrote letters and sent them to Samaria, to the rulers of the city, to the elders, and to the guardians of the sons of Ahab, saying,
2KGS|10|2|"Now then, as soon as this letter comes to you, seeing your master's sons are with you, and there are with you chariots and horses, fortified cities also, and weapons,
2KGS|10|3|select the best and fittest of your master's sons and set him on his father's throne and fight for your master's house."
2KGS|10|4|But they were exceedingly afraid and said, "Behold, the two kings could not stand before him. How then can we stand?"
2KGS|10|5|So he who was over the palace, and he who was over the city, together with the elders and the guardians, sent to Jehu, saying, "We are your servants, and we will do all that you tell us. We will not make anyone king. Do whatever is good in your eyes."
2KGS|10|6|Then he wrote to them a second letter, saying, "If you are on my side, and if you are ready to obey me, take the heads of your master's sons and come to me at Jezreel tomorrow at this time." Now the king's sons, seventy persons, were with the great men of the city, who were bringing them up.
2KGS|10|7|And as soon as the letter came to them, they took the king's sons and slaughtered them, seventy persons, and put their heads in baskets and sent them to him at Jezreel.
2KGS|10|8|When the messenger came and told him, "They have brought the heads of the king's sons," he said, "Lay them in two heaps at the entrance of the gate until the morning."
2KGS|10|9|Then in the morning, when he went out, he stood and said to all the people, "You are innocent. It was I who conspired against my master and killed him, but who struck down all these?
2KGS|10|10|Know then that there shall fall to the earth nothing of the word of the LORD, which the LORD spoke concerning the house of Ahab, for the LORD has done what he said by his servant Elijah."
2KGS|10|11|So Jehu struck down all who remained of the house of Ahab in Jezreel, all his great men and his close friends and his priests, until he left him none remaining.
2KGS|10|12|Then he set out and went to Samaria. On the way, when he was at Beth-eked of the Shepherds,
2KGS|10|13|Jehu met the relatives of Ahaziah king of Judah, and he said, "Who are you?" And they answered, "We are the relatives of Ahaziah, and we came down to visit the royal princes and the sons of the queen mother."
2KGS|10|14|He said, "Take them alive." And they took them alive and slaughtered them at the pit of Beth-eked, forty-two persons, and he spared none of them.
2KGS|10|15|And when he departed from there, he met Jehonadab the son of Rechab coming to meet him. And he greeted him and said to him, "Is your heart true to my heart as mine is to yours?" And Jehonadab answered, "It is." Jehu said, "If it is, give me your hand." So he gave him his hand. And Jehu took him up with him into the chariot.
2KGS|10|16|And he said, "Come with me, and see my zeal for the LORD." So he had him ride in his chariot.
2KGS|10|17|And when he came to Samaria, he struck down all who remained to Ahab in Samaria, till he had wiped them out, according to the word of the LORD that he spoke to Elijah.
2KGS|10|18|Then Jehu assembled all the people and said to them, "Ahab served Baal a little, but Jehu will serve him much.
2KGS|10|19|Now therefore call to me all the prophets of Baal, all his worshipers and all his priests. Let none be missing, for I have a great sacrifice to offer to Baal. Whoever is missing shall not live." But Jehu did it with cunning in order to destroy the worshipers of Baal.
2KGS|10|20|And Jehu ordered, "Sanctify a solemn assembly for Baal." So they proclaimed it.
2KGS|10|21|And Jehu sent throughout all Israel, and all the worshipers of Baal came, so that there was not a man left who did not come. And they entered the house of Baal, and the house of Baal was filled from one end to the other.
2KGS|10|22|He said to him who was in charge of the wardrobe, "Bring out the vestments for all the worshipers of Baal." So he brought out the vestments for them.
2KGS|10|23|Then Jehu went into the house of Baal with Jehonadab the son of Rechab, and he said to the worshipers of Baal, "Search, and see that there is no servant of the LORD here among you, but only the worshipers of Baal."
2KGS|10|24|Then they went in to offer sacrifices and burnt offerings. Now Jehu had stationed eighty men outside and said, "The man who allows any of those whom I give into your hands to escape shall forfeit his life."
2KGS|10|25|So as soon as he had made an end of offering the burnt offering, Jehu said to the guard and to the officers, "Go in and strike them down; let not a man escape." So when they put them to the sword, the guard and the officers cast them out and went into the inner room of the house of Baal,
2KGS|10|26|and they brought out the pillar that was in the house of Baal and burned it.
2KGS|10|27|And they demolished the pillar of Baal, and demolished the house of Baal, and made it a latrine to this day.
2KGS|10|28|Thus Jehu wiped out Baal from Israel.
2KGS|10|29|But Jehu did not turn aside from the sins of Jeroboam the son of Nebat, which he made Israel to sin- that is, the golden calves that were in Bethel and in Dan.
2KGS|10|30|And the LORD said to Jehu, "Because you have done well in carrying out what is right in my eyes, and have done to the house of Ahab according to all that was in my heart, your sons of the fourth generation shall sit on the throne of Israel."
2KGS|10|31|But Jehu was not careful to walk in the law of the LORD the God of Israel with all his heart. He did not turn from the sins of Jeroboam, which he made Israel to sin.
2KGS|10|32|In those days the LORD began to cut off parts of Israel. Hazael defeated them throughout the territory of Israel:
2KGS|10|33|from the Jordan eastward, all the land of Gilead, the Gadites, and the Reubenites, and the Manassites, from Aroer, which is by the Valley of the Arnon, that is, Gilead and Bashan.
2KGS|10|34|Now the rest of the acts of Jehu and all that he did, and all his might, are they not written in the Book of the Chronicles of the Kings of Israel?
2KGS|10|35|So Jehu slept with his fathers, and they buried him in Samaria. And Jehoahaz his son reigned in his place.
2KGS|10|36|The time that Jehu reigned over Israel in Samaria was twenty-eight years.
2KGS|11|1|Now when Athaliah the mother of Ahaziah saw that her son was dead, she arose and destroyed all the royal family.
2KGS|11|2|But Jehosheba, the daughter of King Joram, sister of Ahaziah, took Joash the son of Ahaziah and stole him away from among the king's sons who were being put to death, and she put him and his nurse in a bedroom. Thus they hid him from Athaliah, so that he was not put to death.
2KGS|11|3|And he remained with her six years, hidden in the house of the LORD, while Athaliah reigned over the land.
2KGS|11|4|But in the seventh year Jehoiada sent and brought the captains of the Carites and of the guards, and had them come to him in the house of the LORD. And he made a covenant with them and put them under oath in the house of the LORD, and he showed them the king's son.
2KGS|11|5|And he commanded them, "This is the thing that you shall do: one third of you, those who come off duty on the Sabbath and guard the king's house
2KGS|11|6|(another third being at the gate Sur and a third at the gate behind the guards) shall guard the palace.
2KGS|11|7|And the two divisions of you, which come on duty in force on the Sabbath and guard the house of the LORD on behalf of the king,
2KGS|11|8|shall surround the king, each with his weapons in his hand. And whoever approaches the ranks is to be put to death. Be with the king when he goes out and when he comes in."
2KGS|11|9|The captains did according to all that Jehoiada the priest commanded, and they each brought his men who were to go off duty on the Sabbath, with those who were to come on duty on the Sabbath, and came to Jehoiada the priest.
2KGS|11|10|And the priest gave to the captains the spears and shields that had been King David's, which were in the house of the LORD.
2KGS|11|11|And the guards stood, every man with his weapons in his hand, from the south side of the house to the north side of the house, around the altar and the house on behalf of the king.
2KGS|11|12|Then he brought out the king's son and put the crown on him and gave him the testimony. And they proclaimed him king and anointed him, and they clapped their hands and said, "Long live the king!"
2KGS|11|13|When Athaliah heard the noise of the guard and of the people, she went into the house of the LORD to the people.
2KGS|11|14|And when she looked, there was the king standing by the pillar, according to the custom, and the captains and the trumpeters beside the king, and all the people of the land rejoicing and blowing trumpets. And Athaliah tore her clothes and cried, "Treason! Treason!"
2KGS|11|15|Then Jehoiada the priest commanded the captains who were set over the army, "Bring her out between the ranks, and put to death with the sword anyone who follows her." For the priest said, "Let her not be put to death in the house of the LORD."
2KGS|11|16|So they laid hands on her; and she went through the horses' entrance to the king's house, and there she was put to death.
2KGS|11|17|And Jehoiada made a covenant between the LORD and the king and people, that they should be the LORD's people, and also between the king and the people.
2KGS|11|18|Then all the people of the land went to the house of Baal and tore it down; his altars and his images they broke in pieces, and they killed Mattan the priest of Baal before the altars. And the priest posted watchmen over the house of the LORD.
2KGS|11|19|And he took the captains, the Carites, the guards, and all the people of the land, and they brought the king down from the house of the LORD, marching through the gate of the guards to the king's house. And he took his seat on the throne of the kings.
2KGS|11|20|So all the people of the land rejoiced, and the city was quiet after Athaliah had been put to death with the sword at the king's house.
2KGS|11|21|Jehoash was seven years old when he began to reign.
2KGS|12|1|In the seventh year of Jehu, Jehoash began to reign, and he reigned forty years in Jerusalem. His mother's name was Zibiah of Beersheba.
2KGS|12|2|And Jehoash did what was right in the eyes of the LORD all his days, because Jehoiada the priest instructed him.
2KGS|12|3|Nevertheless, the high places were not taken away; the people continued to sacrifice and make offerings on the high places.
2KGS|12|4|Jehoash said to the priests, "All the money of the holy things that is brought into the house of the LORD, the money for which each man is assessed- the money from the assessment of persons- and the money that a man's heart prompts him to bring into the house of the LORD,
2KGS|12|5|let the priests take, each from his donor, and let them repair the house wherever any need of repairs is discovered."
2KGS|12|6|But by the twenty-third year of King Jehoash, the priests had made no repairs on the house.
2KGS|12|7|Therefore King Jehoash summoned Jehoiada the priest and the other priests and said to them, "Why are you not repairing the house? Now therefore take no more money from your donors, but hand it over for the repair of the house."
2KGS|12|8|So the priests agreed that they should take no more money from the people, and that they should not repair the house.
2KGS|12|9|Then Jehoiada the priest took a chest and bored a hole in the lid of it and set it beside the altar on the right side as one entered the house of the LORD. And the priests who guarded the threshold put in it all the money that was brought into the house of the LORD.
2KGS|12|10|And whenever they saw that there was much money in the chest, the king's secretary and the high priest came up and they bagged and counted the money that was found in the house of the LORD.
2KGS|12|11|Then they would give the money that was weighed out into the hands of the workmen who had the oversight of the house of the LORD. And they paid it out to the carpenters and the builders who worked on the house of the LORD,
2KGS|12|12|and to the masons and the stonecutters, as well as to buy timber and quarried stone for making repairs on the house of the LORD, and for any outlay for the repairs of the house.
2KGS|12|13|But there were not made for the house of the LORD basins of silver, snuffers, bowls, trumpets, or any vessels of gold, or of silver, from the money that was brought into the house of the LORD,
2KGS|12|14|for that was given to the workmen who were repairing the house of the LORD with it.
2KGS|12|15|And they did not ask an accounting from the men into whose hand they delivered the money to pay out to the workmen, for they dealt honestly.
2KGS|12|16|The money from the guilt offerings and the money from the sin offerings was not brought into the house of the LORD; it belonged to the priests.
2KGS|12|17|At that time Hazael king of Syria went up and fought against Gath and took it. But when Hazael set his face to go up against Jerusalem,
2KGS|12|18|Jehoash king of Judah took all the sacred gifts that Jehoshaphat and Jehoram and Ahaziah his fathers, the kings of Judah, had dedicated, and his own sacred gifts, and all the gold that was found in the treasuries of the house of the LORD and of the king's house, and sent these to Hazael king of Syria. Then Hazael went away from Jerusalem.
2KGS|12|19|Now the rest of the acts of Joash and all that he did, are they not written in the Book of the Chronicles of the Kings of Judah?
2KGS|12|20|His servants arose and made a conspiracy and struck down Joash in the house of Millo, on the way that goes down to Silla.
2KGS|12|21|It was Jozacar the son of Shimeath and Jehozabad the son of Shomer, his servants, who struck him down, so that he died. And they buried him with his fathers in the city of David, and Amaziah his son reigned in his place.
2KGS|13|1|In the twenty-third year of Joash the son of Ahaziah, king of Judah, Jehoahaz the son of Jehu began to reign over Israel in Samaria, and he reigned seventeen years.
2KGS|13|2|He did what was evil in the sight of the LORD and followed the sins of Jeroboam the son of Nebat, which he made Israel to sin; he did not depart from them.
2KGS|13|3|And the anger of the LORD was kindled against Israel, and he gave them continually into the hand of Hazael king of Syria and into the hand of Ben-hadad the son of Hazael.
2KGS|13|4|Then Jehoahaz sought the favor of the LORD, and the LORD listened to him, for he saw the oppression of Israel, how the king of Syria oppressed them.
2KGS|13|5|(Therefore the LORD gave Israel a savior, so that they escaped from the hand of the Syrians, and the people of Israel lived in their homes as formerly.
2KGS|13|6|Nevertheless, they did not depart from the sins of the house of Jeroboam, which he made Israel to sin, but walked in them; and the Asherah also remained in Samaria.)
2KGS|13|7|For there was not left to Jehoahaz an army of more than fifty horsemen and ten chariots and ten thousand footmen, for the king of Syria had destroyed them and made them like the dust at threshing.
2KGS|13|8|Now the rest of the acts of Jehoahaz and all that he did, and his might, are they not written in the Book of the Chronicles of the Kings of Israel?
2KGS|13|9|So Jehoahaz slept with his fathers, and they buried him in Samaria, and Joash his son reigned in his place.
2KGS|13|10|In the thirty-seventh year of Joash king of Judah, Jehoash the son of Jehoahaz began to reign over Israel in Samaria, and he reigned sixteen years.
2KGS|13|11|He also did what was evil in the sight of the LORD. He did not depart from all the sins of Jeroboam the son of Nebat, which he made Israel to sin, but he walked in them.
2KGS|13|12|Now the rest of the acts of Joash and all that he did, and the might with which he fought against Amaziah king of Judah, are they not written in the Book of the Chronicles of the Kings of Israel?
2KGS|13|13|So Joash slept with his fathers, and Jeroboam sat on his throne. And Joash was buried in Samaria with the kings of Israel.
2KGS|13|14|Now when Elisha had fallen sick with the illness of which he was to die, Joash king of Israel went down to him and wept before him, crying, "My father, my father! The chariots of Israel and its horsemen!"
2KGS|13|15|And Elisha said to him, "Take a bow and arrows." So he took a bow and arrows.
2KGS|13|16|Then he said to the king of Israel, "Draw the bow," and he drew it. And Elisha laid his hands on the king's hands.
2KGS|13|17|And he said, "Open the window eastward," and he opened it. Then Elisha said, "Shoot," and he shot. And he said, "The LORD's arrow of victory, the arrow of victory over Syria! For you shall fight the Syrians in Aphek until you have made an end of them."
2KGS|13|18|And he said, "Take the arrows," and he took them. And he said to the king of Israel, "Strike the ground with them." And he struck three times and stopped.
2KGS|13|19|Then the man of God was angry with him and said, "You should have struck five or six times; then you would have struck down Syria until you had made an end of it, but now you will strike down Syria only three times."
2KGS|13|20|So Elisha died, and they buried him. Now bands of Moabites used to invade the land in the spring of the year.
2KGS|13|21|And as a man was being buried, behold, a marauding band was seen and the man was thrown into the grave of Elisha, and as soon as the man touched the bones of Elisha, he revived and stood on his feet.
2KGS|13|22|Now Hazael king of Syria oppressed Israel all the days of Jehoahaz.
2KGS|13|23|But the LORD was gracious to them and had compassion on them, and he turned toward them, because of his covenant with Abraham, Isaac, and Jacob, and would not destroy them, nor has he cast them from his presence until now.
2KGS|13|24|When Hazael king of Syria died, Ben-hadad his son became king in his place.
2KGS|13|25|Then Jehoash the son of Jehoahaz took again from Ben-hadad the son of Hazael the cities that he had taken from Jehoahaz his father in war. Three times Joash defeated him and recovered the cities of Israel.
2KGS|14|1|In the second year of Joash the son of Joahaz, king of Israel, Amaziah the son of Joash, king of Judah, began to reign.
2KGS|14|2|He was twenty-five years old when he began to reign, and he reigned twenty-nine years in Jerusalem. His mother's name was Jehoaddin of Jerusalem.
2KGS|14|3|And he did what was right in the eyes of the LORD, yet not like David his father. He did in all things as Joash his father had done.
2KGS|14|4|But the high places were not removed; the people still sacrificed and made offerings on the high places.
2KGS|14|5|And as soon as the royal power was firmly in his hand, he struck down his servants who had struck down the king his father.
2KGS|14|6|But he did not put to death the children of the murderers, according to what is written in the Book of the Law of Moses, where the LORD commanded, "Fathers shall not be put to death because of their children, nor shall children be put to death because of their fathers. But each one shall die for his own sin."
2KGS|14|7|He struck down ten thousand Edomites in the Valley of Salt and took Sela by storm, and called it Joktheel, which is its name to this day.
2KGS|14|8|Then Amaziah sent messengers to Jehoash the son of Jehoahaz, son of Jehu, king of Israel, saying, "Come, let us look one another in the face."
2KGS|14|9|And Jehoash king of Israel sent word to Amaziah king of Judah, "A thistle on Lebanon sent to a cedar on Lebanon, saying, 'Give your daughter to my son for a wife,' and a wild beast of Lebanon passed by and trampled down the thistle.
2KGS|14|10|You have indeed struck down Edom, and your heart has lifted you up. Be content with your glory, and stay at home, for why should you provoke trouble so that you fall, you and Judah with you?"
2KGS|14|11|But Amaziah would not listen. So Jehoash king of Israel went up, and he and Amaziah king of Judah faced one another in battle at Beth-shemesh, which belongs to Judah.
2KGS|14|12|And Judah was defeated by Israel, and every man fled to his home.
2KGS|14|13|And Jehoash king of Israel captured Amaziah king of Judah, the son of Jehoash, son of Ahaziah, at Beth-shemesh, and came to Jerusalem and broke down the wall of Jerusalem for four hundred cubits, from the Ephraim Gate to the Corner Gate.
2KGS|14|14|And he seized all the gold and silver, and all the vessels that were found in the house of the LORD and in the treasuries of the king's house, also hostages, and he returned to Samaria.
2KGS|14|15|Now the rest of the acts of Jehoash that he did, and his might, and how he fought with Amaziah king of Judah, are they not written in the Book of the Chronicles of the Kings of Israel?
2KGS|14|16|And Jehoash slept with his fathers and was buried in Samaria with the kings of Israel, and Jeroboam his son reigned in his place.
2KGS|14|17|Amaziah the son of Joash, king of Judah, lived fifteen years after the death of Jehoash son of Jehoahaz, king of Israel.
2KGS|14|18|Now the rest of the deeds of Amaziah, are they not written in the Book of the Chronicles of the Kings of Judah?
2KGS|14|19|And they made a conspiracy against him in Jerusalem, and he fled to Lachish. But they sent after him to Lachish and put him to death there.
2KGS|14|20|And they brought him on horses; and he was buried in Jerusalem with his fathers in the city of David.
2KGS|14|21|And all the people of Judah took Azariah, who was sixteen years old, and made him king instead of his father Amaziah.
2KGS|14|22|He built Elath and restored it to Judah, after the king slept with his fathers.
2KGS|14|23|In the fifteenth year of Amaziah the son of Joash, king of Judah, Jeroboam the son of Joash, king of Israel, began to reign in Samaria, and he reigned forty-one years.
2KGS|14|24|And he did what was evil in the sight of the LORD. He did not depart from all the sins of Jeroboam the son of Nebat, which he made Israel to sin.
2KGS|14|25|He restored the border of Israel from Lebo-hamath as far as the Sea of the Arabah, according to the word of the LORD, the God of Israel, which he spoke by his servant Jonah the son of Amittai, the prophet, who was from Gath-hepher.
2KGS|14|26|For the LORD saw that the affliction of Israel was very bitter, for there was none left, bond or free, and there was none to help Israel.
2KGS|14|27|But the LORD had not said that he would blot out the name of Israel from under heaven, so he saved them by the hand of Jeroboam the son of Joash.
2KGS|14|28|Now the rest of the acts of Jeroboam and all that he did, and his might, how he fought, and how he restored Damascus and Hamath to Judah in Israel, are they not written in the Book of the Chronicles of the Kings of Israel?
2KGS|14|29|And Jeroboam slept with his fathers, the kings of Israel, and Zechariah his son reigned in his place.
2KGS|15|1|In the twenty-seventh year of Jeroboam king of Israel, Azariah the son of Amaziah, king of Judah, began to reign.
2KGS|15|2|He was sixteen years old when he began to reign, and he reigned fifty-two years in Jerusalem. His mother's name was Jecoliah of Jerusalem.
2KGS|15|3|And he did what was right in the eyes of the LORD, according to all that his father Amaziah had done.
2KGS|15|4|Nevertheless, the high places were not taken away. The people still sacrificed and made offerings on the high places.
2KGS|15|5|And the LORD touched the king, so that he was a leper to the day of his death, and he lived in a separate house. And Jotham the king's son was over the household, governing the people of the land.
2KGS|15|6|Now the rest of the acts of Azariah, and all that he did, are they not written in the Book of the Chronicles of the Kings of Judah?
2KGS|15|7|And Azariah slept with his fathers, and they buried him with his fathers in the city of David, and Jotham his son reigned in his place.
2KGS|15|8|In the thirty-eighth year of Azariah king of Judah, Zechariah the son of Jeroboam reigned over Israel in Samaria six months.
2KGS|15|9|And he did what was evil in the sight of the LORD, as his fathers had done. He did not depart from the sins of Jeroboam the son of Nebat, which he made Israel to sin.
2KGS|15|10|Shallum the son of Jabesh conspired against him and struck him down at Ibleam and put him to death and reigned in his place.
2KGS|15|11|Now the rest of the deeds of Zechariah, behold, they are written in the Book of the Chronicles of the Kings of Israel.
2KGS|15|12|(This was the promise of the LORD that he gave to Jehu, "Your sons shall sit on the throne of Israel to the fourth generation." And so it came to pass.)
2KGS|15|13|Shallum the son of Jabesh began to reign in the thirty-ninth year of Uzziah king of Judah, and he reigned one month in Samaria.
2KGS|15|14|Then Menahem the son of Gadi came up from Tirzah and came to Samaria, and he struck down Shallum the son of Jabesh in Samaria and put him to death and reigned in his place.
2KGS|15|15|Now the rest of the deeds of Shallum, and the conspiracy that he made, behold, they are written in the Book of the Chronicles of the Kings of Israel.
2KGS|15|16|At that time Menahem sacked Tiphsah and all who were in it and its territory from Tirzah on, because they did not open it to him. Therefore he sacked it, and he ripped open all the women in it who were pregnant.
2KGS|15|17|In the thirty-ninth year of Azariah king of Judah, Menahem the son of Gadi began to reign over Israel, and he reigned ten years in Samaria.
2KGS|15|18|And he did what was evil in the sight of the LORD. He did not depart all his days from all the sins of Jeroboam the son of Nebat, which he made Israel to sin.
2KGS|15|19|Pul the king of Assyria came against the land, and Menahem gave Pul a thousand talents of silver, that he might help him to confirm his hold on the royal power.
2KGS|15|20|Menahem exacted the money from Israel, that is, from all the wealthy men, fifty shekels of silver from every man, to give to the king of Assyria. So the king of Assyria turned back and did not stay there in the land.
2KGS|15|21|Now the rest of the deeds of Menahem and all that he did, are they not written in the Book of the Chronicles of the Kings of Israel?
2KGS|15|22|And Menahem slept with his fathers, and Pekahiah his son reigned in his place.
2KGS|15|23|In the fiftieth year of Azariah king of Judah, Pekahiah the son of Menahem began to reign over Israel in Samaria, and he reigned two years.
2KGS|15|24|And he did what was evil in the sight of the LORD. He did not turn away from the sins of Jeroboam the son of Nebat, which he made Israel to sin.
2KGS|15|25|And Pekah the son of Remaliah, his captain, conspired against him with fifty men of the people of Gilead, and struck him down in Samaria, in the citadel of the king's house with Argob and Arieh; he put him to death and reigned in his place.
2KGS|15|26|Now the rest of the deeds of Pekahiah and all that he did, behold, they are written in the Book of the Chronicles of the Kings of Israel.
2KGS|15|27|In the fifty-second year of Azariah king of Judah, Pekah the son of Remaliah began to reign over Israel in Samaria, and he reigned twenty years.
2KGS|15|28|And he did what was evil in the sight of the LORD. He did not depart from the sins of Jeroboam the son of Nebat, which he made Israel to sin.
2KGS|15|29|In the days of Pekah king of Israel, Tiglath-pileser king of Assyria came and captured Ijon, Abel-beth-maacah, Janoah, Kedesh, Hazor, Gilead, and Galilee, all the land of Naphtali, and he carried the people captive to Assyria.
2KGS|15|30|Then Hoshea the son of Elah made a conspiracy against Pekah the son of Remaliah and struck him down and put him to death and reigned in his place, in the twentieth year of Jotham the son of Uzziah.
2KGS|15|31|Now the rest of the acts of Pekah and all that he did, behold, they are written in the Book of the Chronicles of the Kings of Israel.
2KGS|15|32|In the second year of Pekah the son of Remaliah, king of Israel, Jotham the son of Uzziah, king of Judah, began to reign.
2KGS|15|33|He was twenty-five years old when he began to reign, and he reigned sixteen years in Jerusalem. His mother's name was Jerusha the daughter of Zadok.
2KGS|15|34|And he did what was right in the eyes of the LORD, according to all that his father Uzziah had done.
2KGS|15|35|Nevertheless, the high places were not removed. The people still sacrificed and made offerings on the high places. He built the upper gate of the house of the LORD.
2KGS|15|36|Now the rest of the acts of Jotham and all that he did, are they not written in the Book of the Chronicles of the Kings of Judah?
2KGS|15|37|In those days the LORD began to send Rezin the king of Syria and Pekah the son of Remaliah against Judah.
2KGS|15|38|Jotham slept with his fathers and was buried with his fathers in the city of David his father, and Ahaz his son reigned in his place.
2KGS|16|1|In the seventeenth year of Pekah the son of Remaliah, Ahaz the son of Jotham, king of Judah, began to reign.
2KGS|16|2|Ahaz was twenty years old when he began to reign, and he reigned sixteen years in Jerusalem. And he did not do what was right in the eyes of the LORD his God, as his father David had done,
2KGS|16|3|but he walked in the way of the kings of Israel. He even burned his son as an offering, according to the despicable practices of the nations whom the LORD drove out before the people of Israel.
2KGS|16|4|And he sacrificed and made offerings on the high places and on the hills and under every green tree.
2KGS|16|5|Then Rezin king of Syria and Pekah the son of Remaliah, king of Israel, came up to wage war on Jerusalem, and they besieged Ahaz but could not conquer him.
2KGS|16|6|At that time Rezin the king of Syria recovered Elath for Syria and drove the men of Judah from Elath, and the Edomites came to Elath, where they dwell to this day.
2KGS|16|7|So Ahaz sent messengers to Tiglath-pileser king of Assyria, saying, "I am your servant and your son. Come up and rescue me from the hand of the king of Syria and from the hand of the king of Israel, who are attacking me."
2KGS|16|8|Ahaz also took the silver and gold that was found in the house of the LORD and in the treasures of the king's house and sent a present to the king of Assyria.
2KGS|16|9|And the king of Assyria listened to him. The king of Assyria marched up against Damascus and took it, carrying its people captive to Kir, and he killed Rezin.
2KGS|16|10|When King Ahaz went to Damascus to meet Tiglath-pileser king of Assyria, he saw the altar that was at Damascus. And King Ahaz sent to Uriah the priest a model of the altar, and its pattern, exact in all its details.
2KGS|16|11|And Uriah the priest built the altar; in accordance with all that King Ahaz had sent from Damascus, so Uriah the priest made it, before King Ahaz arrived from Damascus.
2KGS|16|12|And when the king came from Damascus, the king viewed the altar. Then the king drew near to the altar and went up on it
2KGS|16|13|and burned his burnt offering and his grain offering and poured his drink offering and threw the blood of his peace offerings on the altar.
2KGS|16|14|And the bronze altar that was before the LORD he removed from the front of the house, from the place between his altar and the house of the LORD, and put it on the north side of his altar.
2KGS|16|15|And King Ahaz commanded Uriah the priest, saying, "On the great altar burn the morning burnt offering and the evening grain offering and the king's burnt offering and his grain offering, with the burnt offering of all the people of the land, and their grain offering and their drink offering. And throw on it all the blood of the burnt offering and all the blood of the sacrifice, but the bronze altar shall be for me to inquire by."
2KGS|16|16|Uriah the priest did all this, as King Ahaz commanded.
2KGS|16|17|And King Ahaz cut off the frames of the stands and removed the basin from them, and he took down the sea from off the bronze oxen that were under it and put it on a stone pedestal.
2KGS|16|18|And the covered way for the Sabbath that had been built inside the house and the outer entrance for the king he caused to go around the house of the LORD, because of the king of Assyria.
2KGS|16|19|Now the rest of the acts of Ahaz that he did, are they not written in the Book of the Chronicles of the Kings of Judah?
2KGS|16|20|And Ahaz slept with his fathers and was buried with his fathers in the city of David, and Hezekiah his son reigned in his place.
2KGS|17|1|In the twelfth year of Ahaz king of Judah, Hoshea the son of Elah began to reign in Samaria over Israel, and he reigned nine years.
2KGS|17|2|And he did what was evil in the sight of the LORD, yet not as the kings of Israel who were before him.
2KGS|17|3|Against him came up Shalmaneser king of Assyria. And Hoshea became his vassal and paid him tribute.
2KGS|17|4|But the king of Assyria found treachery in Hoshea, for he had sent messengers to So, king of Egypt, and offered no tribute to the king of Assyria, as he had done year by year. Therefore the king of Assyria shut him up and bound him in prison.
2KGS|17|5|Then the king of Assyria invaded all the land and came to Samaria, and for three years he besieged it.
2KGS|17|6|In the ninth year of Hoshea, the king of Assyria captured Samaria, and he carried the Israelites away to Assyria and placed them in Halah, and on the Habor, the river of Gozan, and in the cities of the Medes.
2KGS|17|7|And this occurred because the people of Israel had sinned against the LORD their God, who had brought them up out of the land of Egypt from under the hand of Pharaoh king of Egypt, and had feared other gods
2KGS|17|8|and walked in the customs of the nations whom the LORD drove out before the people of Israel, and in the customs that the kings of Israel had practiced.
2KGS|17|9|And the people of Israel did secretly against the LORD their God things that were not right. They built for themselves high places in all their towns, from watchtower to fortified city.
2KGS|17|10|They set up for themselves pillars and Asherim on every high hill and under every green tree,
2KGS|17|11|and there they made offerings on all the high places, as the nations did whom the LORD carried away before them. And they did wicked things, provoking the LORD to anger,
2KGS|17|12|and they served idols, of which the LORD had said to them, "You shall not do this."
2KGS|17|13|Yet the LORD warned Israel and Judah by every prophet and every seer, saying, "Turn from your evil ways and keep my commandments and my statutes, in accordance with all the Law that I commanded your fathers, and that I sent to you by my servants the prophets."
2KGS|17|14|But they would not listen, but were stubborn, as their fathers had been, who did not believe in the LORD their God.
2KGS|17|15|They despised his statutes and his covenant that he made with their fathers and the warnings that he gave them. They went after false idols and became false, and they followed the nations that were around them, concerning whom the LORD had commanded them that they should not do like them.
2KGS|17|16|And they abandoned all the commandments of the LORD their God, and made for themselves metal images of two calves; and they made an Asherah and worshiped all the host of heaven and served Baal.
2KGS|17|17|And they burned their sons and their daughters as offerings and used divination and omens and sold themselves to do evil in the sight of the LORD, provoking him to anger.
2KGS|17|18|Therefore the LORD was very angry with Israel and removed them out of his sight. None was left but the tribe of Judah only.
2KGS|17|19|Judah also did not keep the commandments of the LORD their God, but walked in the customs that Israel had introduced.
2KGS|17|20|And the LORD rejected all the descendants of Israel and afflicted them and gave them into the hand of plunderers, until he had cast them out of his sight.
2KGS|17|21|When he had torn Israel from the house of David, they made Jeroboam the son of Nebat king. And Jeroboam drove Israel from following the LORD and made them commit great sin.
2KGS|17|22|The people of Israel walked in all the sins that Jeroboam did. They did not depart from them,
2KGS|17|23|until the LORD removed Israel out of his sight, as he had spoken by all his servants the prophets. So Israel was exiled from their own land to Assyria until this day.
2KGS|17|24|And the king of Assyria brought people from Babylon, Cuthah, Avva, Hamath, and Sepharvaim, and placed them in the cities of Samaria instead of the people of Israel. And they took possession of Samaria and lived in its cities.
2KGS|17|25|And at the beginning of their dwelling there, they did not fear the LORD. Therefore the LORD sent lions among them, which killed some of them.
2KGS|17|26|So the king of Assyria was told, "The nations that you have carried away and placed in the cities of Samaria do not know the law of the god of the land. Therefore he has sent lions among them, and behold, they are killing them, because they do not know the law of the god of the land."
2KGS|17|27|Then the king of Assyria commanded, "Send there one of the priests whom you carried away from there, and let him go and dwell there and teach them the law of the god of the land."
2KGS|17|28|So one of the priests whom they had carried away from Samaria came and lived in Bethel and taught them how they should fear the LORD.
2KGS|17|29|But every nation still made gods of its own and put them in the shrines of the high places that the Samaritans had made, every nation in the cities in which they lived.
2KGS|17|30|The men of Babylon made Succoth-benoth, the men of Cuth made Nergal, the men of Hamath made Ashima,
2KGS|17|31|and the Avvites made Nibhaz and Tartak; and the Sepharvites burned their children in the fire to Adrammelech and Anammelech, the gods of Sepharvaim.
2KGS|17|32|They also feared the LORD and appointed from among themselves all sorts of people as priests of the high places, who sacrificed for them in the shrines of the high places.
2KGS|17|33|So they feared the LORD but also served their own gods, after the manner of the nations from among whom they had been carried away.
2KGS|17|34|To this day they do according to the former manner. They do not fear the LORD, and they do not follow the statutes or the rules or the law or the commandment that the LORD commanded the children of Jacob, whom he named Israel.
2KGS|17|35|The LORD made a covenant with them and commanded them, "You shall not fear other gods or bow yourselves to them or serve them or sacrifice to them,
2KGS|17|36|but you shall fear the LORD, who brought you out of the land of Egypt with great power and with an outstretched arm. You shall bow yourselves to him, and to him you shall sacrifice.
2KGS|17|37|And the statutes and the rules and the law and the commandment that he wrote for you, you shall always be careful to do. You shall not fear other gods,
2KGS|17|38|and you shall not forget the covenant that I have made with you. You shall not fear other gods,
2KGS|17|39|but you shall fear the LORD your God, and he will deliver you out of the hand of all your enemies."
2KGS|17|40|However, they would not listen, but they did according to their former manner.
2KGS|17|41|So these nations feared the LORD and also served their carved images. Their children did likewise, and their children's children- as their fathers did, so they do to this day.
2KGS|18|1|In the third year of Hoshea son of Elah, king of Israel, Hezekiah the son of Ahaz, king of Judah, began to reign.
2KGS|18|2|He was twenty-five years old when he began to reign, and he reigned twenty-nine years in Jerusalem. His mother's name was Abi the daughter of Zechariah.
2KGS|18|3|And he did what was right in the eyes of the LORD, according to all that David his father had done.
2KGS|18|4|He removed the high places and broke the pillars and cut down the Asherah. And he broke in pieces the bronze serpent that Moses had made, for until those days the people of Israel had made offerings to it (it was called Nehushtan).
2KGS|18|5|He trusted in the LORD the God of Israel, so that there was none like him among all the kings of Judah after him, nor among those who were before him.
2KGS|18|6|For he held fast to the LORD. He did not depart from following him, but kept the commandments that the LORD commanded Moses.
2KGS|18|7|And the LORD was with him; wherever he went out, he prospered. He rebelled against the king of Assyria and would not serve him.
2KGS|18|8|He struck down the Philistines as far as Gaza and its territory, from watchtower to fortified city.
2KGS|18|9|In the fourth year of King Hezekiah, which was the seventh year of Hoshea son of Elah, king of Israel, Shalmaneser king of Assyria came up against Samaria and besieged it,
2KGS|18|10|and at the end of three years he took it. In the sixth year of Hezekiah, which was the ninth year of Hoshea king of Israel, Samaria was taken.
2KGS|18|11|The king of Assyria carried the Israelites away to Assyria and put them in Halah, and on the Habor, the river of Gozan, and in the cities of the Medes,
2KGS|18|12|because they did not obey the voice of the LORD their God but transgressed his covenant, even all that Moses the servant of the LORD commanded. They neither listened nor obeyed.
2KGS|18|13|In the fourteenth year of King Hezekiah, Sennacherib king of Assyria came up against all the fortified cities of Judah and took them.
2KGS|18|14|And Hezekiah king of Judah sent to the king of Assyria at Lachish, saying, "I have done wrong; withdraw from me. Whatever you impose on me I will bear." And the king of Assyria required of Hezekiah king of Judah three hundred talents of silver and thirty talents of gold.
2KGS|18|15|And Hezekiah gave him all the silver that was found in the house of the LORD and in the treasuries of the king's house.
2KGS|18|16|At that time Hezekiah stripped the gold from the doors of the temple of the LORD and from the doorposts that Hezekiah king of Judah had overlaid and gave it to the king of Assyria.
2KGS|18|17|And the king of Assyria sent the Tartan, the Rab-saris, and the Rabshakeh with a great army from Lachish to King Hezekiah at Jerusalem. And they went up and came to Jerusalem. When they arrived, they came and stood by the conduit of the upper pool, which is on the highway to the Washer's Field.
2KGS|18|18|And when they called for the king, there came out to them Eliakim the son of Hilkiah, who was over the household, and Shebnah the secretary, and Joah the son of Asaph, the recorder.
2KGS|18|19|And the Rabshakeh said to them, "Say to Hezekiah, 'Thus says the great king, the king of Assyria: On what do you rest this trust of yours?
2KGS|18|20|Do you think that mere words are strategy and power for war? In whom do you now trust, that you have rebelled against me?
2KGS|18|21|Behold, you are trusting now in Egypt, that broken reed of a staff, which will pierce the hand of any man who leans on it. Such is Pharaoh king of Egypt to all who trust in him.
2KGS|18|22|But if you say to me, "We trust in the LORD our God," is it not he whose high places and altars Hezekiah has removed, saying to Judah and to Jerusalem, "You shall worship before this altar in Jerusalem"?
2KGS|18|23|Come now, make a wager with my master the king of Assyria: I will give you two thousand horses, if you are able on your part to set riders on them.
2KGS|18|24|How then can you repulse a single captain among the least of my master's servants, when you trust in Egypt for chariots and for horsemen?
2KGS|18|25|Moreover, is it without the LORD that I have come up against this place to destroy it? The LORD said to me, Go up against this land, and destroy it.'"
2KGS|18|26|Then Eliakim the son of Hilkiah, and Shebnah, and Joah, said to the Rabshakeh, "Please speak to your servants in Aramaic, for we understand it. Do not speak to us in the language of Judah within the hearing of the people who are on the wall."
2KGS|18|27|But the Rabshakeh said to them, "Has my master sent me to speak these words to your master and to you, and not to the men sitting on the wall, who are doomed with you to eat their own dung and to drink their own urine?"
2KGS|18|28|Then the Rabshakeh stood and called out in a loud voice in the language of Judah: "Hear the word of the great king, the king of Assyria!
2KGS|18|29|Thus says the king: 'Do not let Hezekiah deceive you, for he will not be able to deliver you out of my hand.
2KGS|18|30|Do not let Hezekiah make you trust in the LORD by saying, The LORD will surely deliver us, and this city will not be given into the hand of the king of Assyria.'
2KGS|18|31|Do not listen to Hezekiah, for thus says the king of Assyria: 'Make your peace with me and come out to me. Then each one of you will eat of his own vine, and each one of his own fig tree, and each one of you will drink the water of his own cistern,
2KGS|18|32|until I come and take you away to a land like your own land, a land of grain and wine, a land of bread and vineyards, a land of olive trees and honey, that you may live, and not die. And do not listen to Hezekiah when he misleads you by saying, The LORD will deliver us.
2KGS|18|33|Has any of the gods of the nations ever delivered his land out of the hand of the king of Assyria?
2KGS|18|34|Where are the gods of Hamath and Arpad? Where are the gods of Sepharvaim, Hena, and Ivvah? Have they delivered Samaria out of my hand?
2KGS|18|35|Who among all the gods of the lands have delivered their lands out of my hand, that the LORD should deliver Jerusalem out of my hand?'"
2KGS|18|36|But the people were silent and answered him not a word, for the king's command was, "Do not answer him."
2KGS|18|37|Then Eliakim the son of Hilkiah, who was over the household, and Shebna the secretary, and Joah the son of Asaph, the recorder, came to Hezekiah with their clothes torn and told him the words of the Rabshakeh.
2KGS|19|1|As soon as King Hezekiah heard it, he tore his clothes and covered himself with sackcloth and went into the house of the LORD.
2KGS|19|2|And he sent Eliakim, who was over the household, and Shebna the secretary, and the senior priests, covered with sackcloth, to the prophet Isaiah the son of Amoz.
2KGS|19|3|They said to him, "Thus says Hezekiah, This day is a day of distress, of rebuke, and of disgrace; children have come to the point of birth, and there is no strength to bring them forth.
2KGS|19|4|It may be that the LORD your God heard all the words of the Rabshakeh, whom his master the king of Assyria has sent to mock the living God, and will rebuke the words that the LORD your God has heard; therefore lift up your prayer for the remnant that is left."
2KGS|19|5|When the servants of King Hezekiah came to Isaiah,
2KGS|19|6|Isaiah said to them, "Say to your master, 'Thus says the LORD: Do not be afraid because of the words that you have heard, with which the servants of the king of Assyria have reviled me.
2KGS|19|7|Behold, I will put a spirit in him, so that he shall hear a rumor and return to his own land, and I will make him fall by the sword in his own land.'"
2KGS|19|8|The Rabshakeh returned, and found the king of Assyria fighting against Libnah, for he heard that the king had left Lachish.
2KGS|19|9|Now the king heard concerning Tirhakah king of Cush, "Behold, he has set out to fight against you." So he sent messengers again to Hezekiah, saying,
2KGS|19|10|"Thus shall you speak to Hezekiah king of Judah: 'Do not let your God in whom you trust deceive you by promising that Jerusalem will not be given into the hand of the king of Assyria.
2KGS|19|11|Behold, you have heard what the kings of Assyria have done to all lands, devoting them to destruction. And shall you be delivered?
2KGS|19|12|Have the gods of the nations delivered them, the nations that my fathers destroyed, Gozan, Haran, Rezeph, and the people of Eden who were in Telassar?
2KGS|19|13|Where is the king of Hamath, the king of Arpad, the king of the city of Sepharvaim, the king of Hena, or the king of Ivvah?'"
2KGS|19|14|Hezekiah received the letter from the hand of the messengers and read it; and Hezekiah went up to the house of the LORD and spread it before the LORD.
2KGS|19|15|And Hezekiah prayed before the LORD and said: "O LORD the God of Israel, who is enthroned above the cherubim, you are the God, you alone, of all the kingdoms of the earth; you have made heaven and earth.
2KGS|19|16|Incline your ear, O LORD, and hear; open your eyes, O LORD, and see; and hear the words of Sennacherib, which he has sent to mock the living God.
2KGS|19|17|Truly, O LORD, the kings of Assyria have laid waste the nations and their lands
2KGS|19|18|and have cast their gods into the fire, for they were not gods, but the work of men's hands, wood and stone. Therefore they were destroyed.
2KGS|19|19|So now, O LORD our God, save us, please, from his hand, that all the kingdoms of the earth may know that you, O LORD, are God alone."
2KGS|19|20|Then Isaiah the son of Amoz sent to Hezekiah, saying, "Thus says the LORD, the God of Israel: Your prayer to me about Sennacherib king of Assyria I have heard.
2KGS|19|21|This is the word that the LORD has spoken concerning him: "She despises you, she scorns you- the virgin daughter of Zion; she wags her head behind you- the daughter of Jerusalem.
2KGS|19|22|"Whom have you mocked and reviled? Against whom have you raised your voice and lifted your eyes to the heights? Against the Holy One of Israel!
2KGS|19|23|By your messengers you have mocked the Lord, and you have said, 'With my many chariots I have gone up the heights of the mountains, to the far recesses of Lebanon; I felled its tallest cedars, its choicest cypresses; I entered its farthest lodging place, its most fruitful forest.
2KGS|19|24|I dug wells and drank foreign waters, and I dried up with the sole of my foot all the streams of Egypt.'
2KGS|19|25|"Have you not heard that I determined it long ago? I planned from days of old what now I bring to pass, that you should turn fortified cities into heaps of ruins,
2KGS|19|26|while their inhabitants, shorn of strength, are dismayed and confounded, and have become like plants of the field and like tender grass, like grass on the housetops, blighted before it is grown.
2KGS|19|27|"But I know your sitting down and your going out and coming in, and your raging against me.
2KGS|19|28|Because you have raged against me and your complacency has come into my ears, I will put my hook in your nose and my bit in your mouth, and I will turn you back on the way by which you came.
2KGS|19|29|"And this shall be the sign for you: this year eat what grows of itself, and in the second year what springs of the same. Then in the third year sow and reap and plant vineyards, and eat their fruit.
2KGS|19|30|And the surviving remnant of the house of Judah shall again take root downward and bear fruit upward.
2KGS|19|31|For out of Jerusalem shall go a remnant, and out of Mount Zion a band of survivors. The zeal of the LORD will do this.
2KGS|19|32|"Therefore thus says the LORD concerning the king of Assyria: He shall not come into this city or shoot an arrow there, or come before it with a shield or cast up a siege mound against it.
2KGS|19|33|By the way that he came, by the same he shall return, and he shall not come into this city, declares the LORD.
2KGS|19|34|For I will defend this city to save it, for my own sake and for the sake of my servant David."
2KGS|19|35|And that night the angel of the LORD went out and struck down 185,000 in the camp of the Assyrians. And when people arose early in the morning, behold, these were all dead bodies.
2KGS|19|36|Then Sennacherib king of Assyria departed and went home and lived at Nineveh.
2KGS|19|37|And as he was worshiping in the house of Nisroch his god, Adrammelech and Sharezer, his sons, struck him down with the sword and escaped into the land of Ararat. And Esarhaddon his son reigned in his place.
2KGS|20|1|In those days Hezekiah became sick and was at the point of death. And Isaiah the prophet the son of Amoz came to him and said to him, "Thus says the LORD, 'Set your house in order, for you shall die; you shall not recover.'"
2KGS|20|2|Then Hezekiah turned his face to the wall and prayed to the LORD, saying,
2KGS|20|3|"Now, O LORD, please remember how I have walked before you in faithfulness and with a whole heart, and have done what is good in your sight." And Hezekiah wept bitterly.
2KGS|20|4|And before Isaiah had gone out of the middle court, the word of the LORD came to him:
2KGS|20|5|"Turn back, and say to Hezekiah the leader of my people, Thus says the LORD, the God of David your father: I have heard your prayer; I have seen your tears. Behold, I will heal you. On the third day you shall go up to the house of the LORD,
2KGS|20|6|and I will add fifteen years to your life. I will deliver you and this city out of the hand of the king of Assyria, and I will defend this city for my own sake and for my servant David's sake."
2KGS|20|7|And Isaiah said, "Bring a cake of figs. And let them take and lay it on the boil, that he may recover."
2KGS|20|8|And Hezekiah said to Isaiah, "What shall be the sign that the LORD will heal me, and that I shall go up to the house of the LORD on the third day?"
2KGS|20|9|And Isaiah said, "This shall be the sign to you from the LORD, that the LORD will do the thing that he has promised: shall the shadow go forward ten steps, or go back ten steps?"
2KGS|20|10|And Hezekiah answered, "It is an easy thing for the shadow to lengthen ten steps. Rather let the shadow go back ten steps."
2KGS|20|11|And Isaiah the prophet called to the LORD, and he brought the shadow back ten steps, by which it had gone down on the steps of Ahaz.
2KGS|20|12|At that time Merodach-baladan the son of Baladan, king of Babylon, sent envoys with letters and a present to Hezekiah, for he heard that Hezekiah had been sick.
2KGS|20|13|And Hezekiah welcomed them, and he showed them all his treasure house, the silver, the gold, the spices, the precious oil, his armory, all that was found in his storehouses. There was nothing in his house or in all his realm that Hezekiah did not show them.
2KGS|20|14|Then Isaiah the prophet came to King Hezekiah, and said to him, "What did these men say? And from where did they come to you?" And Hezekiah said, "They have come from a far country, from Babylon."
2KGS|20|15|He said, "What have they seen in your house?" And Hezekiah answered, "They have seen all that is in my house; there is nothing in my storehouses that I did not show them."
2KGS|20|16|Then Isaiah said to Hezekiah, "Hear the word of the LORD:
2KGS|20|17|Behold, the days are coming, when all that is in your house, and that which your fathers have stored up till this day, shall be carried to Babylon. Nothing shall be left, says the LORD.
2KGS|20|18|And some of your own sons, who shall be born to you, shall be taken away, and they shall be eunuchs in the palace of the king of Babylon."
2KGS|20|19|Then said Hezekiah to Isaiah, "The word of the LORD that you have spoken is good." For he thought, "Why not, if there will be peace and security in my days?"
2KGS|20|20|The rest of the deeds of Hezekiah and all his might and how he made the pool and the conduit and brought water into the city, are they not written in the Book of the Chronicles of the Kings of Judah?
2KGS|20|21|And Hezekiah slept with his fathers, and Manasseh his son reigned in his place.
2KGS|21|1|Manasseh was twelve years old when he began to reign, and he reigned fifty-five years in Jerusalem. His mother's name was Hephzibah.
2KGS|21|2|And he did what was evil in the sight of the LORD, according to the despicable practices of the nations whom the LORD drove out before the people of Israel.
2KGS|21|3|For he rebuilt the high places that Hezekiah his father had destroyed, and he erected altars for Baal and made an Asherah, as Ahab king of Israel had done, and worshiped all the host of heaven and served them.
2KGS|21|4|And he built altars in the house of the LORD, of which the LORD had said, "In Jerusalem will I put my name."
2KGS|21|5|And he built altars for all the host of heaven in the two courts of the house of the LORD.
2KGS|21|6|And he burned his son as an offering and used fortune-telling and omens and dealt with mediums and with wizards. He did much evil in the sight of the LORD, provoking him to anger.
2KGS|21|7|And the carved image of Asherah that he had made he set in the house of which the LORD said to David and to Solomon his son, "In this house, and in Jerusalem, which I have chosen out of all the tribes of Israel, I will put my name forever.
2KGS|21|8|And I will not cause the feet of Israel to wander anymore out of the land that I gave to their fathers, if only they will be careful to do according to all that I have commanded them, and according to all the Law that my servant Moses commanded them."
2KGS|21|9|But they did not listen, and Manasseh led them astray to do more evil than the nations had done whom the LORD destroyed before the people of Israel.
2KGS|21|10|And the LORD said by his servants the prophets,
2KGS|21|11|"Because Manasseh king of Judah has committed these abominations and has done things more evil than all that the Amorites did, who were before him, and has made Judah also to sin with his idols,
2KGS|21|12|therefore thus says the LORD, the God of Israel: Behold, I am bringing upon Jerusalem and Judah such disaster that the ears of everyone who hears of it will tingle.
2KGS|21|13|And I will stretch over Jerusalem the measuring line of Samaria, and the plumb line of the house of Ahab, and I will wipe Jerusalem as one wipes a dish, wiping it and turning it upside down.
2KGS|21|14|And I will forsake the remnant of my heritage and give them into the hand of their enemies, and they shall become a prey and a spoil to all their enemies,
2KGS|21|15|because they have done what is evil in my sight and have provoked me to anger, since the day their fathers came out of Egypt, even to this day."
2KGS|21|16|Moreover, Manasseh shed very much innocent blood, till he had filled Jerusalem from one end to another, besides the sin that he made Judah to sin so that they did what was evil in the sight of the LORD.
2KGS|21|17|Now the rest of the acts of Manasseh and all that he did, and the sin that he committed, are they not written in the Book of the Chronicles of the Kings of Judah?
2KGS|21|18|And Manasseh slept with his fathers and was buried in the garden of his house, in the garden of Uzza, and Amon his son reigned in his place.
2KGS|21|19|Amon was twenty-two years old when he began to reign, and he reigned two years in Jerusalem. His mother's name was Meshullemeth the daughter of Haruz of Jotbah.
2KGS|21|20|And he did what was evil in the sight of the LORD, as Manasseh his father had done.
2KGS|21|21|He walked in all the way in which his father walked and served the idols that his father served and worshiped them.
2KGS|21|22|He abandoned the LORD, the God of his fathers, and did not walk in the way of the LORD.
2KGS|21|23|And the servants of Amon conspired against him and put the king to death in his house.
2KGS|21|24|But the people of the land struck down all those who had conspired against King Amon, and the people of the land made Josiah his son king in his place.
2KGS|21|25|Now the rest of the acts of Amon that he did, are they not written in the Book of the Chronicles of the Kings of Judah?
2KGS|21|26|And he was buried in his tomb in the garden of Uzza, and Josiah his son reigned in his place.
2KGS|22|1|Josiah was eight years old when he began to reign, and he reigned thirty-one years in Jerusalem. His mother's name was Jedidah the daughter of Adaiah of Bozkath.
2KGS|22|2|And he did what was right in the eyes of the LORD and walked in all the way of David his father, and he did not turn aside to the right or to the left.
2KGS|22|3|In the eighteenth year of King Josiah, the king sent Shaphan the son of Azaliah, son of Meshullam, the secretary, to the house of the LORD, saying,
2KGS|22|4|"Go up to Hilkiah the high priest, that he may count the money that has been brought into the house of the LORD, which the keepers of the threshold have collected from the people.
2KGS|22|5|And let it be given into the hand of the workmen who have the oversight of the house of the LORD, and let them give it to the workmen who are at the house of the LORD, repairing the house (
2KGS|22|6|that is, to the carpenters, and to the builders, and to the masons), and let them use it for buying timber and quarried stone to repair the house.
2KGS|22|7|But no accounting shall be asked from them for the money that is delivered into their hand, for they deal honestly."
2KGS|22|8|And Hilkiah the high priest said to Shaphan the secretary, "I have found the Book of the Law in the house of the LORD." And Hilkiah gave the book to Shaphan, and he read it.
2KGS|22|9|And Shaphan the secretary came to the king, and reported to the king, "Your servants have emptied out the money that was found in the house and have delivered it into the hand of the workmen who have the oversight of the house of the LORD."
2KGS|22|10|Then Shaphan the secretary told the king, "Hilkiah the priest has given me a book." And Shaphan read it before the king.
2KGS|22|11|When the king heard the words of the Book of the Law, he tore his clothes.
2KGS|22|12|And the king commanded Hilkiah the priest, and Ahikam the son of Shaphan, and Achbor the son of Micaiah, and Shaphan the secretary, and Asaiah the king's servant, saying,
2KGS|22|13|"Go, inquire of the LORD for me, and for the people, and for all Judah, concerning the words of this book that has been found. For great is the wrath of the LORD that is kindled against us, because our fathers have not obeyed the words of this book, to do according to all that is written concerning us."
2KGS|22|14|So Hilkiah the priest, and Ahikam, and Achbor, and Shaphan, and Asaiah went to Huldah the prophetess, the wife of Shallum the son of Tikvah, son of Harhas, keeper of the wardrobe (now she lived in Jerusalem in the Second Quarter), and they talked with her.
2KGS|22|15|And she said to them, "Thus says the LORD, the God of Israel: 'Tell the man who sent you to me,
2KGS|22|16|Thus says the LORD, behold, I will bring disaster upon this place and upon its inhabitants, all the words of the book that the king of Judah has read.
2KGS|22|17|Because they have forsaken me and have made offerings to other gods, that they might provoke me to anger with all the work of their hands, therefore my wrath will be kindled against this place, and it will not be quenched.
2KGS|22|18|But to the king of Judah, who sent you to inquire of the LORD, thus shall you say to him, Thus says the LORD, the God of Israel: Regarding the words that you have heard,
2KGS|22|19|because your heart was penitent, and you humbled yourself before the LORD, when you heard how I spoke against this place and against its inhabitants, that they should become a desolation and a curse, and you have torn your clothes and wept before me, I also have heard you, declares the LORD.
2KGS|22|20|Therefore, behold, I will gather you to your fathers, and you shall be gathered to your grave in peace, and your eyes shall not see all the disaster that I will bring upon this place.'"And they brought back word to the king.
2KGS|23|1|Then the king sent, and all the elders of Judah and Jerusalem were gathered to him.
2KGS|23|2|And the king went up to the house of the LORD, and with him all the men of Judah and all the inhabitants of Jerusalem and the priests and the prophets, all the people, both small and great. And he read in their hearing all the words of the Book of the Covenant that had been found in the house of the LORD.
2KGS|23|3|And the king stood by the pillar and made a covenant before the LORD, to walk after the LORD and to keep his commandments and his testimonies and his statutes with all his heart and all his soul, to perform the words of this covenant that were written in this book. And all the people joined in the covenant.
2KGS|23|4|And the king commanded Hilkiah the high priest and the priests of the second order and the keepers of the threshold to bring out of the temple of the LORD all the vessels made for Baal, for Asherah, and for all the host of heaven. He burned them outside Jerusalem in the fields of the Kidron and carried their ashes to Bethel.
2KGS|23|5|And he deposed the priests whom the kings of Judah had ordained to make offerings in the high places at the cities of Judah and around Jerusalem; those also who burned incense to Baal, to the sun and the moon and the constellations and all the host of the heavens.
2KGS|23|6|And he brought out the Asherah from the house of the LORD, outside Jerusalem, to the brook Kidron, and burned it at the brook Kidron and beat it to dust and cast the dust of it upon the graves of the common people.
2KGS|23|7|And he broke down the houses of the male cult prostitutes who were in the house of the LORD, where the women wove hangings for the Asherah.
2KGS|23|8|And he brought all the priests out of the cities of Judah, and defiled the high places where the priests had made offerings, from Geba to Beersheba. And he broke down the high places of the gates that were at the entrance of the gate of Joshua the governor of the city, which were on one's left at the gate of the city.
2KGS|23|9|However, the priests of the high places did not come up to the altar of the LORD in Jerusalem, but they ate unleavened bread among their brothers.
2KGS|23|10|And he defiled Topheth, which is in the Valley of the Son of Hinnom, that no one might burn his son or his daughter as an offering to Molech.
2KGS|23|11|And he removed the horses that the kings of Judah had dedicated to the sun, at the entrance to the house of the LORD, by the chamber of Nathan-melech the chamberlain, which was in the precincts. And he burned the chariots of the sun with fire.
2KGS|23|12|And the altars on the roof of the upper chamber of Ahaz, which the kings of Judah had made, and the altars that Manasseh had made in the two courts of the house of the LORD, he pulled down and broke in pieces and cast the dust of them into the brook Kidron.
2KGS|23|13|And the king defiled the high places that were east of Jerusalem, to the south of the mount of corruption, which Solomon the king of Israel had built for Ashtoreth the abomination of the Sidonians, and for Chemosh the abomination of Moab, and for Milcom the abomination of the Ammonites.
2KGS|23|14|And he broke in pieces the pillars and cut down the Asherim and filled their places with the bones of men.
2KGS|23|15|Moreover, the altar at Bethel, the high place erected by Jeroboam the son of Nebat, who made Israel to sin, that altar with the high place he pulled down and burned, reducing it to dust. He also burned the Asherah.
2KGS|23|16|And as Josiah turned, he saw the tombs there on the mount. And he sent and took the bones out of the tombs and burned them on the altar and defiled it, according to the word of the LORD that the man of God proclaimed, who had predicted these things.
2KGS|23|17|Then he said, "What is that monument that I see?" And the men of the city told him, "It is the tomb of the man of God who came from Judah and predicted these things that you have done against the altar at Bethel."
2KGS|23|18|And he said, "Let him be; let no man move his bones." So they let his bones alone, with the bones of the prophet who came out of Samaria.
2KGS|23|19|And Josiah removed all the shrines also of the high places that were in the cities of Samaria, which kings of Israel had made, provoking the LORD to anger. He did to them according to all that he had done at Bethel.
2KGS|23|20|And he sacrificed all the priests of the high places who were there, on the altars, and burned human bones on them. Then he returned to Jerusalem.
2KGS|23|21|And the king commanded all the people, "Keep the Passover to the LORD your God, as it is written in this Book of the Covenant."
2KGS|23|22|For no such Passover had been kept since the days of the judges who judged Israel, or during all the days of the kings of Israel or of the kings of Judah.
2KGS|23|23|But in the eighteenth year of King Josiah this Passover was kept to the LORD in Jerusalem.
2KGS|23|24|Moreover, Josiah put away the mediums and the necromancers and the household gods and the idols and all the abominations that were seen in the land of Judah and in Jerusalem, that he might establish the words of the law that were written in the book that Hilkiah the priest found in the house of the LORD.
2KGS|23|25|Before him there was no king like him, who turned to the LORD with all his heart and with all his soul and with all his might, according to all the Law of Moses, nor did any like him arise after him.
2KGS|23|26|Still the LORD did not turn from the burning of his great wrath, by which his anger was kindled against Judah, because of all the provocations with which Manasseh had provoked him.
2KGS|23|27|And the LORD said, "I will remove Judah also out of my sight, as I have removed Israel, and I will cast off this city that I have chosen, Jerusalem, and the house of which I said, My name shall be there."
2KGS|23|28|Now the rest of the acts of Josiah and all that he did, are they not written in the Book of the Chronicles of the Kings of Judah?
2KGS|23|29|In his days Pharaoh Neco king of Egypt went up to the king of Assyria to the river Euphrates. King Josiah went to meet him, and Pharaoh Neco killed him at Megiddo, as soon as he saw him.
2KGS|23|30|And his servants carried him dead in a chariot from Megiddo and brought him to Jerusalem and buried him in his own tomb. And the people of the land took Jehoahaz the son of Josiah, and anointed him, and made him king in his father's place.
2KGS|23|31|Jehoahaz was twenty-three years old when he began to reign, and he reigned three months in Jerusalem. His mother's name was Hamutal the daughter of Jeremiah of Libnah.
2KGS|23|32|And he did what was evil in the sight of the LORD, according to all that his fathers had done.
2KGS|23|33|And Pharaoh Neco put him in bonds at Riblah in the land of Hamath, that he might not reign in Jerusalem, and laid on the land a tribute of a hundred talents of silver and a talent of gold.
2KGS|23|34|And Pharaoh Neco made Eliakim the son of Josiah king in the place of Josiah his father, and changed his name to Jehoiakim. But he took Jehoahaz away, and he came to Egypt and died there.
2KGS|23|35|And Jehoiakim gave the silver and the gold to Pharaoh, but he taxed the land to give the money according to the command of Pharaoh. He exacted the silver and the gold of the people of the land, from everyone according to his assessment, to give it to Pharaoh Neco.
2KGS|23|36|Jehoiakim was twenty-five years old when he began to reign, and he reigned eleven years in Jerusalem. His mother's name was Zebidah the daughter of Pedaiah of Rumah.
2KGS|23|37|And he did what was evil in the sight of the LORD, according to all that his fathers had done.
2KGS|24|1|In his days, Nebuchadnezzar king of Babylon came up, and Jehoiakim became his servant three years. Then he turned and rebelled against him.
2KGS|24|2|And the LORD sent against him bands of the Chaldeans and bands of the Syrians and bands of the Moabites and bands of the Ammonites, and sent them against Judah to destroy it, according to the word of the LORD that he spoke by his servants the prophets.
2KGS|24|3|Surely this came upon Judah at the command of the LORD, to remove them out of his sight, for the sins of Manasseh, according to all that he had done,
2KGS|24|4|and also for the innocent blood that he had shed. For he filled Jerusalem with innocent blood, and the LORD would not pardon.
2KGS|24|5|Now the rest of the deeds of Jehoiakim and all that he did, are they not written in the Book of the Chronicles of the Kings of Judah?
2KGS|24|6|So Jehoiakim slept with his fathers, and Jehoiachin his son reigned in his place.
2KGS|24|7|And the king of Egypt did not come again out of his land, for the king of Babylon had taken all that belonged to the king of Egypt from the Brook of Egypt to the river Euphrates.
2KGS|24|8|Jehoiachin was eighteen years old when he became king, and he reigned three months in Jerusalem. His mother's name was Nehushta the daughter of Elnathan of Jerusalem.
2KGS|24|9|And he did what was evil in the sight of the LORD, according to all that his father had done.
2KGS|24|10|At that time the servants of Nebuchadnezzar king of Babylon came up to Jerusalem, and the city was besieged.
2KGS|24|11|And Nebuchadnezzar king of Babylon came to the city while his servants were besieging it,
2KGS|24|12|and Jehoiachin the king of Judah gave himself up to the king of Babylon, himself and his mother and his servants and his officials and his palace officials. The king of Babylon took him prisoner in the eighth year of his reign
2KGS|24|13|and carried off all the treasures of the house of the LORD and the treasures of the king's house, and cut in pieces all the vessels of gold in the temple of the LORD, which Solomon king of Israel had made, as the LORD had foretold.
2KGS|24|14|He carried away all Jerusalem and all the officials and all the mighty men of valor, 10,000 captives, and all the craftsmen and the smiths. None remained, except the poorest people of the land.
2KGS|24|15|And he carried away Jehoiachin to Babylon. The king's mother, the king's wives, his officials, and the chief men of the land he took into captivity from Jerusalem to Babylon.
2KGS|24|16|And the king of Babylon brought captive to Babylon all the men of valor, 7,000, and the craftsmen and the metal workers, 1,000, all of them strong and fit for war.
2KGS|24|17|And the king of Babylon made Mattaniah, Jehoiachin's uncle, king in his place, and changed his name to Zedekiah.
2KGS|24|18|Zedekiah was twenty-one years old when he became king, and he reigned eleven years in Jerusalem. His mother's name was Hamutal the daughter of Jeremiah of Libnah.
2KGS|24|19|And he did what was evil in the sight of the LORD, according to all that Jehoiakim had done.
2KGS|24|20|For because of the anger of the LORD it came to the point in Jerusalem and Judah that he cast them out from his presence. And Zedekiah rebelled against the king of Babylon.
2KGS|25|1|And in the ninth year of his reign, in the tenth month, on the tenth day of the month, Nebuchadnezzar king of Babylon came with all his army against Jerusalem and laid siege to it. And they built siegeworks all around it.
2KGS|25|2|So the city was besieged till the eleventh year of King Zedekiah.
2KGS|25|3|On the ninth day of the fourth month the famine was so severe in the city that there was no food for the people of the land.
2KGS|25|4|Then a breach was made in the city, and all the men of war fled by night by the way of the gate between the two walls, by the king's garden, though the Chaldeans were around the city. And they went in the direction of the Arabah.
2KGS|25|5|But the army of the Chaldeans pursued the king and overtook him in the plains of Jericho, and all his army was scattered from him.
2KGS|25|6|Then they captured the king and brought him up to the king of Babylon at Riblah, and they passed sentence on him.
2KGS|25|7|They slaughtered the sons of Zedekiah before his eyes, and put out the eyes of Zedekiah and bound him in chains and took him to Babylon.
2KGS|25|8|In the fifth month, on the seventh day of the month- that was the nineteenth year of King Nebuchadnezzar, king of Babylon- Nebuzaradan, the captain of the bodyguard, a servant of the king of Babylon, came to Jerusalem.
2KGS|25|9|And he burned the house of the LORD and the king's house and all the houses of Jerusalem; every great house he burned down.
2KGS|25|10|And all the army of the Chaldeans, who were with the captain of the guard, broke down the walls around Jerusalem.
2KGS|25|11|And the rest of the people who were left in the city and the deserters who had deserted to the king of Babylon, together with the rest of the multitude, Nebuzaradan the captain of the guard carried into exile.
2KGS|25|12|But the captain of the guard left some of the poorest of the land to be vinedressers and plowmen.
2KGS|25|13|And the pillars of bronze that were in the house of the LORD, and the stands and the bronze sea that were in the house of the LORD, the Chaldeans broke in pieces and carried the bronze to Babylon.
2KGS|25|14|And they took away the pots and the shovels and the snuffers and the dishes for incense and all the vessels of bronze used in the temple service,
2KGS|25|15|the fire pans also and the bowls. What was of gold the captain of the guard took away as gold, and what was of silver, as silver.
2KGS|25|16|As for the two pillars, the one sea, and the stands that Solomon had made for the house of the LORD, the bronze of all these vessels was beyond weight.
2KGS|25|17|The height of the one pillar was eighteen cubits, and on it was a capital of bronze. The height of the capital was three cubits. A latticework and pomegranates, all of bronze, were all around the capital. And the second pillar had the same, with the latticework.
2KGS|25|18|And the captain of the guard took Seraiah the chief priest and Zephaniah the second priest and the three keepers of the threshold,
2KGS|25|19|and from the city he took an officer who had been in command of the men of war, and five men of the king's council who were found in the city, and the secretary of the commander of the army who mustered the people of the land, and sixty men of the people of the land who were found in the city.
2KGS|25|20|And Nebuzaradan the captain of the guard took them and brought them to the king of Babylon at Riblah.
2KGS|25|21|And the king of Babylon struck them down and put them to death at Riblah in the land of Hamath. So Judah was taken into exile out of its land.
2KGS|25|22|And over the people who remained in the land of Judah, whom Nebuchadnezzar king of Babylon had left, he appointed Gedaliah the son of Ahikam, son of Shaphan, governor.
2KGS|25|23|Now when all the captains and their men heard that the king of Babylon had appointed Gedaliah governor, they came with their men to Gedaliah at Mizpah, namely, Ishmael the son of Nethaniah, and Johanan the son of Kareah, and Seraiah the son of Tanhumeth the Netophathite, and Jaazaniah the son of the Maacathite.
2KGS|25|24|And Gedaliah swore to them and their men, saying, "Do not be afraid because of the Chaldean officials. Live in the land and serve the king of Babylon, and it shall be well with you."
2KGS|25|25|But in the seventh month, Ishmael the son of Nethaniah, son of Elishama, of the royal family, came with ten men and struck down Gedaliah and put him to death along with the Jews and the Chaldeans who were with him at Mizpah.
2KGS|25|26|Then all the people, both small and great, and the captains of the forces arose and went to Egypt, for they were afraid of the Chaldeans.
2KGS|25|27|And in the thirty-seventh year of the exile of Jehoiachin king of Judah, in the twelfth month, on the twenty-seventh day of the month, Evil-merodach king of Babylon, in the year that he began to reign, graciously freed Jehoiachin king of Judah from prison.
2KGS|25|28|And he spoke kindly to him and gave him a seat above the seats of the kings who were with him in Babylon.
2KGS|25|29|So Jehoiachin put off his prison garments. And every day of his life he dined regularly at the king's table,
2KGS|25|30|and for his allowance, a regular allowance was given him by the king, according to his daily needs, as long as he lived.
