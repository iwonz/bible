JER|1|1|The words of Jeremiah the son of Hilkiah, of the priests that were in Anathoth in the land of Benjamin:
JER|1|2|To whom the word of the LORD came in the days of Josiah the son of Amon king of Judah, in the thirteenth year of his reign.
JER|1|3|It came also in the days of Jehoiakim the son of Josiah king of Judah, unto the end of the eleventh year of Zedekiah the son of Josiah king of Judah, unto the carrying away of Jerusalem captive in the fifth month.
JER|1|4|Then the word of the LORD came unto me, saying,
JER|1|5|Before I formed thee in the belly I knew thee; and before thou camest forth out of the womb I sanctified thee, and I ordained thee a prophet unto the nations.
JER|1|6|Then said I, Ah, Lord GOD! behold, I cannot speak: for I am a child.
JER|1|7|But the LORD said unto me, Say not, I am a child: for thou shalt go to all that I shall send thee, and whatsoever I command thee thou shalt speak.
JER|1|8|Be not afraid of their faces: for I am with thee to deliver thee, saith the LORD.
JER|1|9|Then the LORD put forth his hand, and touched my mouth. And the LORD said unto me, Behold, I have put my words in thy mouth.
JER|1|10|See, I have this day set thee over the nations and over the kingdoms, to root out, and to pull down, and to destroy, and to throw down, to build, and to plant.
JER|1|11|Moreover the word of the LORD came unto me, saying, Jeremiah, what seest thou? And I said, I see a rod of an almond tree.
JER|1|12|Then said the LORD unto me, Thou hast well seen: for I will hasten my word to perform it.
JER|1|13|And the word of the LORD came unto me the second time, saying, What seest thou? And I said, I see a seething pot; and the face thereof is toward the north.
JER|1|14|Then the LORD said unto me, Out of the north an evil shall break forth upon all the inhabitants of the land.
JER|1|15|For, lo, I will call all the families of the kingdoms of the north, saith the LORD; and they shall come, and they shall set every one his throne at the entering of the gates of Jerusalem, and against all the walls thereof round about, and against all the cities of Judah.
JER|1|16|And I will utter my judgments against them touching all their wickedness, who have forsaken me, and have burned incense unto other gods, and worshipped the works of their own hands.
JER|1|17|Thou therefore gird up thy loins, and arise, and speak unto them all that I command thee: be not dismayed at their faces, lest I confound thee before them.
JER|1|18|For, behold, I have made thee this day a defenced city, and an iron pillar, and brasen walls against the whole land, against the kings of Judah, against the princes thereof, against the priests thereof, and against the people of the land.
JER|1|19|And they shall fight against thee; but they shall not prevail against thee; for I am with thee, saith the LORD, to deliver thee.
JER|2|1|Moreover the word of the LORD came to me, saying,
JER|2|2|Go and cry in the ears of Jerusalem, saying, Thus saith the LORD; I remember thee, the kindness of thy youth, the love of thine espousals, when thou wentest after me in the wilderness, in a land that was not sown.
JER|2|3|Israel was holiness unto the LORD, and the firstfruits of his increase: all that devour him shall offend; evil shall come upon them, saith the LORD.
JER|2|4|Hear ye the word of the LORD, O house of Jacob, and all the families of the house of Israel:
JER|2|5|Thus saith the LORD, What iniquity have your fathers found in me, that they are gone far from me, and have walked after vanity, and are become vain?
JER|2|6|Neither said they, Where is the LORD that brought us up out of the land of Egypt, that led us through the wilderness, through a land of deserts and of pits, through a land of drought, and of the shadow of death, through a land that no man passed through, and where no man dwelt?
JER|2|7|And I brought you into a plentiful country, to eat the fruit thereof and the goodness thereof; but when ye entered, ye defiled my land, and made mine heritage an abomination.
JER|2|8|The priests said not, Where is the LORD? and they that handle the law knew me not: the pastors also transgressed against me, and the prophets prophesied by Baal, and walked after things that do not profit.
JER|2|9|Wherefore I will yet plead with you, saith the LORD, and with your children's children will I plead.
JER|2|10|For pass over the isles of Chittim, and see; and send unto Kedar, and consider diligently, and see if there be such a thing.
JER|2|11|Hath a nation changed their gods, which are yet no gods? but my people have changed their glory for that which doth not profit.
JER|2|12|Be astonished, O ye heavens, at this, and be horribly afraid, be ye very desolate, saith the LORD.
JER|2|13|For my people have committed two evils; they have forsaken me the fountain of living waters, and hewed them out cisterns, broken cisterns, that can hold no water.
JER|2|14|Is Israel a servant? is he a homeborn slave? why is he spoiled?
JER|2|15|The young lions roared upon him, and yelled, and they made his land waste: his cities are burned without inhabitant.
JER|2|16|Also the children of Noph and Tahapanes have broken the crown of thy head.
JER|2|17|Hast thou not procured this unto thyself, in that thou hast forsaken the LORD thy God, when he led thee by the way?
JER|2|18|And now what hast thou to do in the way of Egypt, to drink the waters of Sihor? or what hast thou to do in the way of Assyria, to drink the waters of the river?
JER|2|19|Thine own wickedness shall correct thee, and thy backslidings shall reprove thee: know therefore and see that it is an evil thing and bitter, that thou hast forsaken the LORD thy God, and that my fear is not in thee, saith the Lord GOD of hosts.
JER|2|20|For of old time I have broken thy yoke, and burst thy bands; and thou saidst, I will not transgress; when upon every high hill and under every green tree thou wanderest, playing the harlot.
JER|2|21|Yet I had planted thee a noble vine, wholly a right seed: how then art thou turned into the degenerate plant of a strange vine unto me?
JER|2|22|For though thou wash thee with nitre, and take thee much soap, yet thine iniquity is marked before me, saith the Lord GOD.
JER|2|23|How canst thou say, I am not polluted, I have not gone after Baalim? see thy way in the valley, know what thou hast done: thou art a swift dromedary traversing her ways;
JER|2|24|A wild ass used to the wilderness, that snuffeth up the wind at her pleasure; in her occasion who can turn her away? all they that seek her will not weary themselves; in her month they shall find her.
JER|2|25|Withhold thy foot from being unshod, and thy throat from thirst: but thou saidst, There is no hope: no; for I have loved strangers, and after them will I go.
JER|2|26|As the thief is ashamed when he is found, so is the house of Israel ashamed; they, their kings, their princes, and their priests, and their prophets.
JER|2|27|Saying to a stock, Thou art my father; and to a stone, Thou hast brought me forth: for they have turned their back unto me, and not their face: but in the time of their trouble they will say, Arise, and save us.
JER|2|28|But where are thy gods that thou hast made thee? let them arise, if they can save thee in the time of thy trouble: for according to the number of thy cities are thy gods, O Judah.
JER|2|29|Wherefore will ye plead with me? ye all have transgressed against me, saith the LORD.
JER|2|30|In vain have I smitten your children; they received no correction: your own sword hath devoured your prophets, like a destroying lion.
JER|2|31|O generation, see ye the word of the LORD. Have I been a wilderness unto Israel? a land of darkness? wherefore say my people, We are lords; we will come no more unto thee?
JER|2|32|Can a maid forget her ornaments, or a bride her attire? yet my people have forgotten me days without number.
JER|2|33|Why trimmest thou thy way to seek love? therefore hast thou also taught the wicked ones thy ways.
JER|2|34|Also in thy skirts is found the blood of the souls of the poor innocents: I have not found it by secret search, but upon all these.
JER|2|35|Yet thou sayest, Because I am innocent, surely his anger shall turn from me. Behold, I will plead with thee, because thou sayest, I have not sinned.
JER|2|36|Why gaddest thou about so much to change thy way? thou also shalt be ashamed of Egypt, as thou wast ashamed of Assyria.
JER|2|37|Yea, thou shalt go forth from him, and thine hands upon thine head: for the LORD hath rejected thy confidences, and thou shalt not prosper in them.
JER|3|1|They say, If a man put away his wife, and she go from him, and become another man's, shall he return unto her again? shall not that land be greatly polluted? but thou hast played the harlot with many lovers; yet return again to me, saith the LORD.
JER|3|2|Lift up thine eyes unto the high places, and see where thou hast not been lien with. In the ways hast thou sat for them, as the Arabian in the wilderness; and thou hast polluted the land with thy whoredoms and with thy wickedness.
JER|3|3|Therefore the showers have been withholden, and there hath been no latter rain; and thou hadst a whore's forehead, thou refusedst to be ashamed.
JER|3|4|Wilt thou not from this time cry unto me, My father, thou art the guide of my youth?
JER|3|5|Will he reserve his anger for ever? will he keep it to the end? Behold, thou hast spoken and done evil things as thou couldest.
JER|3|6|The LORD said also unto me in the days of Josiah the king, Hast thou seen that which backsliding Israel hath done? she is gone up upon every high mountain and under every green tree, and there hath played the harlot.
JER|3|7|And I said after she had done all these things, Turn thou unto me. But she returned not. And her treacherous sister Judah saw it.
JER|3|8|And I saw, when for all the causes whereby backsliding Israel committed adultery I had put her away, and given her a bill of divorce; yet her treacherous sister Judah feared not, but went and played the harlot also.
JER|3|9|And it came to pass through the lightness of her whoredom, that she defiled the land, and committed adultery with stones and with stocks.
JER|3|10|And yet for all this her treacherous sister Judah hath not turned unto me with her whole heart, but feignedly, saith the LORD.
JER|3|11|And the LORD said unto me, The backsliding Israel hath justified herself more than treacherous Judah.
JER|3|12|Go and proclaim these words toward the north, and say, Return, thou backsliding Israel, saith the LORD; and I will not cause mine anger to fall upon you: for I am merciful, saith the LORD, and I will not keep anger for ever.
JER|3|13|Only acknowledge thine iniquity, that thou hast transgressed against the LORD thy God, and hast scattered thy ways to the strangers under every green tree, and ye have not obeyed my voice, saith the LORD.
JER|3|14|Turn, O backsliding children, saith the LORD; for I am married unto you: and I will take you one of a city, and two of a family, and I will bring you to Zion:
JER|3|15|And I will give you pastors according to mine heart, which shall feed you with knowledge and understanding.
JER|3|16|And it shall come to pass, when ye be multiplied and increased in the land, in those days, saith the LORD, they shall say no more, The ark of the covenant of the LORD: neither shall it come to mind: neither shall they remember it; neither shall they visit it; neither shall that be done any more.
JER|3|17|At that time they shall call Jerusalem the throne of the LORD; and all the nations shall be gathered unto it, to the name of the LORD, to Jerusalem: neither shall they walk any more after the imagination of their evil heart.
JER|3|18|In those days the house of Judah shall walk with the house of Israel, and they shall come together out of the land of the north to the land that I have given for an inheritance unto your fathers.
JER|3|19|But I said, How shall I put thee among the children, and give thee a pleasant land, a goodly heritage of the hosts of nations? and I said, Thou shalt call me, My father; and shalt not turn away from me.
JER|3|20|Surely as a wife treacherously departeth from her husband, so have ye dealt treacherously with me, O house of Israel, saith the LORD.
JER|3|21|A voice was heard upon the high places, weeping and supplications of the children of Israel: for they have perverted their way, and they have forgotten the LORD their God.
JER|3|22|Return, ye backsliding children, and I will heal your backslidings. Behold, we come unto thee; for thou art the LORD our God.
JER|3|23|Truly in vain is salvation hoped for from the hills, and from the multitude of mountains: truly in the LORD our God is the salvation of Israel.
JER|3|24|For shame hath devoured the labour of our fathers from our youth; their flocks and their herds, their sons and their daughters.
JER|3|25|We lie down in our shame, and our confusion covereth us: for we have sinned against the LORD our God, we and our fathers, from our youth even unto this day, and have not obeyed the voice of the LORD our God.
JER|4|1|If thou wilt return, O Israel, saith the LORD, return unto me: and if thou wilt put away thine abominations out of my sight, then shalt thou not remove.
JER|4|2|And thou shalt swear, The LORD liveth, in truth, in judgment, and in righteousness; and the nations shall bless themselves in him, and in him shall they glory.
JER|4|3|For thus saith the LORD to the men of Judah and Jerusalem, Break up your fallow ground, and sow not among thorns.
JER|4|4|Circumcise yourselves to the LORD, and take away the foreskins of your heart, ye men of Judah and inhabitants of Jerusalem: lest my fury come forth like fire, and burn that none can quench it, because of the evil of your doings.
JER|4|5|Declare ye in Judah, and publish in Jerusalem; and say, Blow ye the trumpet in the land: cry, gather together, and say, Assemble yourselves, and let us go into the defenced cities.
JER|4|6|Set up the standard toward Zion: retire, stay not: for I will bring evil from the north, and a great destruction.
JER|4|7|The lion is come up from his thicket, and the destroyer of the Gentiles is on his way; he is gone forth from his place to make thy land desolate; and thy cities shall be laid waste, without an inhabitant.
JER|4|8|For this gird you with sackcloth, lament and howl: for the fierce anger of the LORD is not turned back from us.
JER|4|9|And it shall come to pass at that day, saith the LORD, that the heart of the king shall perish, and the heart of the princes; and the priests shall be astonished, and the prophets shall wonder.
JER|4|10|Then said I, Ah, Lord GOD! surely thou hast greatly deceived this people and Jerusalem, saying, Ye shall have peace; whereas the sword reacheth unto the soul.
JER|4|11|At that time shall it be said to this people and to Jerusalem, A dry wind of the high places in the wilderness toward the daughter of my people, not to fan, nor to cleanse,
JER|4|12|Even a full wind from those places shall come unto me: now also will I give sentence against them.
JER|4|13|Behold, he shall come up as clouds, and his chariots shall be as a whirlwind: his horses are swifter than eagles. Woe unto us! for we are spoiled.
JER|4|14|O Jerusalem, wash thine heart from wickedness, that thou mayest be saved. How long shall thy vain thoughts lodge within thee?
JER|4|15|For a voice declareth from Dan, and publisheth affliction from mount Ephraim.
JER|4|16|Make ye mention to the nations; behold, publish against Jerusalem, that watchers come from a far country, and give out their voice against the cities of Judah.
JER|4|17|As keepers of a field, are they against her round about; because she hath been rebellious against me, saith the LORD.
JER|4|18|Thy way and thy doings have procured these things unto thee; this is thy wickedness, because it is bitter, because it reacheth unto thine heart.
JER|4|19|My bowels, my bowels! I am pained at my very heart; my heart maketh a noise in me; I cannot hold my peace, because thou hast heard, O my soul, the sound of the trumpet, the alarm of war.
JER|4|20|Destruction upon destruction is cried; for the whole land is spoiled: suddenly are my tents spoiled, and my curtains in a moment.
JER|4|21|How long shall I see the standard, and hear the sound of the trumpet?
JER|4|22|For my people is foolish, they have not known me; they are sottish children, and they have none understanding: they are wise to do evil, but to do good they have no knowledge.
JER|4|23|I beheld the earth, and, lo, it was without form, and void; and the heavens, and they had no light.
JER|4|24|I beheld the mountains, and, lo, they trembled, and all the hills moved lightly.
JER|4|25|I beheld, and, lo, there was no man, and all the birds of the heavens were fled.
JER|4|26|I beheld, and, lo, the fruitful place was a wilderness, and all the cities thereof were broken down at the presence of the LORD, and by his fierce anger.
JER|4|27|For thus hath the LORD said, The whole land shall be desolate; yet will I not make a full end.
JER|4|28|For this shall the earth mourn, and the heavens above be black; because I have spoken it, I have purposed it, and will not repent, neither will I turn back from it.
JER|4|29|The whole city shall flee for the noise of the horsemen and bowmen; they shall go into thickets, and climb up upon the rocks: every city shall be forsaken, and not a man dwell therein.
JER|4|30|And when thou art spoiled, what wilt thou do? Though thou clothest thyself with crimson, though thou deckest thee with ornaments of gold, though thou rentest thy face with painting, in vain shalt thou make thyself fair; thy lovers will despise thee, they will seek thy life.
JER|4|31|For I have heard a voice as of a woman in travail, and the anguish as of her that bringeth forth her first child, the voice of the daughter of Zion, that bewaileth herself, that spreadeth her hands, saying, Woe is me now! for my soul is wearied because of murderers.
JER|5|1|Run ye to and fro through the streets of Jerusalem, and see now, and know, and seek in the broad places thereof, if ye can find a man, if there be any that executeth judgment, that seeketh the truth; and I will pardon it.
JER|5|2|And though they say, The LORD liveth; surely they swear falsely.
JER|5|3|O LORD, are not thine eyes upon the truth? thou hast stricken them, but they have not grieved; thou hast consumed them, but they have refused to receive correction: they have made their faces harder than a rock; they have refused to return.
JER|5|4|Therefore I said, Surely these are poor; they are foolish: for they know not the way of the LORD, nor the judgment of their God.
JER|5|5|I will get me unto the great men, and will speak unto them; for they have known the way of the LORD, and the judgment of their God: but these have altogether broken the yoke, and burst the bonds.
JER|5|6|Wherefore a lion out of the forest shall slay them, and a wolf of the evenings shall spoil them, a leopard shall watch over their cities: every one that goeth out thence shall be torn in pieces: because their transgressions are many, and their backslidings are increased.
JER|5|7|How shall I pardon thee for this? thy children have forsaken me, and sworn by them that are no gods: when I had fed them to the full, they then committed adultery, and assembled themselves by troops in the harlots' houses.
JER|5|8|They were as fed horses in the morning: every one neighed after his neighbour's wife.
JER|5|9|Shall I not visit for these things? saith the LORD: and shall not my soul be avenged on such a nation as this?
JER|5|10|Go ye up upon her walls, and destroy; but make not a full end: take away her battlements; for they are not the LORD's.
JER|5|11|For the house of Israel and the house of Judah have dealt very treacherously against me, saith the LORD.
JER|5|12|They have belied the LORD, and said, It is not he; neither shall evil come upon us; neither shall we see sword nor famine:
JER|5|13|And the prophets shall become wind, and the word is not in them: thus shall it be done unto them.
JER|5|14|Wherefore thus saith the LORD God of hosts, Because ye speak this word, behold, I will make my words in thy mouth fire, and this people wood, and it shall devour them.
JER|5|15|Lo, I will bring a nation upon you from far, O house of Israel, saith the LORD: it is a mighty nation, it is an ancient nation, a nation whose language thou knowest not, neither understandest what they say.
JER|5|16|Their quiver is as an open sepulchre, they are all mighty men.
JER|5|17|And they shall eat up thine harvest, and thy bread, which thy sons and thy daughters should eat: they shall eat up thy flocks and thine herds: they shall eat up thy vines and thy fig trees: they shall impoverish thy fenced cities, wherein thou trustedst, with the sword.
JER|5|18|Nevertheless in those days, saith the LORD, I will not make a full end with you.
JER|5|19|And it shall come to pass, when ye shall say, Wherefore doeth the LORD our God all these things unto us? then shalt thou answer them, Like as ye have forsaken me, and served strange gods in your land, so shall ye serve strangers in a land that is not your's.
JER|5|20|Declare this in the house of Jacob, and publish it in Judah, saying,
JER|5|21|Hear now this, O foolish people, and without understanding; which have eyes, and see not; which have ears, and hear not:
JER|5|22|Fear ye not me? saith the LORD: will ye not tremble at my presence, which have placed the sand for the bound of the sea by a perpetual decree, that it cannot pass it: and though the waves thereof toss themselves, yet can they not prevail; though they roar, yet can they not pass over it?
JER|5|23|But this people hath a revolting and a rebellious heart; they are revolted and gone.
JER|5|24|Neither say they in their heart, Let us now fear the LORD our God, that giveth rain, both the former and the latter, in his season: he reserveth unto us the appointed weeks of the harvest.
JER|5|25|Your iniquities have turned away these things, and your sins have withholden good things from you.
JER|5|26|For among my people are found wicked men: they lay wait, as he that setteth snares; they set a trap, they catch men.
JER|5|27|As a cage is full of birds, so are their houses full of deceit: therefore they are become great, and waxen rich.
JER|5|28|They are waxen fat, they shine: yea, they overpass the deeds of the wicked: they judge not the cause, the cause of the fatherless, yet they prosper; and the right of the needy do they not judge.
JER|5|29|Shall I not visit for these things? saith the LORD: shall not my soul be avenged on such a nation as this?
JER|5|30|A wonderful and horrible thing is committed in the land;
JER|5|31|The prophets prophesy falsely, and the priests bear rule by their means; and my people love to have it so: and what will ye do in the end thereof?
JER|6|1|O ye children of Benjamin, gather yourselves to flee out of the midst of Jerusalem, and blow the trumpet in Tekoa, and set up a sign of fire in Bethhaccerem: for evil appeareth out of the north, and great destruction.
JER|6|2|I have likened the daughter of Zion to a comely and delicate woman.
JER|6|3|The shepherds with their flocks shall come unto her; they shall pitch their tents against her round about; they shall feed every one in his place.
JER|6|4|Prepare ye war against her; arise, and let us go up at noon. Woe unto us! for the day goeth away, for the shadows of the evening are stretched out.
JER|6|5|Arise, and let us go by night, and let us destroy her palaces.
JER|6|6|For thus hath the LORD of hosts said, Hew ye down trees, and cast a mount against Jerusalem: this is the city to be visited; she is wholly oppression in the midst of her.
JER|6|7|As a fountain casteth out her waters, so she casteth out her wickedness: violence and spoil is heard in her; before me continually is grief and wounds.
JER|6|8|Be thou instructed, O Jerusalem, lest my soul depart from thee; lest I make thee desolate, a land not inhabited.
JER|6|9|Thus saith the LORD of hosts, They shall throughly glean the remnant of Israel as a vine: turn back thine hand as a grapegatherer into the baskets.
JER|6|10|To whom shall I speak, and give warning, that they may hear? behold, their ear is uncircumcised, and they cannot hearken: behold, the word of the LORD is unto them a reproach; they have no delight in it.
JER|6|11|Therefore I am full of the fury of the LORD; I am weary with holding in: I will pour it out upon the children abroad, and upon the assembly of young men together: for even the husband with the wife shall be taken, the aged with him that is full of days.
JER|6|12|And their houses shall be turned unto others, with their fields and wives together: for I will stretch out my hand upon the inhabitants of the land, saith the LORD.
JER|6|13|For from the least of them even unto the greatest of them every one is given to covetousness; and from the prophet even unto the priest every one dealeth falsely.
JER|6|14|They have healed also the hurt of the daughter of my people slightly, saying, Peace, peace; when there is no peace.
JER|6|15|Were they ashamed when they had committed abomination? nay, they were not at all ashamed, neither could they blush: therefore they shall fall among them that fall: at the time that I visit them they shall be cast down, saith the LORD.
JER|6|16|Thus saith the LORD, Stand ye in the ways, and see, and ask for the old paths, where is the good way, and walk therein, and ye shall find rest for your souls. But they said, We will not walk therein.
JER|6|17|Also I set watchmen over you, saying, Hearken to the sound of the trumpet. But they said, We will not hearken.
JER|6|18|Therefore hear, ye nations, and know, O congregation, what is among them.
JER|6|19|Hear, O earth: behold, I will bring evil upon this people, even the fruit of their thoughts, because they have not hearkened unto my words, nor to my law, but rejected it.
JER|6|20|To what purpose cometh there to me incense from Sheba, and the sweet cane from a far country? your burnt offerings are not acceptable, nor your sacrifices sweet unto me.
JER|6|21|Therefore thus saith the LORD, Behold, I will lay stumblingblocks before this people, and the fathers and the sons together shall fall upon them; the neighbour and his friend shall perish.
JER|6|22|Thus saith the LORD, Behold, a people cometh from the north country, and a great nation shall be raised from the sides of the earth.
JER|6|23|They shall lay hold on bow and spear; they are cruel, and have no mercy; their voice roareth like the sea; and they ride upon horses, set in array as men for war against thee, O daughter of Zion.
JER|6|24|We have heard the fame thereof: our hands wax feeble: anguish hath taken hold of us, and pain, as of a woman in travail.
JER|6|25|Go not forth into the field, nor walk by the way; for the sword of the enemy and fear is on every side.
JER|6|26|O daughter of my people, gird thee with sackcloth, and wallow thyself in ashes: make thee mourning, as for an only son, most bitter lamentation: for the spoiler shall suddenly come upon us.
JER|6|27|I have set thee for a tower and a fortress among my people, that thou mayest know and try their way.
JER|6|28|They are all grievous revolters, walking with slanders: they are brass and iron; they are all corrupters.
JER|6|29|The bellows are burned, the lead is consumed of the fire; the founder melteth in vain: for the wicked are not plucked away.
JER|6|30|Reprobate silver shall men call them, because the LORD hath rejected them.
JER|7|1|The word that came to Jeremiah from the LORD, saying,
JER|7|2|Stand in the gate of the LORD's house, and proclaim there this word, and say, Hear the word of the LORD, all ye of Judah, that enter in at these gates to worship the LORD.
JER|7|3|Thus saith the LORD of hosts, the God of Israel, Amend your ways and your doings, and I will cause you to dwell in this place.
JER|7|4|Trust ye not in lying words, saying, The temple of the LORD, The temple of the LORD, The temple of the LORD, are these.
JER|7|5|For if ye throughly amend your ways and your doings; if ye throughly execute judgment between a man and his neighbour;
JER|7|6|If ye oppress not the stranger, the fatherless, and the widow, and shed not innocent blood in this place, neither walk after other gods to your hurt:
JER|7|7|Then will I cause you to dwell in this place, in the land that I gave to your fathers, for ever and ever.
JER|7|8|Behold, ye trust in lying words, that cannot profit.
JER|7|9|Will ye steal, murder, and commit adultery, and swear falsely, and burn incense unto Baal, and walk after other gods whom ye know not;
JER|7|10|And come and stand before me in this house, which is called by my name, and say, We are delivered to do all these abominations?
JER|7|11|Is this house, which is called by my name, become a den of robbers in your eyes? Behold, even I have seen it, saith the LORD.
JER|7|12|But go ye now unto my place which was in Shiloh, where I set my name at the first, and see what I did to it for the wickedness of my people Israel.
JER|7|13|And now, because ye have done all these works, saith the LORD, and I spake unto you, rising up early and speaking, but ye heard not; and I called you, but ye answered not;
JER|7|14|Therefore will I do unto this house, which is called by my name, wherein ye trust, and unto the place which I gave to you and to your fathers, as I have done to Shiloh.
JER|7|15|And I will cast you out of my sight, as I have cast out all your brethren, even the whole seed of Ephraim.
JER|7|16|Therefore pray not thou for this people, neither lift up cry nor prayer for them, neither make intercession to me: for I will not hear thee.
JER|7|17|Seest thou not what they do in the cities of Judah and in the streets of Jerusalem?
JER|7|18|The children gather wood, and the fathers kindle the fire, and the women knead their dough, to make cakes to the queen of heaven, and to pour out drink offerings unto other gods, that they may provoke me to anger.
JER|7|19|Do they provoke me to anger? saith the LORD: do they not provoke themselves to the confusion of their own faces?
JER|7|20|Therefore thus saith the Lord GOD; Behold, mine anger and my fury shall be poured out upon this place, upon man, and upon beast, and upon the trees of the field, and upon the fruit of the ground; and it shall burn, and shall not be quenched.
JER|7|21|Thus saith the LORD of hosts, the God of Israel; Put your burnt offerings unto your sacrifices, and eat flesh.
JER|7|22|For I spake not unto your fathers, nor commanded them in the day that I brought them out of the land of Egypt, concerning burnt offerings or sacrifices:
JER|7|23|But this thing commanded I them, saying, Obey my voice, and I will be your God, and ye shall be my people: and walk ye in all the ways that I have commanded you, that it may be well unto you.
JER|7|24|But they hearkened not, nor inclined their ear, but walked in the counsels and in the imagination of their evil heart, and went backward, and not forward.
JER|7|25|Since the day that your fathers came forth out of the land of Egypt unto this day I have even sent unto you all my servants the prophets, daily rising up early and sending them:
JER|7|26|Yet they hearkened not unto me, nor inclined their ear, but hardened their neck: they did worse than their fathers.
JER|7|27|Therefore thou shalt speak all these words unto them; but they will not hearken to thee: thou shalt also call unto them; but they will not answer thee.
JER|7|28|But thou shalt say unto them, This is a nation that obeyeth not the voice of the LORD their God, nor receiveth correction: truth is perished, and is cut off from their mouth.
JER|7|29|Cut off thine hair, O Jerusalem, and cast it away, and take up a lamentation on high places; for the LORD hath rejected and forsaken the generation of his wrath.
JER|7|30|For the children of Judah have done evil in my sight, saith the LORD: they have set their abominations in the house which is called by my name, to pollute it.
JER|7|31|And they have built the high places of Tophet, which is in the valley of the son of Hinnom, to burn their sons and their daughters in the fire; which I commanded them not, neither came it into my heart.
JER|7|32|Therefore, behold, the days come, saith the LORD, that it shall no more be called Tophet, nor the valley of the son of Hinnom, but the valley of slaughter: for they shall bury in Tophet, till there be no place.
JER|7|33|And the carcases of this people shall be meat for the fowls of the heaven, and for the beasts of the earth; and none shall fray them away.
JER|7|34|Then will I cause to cease from the cities of Judah, and from the streets of Jerusalem, the voice of mirth, and the voice of gladness, the voice of the bridegroom, and the voice of the bride: for the land shall be desolate.
JER|8|1|At that time, saith the LORD, they shall bring out the bones of the kings of Judah, and the bones of his princes, and the bones of the priests, and the bones of the prophets, and the bones of the inhabitants of Jerusalem, out of their graves:
JER|8|2|And they shall spread them before the sun, and the moon, and all the host of heaven, whom they have loved, and whom they have served, and after whom they have walked, and whom they have sought, and whom they have worshipped: they shall not be gathered, nor be buried; they shall be for dung upon the face of the earth.
JER|8|3|And death shall be chosen rather than life by all the residue of them that remain of this evil family, which remain in all the places whither I have driven them, saith the LORD of hosts.
JER|8|4|Moreover thou shalt say unto them, Thus saith the LORD; Shall they fall, and not arise? shall he turn away, and not return?
JER|8|5|Why then is this people of Jerusalem slidden back by a perpetual backsliding? they hold fast deceit, they refuse to return.
JER|8|6|I hearkened and heard, but they spake not aright: no man repented him of his wickedness, saying, What have I done? every one turned to his course, as the horse rusheth into the battle.
JER|8|7|Yea, the stork in the heaven knoweth her appointed times; and the turtle and the crane and the swallow observe the time of their coming; but my people know not the judgment of the LORD.
JER|8|8|How do ye say, We are wise, and the law of the LORD is with us? Lo, certainly in vain made he it; the pen of the scribes is in vain.
JER|8|9|The wise men are ashamed, they are dismayed and taken: lo, they have rejected the word of the LORD; and what wisdom is in them?
JER|8|10|Therefore will I give their wives unto others, and their fields to them that shall inherit them: for every one from the least even unto the greatest is given to covetousness, from the prophet even unto the priest every one dealeth falsely.
JER|8|11|For they have healed the hurt of the daughter of my people slightly, saying, Peace, peace; when there is no peace.
JER|8|12|Were they ashamed when they had committed abomination? nay, they were not at all ashamed, neither could they blush: therefore shall they fall among them that fall: in the time of their visitation they shall be cast down, saith the LORD.
JER|8|13|I will surely consume them, saith the LORD: there shall be no grapes on the vine, nor figs on the fig tree, and the leaf shall fade; and the things that I have given them shall pass away from them.
JER|8|14|Why do we sit still? assemble yourselves, and let us enter into the defenced cities, and let us be silent there: for the LORD our God hath put us to silence, and given us water of gall to drink, because we have sinned against the LORD.
JER|8|15|We looked for peace, but no good came; and for a time of health, and behold trouble!
JER|8|16|The snorting of his horses was heard from Dan: the whole land trembled at the sound of the neighing of his strong ones; for they are come, and have devoured the land, and all that is in it; the city, and those that dwell therein.
JER|8|17|For, behold, I will send serpents, cockatrices, among you, which will not be charmed, and they shall bite you, saith the LORD.
JER|8|18|When I would comfort myself against sorrow, my heart is faint in me.
JER|8|19|Behold the voice of the cry of the daughter of my people because of them that dwell in a far country: Is not the LORD in Zion? is not her king in her? Why have they provoked me to anger with their graven images, and with strange vanities?
JER|8|20|The harvest is past, the summer is ended, and we are not saved.
JER|8|21|For the hurt of the daughter of my people am I hurt; I am black; astonishment hath taken hold on me.
JER|8|22|Is there no balm in Gilead; is there no physician there? why then is not the health of the daughter of my people recovered?
JER|9|1|Oh that my head were waters, and mine eyes a fountain of tears, that I might weep day and night for the slain of the daughter of my people!
JER|9|2|Oh that I had in the wilderness a lodging place of wayfaring men; that I might leave my people, and go from them! for they be all adulterers, an assembly of treacherous men.
JER|9|3|And they bend their tongues like their bow for lies: but they are not valiant for the truth upon the earth; for they proceed from evil to evil, and they know not me, saith the LORD.
JER|9|4|Take ye heed every one of his neighbour, and trust ye not in any brother: for every brother will utterly supplant, and every neighbour will walk with slanders.
JER|9|5|And they will deceive every one his neighbour, and will not speak the truth: they have taught their tongue to speak lies, and weary themselves to commit iniquity.
JER|9|6|Thine habitation is in the midst of deceit; through deceit they refuse to know me, saith the LORD.
JER|9|7|Therefore thus saith the LORD of hosts, Behold, I will melt them, and try them; for how shall I do for the daughter of my people?
JER|9|8|Their tongue is as an arrow shot out; it speaketh deceit: one speaketh peaceably to his neighbour with his mouth, but in heart he layeth his wait.
JER|9|9|Shall I not visit them for these things? saith the LORD: shall not my soul be avenged on such a nation as this?
JER|9|10|For the mountains will I take up a weeping and wailing, and for the habitations of the wilderness a lamentation, because they are burned up, so that none can pass through them; neither can men hear the voice of the cattle; both the fowl of the heavens and the beast are fled; they are gone.
JER|9|11|And I will make Jerusalem heaps, and a den of dragons; and I will make the cities of Judah desolate, without an inhabitant.
JER|9|12|Who is the wise man, that may understand this? and who is he to whom the mouth of the LORD hath spoken, that he may declare it, for what the land perisheth and is burned up like a wilderness, that none passeth through?
JER|9|13|And the LORD saith, Because they have forsaken my law which I set before them, and have not obeyed my voice, neither walked therein;
JER|9|14|But have walked after the imagination of their own heart, and after Baalim, which their fathers taught them:
JER|9|15|Therefore thus saith the LORD of hosts, the God of Israel; Behold, I will feed them, even this people, with wormwood, and give them water of gall to drink.
JER|9|16|I will scatter them also among the heathen, whom neither they nor their fathers have known: and I will send a sword after them, till I have consumed them.
JER|9|17|Thus saith the LORD of hosts, Consider ye, and call for the mourning women, that they may come; and send for cunning women, that they may come:
JER|9|18|And let them make haste, and take up a wailing for us, that our eyes may run down with tears, and our eyelids gush out with waters.
JER|9|19|For a voice of wailing is heard out of Zion, How are we spoiled! we are greatly confounded, because we have forsaken the land, because our dwellings have cast us out.
JER|9|20|Yet hear the word of the LORD, O ye women, and let your ear receive the word of his mouth, and teach your daughters wailing, and every one her neighbour lamentation.
JER|9|21|For death is come up into our windows, and is entered into our palaces, to cut off the children from without, and the young men from the streets.
JER|9|22|Speak, Thus saith the LORD, Even the carcases of men shall fall as dung upon the open field, and as the handful after the harvestman, and none shall gather them.
JER|9|23|Thus saith the LORD, Let not the wise man glory in his wisdom, neither let the mighty man glory in his might, let not the rich man glory in his riches:
JER|9|24|But let him that glorieth glory in this, that he understandeth and knoweth me, that I am the LORD which exercise lovingkindness, judgment, and righteousness, in the earth: for in these things I delight, saith the LORD.
JER|9|25|Behold, the days come, saith the LORD, that I will punish all them which are circumcised with the uncircumcised;
JER|9|26|Egypt, and Judah, and Edom, and the children of Ammon, and Moab, and all that are in the utmost corners, that dwell in the wilderness: for all these nations are uncircumcised, and all the house of Israel are uncircumcised in the heart.
JER|10|1|Hear ye the word which the LORD speaketh unto you, O house of Israel:
JER|10|2|Thus saith the LORD, Learn not the way of the heathen, and be not dismayed at the signs of heaven; for the heathen are dismayed at them.
JER|10|3|For the customs of the people are vain: for one cutteth a tree out of the forest, the work of the hands of the workman, with the axe.
JER|10|4|They deck it with silver and with gold; they fasten it with nails and with hammers, that it move not.
JER|10|5|They are upright as the palm tree, but speak not: they must needs be borne, because they cannot go. Be not afraid of them; for they cannot do evil, neither also is it in them to do good.
JER|10|6|Forasmuch as there is none like unto thee, O LORD; thou art great, and thy name is great in might.
JER|10|7|Who would not fear thee, O King of nations? for to thee doth it appertain: forasmuch as among all the wise men of the nations, and in all their kingdoms, there is none like unto thee.
JER|10|8|But they are altogether brutish and foolish: the stock is a doctrine of vanities.
JER|10|9|Silver spread into plates is brought from Tarshish, and gold from Uphaz, the work of the workman, and of the hands of the founder: blue and purple is their clothing: they are all the work of cunning men.
JER|10|10|But the LORD is the true God, he is the living God, and an everlasting king: at his wrath the earth shall tremble, and the nations shall not be able to abide his indignation.
JER|10|11|Thus shall ye say unto them, The gods that have not made the heavens and the earth, even they shall perish from the earth, and from under these heavens.
JER|10|12|He hath made the earth by his power, he hath established the world by his wisdom, and hath stretched out the heavens by his discretion.
JER|10|13|When he uttereth his voice, there is a multitude of waters in the heavens, and he causeth the vapours to ascend from the ends of the earth; he maketh lightnings with rain, and bringeth forth the wind out of his treasures.
JER|10|14|Every man is brutish in his knowledge: every founder is confounded by the graven image: for his molten image is falsehood, and there is no breath in them.
JER|10|15|They are vanity, and the work of errors: in the time of their visitation they shall perish.
JER|10|16|The portion of Jacob is not like them: for he is the former of all things; and Israel is the rod of his inheritance: The LORD of hosts is his name.
JER|10|17|Gather up thy wares out of the land, O inhabitant of the fortress.
JER|10|18|For thus saith the LORD, Behold, I will sling out the inhabitants of the land at this once, and will distress them, that they may find it so.
JER|10|19|Woe is me for my hurt! my wound is grievous; but I said, Truly this is a grief, and I must bear it.
JER|10|20|My tabernacle is spoiled, and all my cords are broken: my children are gone forth of me, and they are not: there is none to stretch forth my tent any more, and to set up my curtains.
JER|10|21|For the pastors are become brutish, and have not sought the LORD: therefore they shall not prosper, and all their flocks shall be scattered.
JER|10|22|Behold, the noise of the bruit is come, and a great commotion out of the north country, to make the cities of Judah desolate, and a den of dragons.
JER|10|23|O LORD, I know that the way of man is not in himself: it is not in man that walketh to direct his steps.
JER|10|24|O LORD, correct me, but with judgment; not in thine anger, lest thou bring me to nothing.
JER|10|25|Pour out thy fury upon the heathen that know thee not, and upon the families that call not on thy name: for they have eaten up Jacob, and devoured him, and consumed him, and have made his habitation desolate.
JER|11|1|The word that came to Jeremiah from the LORD saying,
JER|11|2|Hear ye the words of this covenant, and speak unto the men of Judah, and to the inhabitants of Jerusalem;
JER|11|3|And say thou unto them, Thus saith the LORD God of Israel; Cursed be the man that obeyeth not the words of this covenant,
JER|11|4|Which I commanded your fathers in the day that I brought them forth out of the land of Egypt, from the iron furnace, saying, Obey my voice, and do them, according to all which I command you: so shall ye be my people, and I will be your God:
JER|11|5|That I may perform the oath which I have sworn unto your fathers, to give them a land flowing with milk and honey, as it is this day. Then answered I, and said, So be it, O LORD.
JER|11|6|Then the LORD said unto me, Proclaim all these words in the cities of Judah, and in the streets of Jerusalem, saying, Hear ye the words of this covenant, and do them.
JER|11|7|For I earnestly protested unto your fathers in the day that I brought them up out of the land of Egypt, even unto this day, rising early and protesting, saying, Obey my voice.
JER|11|8|Yet they obeyed not, nor inclined their ear, but walked every one in the imagination of their evil heart: therefore I will bring upon them all the words of this covenant, which I commanded them to do: but they did them not.
JER|11|9|And the LORD said unto me, A conspiracy is found among the men of Judah, and among the inhabitants of Jerusalem.
JER|11|10|They are turned back to the iniquities of their forefathers, which refused to hear my words; and they went after other gods to serve them: the house of Israel and the house of Judah have broken my covenant which I made with their fathers.
JER|11|11|Therefore thus saith the LORD, Behold, I will bring evil upon them, which they shall not be able to escape; and though they shall cry unto me, I will not hearken unto them.
JER|11|12|Then shall the cities of Judah and inhabitants of Jerusalem go, and cry unto the gods unto whom they offer incense: but they shall not save them at all in the time of their trouble.
JER|11|13|For according to the number of thy cities were thy gods, O Judah; and according to the number of the streets of Jerusalem have ye set up altars to that shameful thing, even altars to burn incense unto Baal.
JER|11|14|Therefore pray not thou for this people, neither lift up a cry or prayer for them: for I will not hear them in the time that they cry unto me for their trouble.
JER|11|15|What hath my beloved to do in mine house, seeing she hath wrought lewdness with many, and the holy flesh is passed from thee? when thou doest evil, then thou rejoicest.
JER|11|16|The LORD called thy name, A green olive tree, fair, and of goodly fruit: with the noise of a great tumult he hath kindled fire upon it, and the branches of it are broken.
JER|11|17|For the LORD of hosts, that planted thee, hath pronounced evil against thee, for the evil of the house of Israel and of the house of Judah, which they have done against themselves to provoke me to anger in offering incense unto Baal.
JER|11|18|And the LORD hath given me knowledge of it, and I know it: then thou shewedst me their doings.
JER|11|19|But I was like a lamb or an ox that is brought to the slaughter; and I knew not that they had devised devices against me, saying, Let us destroy the tree with the fruit thereof, and let us cut him off from the land of the living, that his name may be no more remembered.
JER|11|20|But, O LORD of hosts, that judgest righteously, that triest the reins and the heart, let me see thy vengeance on them: for unto thee have I revealed my cause.
JER|11|21|Therefore thus saith the LORD of the men of Anathoth, that seek thy life, saying, Prophesy not in the name of the LORD, that thou die not by our hand:
JER|11|22|Therefore thus saith the LORD of hosts, Behold, I will punish them: the young men shall die by the sword; their sons and their daughters shall die by famine:
JER|11|23|And there shall be no remnant of them: for I will bring evil upon the men of Anathoth, even the year of their visitation.
JER|12|1|Righteous art thou, O LORD, when I plead with thee: yet let me talk with thee of thy judgments: Wherefore doth the way of the wicked prosper? wherefore are all they happy that deal very treacherously?
JER|12|2|Thou hast planted them, yea, they have taken root: they grow, yea, they bring forth fruit: thou art near in their mouth, and far from their reins.
JER|12|3|But thou, O LORD, knowest me: thou hast seen me, and tried mine heart toward thee: pull them out like sheep for the slaughter, and prepare them for the day of slaughter.
JER|12|4|How long shall the land mourn, and the herbs of every field wither, for the wickedness of them that dwell therein? the beasts are consumed, and the birds; because they said, He shall not see our last end.
JER|12|5|If thou hast run with the footmen, and they have wearied thee, then how canst thou contend with horses? and if in the land of peace, wherein thou trustedst, they wearied thee, then how wilt thou do in the swelling of Jordan?
JER|12|6|For even thy brethren, and the house of thy father, even they have dealt treacherously with thee; yea, they have called a multitude after thee: believe them not, though they speak fair words unto thee.
JER|12|7|I have forsaken mine house, I have left mine heritage; I have given the dearly beloved of my soul into the hand of her enemies.
JER|12|8|Mine heritage is unto me as a lion in the forest; it crieth out against me: therefore have I hated it.
JER|12|9|Mine heritage is unto me as a speckled bird, the birds round about are against her; come ye, assemble all the beasts of the field, come to devour.
JER|12|10|Many pastors have destroyed my vineyard, they have trodden my portion under foot, they have made my pleasant portion a desolate wilderness.
JER|12|11|They have made it desolate, and being desolate it mourneth unto me; the whole land is made desolate, because no man layeth it to heart.
JER|12|12|The spoilers are come upon all high places through the wilderness: for the sword of the LORD shall devour from the one end of the land even to the other end of the land: no flesh shall have peace.
JER|12|13|They have sown wheat, but shall reap thorns: they have put themselves to pain, but shall not profit: and they shall be ashamed of your revenues because of the fierce anger of the LORD.
JER|12|14|Thus saith the LORD against all mine evil neighbours, that touch the inheritance which I have caused my people Israel to inherit; Behold, I will pluck them out of their land, and pluck out the house of Judah from among them.
JER|12|15|And it shall come to pass, after that I have plucked them out I will return, and have compassion on them, and will bring them again, every man to his heritage, and every man to his land.
JER|12|16|And it shall come to pass, if they will diligently learn the ways of my people, to swear by my name, The LORD liveth; as they taught my people to swear by Baal; then shall they be built in the midst of my people.
JER|12|17|But if they will not obey, I will utterly pluck up and destroy that nation, saith the LORD.
JER|13|1|Thus saith the LORD unto me, Go and get thee a linen girdle, and put it upon thy loins, and put it not in water.
JER|13|2|So I got a girdle according to the word of the LORD, and put it on my loins.
JER|13|3|And the word of the LORD came unto me the second time, saying,
JER|13|4|Take the girdle that thou hast got, which is upon thy loins, and arise, go to Euphrates, and hide it there in a hole of the rock.
JER|13|5|So I went, and hid it by Euphrates, as the LORD commanded me.
JER|13|6|And it came to pass after many days, that the LORD said unto me, Arise, go to Euphrates, and take the girdle from thence, which I commanded thee to hide there.
JER|13|7|Then I went to Euphrates, and digged, and took the girdle from the place where I had hid it: and, behold, the girdle was marred, it was profitable for nothing.
JER|13|8|Then the word of the LORD came unto me, saying,
JER|13|9|Thus saith the LORD, After this manner will I mar the pride of Judah, and the great pride of Jerusalem.
JER|13|10|This evil people, which refuse to hear my words, which walk in the imagination of their heart, and walk after other gods, to serve them, and to worship them, shall even be as this girdle, which is good for nothing.
JER|13|11|For as the girdle cleaveth to the loins of a man, so have I caused to cleave unto me the whole house of Israel and the whole house of Judah, saith the LORD; that they might be unto me for a people, and for a name, and for a praise, and for a glory: but they would not hear.
JER|13|12|Therefore thou shalt speak unto them this word; Thus saith the LORD God of Israel, Every bottle shall be filled with wine: and they shall say unto thee, Do we not certainly know that every bottle shall be filled with wine?
JER|13|13|Then shalt thou say unto them, Thus saith the LORD, Behold, I will fill all the inhabitants of this land, even the kings that sit upon David's throne, and the priests, and the prophets, and all the inhabitants of Jerusalem, with drunkenness.
JER|13|14|And I will dash them one against another, even the fathers and the sons together, saith the LORD: I will not pity, nor spare, nor have mercy, but destroy them.
JER|13|15|Hear ye, and give ear; be not proud: for the LORD hath spoken.
JER|13|16|Give glory to the LORD your God, before he cause darkness, and before your feet stumble upon the dark mountains, and, while ye look for light, he turn it into the shadow of death, and make it gross darkness.
JER|13|17|But if ye will not hear it, my soul shall weep in secret places for your pride; and mine eye shall weep sore, and run down with tears, because the LORD's flock is carried away captive.
JER|13|18|Say unto the king and to the queen, Humble yourselves, sit down: for your principalities shall come down, even the crown of your glory.
JER|13|19|The cities of the south shall be shut up, and none shall open them: Judah shall be carried away captive all of it, it shall be wholly carried away captive.
JER|13|20|Lift up your eyes, and behold them that come from the north: where is the flock that was given thee, thy beautiful flock?
JER|13|21|What wilt thou say when he shall punish thee? for thou hast taught them to be captains, and as chief over thee: shall not sorrows take thee, as a woman in travail?
JER|13|22|And if thou say in thine heart, Wherefore come these things upon me? For the greatness of thine iniquity are thy skirts discovered, and thy heels made bare.
JER|13|23|Can the Ethiopian change his skin, or the leopard his spots? then may ye also do good, that are accustomed to do evil.
JER|13|24|Therefore will I scatter them as the stubble that passeth away by the wind of the wilderness.
JER|13|25|This is thy lot, the portion of thy measures from me, saith the LORD; because thou hast forgotten me, and trusted in falsehood.
JER|13|26|Therefore will I discover thy skirts upon thy face, that thy shame may appear.
JER|13|27|I have seen thine adulteries, and thy neighings, the lewdness of thy whoredom, and thine abominations on the hills in the fields. Woe unto thee, O Jerusalem! wilt thou not be made clean? when shall it once be?
JER|14|1|The word of the LORD that came to Jeremiah concerning the dearth.
JER|14|2|Judah mourneth, and the gates thereof languish; they are black unto the ground; and the cry of Jerusalem is gone up.
JER|14|3|And their nobles have sent their little ones to the waters: they came to the pits, and found no water; they returned with their vessels empty; they were ashamed and confounded, and covered their heads.
JER|14|4|Because the ground is chapt, for there was no rain in the earth, the plowmen were ashamed, they covered their heads.
JER|14|5|Yea, the hind also calved in the field, and forsook it, because there was no grass.
JER|14|6|And the wild asses did stand in the high places, they snuffed up the wind like dragons; their eyes did fail, because there was no grass.
JER|14|7|O LORD, though our iniquities testify against us, do thou it for thy name's sake: for our backslidings are many; we have sinned against thee.
JER|14|8|O the hope of Israel, the saviour thereof in time of trouble, why shouldest thou be as a stranger in the land, and as a wayfaring man that turneth aside to tarry for a night?
JER|14|9|Why shouldest thou be as a man astonied, as a mighty man that cannot save? yet thou, O LORD, art in the midst of us, and we are called by thy name; leave us not.
JER|14|10|Thus saith the LORD unto this people, Thus have they loved to wander, they have not refrained their feet, therefore the LORD doth not accept them; he will now remember their iniquity, and visit their sins.
JER|14|11|Then said the LORD unto me, Pray not for this people for their good.
JER|14|12|When they fast, I will not hear their cry; and when they offer burnt offering and an oblation, I will not accept them: but I will consume them by the sword, and by the famine, and by the pestilence.
JER|14|13|Then said I, Ah, Lord GOD! behold, the prophets say unto them, Ye shall not see the sword, neither shall ye have famine; but I will give you assured peace in this place.
JER|14|14|Then the LORD said unto me, The prophets prophesy lies in my name: I sent them not, neither have I commanded them, neither spake unto them: they prophesy unto you a false vision and divination, and a thing of nought, and the deceit of their heart.
JER|14|15|Therefore thus saith the LORD concerning the prophets that prophesy in my name, and I sent them not, yet they say, Sword and famine shall not be in this land; By sword and famine shall those prophets be consumed.
JER|14|16|And the people to whom they prophesy shall be cast out in the streets of Jerusalem because of the famine and the sword; and they shall have none to bury them, them, their wives, nor their sons, nor their daughters: for I will pour their wickedness upon them.
JER|14|17|Therefore thou shalt say this word unto them; Let mine eyes run down with tears night and day, and let them not cease: for the virgin daughter of my people is broken with a great breach, with a very grievous blow.
JER|14|18|If I go forth into the field, then behold the slain with the sword! and if I enter into the city, then behold them that are sick with famine! yea, both the prophet and the priest go about into a land that they know not.
JER|14|19|Hast thou utterly rejected Judah? hath thy soul lothed Zion? why hast thou smitten us, and there is no healing for us? we looked for peace, and there is no good; and for the time of healing, and behold trouble!
JER|14|20|We acknowledge, O LORD, our wickedness, and the iniquity of our fathers: for we have sinned against thee.
JER|14|21|Do not abhor us, for thy name's sake, do not disgrace the throne of thy glory: remember, break not thy covenant with us.
JER|14|22|Are there any among the vanities of the Gentiles that can cause rain? or can the heavens give showers? art not thou he, O LORD our God? therefore we will wait upon thee: for thou hast made all these things.
JER|15|1|Then said the LORD unto me, Though Moses and Samuel stood before me, yet my mind could not be toward this people: cast them out of my sight, and let them go forth.
JER|15|2|And it shall come to pass, if they say unto thee, Whither shall we go forth? then thou shalt tell them, Thus saith the LORD; Such as are for death, to death; and such as are for the sword, to the sword; and such as are for the famine, to the famine; and such as are for the captivity, to the captivity.
JER|15|3|And I will appoint over them four kinds, saith the LORD: the sword to slay, and the dogs to tear, and the fowls of the heaven, and the beasts of the earth, to devour and destroy.
JER|15|4|And I will cause them to be removed into all kingdoms of the earth, because of Manasseh the son of Hezekiah king of Judah, for that which he did in Jerusalem.
JER|15|5|For who shall have pity upon thee, O Jerusalem? or who shall bemoan thee? or who shall go aside to ask how thou doest?
JER|15|6|Thou hast forsaken me, saith the LORD, thou art gone backward: therefore will I stretch out my hand against thee, and destroy thee; I am weary with repenting.
JER|15|7|And I will fan them with a fan in the gates of the land; I will bereave them of children, I will destroy my people since they return not from their ways.
JER|15|8|Their widows are increased to me above the sand of the seas: I have brought upon them against the mother of the young men a spoiler at noonday: I have caused him to fall upon it suddenly, and terrors upon the city.
JER|15|9|She that hath borne seven languisheth: she hath given up the ghost; her sun is gone down while it was yet day: she hath been ashamed and confounded: and the residue of them will I deliver to the sword before their enemies, saith the LORD.
JER|15|10|Woe is me, my mother, that thou hast borne me a man of strife and a man of contention to the whole earth! I have neither lent on usury, nor men have lent to me on usury; yet every one of them doth curse me.
JER|15|11|The LORD said, Verily it shall be well with thy remnant; verily I will cause the enemy to entreat thee well in the time of evil and in the time of affliction.
JER|15|12|Shall iron break the northern iron and the steel?
JER|15|13|Thy substance and thy treasures will I give to the spoil without price, and that for all thy sins, even in all thy borders.
JER|15|14|And I will make thee to pass with thine enemies into a land which thou knowest not: for a fire is kindled in mine anger, which shall burn upon you.
JER|15|15|O LORD, thou knowest: remember me, and visit me, and revenge me of my persecutors; take me not away in thy longsuffering: know that for thy sake I have suffered rebuke.
JER|15|16|Thy words were found, and I did eat them; and thy word was unto me the joy and rejoicing of mine heart: for I am called by thy name, O LORD God of hosts.
JER|15|17|I sat not in the assembly of the mockers, nor rejoiced; I sat alone because of thy hand: for thou hast filled me with indignation.
JER|15|18|Why is my pain perpetual, and my wound incurable, which refuseth to be healed? wilt thou be altogether unto me as a liar, and as waters that fail?
JER|15|19|Therefore thus saith the LORD, If thou return, then will I bring thee again, and thou shalt stand before me: and if thou take forth the precious from the vile, thou shalt be as my mouth: let them return unto thee; but return not thou unto them.
JER|15|20|And I will make thee unto this people a fenced brasen wall: and they shall fight against thee, but they shall not prevail against thee: for I am with thee to save thee and to deliver thee, saith the LORD.
JER|15|21|And I will deliver thee out of the hand of the wicked, and I will redeem thee out of the hand of the terrible.
JER|16|1|The word of the LORD came also unto me, saying,
JER|16|2|Thou shalt not take thee a wife, neither shalt thou have sons or daughters in this place.
JER|16|3|For thus saith the LORD concerning the sons and concerning the daughters that are born in this place, and concerning their mothers that bare them, and concerning their fathers that begat them in this land;
JER|16|4|They shall die of grievous deaths; they shall not be lamented; neither shall they be buried; but they shall be as dung upon the face of the earth: and they shall be consumed by the sword, and by famine; and their carcases shall be meat for the fowls of heaven, and for the beasts of the earth.
JER|16|5|For thus saith the LORD, Enter not into the house of mourning, neither go to lament nor bemoan them: for I have taken away my peace from this people, saith the LORD, even lovingkindness and mercies.
JER|16|6|Both the great and the small shall die in this land: they shall not be buried, neither shall men lament for them, nor cut themselves, nor make themselves bald for them:
JER|16|7|Neither shall men tear themselves for them in mourning, to comfort them for the dead; neither shall men give them the cup of consolation to drink for their father or for their mother.
JER|16|8|Thou shalt not also go into the house of feasting, to sit with them to eat and to drink.
JER|16|9|For thus saith the LORD of hosts, the God of Israel; Behold, I will cause to cease out of this place in your eyes, and in your days, the voice of mirth, and the voice of gladness, the voice of the bridegroom, and the voice of the bride.
JER|16|10|And it shall come to pass, when thou shalt shew this people all these words, and they shall say unto thee, Wherefore hath the LORD pronounced all this great evil against us? or what is our iniquity? or what is our sin that we have committed against the LORD our God?
JER|16|11|Then shalt thou say unto them, Because your fathers have forsaken me, saith the LORD, and have walked after other gods, and have served them, and have worshipped them, and have forsaken me, and have not kept my law;
JER|16|12|And ye have done worse than your fathers; for, behold, ye walk every one after the imagination of his evil heart, that they may not hearken unto me:
JER|16|13|Therefore will I cast you out of this land into a land that ye know not, neither ye nor your fathers; and there shall ye serve other gods day and night; where I will not shew you favour.
JER|16|14|Therefore, behold, the days come, saith the LORD, that it shall no more be said, The LORD liveth, that brought up the children of Israel out of the land of Egypt;
JER|16|15|But, The LORD liveth, that brought up the children of Israel from the land of the north, and from all the lands whither he had driven them: and I will bring them again into their land that I gave unto their fathers.
JER|16|16|Behold, I will send for many fishers, saith the LORD, and they shall fish them; and after will I send for many hunters, and they shall hunt them from every mountain, and from every hill, and out of the holes of the rocks.
JER|16|17|For mine eyes are upon all their ways: they are not hid from my face, neither is their iniquity hid from mine eyes.
JER|16|18|And first I will recompense their iniquity and their sin double; because they have defiled my land, they have filled mine inheritance with the carcases of their detestable and abominable things.
JER|16|19|O LORD, my strength, and my fortress, and my refuge in the day of affliction, the Gentiles shall come unto thee from the ends of the earth, and shall say, Surely our fathers have inherited lies, vanity, and things wherein there is no profit.
JER|16|20|Shall a man make gods unto himself, and they are no gods?
JER|16|21|Therefore, behold, I will this once cause them to know, I will cause them to know mine hand and my might; and they shall know that my name is The LORD.
JER|17|1|The sin of Judah is written with a pen of iron, and with the point of a diamond: it is graven upon the table of their heart, and upon the horns of your altars;
JER|17|2|Whilst their children remember their altars and their groves by the green trees upon the high hills.
JER|17|3|O my mountain in the field, I will give thy substance and all thy treasures to the spoil, and thy high places for sin, throughout all thy borders.
JER|17|4|And thou, even thyself, shalt discontinue from thine heritage that I gave thee; and I will cause thee to serve thine enemies in the land which thou knowest not: for ye have kindled a fire in mine anger, which shall burn for ever.
JER|17|5|Thus saith the LORD; Cursed be the man that trusteth in man, and maketh flesh his arm, and whose heart departeth from the LORD.
JER|17|6|For he shall be like the heath in the desert, and shall not see when good cometh; but shall inhabit the parched places in the wilderness, in a salt land and not inhabited.
JER|17|7|Blessed is the man that trusteth in the LORD, and whose hope the LORD is.
JER|17|8|For he shall be as a tree planted by the waters, and that spreadeth out her roots by the river, and shall not see when heat cometh, but her leaf shall be green; and shall not be careful in the year of drought, neither shall cease from yielding fruit.
JER|17|9|The heart is deceitful above all things, and desperately wicked: who can know it?
JER|17|10|I the LORD search the heart, I try the reins, even to give every man according to his ways, and according to the fruit of his doings.
JER|17|11|As the partridge sitteth on eggs, and hatcheth them not; so he that getteth riches, and not by right, shall leave them in the midst of his days, and at his end shall be a fool.
JER|17|12|A glorious high throne from the beginning is the place of our sanctuary.
JER|17|13|O LORD, the hope of Israel, all that forsake thee shall be ashamed, and they that depart from me shall be written in the earth, because they have forsaken the LORD, the fountain of living waters.
JER|17|14|Heal me, O LORD, and I shall be healed; save me, and I shall be saved: for thou art my praise.
JER|17|15|Behold, they say unto me, Where is the word of the LORD? let it come now.
JER|17|16|As for me, I have not hastened from being a pastor to follow thee: neither have I desired the woeful day; thou knowest: that which came out of my lips was right before thee.
JER|17|17|Be not a terror unto me: thou art my hope in the day of evil.
JER|17|18|Let them be confounded that persecute me, but let not me be confounded: let them be dismayed, but let not me be dismayed: bring upon them the day of evil, and destroy them with double destruction.
JER|17|19|Thus said the LORD unto me; Go and stand in the gate of the children of the people, whereby the kings of Judah come in, and by the which they go out, and in all the gates of Jerusalem;
JER|17|20|And say unto them, Hear ye the word of the LORD, ye kings of Judah, and all Judah, and all the inhabitants of Jerusalem, that enter in by these gates:
JER|17|21|Thus saith the LORD; Take heed to yourselves, and bear no burden on the sabbath day, nor bring it in by the gates of Jerusalem;
JER|17|22|Neither carry forth a burden out of your houses on the sabbath day, neither do ye any work, but hallow ye the sabbath day, as I commanded your fathers.
JER|17|23|But they obeyed not, neither inclined their ear, but made their neck stiff, that they might not hear, nor receive instruction.
JER|17|24|And it shall come to pass, if ye diligently hearken unto me, saith the LORD, to bring in no burden through the gates of this city on the sabbath day, but hallow the sabbath day, to do no work therein;
JER|17|25|Then shall there enter into the gates of this city kings and princes sitting upon the throne of David, riding in chariots and on horses, they, and their princes, the men of Judah, and the inhabitants of Jerusalem: and this city shall remain for ever.
JER|17|26|And they shall come from the cities of Judah, and from the places about Jerusalem, and from the land of Benjamin, and from the plain, and from the mountains, and from the south, bringing burnt offerings, and sacrifices, and meat offerings, and incense, and bringing sacrifices of praise, unto the house of the LORD.
JER|17|27|But if ye will not hearken unto me to hallow the sabbath day, and not to bear a burden, even entering in at the gates of Jerusalem on the sabbath day; then will I kindle a fire in the gates thereof, and it shall devour the palaces of Jerusalem, and it shall not be quenched.
JER|18|1|The word which came to Jeremiah from the LORD, saying,
JER|18|2|Arise, and go down to the potter's house, and there I will cause thee to hear my words.
JER|18|3|Then I went down to the potter's house, and, behold, he wrought a work on the wheels.
JER|18|4|And the vessel that he made of clay was marred in the hand of the potter: so he made it again another vessel, as seemed good to the potter to make it.
JER|18|5|Then the word of the LORD came to me, saying,
JER|18|6|O house of Israel, cannot I do with you as this potter? saith the LORD. Behold, as the clay is in the potter's hand, so are ye in mine hand, O house of Israel.
JER|18|7|At what instant I shall speak concerning a nation, and concerning a kingdom, to pluck up, and to pull down, and to destroy it;
JER|18|8|If that nation, against whom I have pronounced, turn from their evil, I will repent of the evil that I thought to do unto them.
JER|18|9|And at what instant I shall speak concerning a nation, and concerning a kingdom, to build and to plant it;
JER|18|10|If it do evil in my sight, that it obey not my voice, then I will repent of the good, wherewith I said I would benefit them.
JER|18|11|Now therefore go to, speak to the men of Judah, and to the inhabitants of Jerusalem, saying, Thus saith the LORD; Behold, I frame evil against you, and devise a device against you: return ye now every one from his evil way, and make your ways and your doings good.
JER|18|12|And they said, There is no hope: but we will walk after our own devices, and we will every one do the imagination of his evil heart.
JER|18|13|Therefore thus saith the LORD; Ask ye now among the heathen, who hath heard such things: the virgin of Israel hath done a very horrible thing.
JER|18|14|Will a man leave the snow of Lebanon which cometh from the rock of the field? or shall the cold flowing waters that come from another place be forsaken?
JER|18|15|Because my people hath forgotten me, they have burned incense to vanity, and they have caused them to stumble in their ways from the ancient paths, to walk in paths, in a way not cast up;
JER|18|16|To make their land desolate, and a perpetual hissing; every one that passeth thereby shall be astonished, and wag his head.
JER|18|17|I will scatter them as with an east wind before the enemy; I will shew them the back, and not the face, in the day of their calamity.
JER|18|18|Then said they, Come and let us devise devices against Jeremiah; for the law shall not perish from the priest, nor counsel from the wise, nor the word from the prophet. Come, and let us smite him with the tongue, and let us not give heed to any of his words.
JER|18|19|Give heed to me, O LORD, and hearken to the voice of them that contend with me.
JER|18|20|Shall evil be recompensed for good? for they have digged a pit for my soul. Remember that I stood before thee to speak good for them, and to turn away thy wrath from them.
JER|18|21|Therefore deliver up their children to the famine, and pour out their blood by the force of the sword; and let their wives be bereaved of their children, and be widows; and let their men be put to death; let their young men be slain by the sword in battle.
JER|18|22|Let a cry be heard from their houses, when thou shalt bring a troop suddenly upon them: for they have digged a pit to take me, and hid snares for my feet.
JER|18|23|Yet, LORD, thou knowest all their counsel against me to slay me: forgive not their iniquity, neither blot out their sin from thy sight, but let them be overthrown before thee; deal thus with them in the time of thine anger.
JER|19|1|Thus saith the LORD, Go and get a potter's earthen bottle, and take of the ancients of the people, and of the ancients of the priests;
JER|19|2|And go forth unto the valley of the son of Hinnom, which is by the entry of the east gate, and proclaim there the words that I shall tell thee,
JER|19|3|And say, Hear ye the word of the LORD, O kings of Judah, and inhabitants of Jerusalem; Thus saith the LORD of hosts, the God of Israel; Behold, I will bring evil upon this place, the which whosoever heareth, his ears shall tingle.
JER|19|4|Because they have forsaken me, and have estranged this place, and have burned incense in it unto other gods, whom neither they nor their fathers have known, nor the kings of Judah, and have filled this place with the blood of innocents;
JER|19|5|They have built also the high places of Baal, to burn their sons with fire for burnt offerings unto Baal, which I commanded not, nor spake it, neither came it into my mind:
JER|19|6|Therefore, behold, the days come, saith the LORD, that this place shall no more be called Tophet, nor The valley of the son of Hinnom, but The valley of slaughter.
JER|19|7|And I will make void the counsel of Judah and Jerusalem in this place; and I will cause them to fall by the sword before their enemies, and by the hands of them that seek their lives: and their carcases will I give to be meat for the fowls of the heaven, and for the beasts of the earth.
JER|19|8|And I will make this city desolate, and an hissing; every one that passeth thereby shall be astonished and hiss because of all the plagues thereof.
JER|19|9|And I will cause them to eat the flesh of their sons and the flesh of their daughters, and they shall eat every one the flesh of his friend in the siege and straitness, wherewith their enemies, and they that seek their lives, shall straiten them.
JER|19|10|Then shalt thou break the bottle in the sight of the men that go with thee,
JER|19|11|And shalt say unto them, Thus saith the LORD of hosts; Even so will I break this people and this city, as one breaketh a potter's vessel, that cannot be made whole again: and they shall bury them in Tophet, till there be no place to bury.
JER|19|12|Thus will I do unto this place, saith the LORD, and to the inhabitants thereof, and even make this city as Tophet:
JER|19|13|And the houses of Jerusalem, and the houses of the kings of Judah, shall be defiled as the place of Tophet, because of all the houses upon whose roofs they have burned incense unto all the host of heaven, and have poured out drink offerings unto other gods.
JER|19|14|Then came Jeremiah from Tophet, whither the LORD had sent him to prophesy; and he stood in the court of the LORD's house; and said to all the people,
JER|19|15|Thus saith the LORD of hosts, the God of Israel; Behold, I will bring upon this city and upon all her towns all the evil that I have pronounced against it, because they have hardened their necks, that they might not hear my words.
JER|20|1|Now Pashur the son of Immer the priest, who was also chief governor in the house of the LORD, heard that Jeremiah prophesied these things.
JER|20|2|Then Pashur smote Jeremiah the prophet, and put him in the stocks that were in the high gate of Benjamin, which was by the house of the LORD.
JER|20|3|And it came to pass on the morrow, that Pashur brought forth Jeremiah out of the stocks. Then said Jeremiah unto him, The LORD hath not called thy name Pashur, but Magormissabib.
JER|20|4|For thus saith the LORD, Behold, I will make thee a terror to thyself, and to all thy friends: and they shall fall by the sword of their enemies, and thine eyes shall behold it: and I will give all Judah into the hand of the king of Babylon, and he shall carry them captive into Babylon, and shall slay them with the sword.
JER|20|5|Moreover I will deliver all the strength of this city, and all the labours thereof, and all the precious things thereof, and all the treasures of the kings of Judah will I give into the hand of their enemies, which shall spoil them, and take them, and carry them to Babylon.
JER|20|6|And thou, Pashur, and all that dwell in thine house shall go into captivity: and thou shalt come to Babylon, and there thou shalt die, and shalt be buried there, thou, and all thy friends, to whom thou hast prophesied lies.
JER|20|7|O LORD, thou hast deceived me, and I was deceived; thou art stronger than I, and hast prevailed: I am in derision daily, every one mocketh me.
JER|20|8|For since I spake, I cried out, I cried violence and spoil; because the word of the LORD was made a reproach unto me, and a derision, daily.
JER|20|9|Then I said, I will not make mention of him, nor speak any more in his name. But his word was in mine heart as a burning fire shut up in my bones, and I was weary with forbearing, and I could not stay.
JER|20|10|For I heard the defaming of many, fear on every side. Report, say they, and we will report it. All my familiars watched for my halting, saying, Peradventure he will be enticed, and we shall prevail against him, and we shall take our revenge on him.
JER|20|11|But the LORD is with me as a mighty terrible one: therefore my persecutors shall stumble, and they shall not prevail: they shall be greatly ashamed; for they shall not prosper: their everlasting confusion shall never be forgotten.
JER|20|12|But, O LORD of hosts, that triest the righteous, and seest the reins and the heart, let me see thy vengeance on them: for unto thee have I opened my cause.
JER|20|13|Sing unto the LORD, praise ye the LORD: for he hath delivered the soul of the poor from the hand of evildoers.
JER|20|14|Cursed be the day wherein I was born: let not the day wherein my mother bare me be blessed.
JER|20|15|Cursed be the man who brought tidings to my father, saying, A man child is born unto thee; making him very glad.
JER|20|16|And let that man be as the cities which the LORD overthrew, and repented not: and let him hear the cry in the morning, and the shouting at noontide;
JER|20|17|Because he slew me not from the womb; or that my mother might have been my grave, and her womb to be always great with me.
JER|20|18|Wherefore came I forth out of the womb to see labour and sorrow, that my days should be consumed with shame?
JER|21|1|The word which came unto Jeremiah from the LORD, when king Zedekiah sent unto him Pashur the son of Melchiah, and Zephaniah the son of Maaseiah the priest, saying,
JER|21|2|Enquire, I pray thee, of the LORD for us; for Nebuchadrezzar king of Babylon maketh war against us; if so be that the LORD will deal with us according to all his wondrous works, that he may go up from us.
JER|21|3|Then said Jeremiah unto them, Thus shall ye say to Zedekiah:
JER|21|4|Thus saith the LORD God of Israel; Behold, I will turn back the weapons of war that are in your hands, wherewith ye fight against the king of Babylon, and against the Chaldeans, which besiege you without the walls, and I will assemble them into the midst of this city.
JER|21|5|And I myself will fight against you with an outstretched hand and with a strong arm, even in anger, and in fury, and in great wrath.
JER|21|6|And I will smite the inhabitants of this city, both man and beast: they shall die of a great pestilence.
JER|21|7|And afterward, saith the LORD, I will deliver Zedekiah king of Judah, and his servants, and the people, and such as are left in this city from the pestilence, from the sword, and from the famine, into the hand of Nebuchadrezzar king of Babylon, and into the hand of their enemies, and into the hand of those that seek their life: and he shall smite them with the edge of the sword; he shall not spare them, neither have pity, nor have mercy.
JER|21|8|And unto this people thou shalt say, Thus saith the LORD; Behold, I set before you the way of life, and the way of death.
JER|21|9|He that abideth in this city shall die by the sword, and by the famine, and by the pestilence: but he that goeth out, and falleth to the Chaldeans that besiege you, he shall live, and his life shall be unto him for a prey.
JER|21|10|For I have set my face against this city for evil, and not for good, saith the LORD: it shall be given into the hand of the king of Babylon, and he shall burn it with fire.
JER|21|11|And touching the house of the king of Judah, say, Hear ye the word of the LORD;
JER|21|12|O house of David, thus saith the LORD; Execute judgment in the morning, and deliver him that is spoiled out of the hand of the oppressor, lest my fury go out like fire, and burn that none can quench it, because of the evil of your doings.
JER|21|13|Behold, I am against thee, O inhabitant of the valley, and rock of the plain, saith the LORD; which say, Who shall come down against us? or who shall enter into our habitations?
JER|21|14|But I will punish you according to the fruit of your doings, saith the LORD: and I will kindle a fire in the forest thereof, and it shall devour all things round about it.
JER|22|1|Thus saith the LORD; Go down to the house of the king of Judah, and speak there this word,
JER|22|2|And say, Hear the word of the LORD, O king of Judah, that sittest upon the throne of David, thou, and thy servants, and thy people that enter in by these gates:
JER|22|3|Thus saith the LORD; Execute ye judgment and righteousness, and deliver the spoiled out of the hand of the oppressor: and do no wrong, do no violence to the stranger, the fatherless, nor the widow, neither shed innocent blood in this place.
JER|22|4|For if ye do this thing indeed, then shall there enter in by the gates of this house kings sitting upon the throne of David, riding in chariots and on horses, he, and his servants, and his people.
JER|22|5|But if ye will not hear these words, I swear by myself, saith the LORD, that this house shall become a desolation.
JER|22|6|For thus saith the LORD unto the king's house of Judah; Thou art Gilead unto me, and the head of Lebanon: yet surely I will make thee a wilderness, and cities which are not inhabited.
JER|22|7|And I will prepare destroyers against thee, every one with his weapons: and they shall cut down thy choice cedars, and cast them into the fire.
JER|22|8|And many nations shall pass by this city, and they shall say every man to his neighbour, Wherefore hath the LORD done thus unto this great city?
JER|22|9|Then they shall answer, Because they have forsaken the covenant of the LORD their God, and worshipped other gods, and served them.
JER|22|10|Weep ye not for the dead, neither bemoan him: but weep sore for him that goeth away: for he shall return no more, nor see his native country.
JER|22|11|For thus saith the LORD touching Shallum the son of Josiah king of Judah, which reigned instead of Josiah his father, which went forth out of this place; He shall not return thither any more:
JER|22|12|But he shall die in the place whither they have led him captive, and shall see this land no more.
JER|22|13|Woe unto him that buildeth his house by unrighteousness, and his chambers by wrong; that useth his neighbour's service without wages, and giveth him not for his work;
JER|22|14|That saith, I will build me a wide house and large chambers, and cutteth him out windows; and it is cieled with cedar, and painted with vermilion.
JER|22|15|Shalt thou reign, because thou closest thyself in cedar? did not thy father eat and drink, and do judgment and justice, and then it was well with him?
JER|22|16|He judged the cause of the poor and needy; then it was well with him: was not this to know me? saith the LORD.
JER|22|17|But thine eyes and thine heart are not but for thy covetousness, and for to shed innocent blood, and for oppression, and for violence, to do it.
JER|22|18|Therefore thus saith the LORD concerning Jehoiakim the son of Josiah king of Judah; They shall not lament for him, saying, Ah my brother! or, Ah sister! they shall not lament for him, saying, Ah lord! or, Ah his glory!
JER|22|19|He shall be buried with the burial of an ass, drawn and cast forth beyond the gates of Jerusalem.
JER|22|20|Go up to Lebanon, and cry; and lift up thy voice in Bashan, and cry from the passages: for all thy lovers are destroyed.
JER|22|21|I spake unto thee in thy prosperity; but thou saidst, I will not hear. This hath been thy manner from thy youth, that thou obeyedst not my voice.
JER|22|22|The wind shall eat up all thy pastors, and thy lovers shall go into captivity: surely then shalt thou be ashamed and confounded for all thy wickedness.
JER|22|23|O inhabitant of Lebanon, that makest thy nest in the cedars, how gracious shalt thou be when pangs come upon thee, the pain as of a woman in travail!
JER|22|24|As I live, saith the LORD, though Coniah the son of Jehoiakim king of Judah were the signet upon my right hand, yet would I pluck thee thence;
JER|22|25|And I will give thee into the hand of them that seek thy life, and into the hand of them whose face thou fearest, even into the hand of Nebuchadrezzar king of Babylon, and into the hand of the Chaldeans.
JER|22|26|And I will cast thee out, and thy mother that bare thee, into another country, where ye were not born; and there shall ye die.
JER|22|27|But to the land whereunto they desire to return, thither shall they not return.
JER|22|28|Is this man Coniah a despised broken idol? is he a vessel wherein is no pleasure? wherefore are they cast out, he and his seed, and are cast into a land which they know not?
JER|22|29|O earth, earth, earth, hear the word of the LORD.
JER|22|30|Thus saith the LORD, Write ye this man childless, a man that shall not prosper in his days: for no man of his seed shall prosper, sitting upon the throne of David, and ruling any more in Judah.
JER|23|1|Woe be unto the pastors that destroy and scatter the sheep of my pasture! saith the LORD.
JER|23|2|Therefore thus saith the LORD God of Israel against the pastors that feed my people; Ye have scattered my flock, and driven them away, and have not visited them: behold, I will visit upon you the evil of your doings, saith the LORD.
JER|23|3|And I will gather the remnant of my flock out of all countries whither I have driven them, and will bring them again to their folds; and they shall be fruitful and increase.
JER|23|4|And I will set up shepherds over them which shall feed them: and they shall fear no more, nor be dismayed, neither shall they be lacking, saith the LORD.
JER|23|5|Behold, the days come, saith the LORD, that I will raise unto David a righteous Branch, and a King shall reign and prosper, and shall execute judgment and justice in the earth.
JER|23|6|In his days Judah shall be saved, and Israel shall dwell safely: and this is his name whereby he shall be called, THE LORD OUR RIGHTEOUSNESS.
JER|23|7|Therefore, behold, the days come, saith the LORD, that they shall no more say, The LORD liveth, which brought up the children of Israel out of the land of Egypt;
JER|23|8|But, The LORD liveth, which brought up and which led the seed of the house of Israel out of the north country, and from all countries whither I had driven them; and they shall dwell in their own land.
JER|23|9|Mine heart within me is broken because of the prophets; all my bones shake; I am like a drunken man, and like a man whom wine hath overcome, because of the LORD, and because of the words of his holiness.
JER|23|10|For the land is full of adulterers; for because of swearing the land mourneth; the pleasant places of the wilderness are dried up, and their course is evil, and their force is not right.
JER|23|11|For both prophet and priest are profane; yea, in my house have I found their wickedness, saith the LORD.
JER|23|12|Wherefore their way shall be unto them as slippery ways in the darkness: they shall be driven on, and fall therein: for I will bring evil upon them, even the year of their visitation, saith the LORD.
JER|23|13|And I have seen folly in the prophets of Samaria; they prophesied in Baal, and caused my people Israel to err.
JER|23|14|I have seen also in the prophets of Jerusalem an horrible thing: they commit adultery, and walk in lies: they strengthen also the hands of evildoers, that none doth return from his wickedness; they are all of them unto me as Sodom, and the inhabitants thereof as Gomorrah.
JER|23|15|Therefore thus saith the LORD of hosts concerning the prophets; Behold, I will feed them with wormwood, and make them drink the water of gall: for from the prophets of Jerusalem is profaneness gone forth into all the land.
JER|23|16|Thus saith the LORD of hosts, Hearken not unto the words of the prophets that prophesy unto you: they make you vain: they speak a vision of their own heart, and not out of the mouth of the LORD.
JER|23|17|They say still unto them that despise me, The LORD hath said, Ye shall have peace; and they say unto every one that walketh after the imagination of his own heart, No evil shall come upon you.
JER|23|18|For who hath stood in the counsel of the LORD, and hath perceived and heard his word? who hath marked his word, and heard it?
JER|23|19|Behold, a whirlwind of the LORD is gone forth in fury, even a grievous whirlwind: it shall fall grievously upon the head of the wicked.
JER|23|20|The anger of the LORD shall not return, until he have executed, and till he have performed the thoughts of his heart: in the latter days ye shall consider it perfectly.
JER|23|21|I have not sent these prophets, yet they ran: I have not spoken to them, yet they prophesied.
JER|23|22|But if they had stood in my counsel, and had caused my people to hear my words, then they should have turned them from their evil way, and from the evil of their doings.
JER|23|23|Am I a God at hand, saith the LORD, and not a God afar off?
JER|23|24|Can any hide himself in secret places that I shall not see him? saith the LORD. Do not I fill heaven and earth? saith the LORD.
JER|23|25|I have heard what the prophets said, that prophesy lies in my name, saying, I have dreamed, I have dreamed.
JER|23|26|How long shall this be in the heart of the prophets that prophesy lies? yea, they are prophets of the deceit of their own heart;
JER|23|27|Which think to cause my people to forget my name by their dreams which they tell every man to his neighbour, as their fathers have forgotten my name for Baal.
JER|23|28|The prophet that hath a dream, let him tell a dream; and he that hath my word, let him speak my word faithfully. What is the chaff to the wheat? saith the LORD.
JER|23|29|Is not my word like as a fire? saith the LORD; and like a hammer that breaketh the rock in pieces?
JER|23|30|Therefore, behold, I am against the prophets, saith the LORD, that steal my words every one from his neighbour.
JER|23|31|Behold, I am against the prophets, saith the LORD, that use their tongues, and say, He saith.
JER|23|32|Behold, I am against them that prophesy false dreams, saith the LORD, and do tell them, and cause my people to err by their lies, and by their lightness; yet I sent them not, nor commanded them: therefore they shall not profit this people at all, saith the LORD.
JER|23|33|And when this people, or the prophet, or a priest, shall ask thee, saying, What is the burden of the LORD? thou shalt then say unto them, What burden? I will even forsake you, saith the LORD.
JER|23|34|And as for the prophet, and the priest, and the people, that shall say, The burden of the LORD, I will even punish that man and his house.
JER|23|35|Thus shall ye say every one to his neighbour, and every one to his brother, What hath the LORD answered? and, What hath the LORD spoken?
JER|23|36|And the burden of the LORD shall ye mention no more: for every man's word shall be his burden; for ye have perverted the words of the living God, of the LORD of hosts our God.
JER|23|37|Thus shalt thou say to the prophet, What hath the LORD answered thee? and, What hath the LORD spoken?
JER|23|38|But since ye say, The burden of the LORD; therefore thus saith the LORD; Because ye say this word, The burden of the LORD, and I have sent unto you, saying, Ye shall not say, The burden of the LORD;
JER|23|39|Therefore, behold, I, even I, will utterly forget you, and I will forsake you, and the city that I gave you and your fathers, and cast you out of my presence:
JER|23|40|And I will bring an everlasting reproach upon you, and a perpetual shame, which shall not be forgotten.
JER|24|1|The LORD shewed me, and, behold, two baskets of figs were set before the temple of the LORD, after that Nebuchadrezzar king of Babylon had carried away captive Jeconiah the son of Jehoiakim king of Judah, and the princes of Judah, with the carpenters and smiths, from Jerusalem, and had brought them to Babylon.
JER|24|2|One basket had very good figs, even like the figs that are first ripe: and the other basket had very naughty figs, which could not be eaten, they were so bad.
JER|24|3|Then said the LORD unto me, What seest thou, Jeremiah? And I said, Figs; the good figs, very good; and the evil, very evil, that cannot be eaten, they are so evil.
JER|24|4|Again the word of the LORD came unto me, saying,
JER|24|5|Thus saith the LORD, the God of Israel; Like these good figs, so will I acknowledge them that are carried away captive of Judah, whom I have sent out of this place into the land of the Chaldeans for their good.
JER|24|6|For I will set mine eyes upon them for good, and I will bring them again to this land: and I will build them, and not pull them down; and I will plant them, and not pluck them up.
JER|24|7|And I will give them an heart to know me, that I am the LORD: and they shall be my people, and I will be their God: for they shall return unto me with their whole heart.
JER|24|8|And as the evil figs, which cannot be eaten, they are so evil; surely thus saith the LORD, So will I give Zedekiah the king of Judah, and his princes, and the residue of Jerusalem, that remain in this land, and them that dwell in the land of Egypt:
JER|24|9|And I will deliver them to be removed into all the kingdoms of the earth for their hurt, to be a reproach and a proverb, a taunt and a curse, in all places whither I shall drive them.
JER|24|10|And I will send the sword, the famine, and the pestilence, among them, till they be consumed from off the land that I gave unto them and to their fathers.
JER|25|1|The word that came to Jeremiah concerning all the people of Judah in the fourth year of Jehoiakim the son of Josiah king of Judah, that was the first year of Nebuchadrezzar king of Babylon;
JER|25|2|The which Jeremiah the prophet spake unto all the people of Judah, and to all the inhabitants of Jerusalem, saying,
JER|25|3|From the thirteenth year of Josiah the son of Amon king of Judah, even unto this day, that is the three and twentieth year, the word of the LORD hath come unto me, and I have spoken unto you, rising early and speaking; but ye have not hearkened.
JER|25|4|And the LORD hath sent unto you all his servants the prophets, rising early and sending them; but ye have not hearkened, nor inclined your ear to hear.
JER|25|5|They said, Turn ye again now every one from his evil way, and from the evil of your doings, and dwell in the land that the LORD hath given unto you and to your fathers for ever and ever:
JER|25|6|And go not after other gods to serve them, and to worship them, and provoke me not to anger with the works of your hands; and I will do you no hurt.
JER|25|7|Yet ye have not hearkened unto me, saith the LORD; that ye might provoke me to anger with the works of your hands to your own hurt.
JER|25|8|Therefore thus saith the LORD of hosts; Because ye have not heard my words,
JER|25|9|Behold, I will send and take all the families of the north, saith the LORD, and Nebuchadrezzar the king of Babylon, my servant, and will bring them against this land, and against the inhabitants thereof, and against all these nations round about, and will utterly destroy them, and make them an astonishment, and an hissing, and perpetual desolations.
JER|25|10|Moreover I will take from them the voice of mirth, and the voice of gladness, the voice of the bridegroom, and the voice of the bride, the sound of the millstones, and the light of the candle.
JER|25|11|And this whole land shall be a desolation, and an astonishment; and these nations shall serve the king of Babylon seventy years.
JER|25|12|And it shall come to pass, when seventy years are accomplished, that I will punish the king of Babylon, and that nation, saith the LORD, for their iniquity, and the land of the Chaldeans, and will make it perpetual desolations.
JER|25|13|And I will bring upon that land all my words which I have pronounced against it, even all that is written in this book, which Jeremiah hath prophesied against all the nations.
JER|25|14|For many nations and great kings shall serve themselves of them also: and I will recompense them according to their deeds, and according to the works of their own hands.
JER|25|15|For thus saith the LORD God of Israel unto me; Take the wine cup of this fury at my hand, and cause all the nations, to whom I send thee, to drink it.
JER|25|16|And they shall drink, and be moved, and be mad, because of the sword that I will send among them.
JER|25|17|Then took I the cup at the LORD's hand, and made all the nations to drink, unto whom the LORD had sent me:
JER|25|18|To wit, Jerusalem, and the cities of Judah, and the kings thereof, and the princes thereof, to make them a desolation, an astonishment, an hissing, and a curse; as it is this day;
JER|25|19|Pharaoh king of Egypt, and his servants, and his princes, and all his people;
JER|25|20|And all the mingled people, and all the kings of the land of Uz, and all the kings of the land of the Philistines, and Ashkelon, and Azzah, and Ekron, and the remnant of Ashdod,
JER|25|21|Edom, and Moab, and the children of Ammon,
JER|25|22|And all the kings of Tyrus, and all the kings of Zidon, and the kings of the isles which are beyond the sea,
JER|25|23|Dedan, and Tema, and Buz, and all that are in the utmost corners,
JER|25|24|And all the kings of Arabia, and all the kings of the mingled people that dwell in the desert,
JER|25|25|And all the kings of Zimri, and all the kings of Elam, and all the kings of the Medes,
JER|25|26|And all the kings of the north, far and near, one with another, and all the kingdoms of the world, which are upon the face of the earth: and the king of Sheshach shall drink after them.
JER|25|27|Therefore thou shalt say unto them, Thus saith the LORD of hosts, the God of Israel; Drink ye, and be drunken, and spue, and fall, and rise no more, because of the sword which I will send among you.
JER|25|28|And it shall be, if they refuse to take the cup at thine hand to drink, then shalt thou say unto them, Thus saith the LORD of hosts; Ye shall certainly drink.
JER|25|29|For, lo, I begin to bring evil on the city which is called by my name, and should ye be utterly unpunished? Ye shall not be unpunished: for I will call for a sword upon all the inhabitants of the earth, saith the LORD of hosts.
JER|25|30|Therefore prophesy thou against them all these words, and say unto them, The LORD shall roar from on high, and utter his voice from his holy habitation; he shall mightily roar upon his habitation; he shall give a shout, as they that tread the grapes, against all the inhabitants of the earth.
JER|25|31|A noise shall come even to the ends of the earth; for the LORD hath a controversy with the nations, he will plead with all flesh; he will give them that are wicked to the sword, saith the LORD.
JER|25|32|Thus saith the LORD of hosts, Behold, evil shall go forth from nation to nation, and a great whirlwind shall be raised up from the coasts of the earth.
JER|25|33|And the slain of the LORD shall be at that day from one end of the earth even unto the other end of the earth: they shall not be lamented, neither gathered, nor buried; they shall be dung upon the ground.
JER|25|34|Howl, ye shepherds, and cry; and wallow yourselves in the ashes, ye principal of the flock: for the days of your slaughter and of your dispersions are accomplished; and ye shall fall like a pleasant vessel.
JER|25|35|And the shepherds shall have no way to flee, nor the principal of the flock to escape.
JER|25|36|A voice of the cry of the shepherds, and an howling of the principal of the flock, shall be heard: for the LORD hath spoiled their pasture.
JER|25|37|And the peaceable habitations are cut down because of the fierce anger of the LORD.
JER|25|38|He hath forsaken his covert, as the lion: for their land is desolate because of the fierceness of the oppressor, and because of his fierce anger.
JER|26|1|In the beginning of the reign of Jehoiakim the son of Josiah king of Judah came this word from the LORD, saying,
JER|26|2|Thus saith the LORD; Stand in the court of the LORD's house, and speak unto all the cities of Judah, which come to worship in the LORD's house, all the words that I command thee to speak unto them; diminish not a word:
JER|26|3|If so be they will hearken, and turn every man from his evil way, that I may repent me of the evil, which I purpose to do unto them because of the evil of their doings.
JER|26|4|And thou shalt say unto them, Thus saith the LORD; If ye will not hearken to me, to walk in my law, which I have set before you,
JER|26|5|To hearken to the words of my servants the prophets, whom I sent unto you, both rising up early, and sending them, but ye have not hearkened;
JER|26|6|Then will I make this house like Shiloh, and will make this city a curse to all the nations of the earth.
JER|26|7|So the priests and the prophets and all the people heard Jeremiah speaking these words in the house of the LORD.
JER|26|8|Now it came to pass, when Jeremiah had made an end of speaking all that the LORD had commanded him to speak unto all the people, that the priests and the prophets and all the people took him, saying, Thou shalt surely die.
JER|26|9|Why hast thou prophesied in the name of the LORD, saying, This house shall be like Shiloh, and this city shall be desolate without an inhabitant? And all the people were gathered against Jeremiah in the house of the LORD.
JER|26|10|When the princes of Judah heard these things, then they came up from the king's house unto the house of the LORD, and sat down in the entry of the new gate of the LORD's house.
JER|26|11|Then spake the priests and the prophets unto the princes and to all the people, saying, This man is worthy to die; for he hath prophesied against this city, as ye have heard with your ears.
JER|26|12|Then spake Jeremiah unto all the princes and to all the people, saying, The LORD sent me to prophesy against this house and against this city all the words that ye have heard.
JER|26|13|Therefore now amend your ways and your doings, and obey the voice of the LORD your God; and the LORD will repent him of the evil that he hath pronounced against you.
JER|26|14|As for me, behold, I am in your hand: do with me as seemeth good and meet unto you.
JER|26|15|But know ye for certain, that if ye put me to death, ye shall surely bring innocent blood upon yourselves, and upon this city, and upon the inhabitants thereof: for of a truth the LORD hath sent me unto you to speak all these words in your ears.
JER|26|16|Then said the princes and all the people unto the priests and to the prophets; This man is not worthy to die: for he hath spoken to us in the name of the LORD our God.
JER|26|17|Then rose up certain of the elders of the land, and spake to all the assembly of the people, saying,
JER|26|18|Micah the Morasthite prophesied in the days of Hezekiah king of Judah, and spake to all the people of Judah, saying, Thus saith the LORD of hosts; Zion shall be plowed like a field, and Jerusalem shall become heaps, and the mountain of the house as the high places of a forest.
JER|26|19|Did Hezekiah king of Judah and all Judah put him at all to death? did he not fear the LORD, and besought the LORD, and the LORD repented him of the evil which he had pronounced against them? Thus might we procure great evil against our souls.
JER|26|20|And there was also a man that prophesied in the name of the LORD, Urijah the son of Shemaiah of Kirjathjearim, who prophesied against this city and against this land according to all the words of Jeremiah.
JER|26|21|And when Jehoiakim the king, with all his mighty men, and all the princes, heard his words, the king sought to put him to death: but when Urijah heard it, he was afraid, and fled, and went into Egypt;
JER|26|22|And Jehoiakim the king sent men into Egypt, namely, Elnathan the son of Achbor, and certain men with him into Egypt.
JER|26|23|And they fetched forth Urijah out of Egypt, and brought him unto Jehoiakim the king; who slew him with the sword, and cast his dead body into the graves of the common people.
JER|26|24|Nevertheless the hand of Ahikam the son of Shaphan was with Jeremiah, that they should not give him into the hand of the people to put him to death.
JER|27|1|In the beginning of the reign of Jehoiakim the son of Josiah king of Judah came this word unto Jeremiah from the LORD, saying,
JER|27|2|Thus saith the LORD to me; Make thee bonds and yokes, and put them upon thy neck,
JER|27|3|And send them to the king of Edom, and to the king of Moab, and to the king of the Ammonites, and to the king of Tyrus, and to the king of Zidon, by the hand of the messengers which come to Jerusalem unto Zedekiah king of Judah;
JER|27|4|And command them to say unto their masters, Thus saith the LORD of hosts, the God of Israel; Thus shall ye say unto your masters;
JER|27|5|I have made the earth, the man and the beast that are upon the ground, by my great power and by my outstretched arm, and have given it unto whom it seemed meet unto me.
JER|27|6|And now have I given all these lands into the hand of Nebuchadnezzar the king of Babylon, my servant; and the beasts of the field have I given him also to serve him.
JER|27|7|And all nations shall serve him, and his son, and his son's son, until the very time of his land come: and then many nations and great kings shall serve themselves of him.
JER|27|8|And it shall come to pass, that the nation and kingdom which will not serve the same Nebuchadnezzar the king of Babylon, and that will not put their neck under the yoke of the king of Babylon, that nation will I punish, saith the LORD, with the sword, and with the famine, and with the pestilence, until I have consumed them by his hand.
JER|27|9|Therefore hearken not ye to your prophets, nor to your diviners, nor to your dreamers, nor to your enchanters, nor to your sorcerers, which speak unto you, saying, Ye shall not serve the king of Babylon:
JER|27|10|For they prophesy a lie unto you, to remove you far from your land; and that I should drive you out, and ye should perish.
JER|27|11|But the nations that bring their neck under the yoke of the king of Babylon, and serve him, those will I let remain still in their own land, saith the LORD; and they shall till it, and dwell therein.
JER|27|12|I spake also to Zedekiah king of Judah according to all these words, saying, Bring your necks under the yoke of the king of Babylon, and serve him and his people, and live.
JER|27|13|Why will ye die, thou and thy people, by the sword, by the famine, and by the pestilence, as the LORD hath spoken against the nation that will not serve the king of Babylon?
JER|27|14|Therefore hearken not unto the words of the prophets that speak unto you, saying, Ye shall not serve the king of Babylon: for they prophesy a lie unto you.
JER|27|15|For I have not sent them, saith the LORD, yet they prophesy a lie in my name; that I might drive you out, and that ye might perish, ye, and the prophets that prophesy unto you.
JER|27|16|Also I spake to the priests and to all this people, saying, Thus saith the LORD; Hearken not to the words of your prophets that prophesy unto you, saying, Behold, the vessels of the LORD's house shall now shortly be brought again from Babylon: for they prophesy a lie unto you.
JER|27|17|Hearken not unto them; serve the king of Babylon, and live: wherefore should this city be laid waste?
JER|27|18|But if they be prophets, and if the word of the LORD be with them, let them now make intercession to the LORD of hosts, that the vessels which are left in the house of the LORD, and in the house of the king of Judah, and at Jerusalem, go not to Babylon.
JER|27|19|For thus saith the LORD of hosts concerning the pillars, and concerning the sea, and concerning the bases, and concerning the residue of the vessels that remain in this city.
JER|27|20|Which Nebuchadnezzar king of Babylon took not, when he carried away captive Jeconiah the son of Jehoiakim king of Judah from Jerusalem to Babylon, and all the nobles of Judah and Jerusalem;
JER|27|21|Yea, thus saith the LORD of hosts, the God of Israel, concerning the vessels that remain in the house of the LORD, and in the house of the king of Judah and of Jerusalem;
JER|27|22|They shall be carried to Babylon, and there shall they be until the day that I visit them, saith the LORD; then will I bring them up, and restore them to this place.
JER|28|1|And it came to pass the same year, in the beginning of the reign of Zedekiah king of Judah, in the fourth year, and in the fifth month, that Hananiah the son of Azur the prophet, which was of Gibeon, spake unto me in the house of the LORD, in the presence of the priests and of all the people, saying,
JER|28|2|Thus speaketh the LORD of hosts, the God of Israel, saying, I have broken the yoke of the king of Babylon.
JER|28|3|Within two full years will I bring again into this place all the vessels of the LORD's house, that Nebuchadnezzar king of Babylon took away from this place, and carried them to Babylon:
JER|28|4|And I will bring again to this place Jeconiah the son of Jehoiakim king of Judah, with all the captives of Judah, that went into Babylon, saith the LORD: for I will break the yoke of the king of Babylon.
JER|28|5|Then the prophet Jeremiah said unto the prophet Hananiah in the presence of the priests, and in the presence of all the people that stood in the house of the LORD,
JER|28|6|Even the prophet Jeremiah said, Amen: the LORD do so: the LORD perform thy words which thou hast prophesied, to bring again the vessels of the LORD's house, and all that is carried away captive, from Babylon into this place.
JER|28|7|Nevertheless hear thou now this word that I speak in thine ears, and in the ears of all the people;
JER|28|8|The prophets that have been before me and before thee of old prophesied both against many countries, and against great kingdoms, of war, and of evil, and of pestilence.
JER|28|9|The prophet which prophesieth of peace, when the word of the prophet shall come to pass, then shall the prophet be known, that the LORD hath truly sent him.
JER|28|10|Then Hananiah the prophet took the yoke from off the prophet Jeremiah's neck, and brake it.
JER|28|11|And Hananiah spake in the presence of all the people, saying, Thus saith the LORD; Even so will I break the yoke of Nebuchadnezzar king of Babylon from the neck of all nations within the space of two full years. And the prophet Jeremiah went his way.
JER|28|12|Then the word of the LORD came unto Jeremiah the prophet, after that Hananiah the prophet had broken the yoke from off the neck of the prophet Jeremiah, saying,
JER|28|13|Go and tell Hananiah, saying, Thus saith the LORD; Thou hast broken the yokes of wood; but thou shalt make for them yokes of iron.
JER|28|14|For thus saith the LORD of hosts, the God of Israel; I have put a yoke of iron upon the neck of all these nations, that they may serve Nebuchadnezzar king of Babylon; and they shall serve him: and I have given him the beasts of the field also.
JER|28|15|Then said the prophet Jeremiah unto Hananiah the prophet, Hear now, Hananiah; The LORD hath not sent thee; but thou makest this people to trust in a lie.
JER|28|16|Therefore thus saith the LORD; Behold, I will cast thee from off the face of the earth: this year thou shalt die, because thou hast taught rebellion against the LORD.
JER|28|17|So Hananiah the prophet died the same year in the seventh month.
JER|29|1|Now these are the words of the letter that Jeremiah the prophet sent from Jerusalem unto the residue of the elders which were carried away captives, and to the priests, and to the prophets, and to all the people whom Nebuchadnezzar had carried away captive from Jerusalem to Babylon;
JER|29|2|(After that Jeconiah the king, and the queen, and the eunuchs, the princes of Judah and Jerusalem, and the carpenters, and the smiths, were departed from Jerusalem;)
JER|29|3|By the hand of Elasah the son of Shaphan, and Gemariah the son of Hilkiah, (whom Zedekiah king of Judah sent unto Babylon to Nebuchadnezzar king of Babylon) saying,
JER|29|4|Thus saith the LORD of hosts, the God of Israel, unto all that are carried away captives, whom I have caused to be carried away from Jerusalem unto Babylon;
JER|29|5|Build ye houses, and dwell in them; and plant gardens, and eat the fruit of them;
JER|29|6|Take ye wives, and beget sons and daughters; and take wives for your sons, and give your daughters to husbands, that they may bear sons and daughters; that ye may be increased there, and not diminished.
JER|29|7|And seek the peace of the city whither I have caused you to be carried away captives, and pray unto the LORD for it: for in the peace thereof shall ye have peace.
JER|29|8|For thus saith the LORD of hosts, the God of Israel; Let not your prophets and your diviners, that be in the midst of you, deceive you, neither hearken to your dreams which ye cause to be dreamed.
JER|29|9|For they prophesy falsely unto you in my name: I have not sent them, saith the LORD.
JER|29|10|For thus saith the LORD, That after seventy years be accomplished at Babylon I will visit you, and perform my good word toward you, in causing you to return to this place.
JER|29|11|For I know the thoughts that I think toward you, saith the LORD, thoughts of peace, and not of evil, to give you an expected end.
JER|29|12|Then shall ye call upon me, and ye shall go and pray unto me, and I will hearken unto you.
JER|29|13|And ye shall seek me, and find me, when ye shall search for me with all your heart.
JER|29|14|And I will be found of you, saith the LORD: and I will turn away your captivity, and I will gather you from all the nations, and from all the places whither I have driven you, saith the LORD; and I will bring you again into the place whence I caused you to be carried away captive.
JER|29|15|Because ye have said, The LORD hath raised us up prophets in Babylon;
JER|29|16|Know that thus saith the LORD of the king that sitteth upon the throne of David, and of all the people that dwelleth in this city, and of your brethren that are not gone forth with you into captivity;
JER|29|17|Thus saith the LORD of hosts; Behold, I will send upon them the sword, the famine, and the pestilence, and will make them like vile figs, that cannot be eaten, they are so evil.
JER|29|18|And I will persecute them with the sword, with the famine, and with the pestilence, and will deliver them to be removed to all the kingdoms of the earth, to be a curse, and an astonishment, and an hissing, and a reproach, among all the nations whither I have driven them:
JER|29|19|Because they have not hearkened to my words, saith the LORD, which I sent unto them by my servants the prophets, rising up early and sending them; but ye would not hear, saith the LORD.
JER|29|20|Hear ye therefore the word of the LORD, all ye of the captivity, whom I have sent from Jerusalem to Babylon:
JER|29|21|Thus saith the LORD of hosts, the God of Israel, of Ahab the son of Kolaiah, and of Zedekiah the son of Maaseiah, which prophesy a lie unto you in my name; Behold, I will deliver them into the hand of Nebuchadrezzar king of Babylon; and he shall slay them before your eyes;
JER|29|22|And of them shall be taken up a curse by all the captivity of Judah which are in Babylon, saying, The LORD make thee like Zedekiah and like Ahab, whom the king of Babylon roasted in the fire;
JER|29|23|Because they have committed villany in Israel, and have committed adultery with their neighbours' wives, and have spoken lying words in my name, which I have not commanded them; even I know, and am a witness, saith the LORD.
JER|29|24|Thus shalt thou also speak to Shemaiah the Nehelamite, saying,
JER|29|25|Thus speaketh the LORD of hosts, the God of Israel, saying, Because thou hast sent letters in thy name unto all the people that are at Jerusalem, and to Zephaniah the son of Maaseiah the priest, and to all the priests, saying,
JER|29|26|The LORD hath made thee priest in the stead of Jehoiada the priest, that ye should be officers in the house of the LORD, for every man that is mad, and maketh himself a prophet, that thou shouldest put him in prison, and in the stocks.
JER|29|27|Now therefore why hast thou not reproved Jeremiah of Anathoth, which maketh himself a prophet to you?
JER|29|28|For therefore he sent unto us in Babylon, saying, This captivity is long: build ye houses, and dwell in them; and plant gardens, and eat the fruit of them.
JER|29|29|And Zephaniah the priest read this letter in the ears of Jeremiah the prophet.
JER|29|30|Then came the word of the LORD unto Jeremiah, saying,
JER|29|31|Send to all them of the captivity, saying, Thus saith the LORD concerning Shemaiah the Nehelamite; Because that Shemaiah hath prophesied unto you, and I sent him not, and he caused you to trust in a lie:
JER|29|32|Therefore thus saith the LORD; Behold, I will punish Shemaiah the Nehelamite, and his seed: he shall not have a man to dwell among this people; neither shall he behold the good that I will do for my people, saith the LORD; because he hath taught rebellion against the LORD.
JER|30|1|The word that came to Jeremiah from the LORD, saying,
JER|30|2|Thus speaketh the LORD God of Israel, saying, Write thee all the words that I have spoken unto thee in a book.
JER|30|3|For, lo, the days come, saith the LORD, that I will bring again the captivity of my people Israel and Judah, saith the LORD: and I will cause them to return to the land that I gave to their fathers, and they shall possess it.
JER|30|4|And these are the words that the LORD spake concerning Israel and concerning Judah.
JER|30|5|For thus saith the LORD; We have heard a voice of trembling, of fear, and not of peace.
JER|30|6|Ask ye now, and see whether a man doth travail with child? wherefore do I see every man with his hands on his loins, as a woman in travail, and all faces are turned into paleness?
JER|30|7|Alas! for that day is great, so that none is like it: it is even the time of Jacob's trouble, but he shall be saved out of it.
JER|30|8|For it shall come to pass in that day, saith the LORD of hosts, that I will break his yoke from off thy neck, and will burst thy bonds, and strangers shall no more serve themselves of him:
JER|30|9|But they shall serve the LORD their God, and David their king, whom I will raise up unto them.
JER|30|10|Therefore fear thou not, O my servant Jacob, saith the LORD; neither be dismayed, O Israel: for, lo, I will save thee from afar, and thy seed from the land of their captivity; and Jacob shall return, and shall be in rest, and be quiet, and none shall make him afraid.
JER|30|11|For I am with thee, saith the LORD, to save thee: though I make a full end of all nations whither I have scattered thee, yet I will not make a full end of thee: but I will correct thee in measure, and will not leave thee altogether unpunished.
JER|30|12|For thus saith the LORD, Thy bruise is incurable, and thy wound is grievous.
JER|30|13|There is none to plead thy cause, that thou mayest be bound up: thou hast no healing medicines.
JER|30|14|All thy lovers have forgotten thee; they seek thee not; for I have wounded thee with the wound of an enemy, with the chastisement of a cruel one, for the multitude of thine iniquity; because thy sins were increased.
JER|30|15|Why criest thou for thine affliction? thy sorrow is incurable for the multitude of thine iniquity: because thy sins were increased, I have done these things unto thee.
JER|30|16|Therefore all they that devour thee shall be devoured; and all thine adversaries, every one of them, shall go into captivity; and they that spoil thee shall be a spoil, and all that prey upon thee will I give for a prey.
JER|30|17|For I will restore health unto thee, and I will heal thee of thy wounds, saith the LORD; because they called thee an Outcast, saying, This is Zion, whom no man seeketh after.
JER|30|18|Thus saith the LORD; Behold, I will bring again the captivity of Jacob's tents, and have mercy on his dwellingplaces; and the city shall be builded upon her own heap, and the palace shall remain after the manner thereof.
JER|30|19|And out of them shall proceed thanksgiving and the voice of them that make merry: and I will multiply them, and they shall not be few; I will also glorify them, and they shall not be small.
JER|30|20|Their children also shall be as aforetime, and their congregation shall be established before me, and I will punish all that oppress them.
JER|30|21|And their nobles shall be of themselves, and their governor shall proceed from the midst of them; and I will cause him to draw near, and he shall approach unto me: for who is this that engaged his heart to approach unto me? saith the LORD.
JER|30|22|And ye shall be my people, and I will be your God.
JER|30|23|Behold, the whirlwind of the LORD goeth forth with fury, a continuing whirlwind: it shall fall with pain upon the head of the wicked.
JER|30|24|The fierce anger of the LORD shall not return, until he hath done it, and until he have performed the intents of his heart: in the latter days ye shall consider it.
JER|31|1|At the same time, saith the LORD, will I be the God of all the families of Israel, and they shall be my people.
JER|31|2|Thus saith the LORD, The people which were left of the sword found grace in the wilderness; even Israel, when I went to cause him to rest.
JER|31|3|The LORD hath appeared of old unto me, saying, Yea, I have loved thee with an everlasting love: therefore with lovingkindness have I drawn thee.
JER|31|4|Again I will build thee, and thou shalt be built, O virgin of Israel: thou shalt again be adorned with thy tabrets, and shalt go forth in the dances of them that make merry.
JER|31|5|Thou shalt yet plant vines upon the mountains of Samaria: the planters shall plant, and shall eat them as common things.
JER|31|6|For there shall be a day, that the watchmen upon the mount Ephraim shall cry, Arise ye, and let us go up to Zion unto the LORD our God.
JER|31|7|For thus saith the LORD; Sing with gladness for Jacob, and shout among the chief of the nations: publish ye, praise ye, and say, O LORD, save thy people, the remnant of Israel.
JER|31|8|Behold, I will bring them from the north country, and gather them from the coasts of the earth, and with them the blind and the lame, the woman with child and her that travaileth with child together: a great company shall return thither.
JER|31|9|They shall come with weeping, and with supplications will I lead them: I will cause them to walk by the rivers of waters in a straight way, wherein they shall not stumble: for I am a father to Israel, and Ephraim is my firstborn.
JER|31|10|Hear the word of the LORD, O ye nations, and declare it in the isles afar off, and say, He that scattered Israel will gather him, and keep him, as a shepherd doth his flock.
JER|31|11|For the LORD hath redeemed Jacob, and ransomed him from the hand of him that was stronger than he.
JER|31|12|Therefore they shall come and sing in the height of Zion, and shall flow together to the goodness of the LORD, for wheat, and for wine, and for oil, and for the young of the flock and of the herd: and their soul shall be as a watered garden; and they shall not sorrow any more at all.
JER|31|13|Then shall the virgin rejoice in the dance, both young men and old together: for I will turn their mourning into joy, and will comfort them, and make them rejoice from their sorrow.
JER|31|14|And I will satiate the soul of the priests with fatness, and my people shall be satisfied with my goodness, saith the LORD.
JER|31|15|Thus saith the LORD; A voice was heard in Ramah, lamentation, and bitter weeping; Rahel weeping for her children refused to be comforted for her children, because they were not.
JER|31|16|Thus saith the LORD; Refrain thy voice from weeping, and thine eyes from tears: for thy work shall be rewarded, saith the LORD; and they shall come again from the land of the enemy.
JER|31|17|And there is hope in thine end, saith the LORD, that thy children shall come again to their own border.
JER|31|18|I have surely heard Ephraim bemoaning himself thus; Thou hast chastised me, and I was chastised, as a bullock unaccustomed to the yoke: turn thou me, and I shall be turned; for thou art the LORD my God.
JER|31|19|Surely after that I was turned, I repented; and after that I was instructed, I smote upon my thigh: I was ashamed, yea, even confounded, because I did bear the reproach of my youth.
JER|31|20|Is Ephraim my dear son? is he a pleasant child? for since I spake against him, I do earnestly remember him still: therefore my bowels are troubled for him; I will surely have mercy upon him, saith the LORD.
JER|31|21|Set thee up waymarks, make thee high heaps: set thine heart toward the highway, even the way which thou wentest: turn again, O virgin of Israel, turn again to these thy cities.
JER|31|22|How long wilt thou go about, O thou backsliding daughter? for the LORD hath created a new thing in the earth, A woman shall compass a man.
JER|31|23|Thus saith the LORD of hosts, the God of Israel; As yet they shall use this speech in the land of Judah and in the cities thereof, when I shall bring again their captivity; The LORD bless thee, O habitation of justice, and mountain of holiness.
JER|31|24|And there shall dwell in Judah itself, and in all the cities thereof together, husbandmen, and they that go forth with flocks.
JER|31|25|For I have satiated the weary soul, and I have replenished every sorrowful soul.
JER|31|26|Upon this I awaked, and beheld; and my sleep was sweet unto me.
JER|31|27|Behold, the days come, saith the LORD, that I will sow the house of Israel and the house of Judah with the seed of man, and with the seed of beast.
JER|31|28|And it shall come to pass, that like as I have watched over them, to pluck up, and to break down, and to throw down, and to destroy, and to afflict; so will I watch over them, to build, and to plant, saith the LORD.
JER|31|29|In those days they shall say no more, The fathers have eaten a sour grape, and the children's teeth are set on edge.
JER|31|30|But every one shall die for his own iniquity: every man that eateth the sour grape, his teeth shall be set on edge.
JER|31|31|Behold, the days come, saith the LORD, that I will make a new covenant with the house of Israel, and with the house of Judah:
JER|31|32|Not according to the covenant that I made with their fathers in the day that I took them by the hand to bring them out of the land of Egypt; which my covenant they brake, although I was an husband unto them, saith the LORD:
JER|31|33|But this shall be the covenant that I will make with the house of Israel; After those days, saith the LORD, I will put my law in their inward parts, and write it in their hearts; and will be their God, and they shall be my people.
JER|31|34|And they shall teach no more every man his neighbour, and every man his brother, saying, Know the LORD: for they shall all know me, from the least of them unto the greatest of them, saith the LORD: for I will forgive their iniquity, and I will remember their sin no more.
JER|31|35|Thus saith the LORD, which giveth the sun for a light by day, and the ordinances of the moon and of the stars for a light by night, which divideth the sea when the waves thereof roar; The LORD of hosts is his name:
JER|31|36|If those ordinances depart from before me, saith the LORD, then the seed of Israel also shall cease from being a nation before me for ever.
JER|31|37|Thus saith the LORD; If heaven above can be measured, and the foundations of the earth searched out beneath, I will also cast off all the seed of Israel for all that they have done, saith the LORD.
JER|31|38|Behold, the days come, saith the LORD, that the city shall be built to the LORD from the tower of Hananeel unto the gate of the corner.
JER|31|39|And the measuring line shall yet go forth over against it upon the hill Gareb, and shall compass about to Goath.
JER|31|40|And the whole valley of the dead bodies, and of the ashes, and all the fields unto the brook of Kidron, unto the corner of the horse gate toward the east, shall be holy unto the LORD; it shall not be plucked up, nor thrown down any more for ever.
JER|32|1|The word that came to Jeremiah from the LORD in the tenth year of Zedekiah king of Judah, which was the eighteenth year of Nebuchadrezzar.
JER|32|2|For then the king of Babylon's army besieged Jerusalem: and Jeremiah the prophet was shut up in the court of the prison, which was in the king of Judah's house.
JER|32|3|For Zedekiah king of Judah had shut him up, saying, Wherefore dost thou prophesy, and say, Thus saith the LORD, Behold, I will give this city into the hand of the king of Babylon, and he shall take it;
JER|32|4|And Zedekiah king of Judah shall not escape out of the hand of the Chaldeans, but shall surely be delivered into the hand of the king of Babylon, and shall speak with him mouth to mouth, and his eyes shall behold his eyes;
JER|32|5|And he shall lead Zedekiah to Babylon, and there shall he be until I visit him, saith the LORD: though ye fight with the Chaldeans, ye shall not prosper.
JER|32|6|And Jeremiah said, The word of the LORD came unto me, saying,
JER|32|7|Behold, Hanameel the son of Shallum thine uncle shall come unto thee saying, Buy thee my field that is in Anathoth: for the right of redemption is thine to buy it.
JER|32|8|So Hanameel mine uncle's son came to me in the court of the prison according to the word of the LORD, and said unto me, Buy my field, I pray thee, that is in Anathoth, which is in the country of Benjamin: for the right of inheritance is thine, and the redemption is thine; buy it for thyself. Then I knew that this was the word of the LORD.
JER|32|9|And I bought the field of Hanameel my uncle's son, that was in Anathoth, and weighed him the money, even seventeen shekels of silver.
JER|32|10|And I subscribed the evidence, and sealed it, and took witnesses, and weighed him the money in the balances.
JER|32|11|So I took the evidence of the purchase, both that which was sealed according to the law and custom, and that which was open:
JER|32|12|And I gave the evidence of the purchase unto Baruch the son of Neriah, the son of Maaseiah, in the sight of Hanameel mine uncle's son, and in the presence of the witnesses that subscribed the book of the purchase, before all the Jews that sat in the court of the prison.
JER|32|13|And I charged Baruch before them, saying,
JER|32|14|Thus saith the LORD of hosts, the God of Israel; Take these evidences, this evidence of the purchase, both which is sealed, and this evidence which is open; and put them in an earthen vessel, that they may continue many days.
JER|32|15|For thus saith the LORD of hosts, the God of Israel; Houses and fields and vineyards shall be possessed again in this land.
JER|32|16|Now when I had delivered the evidence of the purchase unto Baruch the son of Neriah, I prayed unto the LORD, saying,
JER|32|17|Ah Lord GOD! behold, thou hast made the heaven and the earth by thy great power and stretched out arm, and there is nothing too hard for thee:
JER|32|18|Thou shewest lovingkindness unto thousands, and recompensest the iniquity of the fathers into the bosom of their children after them: the Great, the Mighty God, the LORD of hosts, is his name,
JER|32|19|Great in counsel, and mighty in work: for thine eyes are open upon all the ways of the sons of men: to give every one according to his ways, and according to the fruit of his doings:
JER|32|20|Which hast set signs and wonders in the land of Egypt, even unto this day, and in Israel, and among other men; and hast made thee a name, as at this day;
JER|32|21|And hast brought forth thy people Israel out of the land of Egypt with signs, and with wonders, and with a strong hand, and with a stretched out arm, and with great terror;
JER|32|22|And hast given them this land, which thou didst swear to their fathers to give them, a land flowing with milk and honey;
JER|32|23|And they came in, and possessed it; but they obeyed not thy voice, neither walked in thy law; they have done nothing of all that thou commandedst them to do: therefore thou hast caused all this evil to come upon them:
JER|32|24|Behold the mounts, they are come unto the city to take it; and the city is given into the hand of the Chaldeans, that fight against it, because of the sword, and of the famine, and of the pestilence: and what thou hast spoken is come to pass; and, behold, thou seest it.
JER|32|25|And thou hast said unto me, O Lord GOD, Buy thee the field for money, and take witnesses; for the city is given into the hand of the Chaldeans.
JER|32|26|Then came the word of the LORD unto Jeremiah, saying,
JER|32|27|Behold, I am the LORD, the God of all flesh: is there any thing too hard for me?
JER|32|28|Therefore thus saith the LORD; Behold, I will give this city into the hand of the Chaldeans, and into the hand of Nebuchadrezzar king of Babylon, and he shall take it:
JER|32|29|And the Chaldeans, that fight against this city, shall come and set fire on this city, and burn it with the houses, upon whose roofs they have offered incense unto Baal, and poured out drink offerings unto other gods, to provoke me to anger.
JER|32|30|For the children of Israel and the children of Judah have only done evil before me from their youth: for the children of Israel have only provoked me to anger with the work of their hands, saith the LORD.
JER|32|31|For this city hath been to me as a provocation of mine anger and of my fury from the day that they built it even unto this day; that I should remove it from before my face,
JER|32|32|Because of all the evil of the children of Israel and of the children of Judah, which they have done to provoke me to anger, they, their kings, their princes, their priests, and their prophets, and the men of Judah, and the inhabitants of Jerusalem.
JER|32|33|And they have turned unto me the back, and not the face: though I taught them, rising up early and teaching them, yet they have not hearkened to receive instruction.
JER|32|34|But they set their abominations in the house, which is called by my name, to defile it.
JER|32|35|And they built the high places of Baal, which are in the valley of the son of Hinnom, to cause their sons and their daughters to pass through the fire unto Molech; which I commanded them not, neither came it into my mind, that they should do this abomination, to cause Judah to sin.
JER|32|36|And now therefore thus saith the LORD, the God of Israel, concerning this city, whereof ye say, It shall be delivered into the hand of the king of Babylon by the sword, and by the famine, and by the pestilence;
JER|32|37|Behold, I will gather them out of all countries, whither I have driven them in mine anger, and in my fury, and in great wrath; and I will bring them again unto this place, and I will cause them to dwell safely:
JER|32|38|And they shall be my people, and I will be their God:
JER|32|39|And I will give them one heart, and one way, that they may fear me for ever, for the good of them, and of their children after them:
JER|32|40|And I will make an everlasting covenant with them, that I will not turn away from them, to do them good; but I will put my fear in their hearts, that they shall not depart from me.
JER|32|41|Yea, I will rejoice over them to do them good, and I will plant them in this land assuredly with my whole heart and with my whole soul.
JER|32|42|For thus saith the LORD; Like as I have brought all this great evil upon this people, so will I bring upon them all the good that I have promised them.
JER|32|43|And fields shall be bought in this land, whereof ye say, It is desolate without man or beast; it is given into the hand of the Chaldeans.
JER|32|44|Men shall buy fields for money, and subscribe evidences, and seal them, and take witnesses in the land of Benjamin, and in the places about Jerusalem, and in the cities of Judah, and in the cities of the mountains, and in the cities of the valley, and in the cities of the south: for I will cause their captivity to return, saith the LORD.
JER|33|1|Moreover the word of the LORD came unto Jeremiah the second time, while he was yet shut up in the court of the prison, saying,
JER|33|2|Thus saith the LORD the maker thereof, the LORD that formed it, to establish it; the LORD is his name;
JER|33|3|Call unto me, and I will answer thee, and shew thee great and mighty things, which thou knowest not.
JER|33|4|For thus saith the LORD, the God of Israel, concerning the houses of this city, and concerning the houses of the kings of Judah, which are thrown down by the mounts, and by the sword;
JER|33|5|They come to fight with the Chaldeans, but it is to fill them with the dead bodies of men, whom I have slain in mine anger and in my fury, and for all whose wickedness I have hid my face from this city.
JER|33|6|Behold, I will bring it health and cure, and I will cure them, and will reveal unto them the abundance of peace and truth.
JER|33|7|And I will cause the captivity of Judah and the captivity of Israel to return, and will build them, as at the first.
JER|33|8|And I will cleanse them from all their iniquity, whereby they have sinned against me; and I will pardon all their iniquities, whereby they have sinned, and whereby they have transgressed against me.
JER|33|9|And it shall be to me a name of joy, a praise and an honour before all the nations of the earth, which shall hear all the good that I do unto them: and they shall fear and tremble for all the goodness and for all the prosperity that I procure unto it.
JER|33|10|Thus saith the LORD; Again there shall be heard in this place, which ye say shall be desolate without man and without beast, even in the cities of Judah, and in the streets of Jerusalem, that are desolate, without man, and without inhabitant, and without beast,
JER|33|11|The voice of joy, and the voice of gladness, the voice of the bridegroom, and the voice of the bride, the voice of them that shall say, Praise the LORD of hosts: for the LORD is good; for his mercy endureth for ever: and of them that shall bring the sacrifice of praise into the house of the LORD. For I will cause to return the captivity of the land, as at the first, saith the LORD.
JER|33|12|Thus saith the LORD of hosts; Again in this place, which is desolate without man and without beast, and in all the cities thereof, shall be an habitation of shepherds causing their flocks to lie down.
JER|33|13|In the cities of the mountains, in the cities of the vale, and in the cities of the south, and in the land of Benjamin, and in the places about Jerusalem, and in the cities of Judah, shall the flocks pass again under the hands of him that telleth them, saith the LORD.
JER|33|14|Behold, the days come, saith the LORD, that I will perform that good thing which I have promised unto the house of Israel and to the house of Judah.
JER|33|15|In those days, and at that time, will I cause the Branch of righteousness to grow up unto David; and he shall execute judgment and righteousness in the land.
JER|33|16|In those days shall Judah be saved, and Jerusalem shall dwell safely: and this is the name wherewith she shall be called, The LORD our righteousness.
JER|33|17|For thus saith the LORD; David shall never want a man to sit upon the throne of the house of Israel;
JER|33|18|Neither shall the priests the Levites want a man before me to offer burnt offerings, and to kindle meat offerings, and to do sacrifice continually.
JER|33|19|And the word of the LORD came unto Jeremiah, saying,
JER|33|20|Thus saith the LORD; If ye can break my covenant of the day, and my covenant of the night, and that there should not be day and night in their season;
JER|33|21|Then may also my covenant be broken with David my servant, that he should not have a son to reign upon his throne; and with the Levites the priests, my ministers.
JER|33|22|As the host of heaven cannot be numbered, neither the sand of the sea measured: so will I multiply the seed of David my servant, and the Levites that minister unto me.
JER|33|23|Moreover the word of the LORD came to Jeremiah, saying,
JER|33|24|Considerest thou not what this people have spoken, saying, The two families which the LORD hath chosen, he hath even cast them off? thus they have despised my people, that they should be no more a nation before them.
JER|33|25|Thus saith the LORD; If my covenant be not with day and night, and if I have not appointed the ordinances of heaven and earth;
JER|33|26|Then will I cast away the seed of Jacob and David my servant, so that I will not take any of his seed to be rulers over the seed of Abraham, Isaac, and Jacob: for I will cause their captivity to return, and have mercy on them.
JER|34|1|The word which came unto Jeremiah from the LORD, when Nebuchadnezzar king of Babylon, and all his army, and all the kingdoms of the earth of his dominion, and all the people, fought against Jerusalem, and against all the cities thereof, saying,
JER|34|2|Thus saith the LORD, the God of Israel; Go and speak to Zedekiah king of Judah, and tell him, Thus saith the LORD; Behold, I will give this city into the hand of the king of Babylon, and he shall burn it with fire:
JER|34|3|And thou shalt not escape out of his hand, but shalt surely be taken, and delivered into his hand; and thine eyes shall behold the eyes of the king of Babylon, and he shall speak with thee mouth to mouth, and thou shalt go to Babylon.
JER|34|4|Yet hear the word of the LORD, O Zedekiah king of Judah; Thus saith the LORD of thee, Thou shalt not die by the sword:
JER|34|5|But thou shalt die in peace: and with the burnings of thy fathers, the former kings which were before thee, so shall they burn odours for thee; and they will lament thee, saying, Ah lord! for I have pronounced the word, saith the LORD.
JER|34|6|Then Jeremiah the prophet spake all these words unto Zedekiah king of Judah in Jerusalem,
JER|34|7|When the king of Babylon's army fought against Jerusalem, and against all the cities of Judah that were left, against Lachish, and against Azekah: for these defenced cities remained of the cities of Judah.
JER|34|8|This is the word that came unto Jeremiah from the LORD, after that the king Zedekiah had made a covenant with all the people which were at Jerusalem, to proclaim liberty unto them;
JER|34|9|That every man should let his manservant, and every man his maidservant, being an Hebrew or an Hebrewess, go free; that none should serve himself of them, to wit, of a Jew his brother.
JER|34|10|Now when all the princes, and all the people, which had entered into the covenant, heard that every one should let his manservant, and every one his maidservant, go free, that none should serve themselves of them any more, then they obeyed, and let them go.
JER|34|11|But afterward they turned, and caused the servants and the handmaids, whom they had let go free, to return, and brought them into subjection for servants and for handmaids.
JER|34|12|Therefore the word of the LORD came to Jeremiah from the LORD, saying,
JER|34|13|Thus saith the LORD, the God of Israel; I made a covenant with your fathers in the day that I brought them forth out of the land of Egypt, out of the house of bondmen, saying,
JER|34|14|At the end of seven years let ye go every man his brother an Hebrew, which hath been sold unto thee; and when he hath served thee six years, thou shalt let him go free from thee: but your fathers hearkened not unto me, neither inclined their ear.
JER|34|15|And ye were now turned, and had done right in my sight, in proclaiming liberty every man to his neighbour; and ye had made a covenant before me in the house which is called by my name:
JER|34|16|But ye turned and polluted my name, and caused every man his servant, and every man his handmaid, whom he had set at liberty at their pleasure, to return, and brought them into subjection, to be unto you for servants and for handmaids.
JER|34|17|Therefore thus saith the LORD; Ye have not hearkened unto me, in proclaiming liberty, every one to his brother, and every man to his neighbour: behold, I proclaim a liberty for you, saith the LORD, to the sword, to the pestilence, and to the famine; and I will make you to be removed into all the kingdoms of the earth.
JER|34|18|And I will give the men that have transgressed my covenant, which have not performed the words of the covenant which they had made before me, when they cut the calf in twain, and passed between the parts thereof,
JER|34|19|The princes of Judah, and the princes of Jerusalem, the eunuchs, and the priests, and all the people of the land, which passed between the parts of the calf;
JER|34|20|I will even give them into the hand of their enemies, and into the hand of them that seek their life: and their dead bodies shall be for meat unto the fowls of the heaven, and to the beasts of the earth.
JER|34|21|And Zedekiah king of Judah and his princes will I give into the hand of their enemies, and into the hand of them that seek their life, and into the hand of the king of Babylon's army, which are gone up from you.
JER|34|22|Behold, I will command, saith the LORD, and cause them to return to this city; and they shall fight against it, and take it, and burn it with fire: and I will make the cities of Judah a desolation without an inhabitant.
JER|35|1|The word which came unto Jeremiah from the LORD in the days of Jehoiakim the son of Josiah king of Judah, saying,
JER|35|2|Go unto the house of the Rechabites, and speak unto them, and bring them into the house of the LORD, into one of the chambers, and give them wine to drink.
JER|35|3|Then I took Jaazaniah the son of Jeremiah, the son of Habaziniah, and his brethren, and all his sons, and the whole house of the Rechabites;
JER|35|4|And I brought them into the house of the LORD, into the chamber of the sons of Hanan, the son of Igdaliah, a man of God, which was by the chamber of the princes, which was above the chamber of Maaseiah the son of Shallum, the keeper of the door:
JER|35|5|And I set before the sons of the house of the Rechabites pots full of wine, and cups, and I said unto them, Drink ye wine.
JER|35|6|But they said, We will drink no wine: for Jonadab the son of Rechab our father commanded us, saying, Ye shall drink no wine, neither ye, nor your sons for ever:
JER|35|7|Neither shall ye build house, nor sow seed, nor plant vineyard, nor have any: but all your days ye shall dwell in tents; that ye may live many days in the land where ye be strangers.
JER|35|8|Thus have we obeyed the voice of Jonadab the son of Rechab our father in all that he hath charged us, to drink no wine all our days, we, our wives, our sons, nor our daughters;
JER|35|9|Nor to build houses for us to dwell in: neither have we vineyard, nor field, nor seed:
JER|35|10|But we have dwelt in tents, and have obeyed, and done according to all that Jonadab our father commanded us.
JER|35|11|But it came to pass, when Nebuchadrezzar king of Babylon came up into the land, that we said, Come, and let us go to Jerusalem for fear of the army of the Chaldeans, and for fear of the army of the Syrians: so we dwell at Jerusalem.
JER|35|12|Then came the word of the LORD unto Jeremiah, saying,
JER|35|13|Thus saith the LORD of hosts, the God of Israel; Go and tell the men of Judah and the inhabitants of Jerusalem, Will ye not receive instruction to hearken to my words? saith the LORD.
JER|35|14|The words of Jonadab the son of Rechab, that he commanded his sons not to drink wine, are performed; for unto this day they drink none, but obey their father's commandment: notwithstanding I have spoken unto you, rising early and speaking; but ye hearkened not unto me.
JER|35|15|I have sent also unto you all my servants the prophets, rising up early and sending them, saying, Return ye now every man from his evil way, and amend your doings, and go not after other gods to serve them, and ye shall dwell in the land which I have given to you and to your fathers: but ye have not inclined your ear, nor hearkened unto me.
JER|35|16|Because the sons of Jonadab the son of Rechab have performed the commandment of their father, which he commanded them; but this people hath not hearkened unto me:
JER|35|17|Therefore thus saith the LORD God of hosts, the God of Israel; Behold, I will bring upon Judah and upon all the inhabitants of Jerusalem all the evil that I have pronounced against them: because I have spoken unto them, but they have not heard; and I have called unto them, but they have not answered.
JER|35|18|And Jeremiah said unto the house of the Rechabites, Thus saith the LORD of hosts, the God of Israel; Because ye have obeyed the commandment of Jonadab your father, and kept all his precepts, and done according unto all that he hath commanded you:
JER|35|19|Therefore thus saith the LORD of hosts, the God of Israel; Jonadab the son of Rechab shall not want a man to stand before me for ever.
JER|36|1|And it came to pass in the fourth year of Jehoiakim the son of Josiah king of Judah, that this word came unto Jeremiah from the LORD, saying,
JER|36|2|Take thee a roll of a book, and write therein all the words that I have spoken unto thee against Israel, and against Judah, and against all the nations, from the day I spake unto thee, from the days of Josiah, even unto this day.
JER|36|3|It may be that the house of Judah will hear all the evil which I purpose to do unto them; that they may return every man from his evil way; that I may forgive their iniquity and their sin.
JER|36|4|Then Jeremiah called Baruch the son of Neriah: and Baruch wrote from the mouth of Jeremiah all the words of the LORD, which he had spoken unto him, upon a roll of a book.
JER|36|5|And Jeremiah commanded Baruch, saying, I am shut up; I cannot go into the house of the LORD:
JER|36|6|Therefore go thou, and read in the roll, which thou hast written from my mouth, the words of the LORD in the ears of the people in the LORD's house upon the fasting day: and also thou shalt read them in the ears of all Judah that come out of their cities.
JER|36|7|It may be they will present their supplication before the LORD, and will return every one from his evil way: for great is the anger and the fury that the LORD hath pronounced against this people.
JER|36|8|And Baruch the son of Neriah did according to all that Jeremiah the prophet commanded him, reading in the book the words of the LORD in the LORD's house.
JER|36|9|And it came to pass in the fifth year of Jehoiakim the son of Josiah king of Judah, in the ninth month, that they proclaimed a fast before the LORD to all the people in Jerusalem, and to all the people that came from the cities of Judah unto Jerusalem.
JER|36|10|Then read Baruch in the book the words of Jeremiah in the house of the LORD, in the chamber of Gemariah the son of Shaphan the scribe, in the higher court, at the entry of the new gate of the LORD's house, in the ears of all the people.
JER|36|11|When Michaiah the son of Gemariah, the son of Shaphan, had heard out of the book all the words of the LORD,
JER|36|12|Then he went down into the king's house, into the scribe's chamber: and, lo, all the princes sat there, even Elishama the scribe, and Delaiah the son of Shemaiah, and Elnathan the son of Achbor, and Gemariah the son of Shaphan, and Zedekiah the son of Hananiah, and all the princes.
JER|36|13|Then Michaiah declared unto them all the words that he had heard, when Baruch read the book in the ears of the people.
JER|36|14|Therefore all the princes sent Jehudi the son of Nethaniah, the son of Shelemiah, the son of Cushi, unto Baruch, saying, Take in thine hand the roll wherein thou hast read in the ears of the people, and come. So Baruch the son of Neriah took the roll in his hand, and came unto them.
JER|36|15|And they said unto him, Sit down now, and read it in our ears. So Baruch read it in their ears.
JER|36|16|Now it came to pass, when they had heard all the words, they were afraid both one and other, and said unto Baruch, We will surely tell the king of all these words.
JER|36|17|And they asked Baruch, saying, Tell us now, How didst thou write all these words at his mouth?
JER|36|18|Then Baruch answered them, He pronounced all these words unto me with his mouth, and I wrote them with ink in the book.
JER|36|19|Then said the princes unto Baruch, Go, hide thee, thou and Jeremiah; and let no man know where ye be.
JER|36|20|And they went in to the king into the court, but they laid up the roll in the chamber of Elishama the scribe, and told all the words in the ears of the king.
JER|36|21|So the king sent Jehudi to fetch the roll: and he took it out of Elishama the scribe's chamber. And Jehudi read it in the ears of the king, and in the ears of all the princes which stood beside the king.
JER|36|22|Now the king sat in the winterhouse in the ninth month: and there was a fire on the hearth burning before him.
JER|36|23|And it came to pass, that when Jehudi had read three or four leaves, he cut it with the penknife, and cast it into the fire that was on the hearth, until all the roll was consumed in the fire that was on the hearth.
JER|36|24|Yet they were not afraid, nor rent their garments, neither the king, nor any of his servants that heard all these words.
JER|36|25|Nevertheless Elnathan and Delaiah and Gemariah had made intercession to the king that he would not burn the roll: but he would not hear them.
JER|36|26|But the king commanded Jerahmeel the son of Hammelech, and Seraiah the son of Azriel, and Shelemiah the son of Abdeel, to take Baruch the scribe and Jeremiah the prophet: but the LORD hid them.
JER|36|27|Then the word of the LORD came to Jeremiah, after that the king had burned the roll, and the words which Baruch wrote at the mouth of Jeremiah, saying,
JER|36|28|Take thee again another roll, and write in it all the former words that were in the first roll, which Jehoiakim the king of Judah hath burned.
JER|36|29|And thou shalt say to Jehoiakim king of Judah, Thus saith the LORD; Thou hast burned this roll, saying, Why hast thou written therein, saying, The king of Babylon shall certainly come and destroy this land, and shall cause to cease from thence man and beast?
JER|36|30|Therefore thus saith the LORD of Jehoiakim king of Judah; He shall have none to sit upon the throne of David: and his dead body shall be cast out in the day to the heat, and in the night to the frost.
JER|36|31|And I will punish him and his seed and his servants for their iniquity; and I will bring upon them, and upon the inhabitants of Jerusalem, and upon the men of Judah, all the evil that I have pronounced against them; but they hearkened not.
JER|36|32|Then took Jeremiah another roll, and gave it to Baruch the scribe, the son of Neriah; who wrote therein from the mouth of Jeremiah all the words of the book which Jehoiakim king of Judah had burned in the fire: and there were added besides unto them many like words.
JER|37|1|And king Zedekiah the son of Josiah reigned instead of Coniah the son of Jehoiakim, whom Nebuchadrezzar king of Babylon made king in the land of Judah.
JER|37|2|But neither he, nor his servants, nor the people of the land, did hearken unto the words of the LORD, which he spake by the prophet Jeremiah.
JER|37|3|And Zedekiah the king sent Jehucal the son of Shelemiah and Zephaniah the son of Maaseiah the priest to the prophet Jeremiah, saying, Pray now unto the LORD our God for us.
JER|37|4|Now Jeremiah came in and went out among the people: for they had not put him into prison.
JER|37|5|Then Pharaoh's army was come forth out of Egypt: and when the Chaldeans that besieged Jerusalem heard tidings of them, they departed from Jerusalem.
JER|37|6|Then came the word of the LORD unto the prophet Jeremiah saying,
JER|37|7|Thus saith the LORD, the God of Israel; Thus shall ye say to the king of Judah, that sent you unto me to enquire of me; Behold, Pharaoh's army, which is come forth to help you, shall return to Egypt into their own land.
JER|37|8|And the Chaldeans shall come again, and fight against this city, and take it, and burn it with fire.
JER|37|9|Thus saith the LORD; Deceive not yourselves, saying, The Chaldeans shall surely depart from us: for they shall not depart.
JER|37|10|For though ye had smitten the whole army of the Chaldeans that fight against you, and there remained but wounded men among them, yet should they rise up every man in his tent, and burn this city with fire.
JER|37|11|And it came to pass, that when the army of the Chaldeans was broken up from Jerusalem for fear of Pharaoh's army,
JER|37|12|Then Jeremiah went forth out of Jerusalem to go into the land of Benjamin, to separate himself thence in the midst of the people.
JER|37|13|And when he was in the gate of Benjamin, a captain of the ward was there, whose name was Irijah, the son of Shelemiah, the son of Hananiah; and he took Jeremiah the prophet, saying, Thou fallest away to the Chaldeans.
JER|37|14|Then said Jeremiah, It is false; I fall not away to the Chaldeans. But he hearkened not to him: so Irijah took Jeremiah, and brought him to the princes.
JER|37|15|Wherefore the princes were wroth with Jeremiah, and smote him, and put him in prison in the house of Jonathan the scribe: for they had made that the prison.
JER|37|16|When Jeremiah was entered into the dungeon, and into the cabins, and Jeremiah had remained there many days;
JER|37|17|Then Zedekiah the king sent, and took him out: and the king asked him secretly in his house, and said, Is there any word from the LORD? And Jeremiah said, There is: for, said he, thou shalt be delivered into the hand of the king of Babylon.
JER|37|18|Moreover Jeremiah said unto king Zedekiah, What have I offended against thee, or against thy servants, or against this people, that ye have put me in prison?
JER|37|19|Where are now your prophets which prophesied unto you, saying, The king of Babylon shall not come against you, nor against this land?
JER|37|20|Therefore hear now, I pray thee, O my lord the king: let my supplication, I pray thee, be accepted before thee; that thou cause me not to return to the house of Jonathan the scribe, lest I die there.
JER|37|21|Then Zedekiah the king commanded that they should commit Jeremiah into the court of the prison, and that they should give him daily a piece of bread out of the bakers' street, until all the bread in the city were spent. Thus Jeremiah remained in the court of the prison.
JER|38|1|Then Shephatiah the son of Mattan, and Gedaliah the son of Pashur, and Jucal the son of Shelemiah, and Pashur the son of Malchiah, heard the words that Jeremiah had spoken unto all the people, saying,
JER|38|2|Thus saith the LORD, He that remaineth in this city shall die by the sword, by the famine, and by the pestilence: but he that goeth forth to the Chaldeans shall live; for he shall have his life for a prey, and shall live.
JER|38|3|Thus saith the LORD, This city shall surely be given into the hand of the king of Babylon's army, which shall take it.
JER|38|4|Therefore the princes said unto the king, We beseech thee, let this man be put to death: for thus he weakeneth the hands of the men of war that remain in this city, and the hands of all the people, in speaking such words unto them: for this man seeketh not the welfare of this people, but the hurt.
JER|38|5|Then Zedekiah the king said, Behold, he is in your hand: for the king is not he that can do any thing against you.
JER|38|6|Then took they Jeremiah, and cast him into the dungeon of Malchiah the son of Hammelech, that was in the court of the prison: and they let down Jeremiah with cords. And in the dungeon there was no water, but mire: so Jeremiah sunk in the mire.
JER|38|7|Now when Ebedmelech the Ethiopian, one of the eunuchs which was in the king's house, heard that they had put Jeremiah in the dungeon; the king then sitting in the gate of Benjamin;
JER|38|8|Ebedmelech went forth out of the king's house, and spake to the king saying,
JER|38|9|My lord the king, these men have done evil in all that they have done to Jeremiah the prophet, whom they have cast into the dungeon; and he is like to die for hunger in the place where he is: for there is no more bread in the city.
JER|38|10|Then the king commanded Ebedmelech the Ethiopian, saying, Take from hence thirty men with thee, and take up Jeremiah the prophet out of the dungeon, before he die.
JER|38|11|So Ebedmelech took the men with him, and went into the house of the king under the treasury, and took thence old cast clouts and old rotten rags, and let them down by cords into the dungeon to Jeremiah.
JER|38|12|And Ebedmelech the Ethiopian said unto Jeremiah, Put now these old cast clouts and rotten rags under thine armholes under the cords. And Jeremiah did so.
JER|38|13|So they drew up Jeremiah with cords, and took him up out of the dungeon: and Jeremiah remained in the court of the prison.
JER|38|14|Then Zedekiah the king sent, and took Jeremiah the prophet unto him into the third entry that is in the house of the LORD: and the king said unto Jeremiah, I will ask thee a thing; hide nothing from me.
JER|38|15|Then Jeremiah said unto Zedekiah, If I declare it unto thee, wilt thou not surely put me to death? and if I give thee counsel, wilt thou not hearken unto me?
JER|38|16|So Zedekiah the king sware secretly unto Jeremiah, saying, As the LORD liveth, that made us this soul, I will not put thee to death, neither will I give thee into the hand of these men that seek thy life.
JER|38|17|Then said Jeremiah unto Zedekiah, Thus saith the LORD, the God of hosts, the God of Israel; If thou wilt assuredly go forth unto the king of Babylon's princes, then thy soul shall live, and this city shall not be burned with fire; and thou shalt live, and thine house:
JER|38|18|But if thou wilt not go forth to the king of Babylon's princes, then shall this city be given into the hand of the Chaldeans, and they shall burn it with fire, and thou shalt not escape out of their hand.
JER|38|19|And Zedekiah the king said unto Jeremiah, I am afraid of the Jews that are fallen to the Chaldeans, lest they deliver me into their hand, and they mock me.
JER|38|20|But Jeremiah said, They shall not deliver thee. Obey, I beseech thee, the voice of the LORD, which I speak unto thee: so it shall be well unto thee, and thy soul shall live.
JER|38|21|But if thou refuse to go forth, this is the word that the LORD hath shewed me:
JER|38|22|And, behold, all the women that are left in the king of Judah's house shall be brought forth to the king of Babylon's princes, and those women shall say, Thy friends have set thee on, and have prevailed against thee: thy feet are sunk in the mire, and they are turned away back.
JER|38|23|So they shall bring out all thy wives and thy children to the Chaldeans: and thou shalt not escape out of their hand, but shalt be taken by the hand of the king of Babylon: and thou shalt cause this city to be burned with fire.
JER|38|24|Then said Zedekiah unto Jeremiah, Let no man know of these words, and thou shalt not die.
JER|38|25|But if the princes hear that I have talked with thee, and they come unto thee, and say unto thee, Declare unto us now what thou hast said unto the king, hide it not from us, and we will not put thee to death; also what the king said unto thee:
JER|38|26|Then thou shalt say unto them, I presented my supplication before the king, that he would not cause me to return to Jonathan's house, to die there.
JER|38|27|Then came all the princes unto Jeremiah, and asked him: and he told them according to all these words that the king had commanded. So they left off speaking with him; for the matter was not perceived.
JER|38|28|So Jeremiah abode in the court of the prison until the day that Jerusalem was taken: and he was there when Jerusalem was taken.
JER|39|1|In the ninth year of Zedekiah king of Judah, in the tenth month, came Nebuchadrezzar king of Babylon and all his army against Jerusalem, and they besieged it.
JER|39|2|And in the eleventh year of Zedekiah, in the fourth month, the ninth day of the month, the city was broken up.
JER|39|3|And all the princes of the king of Babylon came in, and sat in the middle gate, even Nergalsharezer, Samgarnebo, Sarsechim, Rabsaris, Nergalsharezer, Rabmag, with all the residue of the princes of the king of Babylon.
JER|39|4|And it came to pass, that when Zedekiah the king of Judah saw them, and all the men of war, then they fled, and went forth out of the city by night, by the way of the king's garden, by the gate betwixt the two walls: and he went out the way of the plain.
JER|39|5|But the Chaldeans' army pursued after them, and overtook Zedekiah in the plains of Jericho: and when they had taken him, they brought him up to Nebuchadnezzar king of Babylon to Riblah in the land of Hamath, where he gave judgment upon him.
JER|39|6|Then the king of Babylon slew the sons of Zedekiah in Riblah before his eyes: also the king of Babylon slew all the nobles of Judah.
JER|39|7|Moreover he put out Zedekiah's eyes, and bound him with chains, to carry him to Babylon.
JER|39|8|And the Chaldeans burned the king's house, and the houses of the people, with fire, and brake down the walls of Jerusalem.
JER|39|9|Then Nebuzaradan the captain of the guard carried away captive into Babylon the remnant of the people that remained in the city, and those that fell away, that fell to him, with the rest of the people that remained.
JER|39|10|But Nebuzaradan the captain of the guard left of the poor of the people, which had nothing, in the land of Judah, and gave them vineyards and fields at the same time.
JER|39|11|Now Nebuchadrezzar king of Babylon gave charge concerning Jeremiah to Nebuzaradan the captain of the guard, saying,
JER|39|12|Take him, and look well to him, and do him no harm; but do unto him even as he shall say unto thee.
JER|39|13|So Nebuzaradan the captain of the guard sent, and Nebushasban, Rabsaris, and Nergalsharezer, Rabmag, and all the king of Babylon's princes;
JER|39|14|Even they sent, and took Jeremiah out of the court of the prison, and committed him unto Gedaliah the son of Ahikam the son of Shaphan, that he should carry him home: so he dwelt among the people.
JER|39|15|Now the word of the LORD came unto Jeremiah, while he was shut up in the court of the prison, saying,
JER|39|16|Go and speak to Ebedmelech the Ethiopian, saying, Thus saith the LORD of hosts, the God of Israel; Behold, I will bring my words upon this city for evil, and not for good; and they shall be accomplished in that day before thee.
JER|39|17|But I will deliver thee in that day, saith the LORD: and thou shalt not be given into the hand of the men of whom thou art afraid.
JER|39|18|For I will surely deliver thee, and thou shalt not fall by the sword, but thy life shall be for a prey unto thee: because thou hast put thy trust in me, saith the LORD.
JER|40|1|The word that came to Jeremiah from the LORD, after that Nebuzaradan the captain of the guard had let him go from Ramah, when he had taken him being bound in chains among all that were carried away captive of Jerusalem and Judah, which were carried away captive unto Babylon.
JER|40|2|And the captain of the guard took Jeremiah, and said unto him, The LORD thy God hath pronounced this evil upon this place.
JER|40|3|Now the LORD hath brought it, and done according as he hath said: because ye have sinned against the LORD, and have not obeyed his voice, therefore this thing is come upon you.
JER|40|4|And now, behold, I loose thee this day from the chains which were upon thine hand. If it seem good unto thee to come with me into Babylon, come; and I will look well unto thee: but if it seem ill unto thee to come with me into Babylon, forbear: behold, all the land is before thee: whither it seemeth good and convenient for thee to go, thither go.
JER|40|5|Now while he was not yet gone back, he said, Go back also to Gedaliah the son of Ahikam the son of Shaphan, whom the king of Babylon hath made governor over the cities of Judah, and dwell with him among the people: or go wheresoever it seemeth convenient unto thee to go. So the captain of the guard gave him victuals and a reward, and let him go.
JER|40|6|Then went Jeremiah unto Gedaliah the son of Ahikam to Mizpah; and dwelt with him among the people that were left in the land.
JER|40|7|Now when all the captains of the forces which were in the fields, even they and their men, heard that the king of Babylon had made Gedaliah the son of Ahikam governor in the land, and had committed unto him men, and women, and children, and of the poor of the land, of them that were not carried away captive to Babylon;
JER|40|8|Then they came to Gedaliah to Mizpah, even Ishmael the son of Nethaniah, and Johanan and Jonathan the sons of Kareah, and Seraiah the son of Tanhumeth, and the sons of Ephai the Netophathite, and Jezaniah the son of a Maachathite, they and their men.
JER|40|9|And Gedaliah the son of Ahikam the son of Shaphan sware unto them and to their men, saying, Fear not to serve the Chaldeans: dwell in the land, and serve the king of Babylon, and it shall be well with you.
JER|40|10|As for me, behold, I will dwell at Mizpah, to serve the Chaldeans, which will come unto us: but ye, gather ye wine, and summer fruits, and oil, and put them in your vessels, and dwell in your cities that ye have taken.
JER|40|11|Likewise when all the Jews that were in Moab, and among the Ammonites, and in Edom, and that were in all the countries, heard that the king of Babylon had left a remnant of Judah, and that he had set over them Gedaliah the son of Ahikam the son of Shaphan;
JER|40|12|Even all the Jews returned out of all places whither they were driven, and came to the land of Judah, to Gedaliah, unto Mizpah, and gathered wine and summer fruits very much.
JER|40|13|Moreover Johanan the son of Kareah, and all the captains of the forces that were in the fields, came to Gedaliah to Mizpah,
JER|40|14|And said unto him, Dost thou certainly know that Baalis the king of the Ammonites hath sent Ishmael the son of Nethaniah to slay thee? But Gedaliah the son of Ahikam believed them not.
JER|40|15|Then Johanan the son of Kareah spake to Gedaliah in Mizpah secretly saying, Let me go, I pray thee, and I will slay Ishmael the son of Nethaniah, and no man shall know it: wherefore should he slay thee, that all the Jews which are gathered unto thee should be scattered, and the remnant in Judah perish?
JER|40|16|But Gedaliah the son of Ahikam said unto Johanan the son of Kareah, Thou shalt not do this thing: for thou speakest falsely of Ishmael.
JER|41|1|Now it came to pass in the seventh month, that Ishmael the son of Nethaniah the son of Elishama, of the seed royal, and the princes of the king, even ten men with him, came unto Gedaliah the son of Ahikam to Mizpah; and there they did eat bread together in Mizpah.
JER|41|2|Then arose Ishmael the son of Nethaniah, and the ten men that were with him, and smote Gedaliah the son of Ahikam the son of Shaphan with the sword, and slew him, whom the king of Babylon had made governor over the land.
JER|41|3|Ishmael also slew all the Jews that were with him, even with Gedaliah, at Mizpah, and the Chaldeans that were found there, and the men of war.
JER|41|4|And it came to pass the second day after he had slain Gedaliah, and no man knew it,
JER|41|5|That there came certain from Shechem, from Shiloh, and from Samaria, even fourscore men, having their beards shaven, and their clothes rent, and having cut themselves, with offerings and incense in their hand, to bring them to the house of the LORD.
JER|41|6|And Ishmael the son of Nethaniah went forth from Mizpah to meet them, weeping all along as he went: and it came to pass, as he met them, he said unto them, Come to Gedaliah the son of Ahikam.
JER|41|7|And it was so, when they came into the midst of the city, that Ishmael the son of Nethaniah slew them, and cast them into the midst of the pit, he, and the men that were with him.
JER|41|8|But ten men were found among them that said unto Ishmael, Slay us not: for we have treasures in the field, of wheat, and of barley, and of oil, and of honey. So he forbare, and slew them not among their brethren.
JER|41|9|Now the pit wherein Ishmael had cast all the dead bodies of the men, whom he had slain because of Gedaliah, was it which Asa the king had made for fear of Baasha king of Israel: and Ishmael the son of Nethaniah filled it with them that were slain.
JER|41|10|Then Ishmael carried away captive all the residue of the people that were in Mizpah, even the king's daughters, and all the people that remained in Mizpah, whom Nebuzaradan the captain of the guard had committed to Gedaliah the son of Ahikam: and Ishmael the son of Nethaniah carried them away captive, and departed to go over to the Ammonites.
JER|41|11|But when Johanan the son of Kareah, and all the captains of the forces that were with him, heard of all the evil that Ishmael the son of Nethaniah had done,
JER|41|12|Then they took all the men, and went to fight with Ishmael the son of Nethaniah, and found him by the great waters that are in Gibeon.
JER|41|13|Now it came to pass, that when all the people which were with Ishmael saw Johanan the son of Kareah, and all the captains of the forces that were with him, then they were glad.
JER|41|14|So all the people that Ishmael had carried away captive from Mizpah cast about and returned, and went unto Johanan the son of Kareah.
JER|41|15|But Ishmael the son of Nethaniah escaped from Johanan with eight men, and went to the Ammonites.
JER|41|16|Then took Johanan the son of Kareah, and all the captains of the forces that were with him, all the remnant of the people whom he had recovered from Ishmael the son of Nethaniah, from Mizpah, after that he had slain Gedaliah the son of Ahikam, even mighty men of war, and the women, and the children, and the eunuchs, whom he had brought again from Gibeon:
JER|41|17|And they departed, and dwelt in the habitation of Chimham, which is by Bethlehem, to go to enter into Egypt,
JER|41|18|Because of the Chaldeans: for they were afraid of them, because Ishmael the son of Nethaniah had slain Gedaliah the son of Ahikam, whom the king of Babylon made governor in the land.
JER|42|1|Then all the captains of the forces, and Johanan the son of Kareah, and Jezaniah the son of Hoshaiah, and all the people from the least even unto the greatest, came near,
JER|42|2|And said unto Jeremiah the prophet, Let, we beseech thee, our supplication be accepted before thee, and pray for us unto the LORD thy God, even for all this remnant; (for we are left but a few of many, as thine eyes do behold us:)
JER|42|3|That the LORD thy God may shew us the way wherein we may walk, and the thing that we may do.
JER|42|4|Then Jeremiah the prophet said unto them, I have heard you; behold, I will pray unto the LORD your God according to your words; and it shall come to pass, that whatsoever thing the LORD shall answer you, I will declare it unto you; I will keep nothing back from you.
JER|42|5|Then they said to Jeremiah, The LORD be a true and faithful witness between us, if we do not even according to all things for the which the LORD thy God shall send thee to us.
JER|42|6|Whether it be good, or whether it be evil, we will obey the voice of the LORD our God, to whom we send thee; that it may be well with us, when we obey the voice of the LORD our God.
JER|42|7|And it came to pass after ten days, that the word of the LORD came unto Jeremiah.
JER|42|8|Then called he Johanan the son of Kareah, and all the captains of the forces which were with him, and all the people from the least even to the greatest,
JER|42|9|And said unto them, Thus saith the LORD, the God of Israel, unto whom ye sent me to present your supplication before him;
JER|42|10|If ye will still abide in this land, then will I build you, and not pull you down, and I will plant you, and not pluck you up: for I repent me of the evil that I have done unto you.
JER|42|11|Be not afraid of the king of Babylon, of whom ye are afraid; be not afraid of him, saith the LORD: for I am with you to save you, and to deliver you from his hand.
JER|42|12|And I will shew mercies unto you, that he may have mercy upon you, and cause you to return to your own land.
JER|42|13|But if ye say, We will not dwell in this land, neither obey the voice of the LORD your God,
JER|42|14|Saying, No; but we will go into the land of Egypt, where we shall see no war, nor hear the sound of the trumpet, nor have hunger of bread; and there will we dwell:
JER|42|15|And now therefore hear the word of the LORD, ye remnant of Judah; Thus saith the LORD of hosts, the God of Israel; If ye wholly set your faces to enter into Egypt, and go to sojourn there;
JER|42|16|Then it shall come to pass, that the sword, which ye feared, shall overtake you there in the land of Egypt, and the famine, whereof ye were afraid, shall follow close after you there in Egypt; and there ye shall die.
JER|42|17|So shall it be with all the men that set their faces to go into Egypt to sojourn there; they shall die by the sword, by the famine, and by the pestilence: and none of them shall remain or escape from the evil that I will bring upon them.
JER|42|18|For thus saith the LORD of hosts, the God of Israel; As mine anger and my fury hath been poured forth upon the inhabitants of Jerusalem; so shall my fury be poured forth upon you, when ye shall enter into Egypt: and ye shall be an execration, and an astonishment, and a curse, and a reproach; and ye shall see this place no more.
JER|42|19|The LORD hath said concerning you, O ye remnant of Judah; Go ye not into Egypt: know certainly that I have admonished you this day.
JER|42|20|For ye dissembled in your hearts, when ye sent me unto the LORD your God, saying, Pray for us unto the LORD our God; and according unto all that the LORD our God shall say, so declare unto us, and we will do it.
JER|42|21|And now I have this day declared it to you; but ye have not obeyed the voice of the LORD your God, nor any thing for the which he hath sent me unto you.
JER|42|22|Now therefore know certainly that ye shall die by the sword, by the famine, and by the pestilence, in the place whither ye desire to go and to sojourn.
JER|43|1|And it came to pass, that when Jeremiah had made an end of speaking unto all the people all the words of the LORD their God, for which the LORD their God had sent him to them, even all these words,
JER|43|2|Then spake Azariah the son of Hoshaiah, and Johanan the son of Kareah, and all the proud men, saying unto Jeremiah, Thou speakest falsely: the LORD our God hath not sent thee to say, Go not into Egypt to sojourn there:
JER|43|3|But Baruch the son of Neriah setteth thee on against us, for to deliver us into the hand of the Chaldeans, that they might put us to death, and carry us away captives into Babylon.
JER|43|4|So Johanan the son of Kareah, and all the captains of the forces, and all the people, obeyed not the voice of the LORD, to dwell in the land of Judah.
JER|43|5|But Johanan the son of Kareah, and all the captains of the forces, took all the remnant of Judah, that were returned from all nations, whither they had been driven, to dwell in the land of Judah;
JER|43|6|Even men, and women, and children, and the king's daughters, and every person that Nebuzaradan the captain of the guard had left with Gedaliah the son of Ahikam the son of Shaphan, and Jeremiah the prophet, and Baruch the son of Neriah.
JER|43|7|So they came into the land of Egypt: for they obeyed not the voice of the LORD: thus came they even to Tahpanhes.
JER|43|8|Then came the word of the LORD unto Jeremiah in Tahpanhes, saying,
JER|43|9|Take great stones in thine hand, and hide them in the clay in the brickkiln, which is at the entry of Pharaoh's house in Tahpanhes, in the sight of the men of Judah;
JER|43|10|And say unto them, Thus saith the LORD of hosts, the God of Israel; Behold, I will send and take Nebuchadrezzar the king of Babylon, my servant, and will set his throne upon these stones that I have hid; and he shall spread his royal pavilion over them.
JER|43|11|And when he cometh, he shall smite the land of Egypt, and deliver such as are for death to death; and such as are for captivity to captivity; and such as are for the sword to the sword.
JER|43|12|And I will kindle a fire in the houses of the gods of Egypt; and he shall burn them, and carry them away captives: and he shall array himself with the land of Egypt, as a shepherd putteth on his garment; and he shall go forth from thence in peace.
JER|43|13|He shall break also the images of Bethshemesh, that is in the land of Egypt; and the houses of the gods of the Egyptians shall he burn with fire.
JER|44|1|The word that came to Jeremiah concerning all the Jews which dwell in the land of Egypt, which dwell at Migdol, and at Tahpanhes, and at Noph, and in the country of Pathros, saying,
JER|44|2|Thus saith the LORD of hosts, the God of Israel; Ye have seen all the evil that I have brought upon Jerusalem, and upon all the cities of Judah; and, behold, this day they are a desolation, and no man dwelleth therein,
JER|44|3|Because of their wickedness which they have committed to provoke me to anger, in that they went to burn incense, and to serve other gods, whom they knew not, neither they, ye, nor your fathers.
JER|44|4|Howbeit I sent unto you all my servants the prophets, rising early and sending them, saying, Oh, do not this abominable thing that I hate.
JER|44|5|But they hearkened not, nor inclined their ear to turn from their wickedness, to burn no incense unto other gods.
JER|44|6|Wherefore my fury and mine anger was poured forth, and was kindled in the cities of Judah and in the streets of Jerusalem; and they are wasted and desolate, as at this day.
JER|44|7|Therefore now thus saith the LORD, the God of hosts, the God of Israel; Wherefore commit ye this great evil against your souls, to cut off from you man and woman, child and suckling, out of Judah, to leave you none to remain;
JER|44|8|In that ye provoke me unto wrath with the works of your hands, burning incense unto other gods in the land of Egypt, whither ye be gone to dwell, that ye might cut yourselves off, and that ye might be a curse and a reproach among all the nations of the earth?
JER|44|9|Have ye forgotten the wickedness of your fathers, and the wickedness of the kings of Judah, and the wickedness of their wives, and your own wickedness, and the wickedness of your wives, which they have committed in the land of Judah, and in the streets of Jerusalem?
JER|44|10|They are not humbled even unto this day, neither have they feared, nor walked in my law, nor in my statutes, that I set before you and before your fathers.
JER|44|11|Therefore thus saith the LORD of hosts, the God of Israel; Behold, I will set my face against you for evil, and to cut off all Judah.
JER|44|12|And I will take the remnant of Judah, that have set their faces to go into the land of Egypt to sojourn there, and they shall all be consumed, and fall in the land of Egypt; they shall even be consumed by the sword and by the famine: they shall die, from the least even unto the greatest, by the sword and by the famine: and they shall be an execration, and an astonishment, and a curse, and a reproach.
JER|44|13|For I will punish them that dwell in the land of Egypt, as I have punished Jerusalem, by the sword, by the famine, and by the pestilence:
JER|44|14|So that none of the remnant of Judah, which are gone into the land of Egypt to sojourn there, shall escape or remain, that they should return into the land of Judah, to the which they have a desire to return to dwell there: for none shall return but such as shall escape.
JER|44|15|Then all the men which knew that their wives had burned incense unto other gods, and all the women that stood by, a great multitude, even all the people that dwelt in the land of Egypt, in Pathros, answered Jeremiah, saying,
JER|44|16|As for the word that thou hast spoken unto us in the name of the LORD, we will not hearken unto thee.
JER|44|17|But we will certainly do whatsoever thing goeth forth out of our own mouth, to burn incense unto the queen of heaven, and to pour out drink offerings unto her, as we have done, we, and our fathers, our kings, and our princes, in the cities of Judah, and in the streets of Jerusalem: for then had we plenty of victuals, and were well, and saw no evil.
JER|44|18|But since we left off to burn incense to the queen of heaven, and to pour out drink offerings unto her, we have wanted all things, and have been consumed by the sword and by the famine.
JER|44|19|And when we burned incense to the queen of heaven, and poured out drink offerings unto her, did we make her cakes to worship her, and pour out drink offerings unto her, without our men?
JER|44|20|Then Jeremiah said unto all the people, to the men, and to the women, and to all the people which had given him that answer, saying,
JER|44|21|The incense that ye burned in the cities of Judah, and in the streets of Jerusalem, ye, and your fathers, your kings, and your princes, and the people of the land, did not the LORD remember them, and came it not into his mind?
JER|44|22|So that the LORD could no longer bear, because of the evil of your doings, and because of the abominations which ye have committed; therefore is your land a desolation, and an astonishment, and a curse, without an inhabitant, as at this day.
JER|44|23|Because ye have burned incense, and because ye have sinned against the LORD, and have not obeyed the voice of the LORD, nor walked in his law, nor in his statutes, nor in his testimonies; therefore this evil is happened unto you, as at this day.
JER|44|24|Moreover Jeremiah said unto all the people, and to all the women, Hear the word of the LORD, all Judah that are in the land of Egypt:
JER|44|25|Thus saith the LORD of hosts, the God of Israel, saying; Ye and your wives have both spoken with your mouths, and fulfilled with your hand, saying, We will surely perform our vows that we have vowed, to burn incense to the queen of heaven, and to pour out drink offerings unto her: ye will surely accomplish your vows, and surely perform your vows.
JER|44|26|Therefore hear ye the word of the LORD, all Judah that dwell in the land of Egypt; Behold, I have sworn by my great name, saith the LORD, that my name shall no more be named in the mouth of any man of Judah in all the land of Egypt, saying, The Lord GOD liveth.
JER|44|27|Behold, I will watch over them for evil, and not for good: and all the men of Judah that are in the land of Egypt shall be consumed by the sword and by the famine, until there be an end of them.
JER|44|28|Yet a small number that escape the sword shall return out of the land of Egypt into the land of Judah, and all the remnant of Judah, that are gone into the land of Egypt to sojourn there, shall know whose words shall stand, mine, or their's.
JER|44|29|And this shall be a sign unto you, saith the LORD, that I will punish you in this place, that ye may know that my words shall surely stand against you for evil:
JER|44|30|Thus saith the LORD; Behold, I will give Pharaohhophra king of Egypt into the hand of his enemies, and into the hand of them that seek his life; as I gave Zedekiah king of Judah into the hand of Nebuchadrezzar king of Babylon, his enemy, and that sought his life.
JER|45|1|The word that Jeremiah the prophet spake unto Baruch the son of Neriah, when he had written these words in a book at the mouth of Jeremiah, in the fourth year of Jehoiakim the son of Josiah king of Judah, saying,
JER|45|2|Thus saith the LORD, the God of Israel, unto thee, O Baruch:
JER|45|3|Thou didst say, Woe is me now! for the LORD hath added grief to my sorrow; I fainted in my sighing, and I find no rest.
JER|45|4|Thus shalt thou say unto him, The LORD saith thus; Behold, that which I have built will I break down, and that which I have planted I will pluck up, even this whole land.
JER|45|5|And seekest thou great things for thyself? seek them not: for, behold, I will bring evil upon all flesh, saith the LORD: but thy life will I give unto thee for a prey in all places whither thou goest.
JER|46|1|The word of the LORD which came to Jeremiah the prophet against the Gentiles;
JER|46|2|Against Egypt, against the army of Pharaohnecho king of Egypt, which was by the river Euphrates in Carchemish, which Nebuchadrezzar king of Babylon smote in the fourth year of Jehoiakim the son of Josiah king of Judah.
JER|46|3|Order ye the buckler and shield, and draw near to battle.
JER|46|4|Harness the horses; and get up, ye horsemen, and stand forth with your helmets; furbish the spears, and put on the brigandines.
JER|46|5|Wherefore have I seen them dismayed and turned away back? and their mighty ones are beaten down, and are fled apace, and look not back: for fear was round about, saith the LORD.
JER|46|6|Let not the swift flee away, nor the mighty man escape; they shall stumble, and fall toward the north by the river Euphrates.
JER|46|7|Who is this that cometh up as a flood, whose waters are moved as the rivers?
JER|46|8|Egypt riseth up like a flood, and his waters are moved like the rivers; and he saith, I will go up, and will cover the earth; I will destroy the city and the inhabitants thereof.
JER|46|9|Come up, ye horses; and rage, ye chariots; and let the mighty men come forth; the Ethiopians and the Libyans, that handle the shield; and the Lydians, that handle and bend the bow.
JER|46|10|For this is the day of the Lord GOD of hosts, a day of vengeance, that he may avenge him of his adversaries: and the sword shall devour, and it shall be satiate and made drunk with their blood: for the Lord GOD of hosts hath a sacrifice in the north country by the river Euphrates.
JER|46|11|Go up into Gilead, and take balm, O virgin, the daughter of Egypt: in vain shalt thou use many medicines; for thou shalt not be cured.
JER|46|12|The nations have heard of thy shame, and thy cry hath filled the land: for the mighty man hath stumbled against the mighty, and they are fallen both together.
JER|46|13|The word that the LORD spake to Jeremiah the prophet, how Nebuchadrezzar king of Babylon should come and smite the land of Egypt.
JER|46|14|Declare ye in Egypt, and publish in Migdol, and publish in Noph and in Tahpanhes: say ye, Stand fast, and prepare thee; for the sword shall devour round about thee.
JER|46|15|Why are thy valiant men swept away? they stood not, because the LORD did drive them.
JER|46|16|He made many to fall, yea, one fell upon another: and they said, Arise, and let us go again to our own people, and to the land of our nativity, from the oppressing sword.
JER|46|17|They did cry there, Pharaoh king of Egypt is but a noise; he hath passed the time appointed.
JER|46|18|As I live, saith the King, whose name is the LORD of hosts, Surely as Tabor is among the mountains, and as Carmel by the sea, so shall he come.
JER|46|19|O thou daughter dwelling in Egypt, furnish thyself to go into captivity: for Noph shall be waste and desolate without an inhabitant.
JER|46|20|Egypt is like a very fair heifer, but destruction cometh; it cometh out of the north.
JER|46|21|Also her hired men are in the midst of her like fatted bullocks; for they also are turned back, and are fled away together: they did not stand, because the day of their calamity was come upon them, and the time of their visitation.
JER|46|22|The voice thereof shall go like a serpent; for they shall march with an army, and come against her with axes, as hewers of wood.
JER|46|23|They shall cut down her forest, saith the LORD, though it cannot be searched; because they are more than the grasshoppers, and are innumerable.
JER|46|24|The daughter of Egypt shall be confounded; she shall be delivered into the hand of the people of the north.
JER|46|25|The LORD of hosts, the God of Israel, saith; Behold, I will punish the multitude of No, and Pharaoh, and Egypt, with their gods, and their kings; even Pharaoh, and all them that trust in him:
JER|46|26|And I will deliver them into the hand of those that seek their lives, and into the hand of Nebuchadrezzar king of Babylon, and into the hand of his servants: and afterward it shall be inhabited, as in the days of old, saith the LORD.
JER|46|27|But fear not thou, O my servant Jacob, and be not dismayed, O Israel: for, behold, I will save thee from afar off, and thy seed from the land of their captivity; and Jacob shall return, and be in rest and at ease, and none shall make him afraid.
JER|46|28|Fear thou not, O Jacob my servant, saith the LORD: for I am with thee; for I will make a full end of all the nations whither I have driven thee: but I will not make a full end of thee, but correct thee in measure; yet will I not leave thee wholly unpunished.
JER|47|1|The word of the LORD that came to Jeremiah the prophet against the Philistines, before that Pharaoh smote Gaza.
JER|47|2|Thus saith the LORD; Behold, waters rise up out of the north, and shall be an overflowing flood, and shall overflow the land, and all that is therein; the city, and them that dwell therein: then the men shall cry, and all the inhabitants of the land shall howl.
JER|47|3|At the noise of the stamping of the hoofs of his strong horses, at the rushing of his chariots, and at the rumbling of his wheels, the fathers shall not look back to their children for feebleness of hands;
JER|47|4|Because of the day that cometh to spoil all the Philistines, and to cut off from Tyrus and Zidon every helper that remaineth: for the LORD will spoil the Philistines, the remnant of the country of Caphtor.
JER|47|5|Baldness is come upon Gaza; Ashkelon is cut off with the remnant of their valley: how long wilt thou cut thyself?
JER|47|6|O thou sword of the LORD, how long will it be ere thou be quiet? put up thyself into thy scabbard, rest, and be still.
JER|47|7|How can it be quiet, seeing the LORD hath given it a charge against Ashkelon, and against the sea shore? there hath he appointed it.
JER|48|1|Against Moab thus saith the LORD of hosts, the God of Israel; Woe unto Nebo! for it is spoiled: Kiriathaim is confounded and taken: Misgab is confounded and dismayed.
JER|48|2|There shall be no more praise of Moab: in Heshbon they have devised evil against it; come, and let us cut it off from being a nation. Also thou shalt be cut down, O Madmen; the sword shall pursue thee.
JER|48|3|A voice of crying shall be from Horonaim, spoiling and great destruction.
JER|48|4|Moab is destroyed; her little ones have caused a cry to be heard.
JER|48|5|For in the going up of Luhith continual weeping shall go up; for in the going down of Horonaim the enemies have heard a cry of destruction.
JER|48|6|Flee, save your lives, and be like the heath in the wilderness.
JER|48|7|For because thou hast trusted in thy works and in thy treasures, thou shalt also be taken: and Chemosh shall go forth into captivity with his priests and his princes together.
JER|48|8|And the spoiler shall come upon every city, and no city shall escape: the valley also shall perish, and the plain shall be destroyed, as the LORD hath spoken.
JER|48|9|Give wings unto Moab, that it may flee and get away: for the cities thereof shall be desolate, without any to dwell therein.
JER|48|10|Cursed be he that doeth the work of the LORD deceitfully, and cursed be he that keepeth back his sword from blood.
JER|48|11|Moab hath been at ease from his youth, and he hath settled on his lees, and hath not been emptied from vessel to vessel, neither hath he gone into captivity: therefore his taste remained in him, and his scent is not changed.
JER|48|12|Therefore, behold, the days come, saith the LORD, that I will send unto him wanderers, that shall cause him to wander, and shall empty his vessels, and break their bottles.
JER|48|13|And Moab shall be ashamed of Chemosh, as the house of Israel was ashamed of Bethel their confidence.
JER|48|14|How say ye, We are mighty and strong men for the war?
JER|48|15|Moab is spoiled, and gone up out of her cities, and his chosen young men are gone down to the slaughter, saith the King, whose name is the LORD of hosts.
JER|48|16|The calamity of Moab is near to come, and his affliction hasteth fast.
JER|48|17|All ye that are about him, bemoan him; and all ye that know his name, say, How is the strong staff broken, and the beautiful rod!
JER|48|18|Thou daughter that dost inhabit Dibon, come down from thy glory, and sit in thirst; for the spoiler of Moab shall come upon thee, and he shall destroy thy strong holds.
JER|48|19|O inhabitant of Aroer, stand by the way, and espy; ask him that fleeth, and her that escapeth, and say, What is done?
JER|48|20|Moab is confounded; for it is broken down: howl and cry; tell ye it in Arnon, that Moab is spoiled,
JER|48|21|And judgment is come upon the plain country; upon Holon, and upon Jahazah, and upon Mephaath,
JER|48|22|And upon Dibon, and upon Nebo, and upon Bethdiblathaim,
JER|48|23|And upon Kiriathaim, and upon Bethgamul, and upon Bethmeon,
JER|48|24|And upon Kerioth, and upon Bozrah, and upon all the cities of the land of Moab, far or near.
JER|48|25|The horn of Moab is cut off, and his arm is broken, saith the LORD.
JER|48|26|Make ye him drunken: for he magnified himself against the LORD: Moab also shall wallow in his vomit, and he also shall be in derision.
JER|48|27|For was not Israel a derision unto thee? was he found among thieves? for since thou spakest of him, thou skippedst for joy.
JER|48|28|O ye that dwell in Moab, leave the cities, and dwell in the rock, and be like the dove that maketh her nest in the sides of the hole's mouth.
JER|48|29|We have heard the pride of Moab, (he is exceeding proud) his loftiness, and his arrogancy, and his pride, and the haughtiness of his heart.
JER|48|30|I know his wrath, saith the LORD; but it shall not be so; his lies shall not so effect it.
JER|48|31|Therefore will I howl for Moab, and I will cry out for all Moab; mine heart shall mourn for the men of Kirheres.
JER|48|32|O vine of Sibmah, I will weep for thee with the weeping of Jazer: thy plants are gone over the sea, they reach even to the sea of Jazer: the spoiler is fallen upon thy summer fruits and upon thy vintage.
JER|48|33|And joy and gladness is taken from the plentiful field, and from the land of Moab, and I have caused wine to fail from the winepresses: none shall tread with shouting; their shouting shall be no shouting.
JER|48|34|From the cry of Heshbon even unto Elealeh, and even unto Jahaz, have they uttered their voice, from Zoar even unto Horonaim, as an heifer of three years old: for the waters also of Nimrim shall be desolate.
JER|48|35|Moreover I will cause to cease in Moab, saith the LORD, him that offereth in the high places, and him that burneth incense to his gods.
JER|48|36|Therefore mine heart shall sound for Moab like pipes, and mine heart shall sound like pipes for the men of Kirheres: because the riches that he hath gotten are perished.
JER|48|37|For every head shall be bald, and every beard clipped: upon all the hands shall be cuttings, and upon the loins sackcloth.
JER|48|38|There shall be lamentation generally upon all the housetops of Moab, and in the streets thereof: for I have broken Moab like a vessel wherein is no pleasure, saith the LORD.
JER|48|39|They shall howl, saying, How is it broken down! how hath Moab turned the back with shame! so shall Moab be a derision and a dismaying to all them about him.
JER|48|40|For thus saith the LORD; Behold, he shall fly as an eagle, and shall spread his wings over Moab.
JER|48|41|Kerioth is taken, and the strong holds are surprised, and the mighty men's hearts in Moab at that day shall be as the heart of a woman in her pangs.
JER|48|42|And Moab shall be destroyed from being a people, because he hath magnified himself against the LORD.
JER|48|43|Fear, and the pit, and the snare, shall be upon thee, O inhabitant of Moab, saith the LORD.
JER|48|44|He that fleeth from the fear shall fall into the pit; and he that getteth up out of the pit shall be taken in the snare: for I will bring upon it, even upon Moab, the year of their visitation, saith the LORD.
JER|48|45|They that fled stood under the shadow of Heshbon because of the force: but a fire shall come forth out of Heshbon, and a flame from the midst of Sihon, and shall devour the corner of Moab, and the crown of the head of the tumultuous ones.
JER|48|46|Woe be unto thee, O Moab! the people of Chemosh perisheth: for thy sons are taken captives, and thy daughters captives.
JER|48|47|Yet will I bring again the captivity of Moab in the latter days, saith the LORD. Thus far is the judgment of Moab.
JER|49|1|Concerning the Ammonites, thus saith the LORD; Hath Israel no sons? hath he no heir? why then doth their king inherit Gad, and his people dwell in his cities?
JER|49|2|Therefore, behold, the days come, saith the LORD, that I will cause an alarm of war to be heard in Rabbah of the Ammonites; and it shall be a desolate heap, and her daughters shall be burned with fire: then shall Israel be heir unto them that were his heirs, saith the LORD.
JER|49|3|Howl, O Heshbon, for Ai is spoiled: cry, ye daughters of Rabbah, gird you with sackcloth; lament, and run to and fro by the hedges; for their king shall go into captivity, and his priests and his princes together.
JER|49|4|Wherefore gloriest thou in the valleys, thy flowing valley, O backsliding daughter? that trusted in her treasures, saying, Who shall come unto me?
JER|49|5|Behold, I will bring a fear upon thee, saith the Lord GOD of hosts, from all those that be about thee; and ye shall be driven out every man right forth; and none shall gather up him that wandereth.
JER|49|6|And afterward I will bring again the captivity of the children of Ammon, saith the LORD.
JER|49|7|Concerning Edom, thus saith the LORD of hosts; Is wisdom no more in Teman? is counsel perished from the prudent? is their wisdom vanished?
JER|49|8|Flee ye, turn back, dwell deep, O inhabitants of Dedan; for I will bring the calamity of Esau upon him, the time that I will visit him.
JER|49|9|If grapegatherers come to thee, would they not leave some gleaning grapes? if thieves by night, they will destroy till they have enough.
JER|49|10|But I have made Esau bare, I have uncovered his secret places, and he shall not be able to hide himself: his seed is spoiled, and his brethren, and his neighbours, and he is not.
JER|49|11|Leave thy fatherless children, I will preserve them alive; and let thy widows trust in me.
JER|49|12|For thus saith the LORD; Behold, they whose judgment was not to drink of the cup have assuredly drunken; and art thou he that shall altogether go unpunished? thou shalt not go unpunished, but thou shalt surely drink of it.
JER|49|13|For I have sworn by myself, saith the LORD, that Bozrah shall become a desolation, a reproach, a waste, and a curse; and all the cities thereof shall be perpetual wastes.
JER|49|14|I have heard a rumour from the LORD, and an ambassador is sent unto the heathen, saying, Gather ye together, and come against her, and rise up to the battle.
JER|49|15|For, lo, I will make thee small among the heathen, and despised among men.
JER|49|16|Thy terribleness hath deceived thee, and the pride of thine heart, O thou that dwellest in the clefts of the rock, that holdest the height of the hill: though thou shouldest make thy nest as high as the eagle, I will bring thee down from thence, saith the LORD.
JER|49|17|Also Edom shall be a desolation: every one that goeth by it shall be astonished, and shall hiss at all the plagues thereof.
JER|49|18|As in the overthrow of Sodom and Gomorrah and the neighbour cities thereof, saith the LORD, no man shall abide there, neither shall a son of man dwell in it.
JER|49|19|Behold, he shall come up like a lion from the swelling of Jordan against the habitation of the strong: but I will suddenly make him run away from her: and who is a chosen man, that I may appoint over her? for who is like me? and who will appoint me the time? and who is that shepherd that will stand before me?
JER|49|20|Therefore hear the counsel of the LORD, that he hath taken against Edom; and his purposes, that he hath purposed against the inhabitants of Teman: Surely the least of the flock shall draw them out: surely he shall make their habitations desolate with them.
JER|49|21|The earth is moved at the noise of their fall, at the cry the noise thereof was heard in the Red sea.
JER|49|22|Behold, he shall come up and fly as the eagle, and spread his wings over Bozrah: and at that day shall the heart of the mighty men of Edom be as the heart of a woman in her pangs.
JER|49|23|Concerning Damascus. Hamath is confounded, and Arpad: for they have heard evil tidings: they are fainthearted; there is sorrow on the sea; it cannot be quiet.
JER|49|24|Damascus is waxed feeble, and turneth herself to flee, and fear hath seized on her: anguish and sorrows have taken her, as a woman in travail.
JER|49|25|How is the city of praise not left, the city of my joy!
JER|49|26|Therefore her young men shall fall in her streets, and all the men of war shall be cut off in that day, saith the LORD of hosts.
JER|49|27|And I will kindle a fire in the wall of Damascus, and it shall consume the palaces of Benhadad.
JER|49|28|Concerning Kedar, and concerning the kingdoms of Hazor, which Nebuchadrezzar king of Babylon shall smite, thus saith the LORD; Arise ye, go up to Kedar, and spoil the men of the east.
JER|49|29|Their tents and their flocks shall they take away: they shall take to themselves their curtains, and all their vessels, and their camels; and they shall cry unto them, Fear is on every side.
JER|49|30|Flee, get you far off, dwell deep, O ye inhabitants of Hazor, saith the LORD; for Nebuchadrezzar king of Babylon hath taken counsel against you, and hath conceived a purpose against you.
JER|49|31|Arise, get you up unto the wealthy nation, that dwelleth without care, saith the LORD, which have neither gates nor bars, which dwell alone.
JER|49|32|And their camels shall be a booty, and the multitude of their cattle a spoil: and I will scatter into all winds them that are in the utmost corners; and I will bring their calamity from all sides thereof, saith the LORD.
JER|49|33|And Hazor shall be a dwelling for dragons, and a desolation for ever: there shall no man abide there, nor any son of man dwell in it.
JER|49|34|The word of the LORD that came to Jeremiah the prophet against Elam in the beginning of the reign of Zedekiah king of Judah, saying,
JER|49|35|Thus saith the LORD of hosts; Behold, I will break the bow of Elam, the chief of their might.
JER|49|36|And upon Elam will I bring the four winds from the four quarters of heaven, and will scatter them toward all those winds; and there shall be no nation whither the outcasts of Elam shall not come.
JER|49|37|For I will cause Elam to be dismayed before their enemies, and before them that seek their life: and I will bring evil upon them, even my fierce anger, saith the LORD; and I will send the sword after them, till I have consumed them:
JER|49|38|And I will set my throne in Elam, and will destroy from thence the king and the princes, saith the LORD.
JER|49|39|But it shall come to pass in the latter days, that I will bring again the captivity of Elam, saith the LORD.
JER|50|1|The word that the LORD spake against Babylon and against the land of the Chaldeans by Jeremiah the prophet.
JER|50|2|Declare ye among the nations, and publish, and set up a standard; publish, and conceal not: say, Babylon is taken, Bel is confounded, Merodach is broken in pieces; her idols are confounded, her images are broken in pieces.
JER|50|3|For out of the north there cometh up a nation against her, which shall make her land desolate, and none shall dwell therein: they shall remove, they shall depart, both man and beast.
JER|50|4|In those days, and in that time, saith the LORD, the children of Israel shall come, they and the children of Judah together, going and weeping: they shall go, and seek the LORD their God.
JER|50|5|They shall ask the way to Zion with their faces thitherward, saying, Come, and let us join ourselves to the LORD in a perpetual covenant that shall not be forgotten.
JER|50|6|My people hath been lost sheep: their shepherds have caused them to go astray, they have turned them away on the mountains: they have gone from mountain to hill, they have forgotten their restingplace.
JER|50|7|All that found them have devoured them: and their adversaries said, We offend not, because they have sinned against the LORD, the habitation of justice, even the LORD, the hope of their fathers.
JER|50|8|Remove out of the midst of Babylon, and go forth out of the land of the Chaldeans, and be as the he goats before the flocks.
JER|50|9|For, lo, I will raise and cause to come up against Babylon an assembly of great nations from the north country: and they shall set themselves in array against her; from thence she shall be taken: their arrows shall be as of a mighty expert man; none shall return in vain.
JER|50|10|And Chaldea shall be a spoil: all that spoil her shall be satisfied, saith the LORD.
JER|50|11|Because ye were glad, because ye rejoiced, O ye destroyers of mine heritage, because ye are grown fat as the heifer at grass, and bellow as bulls;
JER|50|12|Your mother shall be sore confounded; she that bare you shall be ashamed: behold, the hindermost of the nations shall be a wilderness, a dry land, and a desert.
JER|50|13|Because of the wrath of the LORD it shall not be inhabited, but it shall be wholly desolate: every one that goeth by Babylon shall be astonished, and hiss at all her plagues.
JER|50|14|Put yourselves in array against Babylon round about: all ye that bend the bow, shoot at her, spare no arrows: for she hath sinned against the LORD.
JER|50|15|Shout against her round about: she hath given her hand: her foundations are fallen, her walls are thrown down: for it is the vengeance of the LORD: take vengeance upon her; as she hath done, do unto her.
JER|50|16|Cut off the sower from Babylon, and him that handleth the sickle in the time of harvest: for fear of the oppressing sword they shall turn every one to his people, and they shall flee every one to his own land.
JER|50|17|Israel is a scattered sheep; the lions have driven him away: first the king of Assyria hath devoured him; and last this Nebuchadrezzar king of Babylon hath broken his bones.
JER|50|18|Therefore thus saith the LORD of hosts, the God of Israel; Behold, I will punish the king of Babylon and his land, as I have punished the king of Assyria.
JER|50|19|And I will bring Israel again to his habitation, and he shall feed on Carmel and Bashan, and his soul shall be satisfied upon mount Ephraim and Gilead.
JER|50|20|In those days, and in that time, saith the LORD, the iniquity of Israel shall be sought for, and there shall be none; and the sins of Judah, and they shall not be found: for I will pardon them whom I reserve.
JER|50|21|Go up against the land of Merathaim, even against it, and against the inhabitants of Pekod: waste and utterly destroy after them, saith the LORD, and do according to all that I have commanded thee.
JER|50|22|A sound of battle is in the land, and of great destruction.
JER|50|23|How is the hammer of the whole earth cut asunder and broken! how is Babylon become a desolation among the nations!
JER|50|24|I have laid a snare for thee, and thou art also taken, O Babylon, and thou wast not aware: thou art found, and also caught, because thou hast striven against the LORD.
JER|50|25|The LORD hath opened his armoury, and hath brought forth the weapons of his indignation: for this is the work of the Lord GOD of hosts in the land of the Chaldeans.
JER|50|26|Come against her from the utmost border, open her storehouses: cast her up as heaps, and destroy her utterly: let nothing of her be left.
JER|50|27|Slay all her bullocks; let them go down to the slaughter: woe unto them! for their day is come, the time of their visitation.
JER|50|28|The voice of them that flee and escape out of the land of Babylon, to declare in Zion the vengeance of the LORD our God, the vengeance of his temple.
JER|50|29|Call together the archers against Babylon: all ye that bend the bow, camp against it round about; let none thereof escape: recompense her according to her work; according to all that she hath done, do unto her: for she hath been proud against the LORD, against the Holy One of Israel.
JER|50|30|Therefore shall her young men fall in the streets, and all her men of war shall be cut off in that day, saith the LORD.
JER|50|31|Behold, I am against thee, O thou most proud, saith the Lord GOD of hosts: for thy day is come, the time that I will visit thee.
JER|50|32|And the most proud shall stumble and fall, and none shall raise him up: and I will kindle a fire in his cities, and it shall devour all round about him.
JER|50|33|Thus saith the LORD of hosts; The children of Israel and the children of Judah were oppressed together: and all that took them captives held them fast; they refused to let them go.
JER|50|34|Their Redeemer is strong; the LORD of hosts is his name: he shall throughly plead their cause, that he may give rest to the land, and disquiet the inhabitants of Babylon.
JER|50|35|A sword is upon the Chaldeans, saith the LORD, and upon the inhabitants of Babylon, and upon her princes, and upon her wise men.
JER|50|36|A sword is upon the liars; and they shall dote: a sword is upon her mighty men; and they shall be dismayed.
JER|50|37|A sword is upon their horses, and upon their chariots, and upon all the mingled people that are in the midst of her; and they shall become as women: a sword is upon her treasures; and they shall be robbed.
JER|50|38|A drought is upon her waters; and they shall be dried up: for it is the land of graven images, and they are mad upon their idols.
JER|50|39|Therefore the wild beasts of the desert with the wild beasts of the islands shall dwell there, and the owls shall dwell therein: and it shall be no more inhabited for ever; neither shall it be dwelt in from generation to generation.
JER|50|40|As God overthrew Sodom and Gomorrah and the neighbour cities thereof, saith the LORD; so shall no man abide there, neither shall any son of man dwell therein.
JER|50|41|Behold, a people shall come from the north, and a great nation, and many kings shall be raised up from the coasts of the earth.
JER|50|42|They shall hold the bow and the lance: they are cruel, and will not shew mercy: their voice shall roar like the sea, and they shall ride upon horses, every one put in array, like a man to the battle, against thee, O daughter of Babylon.
JER|50|43|The king of Babylon hath heard the report of them, and his hands waxed feeble: anguish took hold of him, and pangs as of a woman in travail.
JER|50|44|Behold, he shall come up like a lion from the swelling of Jordan unto the habitation of the strong: but I will make them suddenly run away from her: and who is a chosen man, that I may appoint over her? for who is like me? and who will appoint me the time? and who is that shepherd that will stand before me?
JER|50|45|Therefore hear ye the counsel of the LORD, that he hath taken against Babylon; and his purposes, that he hath purposed against the land of the Chaldeans: Surely the least of the flock shall draw them out: surely he shall make their habitation desolate with them.
JER|50|46|At the noise of the taking of Babylon the earth is moved, and the cry is heard among the nations.
JER|51|1|Thus saith the LORD; Behold, I will raise up against Babylon, and against them that dwell in the midst of them that rise up against me, a destroying wind;
JER|51|2|And will send unto Babylon fanners, that shall fan her, and shall empty her land: for in the day of trouble they shall be against her round about.
JER|51|3|Against him that bendeth let the archer bend his bow, and against him that lifteth himself up in his brigandine: and spare ye not her young men; destroy ye utterly all her host.
JER|51|4|Thus the slain shall fall in the land of the Chaldeans, and they that are thrust through in her streets.
JER|51|5|For Israel hath not been forsaken, nor Judah of his God, of the LORD of hosts; though their land was filled with sin against the Holy One of Israel.
JER|51|6|Flee out of the midst of Babylon, and deliver every man his soul: be not cut off in her iniquity; for this is the time of the LORD's vengeance; he will render unto her a recompence.
JER|51|7|Babylon hath been a golden cup in the LORD's hand, that made all the earth drunken: the nations have drunken of her wine; therefore the nations are mad.
JER|51|8|Babylon is suddenly fallen and destroyed: howl for her; take balm for her pain, if so be she may be healed.
JER|51|9|We would have healed Babylon, but she is not healed: forsake her, and let us go every one into his own country: for her judgment reacheth unto heaven, and is lifted up even to the skies.
JER|51|10|The LORD hath brought forth our righteousness: come, and let us declare in Zion the work of the LORD our God.
JER|51|11|Make bright the arrows; gather the shields: the LORD hath raised up the spirit of the kings of the Medes: for his device is against Babylon, to destroy it; because it is the vengeance of the LORD, the vengeance of his temple.
JER|51|12|Set up the standard upon the walls of Babylon, make the watch strong, set up the watchmen, prepare the ambushes: for the LORD hath both devised and done that which he spake against the inhabitants of Babylon.
JER|51|13|O thou that dwellest upon many waters, abundant in treasures, thine end is come, and the measure of thy covetousness.
JER|51|14|The LORD of hosts hath sworn by himself, saying, Surely I will fill thee with men, as with caterpillers; and they shall lift up a shout against thee.
JER|51|15|He hath made the earth by his power, he hath established the world by his wisdom, and hath stretched out the heaven by his understanding.
JER|51|16|When he uttereth his voice, there is a multitude of waters in the heavens; and he causeth the vapours to ascend from the ends of the earth: he maketh lightnings with rain, and bringeth forth the wind out of his treasures.
JER|51|17|Every man is brutish by his knowledge; every founder is confounded by the graven image: for his molten image is falsehood, and there is no breath in them.
JER|51|18|They are vanity, the work of errors: in the time of their visitation they shall perish.
JER|51|19|The portion of Jacob is not like them; for he is the former of all things: and Israel is the rod of his inheritance: the LORD of hosts is his name.
JER|51|20|Thou art my battle axe and weapons of war: for with thee will I break in pieces the nations, and with thee will I destroy kingdoms;
JER|51|21|And with thee will I break in pieces the horse and his rider; and with thee will I break in pieces the chariot and his rider;
JER|51|22|With thee also will I break in pieces man and woman; and with thee will I break in pieces old and young; and with thee will I break in pieces the young man and the maid;
JER|51|23|I will also break in pieces with thee the shepherd and his flock; and with thee will I break in pieces the husbandman and his yoke of oxen; and with thee will I break in pieces captains and rulers.
JER|51|24|And I will render unto Babylon and to all the inhabitants of Chaldea all their evil that they have done in Zion in your sight, saith the LORD.
JER|51|25|Behold, I am against thee, O destroying mountain, saith the LORD, which destroyest all the earth: and I will stretch out mine hand upon thee, and roll thee down from the rocks, and will make thee a burnt mountain.
JER|51|26|And they shall not take of thee a stone for a corner, nor a stone for foundations; but thou shalt be desolate for ever, saith the LORD.
JER|51|27|Set ye up a standard in the land, blow the trumpet among the nations, prepare the nations against her, call together against her the kingdoms of Ararat, Minni, and Ashchenaz; appoint a captain against her; cause the horses to come up as the rough caterpillers.
JER|51|28|Prepare against her the nations with the kings of the Medes, the captains thereof, and all the rulers thereof, and all the land of his dominion.
JER|51|29|And the land shall tremble and sorrow: for every purpose of the LORD shall be performed against Babylon, to make the land of Babylon a desolation without an inhabitant.
JER|51|30|The mighty men of Babylon have forborn to fight, they have remained in their holds: their might hath failed; they became as women: they have burned her dwellingplaces; her bars are broken.
JER|51|31|One post shall run to meet another, and one messenger to meet another, to shew the king of Babylon that his city is taken at one end,
JER|51|32|And that the passages are stopped, and the reeds they have burned with fire, and the men of war are affrighted.
JER|51|33|For thus saith the LORD of hosts, the God of Israel; The daughter of Babylon is like a threshingfloor, it is time to thresh her: yet a little while, and the time of her harvest shall come.
JER|51|34|Nebuchadrezzar the king of Babylon hath devoured me, he hath crushed me, he hath made me an empty vessel, he hath swallowed me up like a dragon, he hath filled his belly with my delicates, he hath cast me out.
JER|51|35|The violence done to me and to my flesh be upon Babylon, shall the inhabitant of Zion say; and my blood upon the inhabitants of Chaldea, shall Jerusalem say.
JER|51|36|Therefore thus saith the LORD; Behold, I will plead thy cause, and take vengeance for thee; and I will dry up her sea, and make her springs dry.
JER|51|37|And Babylon shall become heaps, a dwellingplace for dragons, an astonishment, and an hissing, without an inhabitant.
JER|51|38|They shall roar together like lions: they shall yell as lions' whelps.
JER|51|39|In their heat I will make their feasts, and I will make them drunken, that they may rejoice, and sleep a perpetual sleep, and not wake, saith the LORD.
JER|51|40|I will bring them down like lambs to the slaughter, like rams with he goats.
JER|51|41|How is Sheshach taken! and how is the praise of the whole earth surprised! how is Babylon become an astonishment among the nations!
JER|51|42|The sea is come up upon Babylon: she is covered with the multitude of the waves thereof.
JER|51|43|Her cities are a desolation, a dry land, and a wilderness, a land wherein no man dwelleth, neither doth any son of man pass thereby.
JER|51|44|And I will punish Bel in Babylon, and I will bring forth out of his mouth that which he hath swallowed up: and the nations shall not flow together any more unto him: yea, the wall of Babylon shall fall.
JER|51|45|My people, go ye out of the midst of her, and deliver ye every man his soul from the fierce anger of the LORD.
JER|51|46|And lest your heart faint, and ye fear for the rumour that shall be heard in the land; a rumour shall both come one year, and after that in another year shall come a rumour, and violence in the land, ruler against ruler.
JER|51|47|Therefore, behold, the days come, that I will do judgment upon the graven images of Babylon: and her whole land shall be confounded, and all her slain shall fall in the midst of her.
JER|51|48|Then the heaven and the earth, and all that is therein, shall sing for Babylon: for the spoilers shall come unto her from the north, saith the LORD.
JER|51|49|As Babylon hath caused the slain of Israel to fall, so at Babylon shall fall the slain of all the earth.
JER|51|50|Ye that have escaped the sword, go away, stand not still: remember the LORD afar off, and let Jerusalem come into your mind.
JER|51|51|We are confounded, because we have heard reproach: shame hath covered our faces: for strangers are come into the sanctuaries of the LORD's house.
JER|51|52|Wherefore, behold, the days come, saith the LORD, that I will do judgment upon her graven images: and through all her land the wounded shall groan.
JER|51|53|Though Babylon should mount up to heaven, and though she should fortify the height of her strength, yet from me shall spoilers come unto her, saith the LORD.
JER|51|54|A sound of a cry cometh from Babylon, and great destruction from the land of the Chaldeans:
JER|51|55|Because the LORD hath spoiled Babylon, and destroyed out of her the great voice; when her waves do roar like great waters, a noise of their voice is uttered:
JER|51|56|Because the spoiler is come upon her, even upon Babylon, and her mighty men are taken, every one of their bows is broken: for the LORD God of recompences shall surely requite.
JER|51|57|And I will make drunk her princes, and her wise men, her captains, and her rulers, and her mighty men: and they shall sleep a perpetual sleep, and not wake, saith the King, whose name is the LORD of hosts.
JER|51|58|Thus saith the LORD of hosts; The broad walls of Babylon shall be utterly broken, and her high gates shall be burned with fire; and the people shall labour in vain, and the folk in the fire, and they shall be weary.
JER|51|59|The word which Jeremiah the prophet commanded Seraiah the son of Neriah, the son of Maaseiah, when he went with Zedekiah the king of Judah into Babylon in the fourth year of his reign. And this Seraiah was a quiet prince.
JER|51|60|So Jeremiah wrote in a book all the evil that should come upon Babylon, even all these words that are written against Babylon.
JER|51|61|And Jeremiah said to Seraiah, When thou comest to Babylon, and shalt see, and shalt read all these words;
JER|51|62|Then shalt thou say, O LORD, thou hast spoken against this place, to cut it off, that none shall remain in it, neither man nor beast, but that it shall be desolate for ever.
JER|51|63|And it shall be, when thou hast made an end of reading this book, that thou shalt bind a stone to it, and cast it into the midst of Euphrates:
JER|51|64|And thou shalt say, Thus shall Babylon sink, and shall not rise from the evil that I will bring upon her: and they shall be weary. Thus far are the words of Jeremiah.
JER|52|1|Zedekiah was one and twenty years old when he began to reign, and he reigned eleven years in Jerusalem. And his mother's name was Hamutal the daughter of Jeremiah of Libnah.
JER|52|2|And he did that which was evil in the eyes of the LORD, according to all that Jehoiakim had done.
JER|52|3|For through the anger of the LORD it came to pass in Jerusalem and Judah, till he had cast them out from his presence, that Zedekiah rebelled against the king of Babylon.
JER|52|4|And it came to pass in the ninth year of his reign, in the tenth month, in the tenth day of the month, that Nebuchadrezzar king of Babylon came, he and all his army, against Jerusalem, and pitched against it, and built forts against it round about.
JER|52|5|So the city was besieged unto the eleventh year of king Zedekiah.
JER|52|6|And in the fourth month, in the ninth day of the month, the famine was sore in the city, so that there was no bread for the people of the land.
JER|52|7|Then the city was broken up, and all the men of war fled, and went forth out of the city by night by the way of the gate between the two walls, which was by the king's garden; (now the Chaldeans were by the city round about:) and they went by the way of the plain.
JER|52|8|But the army of the Chaldeans pursued after the king, and overtook Zedekiah in the plains of Jericho; and all his army was scattered from him.
JER|52|9|Then they took the king, and carried him up unto the king of Babylon to Riblah in the land of Hamath; where he gave judgment upon him.
JER|52|10|And the king of Babylon slew the sons of Zedekiah before his eyes: he slew also all the princes of Judah in Riblah.
JER|52|11|Then he put out the eyes of Zedekiah; and the king of Babylon bound him in chains, and carried him to Babylon, and put him in prison till the day of his death.
JER|52|12|Now in the fifth month, in the tenth day of the month, which was the nineteenth year of Nebuchadrezzar king of Babylon, came Nebuzaradan, captain of the guard, which served the king of Babylon, into Jerusalem,
JER|52|13|And burned the house of the LORD, and the king's house; and all the houses of Jerusalem, and all the houses of the great men, burned he with fire:
JER|52|14|And all the army of the Chaldeans, that were with the captain of the guard, brake down all the walls of Jerusalem round about.
JER|52|15|Then Nebuzaradan the captain of the guard carried away captive certain of the poor of the people, and the residue of the people that remained in the city, and those that fell away, that fell to the king of Babylon, and the rest of the multitude.
JER|52|16|But Nebuzaradan the captain of the guard left certain of the poor of the land for vinedressers and for husbandmen.
JER|52|17|Also the pillars of brass that were in the house of the LORD, and the bases, and the brasen sea that was in the house of the LORD, the Chaldeans brake, and carried all the brass of them to Babylon.
JER|52|18|The caldrons also, and the shovels, and the snuffers, and the bowls, and the spoons, and all the vessels of brass wherewith they ministered, took they away.
JER|52|19|And the basons, and the firepans, and the bowls, and the caldrons, and the candlesticks, and the spoons, and the cups; that which was of gold in gold, and that which was of silver in silver, took the captain of the guard away.
JER|52|20|The two pillars, one sea, and twelve brasen bulls that were under the bases, which king Solomon had made in the house of the LORD: the brass of all these vessels was without weight.
JER|52|21|And concerning the pillars, the height of one pillar was eighteen cubits; and a fillet of twelve cubits did compass it; and the thickness thereof was four fingers: it was hollow.
JER|52|22|And a chapiter of brass was upon it; and the height of one chapiter was five cubits, with network and pomegranates upon the chapiters round about, all of brass. The second pillar also and the pomegranates were like unto these.
JER|52|23|And there were ninety and six pomegranates on a side; and all the pomegranates upon the network were an hundred round about.
JER|52|24|And the captain of the guard took Seraiah the chief priest, and Zephaniah the second priest, and the three keepers of the door:
JER|52|25|He took also out of the city an eunuch, which had the charge of the men of war; and seven men of them that were near the king's person, which were found in the city; and the principal scribe of the host, who mustered the people of the land; and threescore men of the people of the land, that were found in the midst of the city.
JER|52|26|So Nebuzaradan the captain of the guard took them, and brought them to the king of Babylon to Riblah.
JER|52|27|And the king of Babylon smote them, and put them to death in Riblah in the land of Hamath. Thus Judah was carried away captive out of his own land.
JER|52|28|This is the people whom Nebuchadrezzar carried away captive: in the seventh year three thousand Jews and three and twenty:
JER|52|29|In the eighteenth year of Nebuchadrezzar he carried away captive from Jerusalem eight hundred thirty and two persons:
JER|52|30|In the three and twentieth year of Nebuchadrezzar Nebuzaradan the captain of the guard carried away captive of the Jews seven hundred forty and five persons: all the persons were four thousand and six hundred.
JER|52|31|And it came to pass in the seven and thirtieth year of the captivity of Jehoiachin king of Judah, in the twelfth month, in the five and twentieth day of the month, that Evilmerodach king of Babylon in the first year of his reign lifted up the head of Jehoiachin king of Judah, and brought him forth out of prison.
JER|52|32|And spake kindly unto him, and set his throne above the throne of the kings that were with him in Babylon,
JER|52|33|And changed his prison garments: and he did continually eat bread before him all the days of his life.
JER|52|34|And for his diet, there was a continual diet given him of the king of Babylon, every day a portion until the day of his death, all the days of his life.
