2JOHN|1|1|我作长老的写信给蒙拣选的夫人 和她的儿女，就是我真心所爱的；不但我爱，也是一切认识真理的人所爱的，
2JOHN|1|2|这是因为真理住在我们里面，也必与我们同在直到永远。
2JOHN|1|3|愿恩惠、怜悯、平安 从父上帝和他儿子耶稣基督，在真理和爱中必与我们同在。
2JOHN|1|4|我非常欢喜见你的儿女，有照我们从父所受之命令遵行真理的。
2JOHN|1|5|夫人哪，我现在请求你，我们大家要彼此相爱。我写给你的，并不是一条新命令，而是我们从起初就有的。
2JOHN|1|6|这就是爱，就是照他的命令行事；这就是命令，你们要照这命令行，正如你们从起初所听见的。
2JOHN|1|7|有许多迷惑人的已经来到世上，他们不宣认耶稣基督是成了肉身来的；这样的人是迷惑人的，是敌基督的。
2JOHN|1|8|你们要小心，不要失去你们 所完成的工作，而要得到充足的赏赐。
2JOHN|1|9|凡越过基督的教导而不持守的，就没有上帝；凡持守这教导的，就有父又有子。
2JOHN|1|10|若有人到你们那里而不传这教导，不要接他到家里，也不要向他问安；
2JOHN|1|11|因为向他问安的，就在他的恶行上有份。
2JOHN|1|12|我还有许多事要写给你们，却不愿意用纸用墨，但盼望到你们那里，与你们面对面谈论，使我们的喜乐得以满足。
2JOHN|1|13|你那蒙拣选的姊妹的儿女向你问安。
