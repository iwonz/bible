1SAM|1|1|Fuit vir unus de Ramathaim Suphita de monte Ephraim, et nomen eius Elcana filius Ieroham filii Eliu filii Thohu filii Suph, Ephrathaeus.
1SAM|1|2|Et habuit duas uxores: nomen uni Anna et nomen secundae Phenenna. Fueruntque Phenennae filii, Annae autem non erant liberi.
1SAM|1|3|Et ascendebat vir ille de civitate sua singulis annis, ut adoraret et sacrificaret Domino exercituum in Silo. Erant autem ibi duo filii Heli, Ophni et Phinees, sacerdotes Domini.
1SAM|1|4|Venit ergo dies, et immolavit Elcana dabatque Phenennae uxori suae et cunctis filiis eius et filiabus partes;
1SAM|1|5|Annae autem dabat unam partem electam, quia Annam diligebat; Dominus autem concluserat vulvam eius.
1SAM|1|6|Affligebat quoque eam aemula eius et vehementer angebat, ut conturbaret eam, quod conclusisset Dominus vulvam eius.
1SAM|1|7|Sicque faciebat per singulos annos, cum, redeunte tempore, ascenderent templum Domini, et sic provocabat eam. Porro illa flebat et non capiebat cibum.
1SAM|1|8|Dixit ergo ei Elcana vir suus: " Anna, cur fles et quare non comedis? Et quam ob rem affligitur cor tuum? Numquid non ego melior sum tibi quam decem filii? ".
1SAM|1|9|Surrexit autem Anna, postquam comederant et biberant in Silo, et Heli sacerdote sedente super sellam ante postes templi Domini.
1SAM|1|10|Cum esset Anna amaro animo, oravit Dominum flens largiter
1SAM|1|11|et votum vovit dicens: " Domine exercituum, si respiciens videris afflictionem famulae tuae et recordatus mei fueris nec oblitus ancillae tuae dederisque servae tuae sexum virilem, dabo eum Domino omnes dies vitae eius, et novacula non ascendet super caput eius ".
1SAM|1|12|Factum est ergo, cum illa multiplicaret preces coram Domino, ut Heli observaret os eius.
1SAM|1|13|Porro Anna loquebatur in corde suo; tantumque labia illius movebantur, et vox penitus non audiebatur. Aestimavit igitur eam Heli temulentam
1SAM|1|14|dixitque ei: " Usquequo ebria eris? Digere paulisper vinum, quo mades!.
1SAM|1|15|Respondens Anna: " Nequaquam, inquit, domine mi; nam mulier infelix nimis ego sum: vinumque et omne, quod inebriare potest, non bibi, sed effudi animam meam in conspectu Domini.
1SAM|1|16|Ne reputes ancillam tuam quasi unam de filiabus Belial, quia ex multitudine doloris et maeroris mei locuta sum usque in praesens ".
1SAM|1|17|Tunc Heli ait ei: " Vade in pace, et Deus Israel det tibi petitionem, quam rogasti eum ".
1SAM|1|18|Et illa dixit: " Utinam inveniat ancilla tua gratiam in oculis tuis ". Et abiit mulier in viam suam et comedit; vultusque illius non fuerunt amplius sicut prius.
1SAM|1|19|Et surrexerunt mane et adoraverunt coram Domino.Reversique sunt et venerunt in domum suam in Rama. Cognovit autem Elcana Annam uxorem suam, et recordatus est eius Dominus.
1SAM|1|20|Et factum est post circulum dierum concepit Anna et peperit filium vocavitque nomen eius Samuel, eo quod a Domino postulasset eum.
1SAM|1|21|Ascendit autem vir Elcana et omnis domus eius, ut immolaret Domino hostiam annuam et votum suum.
1SAM|1|22|Et Anna non ascendit; dixit enim viro suo: " Non vadam, donec ablactetur infans, et ducam eum, et appareat ante conspectum Domini et maneat ibi iugiter ".
1SAM|1|23|Et ait ei Elcana vir suus: " Fac, quod bonum tibi videtur, et mane, donec ablactes eum; precorque, ut impleat Dominus verbum suum ". Mansit ergo mulier et lactavit filium suum, donec amoveret eum a lacte.
1SAM|1|24|Et adduxit eum secum, postquam ablactaverat, cum vitulo trium annorum et tribus modiis farinae et utre vini; et adduxit eum ad domum Domini in Silo. Puer autem erat adhuc infantulus.
1SAM|1|25|Et immolaverunt vitulum et obtulerunt puerum Heli,
1SAM|1|26|et ait Anna: " Obsecro, mi domine; vivit anima tua, domine, ego sum illa mulier, quae steti coram te hic orans Dominum.
1SAM|1|27|Pro puero isto oravi, et dedit mihi Dominus petitionem meam, quam postulavi eum.
1SAM|1|28|Idcirco et ego commodavi eum Domino; cunctis diebus, quibus vivet, postulatus erit pro Domino ".Et adoraverunt ibi Dominum.
1SAM|2|1|Et oravit Anna et ait: Exsultavit cor meum in Do mino,exaltatum est cornu meum in Deo meo;dilatatum est os meum super inimicos meos,quoniam laetata sum in salutari tuo.
1SAM|2|2|Non est sanctus ut est Dominus;neque enim est alius extra te,et non est fortis sicut Deus noster.
1SAM|2|3|Nolite multiplicare loqui sublimia gloriantes.Recedant superba de ore vestro,quia Deus scientiarum Dominus est, et ab eo ponderantur actiones.
1SAM|2|4|Arcus fortium confractus est,et infirmi accincti sunt robore.
1SAM|2|5|Saturati prius pro pane se locaverunt,et famelici non eguerunt amplius.Sterilis peperit plurimos,et, quae multos habebat filios, emarcuit.
1SAM|2|6|Dominus mortificat et vivificat,deducit ad infernum et reducit.
1SAM|2|7|Dominus pauperem facit et ditat,humiliat et sublevat;
1SAM|2|8|suscitat de pulvere egenumet de stercore elevat pauperem,ut sedeat cum principibuset solium gloriae teneat.Domini enim sunt cardines terrae, et posuit super eos orbem.
1SAM|2|9|Pedes sanctorum suorum servabit,et impii in tenebris conticescent,quia non in fortitudine sua roborabitur vir.
1SAM|2|10|Dominus conteret adversarios suos;super ipsos in caelis tonabit.Dominus iudicabit fines terraeet dabit imperium regi suoet sublimabit cornu christi sui ".
1SAM|2|11|Et abiit Elcana in Rama in domum suam. Puer autem erat minister in conspectu Domini ante faciem Heli sacerdotis.
1SAM|2|12|Porro filii Heli filii Belial nescientes Dominum
1SAM|2|13|neque officium sacerdotum ad populum, sed, quicumque immolasset victimam, veniebat puer sacerdotis, dum coquerentur carnes, et habebat fuscinulam tridentem in manu sua
1SAM|2|14|et mittebat eam in lebetem vel in caldariam aut in ollam sive in cacabum et omne, quod levabat fuscinula, tollebat sacerdos sibi. Sic faciebant universo Israeli venienti in Silo.
1SAM|2|15|Etiam, antequam adolerent adipem, veniebat puer sacerdotis et dicebat immolanti: " Da mihi carnem, ut coquam sacerdoti; non enim accipiet a te carnem coctam sed crudam ".
1SAM|2|16|Dicebatque illi immolans: " Incendatur primum iuxta morem hodie adeps, et tolle tibi, quantumcumque desiderat anima tua ". Qui respondens aiebat ei: " Nequaquam; nunc enim dabis, alioquin tollam vi ".
1SAM|2|17|Erat ergo peccatum puerorum grande nimis coram Domino, quia detrahebant sacrificio Domini.
1SAM|2|18|Samuel autem ministrabat ante faciem Domini, puer accinctus ephod lineo.
1SAM|2|19|Et tunicam parvam faciebat ei mater sua, quam afferebat ei singulis annis ascendens cum viro suo, ut immolaret hostiam annuam.
1SAM|2|20|Et benedicebat Heli Elcanae et uxori eius dicebatque: " Reddat tibi Dominus semen de muliere hac pro petitione, quae postulata est pro Domino. Et abierunt in locum suum.
1SAM|2|21|Visitavit ergo Dominus Annam, et concepit et peperit tres filios et duas filias. Et crevit puer Samuel apud Dominum.
1SAM|2|22|Heli autem erat senex valde et audivit omnia, quae faciebant filii sui universo Israeli et quomodo dormiebant cum mulieribus, quae ministrabant ad ostium tabernaculi,
1SAM|2|23|et dixit eis: " Quare facitis res huiuscemodi, quas ego audio, res pessimas, ab omni populo?
1SAM|2|24|Nolite, filii mei; non enim est bona fama, quam ego audio, ut transgredi faciatis populum Domini.
1SAM|2|25|Si peccaverit vir in virum,arbiter ei potest esse Deus;si autem in Dominum peccaverit vir,quis intercedet pro eo? ".Et non audierunt vocem patris sui, quia voluit Dominus occidere eos.
1SAM|2|26|Puer autem Samuel proficiebat atque crescebat et placebat tam Domino quam hominibus.
1SAM|2|27|Venit autem vir Dei ad Heli et ait ad eum: " Haec dicit Dominus: Numquid non aperte revelatus sum domui patris tui, cum esset in Aegypto in domo pharaonis?
1SAM|2|28|Et elegi eum ex omnibus tribubus Israel mihi in sacerdotem, ut ascenderet ad altare meum et adoleret mihi incensum et portaret ephod coram me; et dedi domui patris tui omnia de sacrificiis filiorum Israel.
1SAM|2|29|Quare calce abicitis victimam meam et munera mea, quae praecepi, ut offerrentur in templo, et magis honorasti filios tuos quam me, ut impinguaremini primitiis omnis sacrificii Israel populi mei?
1SAM|2|30|Propterea ait Dominus, Deus Israel: Loquens locutus sum, ut domus tua et domus patris tui ministraret in conspectu meo usque in sempiternum. Nunc autem, dicit Dominus, absit hoc a me. Sed quicumque glorificaverit me, glorificabo eum; qui autem contemnunt me, erunt ignobiles.
1SAM|2|31|Ecce dies veniunt, et praecidam brachium tuum et brachium domus patris tui, ut non sit senex in domo tua.
1SAM|2|32|Et videbis aemulum tuum in templo in universis prosperis Israel; et non erit senex in domo tua omnibus diebus.
1SAM|2|33|Verumtamen non auferam penitus virum ex te ab altari meo; sed ut deficiant oculi tui, et tabescat anima tua, et pars magna domus tuae morietur, cum ad virilem aetatem venerit.
1SAM|2|34|Hoc autem erit tibi signum, quod venturum est duobus filiis tuis Ophni et Phinees: in die uno morientur ambo.
1SAM|2|35|Et suscitabo mihi sacerdotem fidelem, qui iuxta cor meum et animam meam faciat; et aedificabo ei domum fidelem, et ambulabit coram christo meo cunctis diebus.
1SAM|2|36|Futurum est autem ut quicumque remanserit in domo tua, veniat, ut procidat ante illum pro nummo argenteo et torta panis dicatque: "Dimitte me, obsecro, ad unam partem sacerdotalem, ut comedam buccellam panis" ".
1SAM|3|1|Puer autem Samuel ministrabat Domino coram Heli. Et sermo Domini erat pretiosus in diebus illis: non erat visio frequens.
1SAM|3|2|Factum est ergo in die quadam, Heli iacebat in loco suo, et oculi eius caligaverant, nec poterat videre.
1SAM|3|3|Lucerna Dei nondum exstincta erat, et Samuel dormiebat in templo Domini, ubi erat arca Dei.
1SAM|3|4|Et vocavit Dominus Samuel, qui respondens ait: " Ecce ego ".
1SAM|3|5|Et cucurrit ad Heli et dixit: " Ecce ego; vocasti enim me ". Qui dixit: Non vocavi. Revertere; dormi! ". Et abiit et dormivit.
1SAM|3|6|Et Dominus rursum vocavit Samuel. Consurgensque Samuel abiit ad Heli et dixit: " Ecce ego, quia vocasti me ". Qui respondit: " Non vocavi te, fili mi. Revertere et dormi! ".
1SAM|3|7|Porro Samuel necdum sciebat Dominum, neque revelatus fuerat ei sermo Domini.
1SAM|3|8|Et Dominus rursum vocavit Samuel tertio, qui consurgens abiit ad Heli
1SAM|3|9|et ait: " Ecce ego, quia vocasti me ". Intellexit igitur Heli quia Dominus vocaret puerum, et ait ad Samuel: " Vade et dormi; et, si deinceps vocaverit te, dices: " Loquere, Domine, quia audit servus tuus" ". Abiit ergo Samuel et dormivit in loco suo.
1SAM|3|10|Et venit Dominus et stetit et vocavit, sicut vocaverat prius: " Samuel, Samuel ". Et ait Samuel: " Loquere, quia audit servus tuus ".
1SAM|3|11|Et dixit Dominus ad Samuel: " Ecce ego facio verbum in Israel, quod quicumque audierit, tinnient ambae aures eius.
1SAM|3|12|In die illo suscitabo adversum Heli omnia, quae locutus sum super domum eius: incipiam et complebo.
1SAM|3|13|Praedixi enim ei quod iudicaturus essem domum eius in aeternum propter iniquitatem, eo quod noverat filios suos contemnere Deum et non corripuit eos.
1SAM|3|14|Idcirco iuravi domui Heli quod non expietur iniquitas domus eius victimis et muneribus usque in aeternum ".
1SAM|3|15|Dormivit autem Samuel usque mane aperuitque ostia domus Domini. Et Samuel timebat indicare visionem Heli.
1SAM|3|16|Vocavit ergo Heli Samuelem et dixit: " Samuel, fili mi ". Qui respondens ait: " Praesto sum ".
1SAM|3|17|Et interrogavit eum: " Quis est sermo, quem locutus est ad te? Oro te, ne celaveris me. Haec faciat tibi Deus et haec addat, si absconderis a me sermonem ex omnibus verbis, quae dicta sunt tibi ".
1SAM|3|18|Indicavit itaque ei Samuel universos sermones et non abscondit ab eo. Et ille respondit: " Dominus est! Quod bonum est in oculis suis, faciat ".
1SAM|3|19|Crevit autem Samuel, et Dominus erat cum eo, et non cecidit ex omnibus verbis eius in terram.
1SAM|3|20|Et cognovit universus Israel a Dan usque Bersabee quod constitutus esset Samuel propheta Domini.
1SAM|3|21|Et addidit Dominus ut appareret in Silo, quoniam revelatus fuerat Dominus Samueli in Silo iuxta verbum Domini. Et evenit sermo Samuelis universo Israeli.
1SAM|4|1|Et factum est in diebus illis, convenerunt Philisthim in pu gnam; et egressus est Israel obviam Philisthim in proelium et castrametatus est iuxta Abenezer. Porro Philisthim venerunt in Aphec
1SAM|4|2|et instruxerunt aciem contra Israel. Crescente autem certamine, terga vertit Israel Philisthaeis; et caesi sunt in illo certamine passim per agros quasi quattuor milia virorum.
1SAM|4|3|Et reversus est populus ad castra, dixeruntque maiores natu de Israel: " Quare percussit nos Dominus hodie coram Philisthim? Afferamus ad nos de Silo arcam foederis Domini, et veniat in medium nostri, ut salvet nos de manu inimicorum nostrorum ".
1SAM|4|4|Misit ergo populus in Silo, et tulerunt inde arcam foederis Domini exercituum sedentis super cherubim; erantque duo filii Heli cum arca foederis Dei, Ophni et Phinees.
1SAM|4|5|Cumque venisset arca foederis Domini in castra, vociferatus est omnis Israel clamore grandi, et personuit terra.
1SAM|4|6|Et audierunt Philisthim vocem clamoris dixeruntque: " Quaenam est haec vox clamoris magni in castris Hebraeorum? ". Et cognoverunt quod arca Domini venisset in castra.
1SAM|4|7|Timueruntque Philisthim dicentes: " Venit Deus in castra! ". Et ingemuerunt dicentes:
1SAM|4|8|" Vae nobis! Non enim fuit tanta exsultatio heri et nudiustertius. Vae nobis! Quis nos servabit de manu deorum sublimium istorum? Hi sunt dii, qui percusserunt Aegyptum omni plaga in deserto.
1SAM|4|9|Confortamini et estote viri, Philisthim, ne serviatis Hebraeis, sicut illi servierunt vobis. Estote viri et bellate! ".
1SAM|4|10|Pugnaverunt ergo Philisthim, et caesus est Israel, et fugit unusquisque in tabernaculum suum; et facta est plaga magna nimis, et ceciderunt de Israel triginta milia peditum.
1SAM|4|11|Et arca Dei capta est; duoque filii Heli mortui sunt, Ophni et Phinees.
1SAM|4|12|Currens autem vir de Beniamin ex acie venit in Silo in die illo scissa veste et conspersus pulvere caput.
1SAM|4|13|Cumque ille venisset, Heli sedebat super sellam iuxta portam aspectans viam; erat enim cor eius pavens pro arca Dei. Vir autem ille, postquam ingressus est, nuntiavit urbi; et ululavit omnis civitas.
1SAM|4|14|Et audivit Heli sonitum clamoris dixitque: " Quis est hic sonitus tumultus huius? ". At ille festinavit et venit et nuntiavit Heli.
1SAM|4|15|Heli autem erat nonaginta et octo annorum, et oculi eius caligaverant, et videre non poterat.
1SAM|4|16|Et dixit ad Heli: " Ego sum qui veni de proelio et ego qui de acie fugi hodie ". Cui ille ait: " Quid actum est, fili mi? ".
1SAM|4|17|Respondens autem, qui nuntiabat: " Fugit, inquit, Israel coram Philisthim, et ruina magna facta est in populo; insuper et duo filii tui mortui sunt, Ophni et Phinees, et arca Dei capta est ".
1SAM|4|18|Cumque ille nominasset arcam Dei, cecidit de sella retrorsum iuxta ostium et, fractis cervicibus, mortuus est; senex enim erat vir et gravis. Et ipse iudicavit Israel quadraginta annis.
1SAM|4|19|Nurus autem eius, uxor Phinees, praegnans erat vicinaque partui. Et, audito nuntio quod capta esset arca Dei et mortuus socer suus et vir suus, incurvavit se et peperit; irruerant enim in eam dolores subiti.
1SAM|4|20|In ipso autem momento mortis eius dixerunt ei, quae stabant circa eam: Ne timeas, quia filium peperisti ". Quae non respondit eis neque animadvertit.
1SAM|4|21|Et vocavit puerum Ichabod dicens: " Translata est gloria de Israel! ", quia capta est arca Dei et pro socero suo et pro viro suo.
1SAM|4|22|Et ait: " Translata est gloria ab Israel, eo quod capta est arca Dei!.
1SAM|5|1|Philisthim autem tulerunt arcam Dei et asportaverunt eam a Abenezer in Azotum.
1SAM|5|2|Tulerunt Philisthim arcam Dei et intulerunt eam in templum Dagon et statuerunt eam iuxta Dagon.
1SAM|5|3|Cumque surrexissent Azotii altera die, ecce Dagon iacebat pronus in terram ante arcam Domini; et tulerunt Dagon et restituerunt eum in loco suo.
1SAM|5|4|Rursumque mane die altera consurgentes invenerunt Dagon iacentem super faciem suam in terram coram arca Domini; caput autem Dagon et duae palmae manuum eius abscisae erant super limen:
1SAM|5|5|porro Dagon truncus solus remanserat in loco suo. Propter hanc causam non calcant sacerdotes Dagon et omnes, qui ingrediuntur templum eius, super limen Dagon in Azoto usque in hodiernum diem.
1SAM|5|6|Aggravata est autem manus Domini super Azotios, et demolitus est eos et percussit eos tumoribus, Azotum et fines eius.
1SAM|5|7|Videntes autem viri Azotii huiuscemodi plagam dixerunt: " Non maneat arca Dei Israel apud nos, quoniam dura est manus eius super nos et super Dagon deum nostrum ".
1SAM|5|8|Et mittentes congregaverunt omnes principes Philisthinorum ad se et dixerunt: " Quid faciemus de arca Dei Israel? ". Responderuntque: " In Geth circumducatur arca Dei Israel ". Et circumduxerunt arcam Dei Israel.
1SAM|5|9|Postquam autem circumduxerunt eam, facta est manus Domini super civitatem, pavor magnus nimis; et percussit viros urbis a parvo usque ad maiorem, et eruperunt eis tumores.
1SAM|5|10|Miserunt ergo arcam Dei in Accaron.Cumque venisset arca Dei in Accaron, exclamaverunt Accaronitae dicentes: " Adduxerunt ad nos arcam Dei Israel, ut interficiat nos et populum nostrum!.
1SAM|5|11|Miserunt itaque et congregaverunt omnes principes Philisthinorum et dixerunt: " Dimittite arcam Dei Israel, et revertatur in locum suum et non interficiat nos cum populo nostro ".
1SAM|5|12|Fiebat enim pavor mortis in tota civitate, et gravissima valde manus Dei. Viri quoque, qui mortui non fuerant, percutiebantur tumoribus, et ascendebat ululatus civitatis in caelum.
1SAM|6|1|Fuit ergo arca Domini in regio ne Philisthinorum septem mensi bus;
1SAM|6|2|et vocaverunt Philisthim sacerdotes et divinos dicentes: " Quid faciemus de arca Domini? Indicate nobis quomodo remittemus eam in locum suum ".Qui dixerunt:
1SAM|6|3|" Si remittitis arcam Dei Israel, nolite dimittere eam vacuam, sed, quod debetis, reddite ei pro peccato, et tunc curabimini; scietis quare non recedat manus eius a vobis ".
1SAM|6|4|Qui dixerunt: " Quid est quod pro delicto reddere debeamus ei? ". Responderuntque illi:
1SAM|6|5|" Iuxta numerum principum Philisthinorum quinque tumores aureos facietis et quinque mures aureos, quia plaga una fuit omnibus vobis et principibus vestris. Facietisque similitudines tumorum vestrorum et similitudines murium, qui demoliti sunt terram, et dabitis Deo Israel gloriam, si forte relevet manum suam a vobis et a diis vestris et a terra vestra.
1SAM|6|6|Quare gravatis corda vestra, sicut aggravavit Aegyptus et pharao cor suum? Nonne, postquam percussit eos, tunc dimiserunt eos, et abierunt?
1SAM|6|7|Nunc ergo arripite et facite plaustrum novum unum et duas vaccas fetas, quibus non est impositum iugum, iungite in plaustro; et recludite vitulos earum domi.
1SAM|6|8|Tolletisque arcam Domini et ponetis in plaustro; et similitudines aureas, quas exsolvistis ei pro delicto, ponetis in capsella ad latus eius et dimittite eam, ut vadat,
1SAM|6|9|et aspicietis. Et siquidem per viam finium suorum ascenderit contra Bethsames, ipse fecit nobis hoc malum grande; sin autem minime, sciemus quia nequaquam manus eius tetigit nos, sed casu accidit ".
1SAM|6|10|Fecerunt ergo illi hoc modo et tollentes duas vaccas, quae lactabant vitulos, iunxerunt ad plaustrum vitulosque earum concluserunt domi;
1SAM|6|11|et posuerunt arcam Dei super plaustrum et capsellam, quae habebat mures aureos et similitudines tumorum.
1SAM|6|12|Ibant autem in directum vaccae per viam, quae ducit Bethsames, et itinere uno gradiebantur pergentes et mugientes et non declinabant neque ad dextram neque ad sinistram. Sed et principes Philisthim sequebantur usque ad terminos Bethsames.
1SAM|6|13|Porro Bethsamitae metebant triticum in valle; et elevantes oculos viderunt arcam et gavisi sunt, cum vidissent.
1SAM|6|14|Et plaustrum venit in agrum Iosue Bethsamitae et stetit ibi. Erat autem ibi lapis magnus; et conciderunt ligna plaustri vaccasque imposuerunt super ea holocaustum Domino.
1SAM|6|15|Levitae autem deposuerunt arcam Dei et capsellam, quae erat iuxta eam, in qua erant similitudines aureae; et posuerunt super lapidem grandem. Viri autem Bethsamitae obtulerunt holocausta et immolaverunt victimas in die illa Domino.
1SAM|6|16|Et quinque principes Philisthinorum viderunt et reversi sunt in Accaron in die illa.
1SAM|6|17|Hi sunt autem tumores aurei, quos reddiderunt Philisthim pro delicto Domino: Azotus unum, Gaza unum, Ascalon unum, Geth unum, Accaron unum;
1SAM|6|18|et mures aureos secundum numerum urbium Philisthim quinque principum, ab urbe murata usque ad villam, quae erat absque muro; et lapis ille magnus, super quem posuerunt arcam Domini, testis est usque in hunc diem in agro Iosue Bethsamitis.
1SAM|6|19|Filii autem Iechoniae non sunt gavisi super viros Bethsamites quia viderant arcam Domini; et percussit Dominus de populo septuaginta viros. Luxitque populus eo quod Dominus percussisset plebem plaga magna;
1SAM|6|20|et dixerunt viri Bethsamitae: " Quis poterit stare in conspectu Domini, Dei sancti huius? Et ad quem ascendet a nobis? ".
1SAM|6|21|Miseruntque nuntios ad habitatores Cariathiarim dicentes: " Reduxerunt Philisthim arcam Domini. Descendite et ducite eam sursum ad vos ".
1SAM|7|1|Venerunt ergo viri Cariathiarim et duxerunt arcam Domini sursum et intulerunt eam in domum Abinadab in colle; Eleazarum autem filium eius sanctificaverunt, ut custodiret arcam Domini.
1SAM|7|2|Et factum est, ex qua die mansit arca Domini in Cariathiarim, multiplicati sunt dies; erat quippe iam annus vicesimus, et ingemuit omnis domus Israel post Dominum.
1SAM|7|3|Ait autem Samuel ad universam domum Israel dicens: " Si in toto corde vestro revertimini ad Dominum, auferte deos alienos de medio vestri et Astharoth et praeparate corda vestra Domino et servite ei soli, et eruet vos de manu Philisthim ".
1SAM|7|4|Abstulerunt ergo filii Israel Baalim et Astharoth et servierunt Domino soli.
1SAM|7|5|Dixit autem Samuel: " Congregate universum Israel in Maspha, ut orem pro vobis Dominum ".
1SAM|7|6|Et convenerunt in Maspha hauseruntque aquam et effuderunt in conspectu Domini et ieiunaverunt in die illa et dixerunt ibi: " Peccavimus Domino ". Iudicavitque Samuel filios Israel in Maspha.
1SAM|7|7|Et audierunt Philisthim quod congregati essent filii Israel in Maspha, et ascenderunt principes Philisthinorum ad Israel. Quod cum audissent filii Israel, timuerunt a facie Philisthinorum
1SAM|7|8|dixeruntque ad Samuel: " Ne cesses pro nobis clamare ad Dominum Deum nostrum, ut salvet nos de manu Philisthinorum ".
1SAM|7|9|Tulit ergo Samuel agnum lactantem unum et obtulit illum holocaustum integrum Domino; et clamavit Samuel ad Dominum pro Israel, et exaudivit eum Dominus.
1SAM|7|10|Factum est autem cum Samuel offerret holocaustum, Philisthim iniere proelium contra Israel. Intonuit autem Dominus fragore magno in die illa super Philisthim et exterruit eos, et caesi sunt a facie Israel.
1SAM|7|11|Egressique viri Israel de Maspha persecuti sunt Philisthaeos et percusserunt eos usque ad locum, qui erat subter Bethchar.
1SAM|7|12|Tulit autem Samuel lapidem unum et posuit eum inter Maspha et inter Sen et vocavit nomen loci illius Abenezer (id est Lapis adiutorii) dixitque: " Hucusque auxiliatus est nobis Dominus ".
1SAM|7|13|Et humiliati sunt Philisthim nec apposuerunt ultra ut venirent in terminos Israel. Facta est itaque manus Domini super Philisthaeos cunctis diebus Samuel.
1SAM|7|14|Et redditae sunt urbes, quas tulerant Philisthim ab Israel, Israeli ab Accaron usque Geth; et terminos earum liberavit Israel de manu Philisthinorum. Eratque pax inter Israel et Amorraeum.
1SAM|7|15|Iudicabat quoque Samuel Israel cunctis diebus vitae suae
1SAM|7|16|et ibat per singulos annos circumiens Bethel et Galgala et Maspha et iudicabat Israelem in supradictis locis. Revertebaturque in Rama; ibi enim erat domus eius, et ibi iudicabat Israelem. Aedificavit etiam ibi altare Domino.
1SAM|8|1|Factum est autem cum senuis set, Samuel posuit filios suos iu dices Israel.
1SAM|8|2|Fuitque nomen filii eius primogeniti Ioel et nomen secundi Abia; iudicabant in Bersabee.
1SAM|8|3|Et non ambulaverunt filii illius in viis eius, sed declinaverunt post avaritiam acceperuntque munera et perverterunt iudicium.
1SAM|8|4|Congregati ergo universi maiores natu Israel venerunt ad Samuel in Rama
1SAM|8|5|dixeruntque ei: " Ecce tu senuisti, et filii tui non ambulant in viis tuis; nunc ergo constitue nobis regem, ut iudicet nos, sicut universae habent nationes ".
1SAM|8|6|Displicuitque sermo in oculis Samuelis, eo quod dixissent: " Da nobis regem, ut iudicet nos ". Et oravit Samuel ad Dominum.
1SAM|8|7|Dixit autem Dominus ad Samuel: " Audi vocem populi in omnibus, quae loquuntur tibi; non enim te abiecerunt, sed me abiecerunt, ne regnem super eos.
1SAM|8|8|Iuxta omnia opera sua, quae fecerunt a die, qua eduxi eos de Aegypto, usque ad diem hanc, sicut dereliquerunt me et servierunt diis alienis, sic faciunt etiam tibi.
1SAM|8|9|Nunc ergo audi vocem eorum; verumtamen contestare eos et praedic eis ius regis, qui regnaturus est super eos ".
1SAM|8|10|Dixit itaque Samuel omnia verba Domini ad populum, qui petierat a se regem,
1SAM|8|11|et ait: " Hoc erit ius regis, qui imperaturus est vobis: Filios vestros tollet et ponet in curribus suis facietque sibi equites, et current ante quadrigas eius;
1SAM|8|12|et constituet sibi tribunos et centuriones et aratores agrorum suorum et messores segetum et fabros armorum et curruum suorum.
1SAM|8|13|Filias quoque vestras faciet sibi unguentarias et focarias et panificas.
1SAM|8|14|Agros quoque vestros et vineas et oliveta optima tollet et dabit servis suis.
1SAM|8|15|Sed et segetes vestras et vinearum reditus addecimabit, ut det eunuchis et famulis suis.
1SAM|8|16|Servos etiam vestros et ancillas et boves vestros optimos et asinos auferet et ponet in opere suo.
1SAM|8|17|Greges vestros addecimabit, vosque eritis ei servi.
1SAM|8|18|Et clamabitis in die illa a facie regis vestri, quem elegistis vobis, et non exaudiet vos Dominus in die illa ".
1SAM|8|19|Noluit autem populus audire vocem Samuel, sed dixerunt: " Nequaquam: rex enim erit super nos,
1SAM|8|20|et erimus nos quoque sicut omnes gentes; et iudicabit nos rex noster et egredietur ante nos et pugnabit bella nostra pro nobis ".
1SAM|8|21|Et audivit Samuel omnia verba populi et locutus est ea in auribus Domini.
1SAM|8|22|Dixit autem Dominus ad Samuel: " Audi vocem eorum et constitue super eos regem ". Et ait Samuel ad viros Israel: " Vadat unusquisque in civitatem suam ".
1SAM|9|1|Et erat vir de Beniamin nomine Cis filius Abiel filii Seror filii Be chorath filii Aphia, Beniaminita vir potens.
1SAM|9|2|Et erat ei filius vocabulo Saul electus et bonus, et non erat vir de filiis Israel melior illo; ab umero et sursum eminebat super omnem populum.
1SAM|9|3|Perierant autem asinae Cis patris Saul, et dixit Cis ad Saul filium suum: " Tolle tecum unum de pueris et consurgens vade et quaere asinas ". Qui cum transissent per montem Ephraim
1SAM|9|4|et per terram Salisa et non invenissent, transierunt etiam per terram Salim, et non erant, sed et per terram Iemini et minime reppererunt.
1SAM|9|5|Cum autem venissent in terram Suph, dixit Saul ad puerum suum, qui erat cum eo: " Veni, et revertamur, ne forte dimiserit pater meus asinas et sollicitus sit pro nobis ".
1SAM|9|6|Qui ait ei: " Ecce est vir Dei in civitate hac, vir nobilis. Omne quod loquitur, absque ambiguitate venit. Nunc ergo eamus illuc, si forte indicet nobis de via nostra, propter quam venimus ".
1SAM|9|7|Dixitque Saul ad puerum suum: " Ecce ibimus; quid feremus ad virum? Panis defecit in sitarciis nostris, et sportulam non habemus, ut demus homini Dei. Quid habemus? ".
1SAM|9|8|Rursum puer respondit Sauli et ait: " Ecce inventa est in manu mea quarta pars sicli argenti; demus homini Dei, ut indicet nobis viam nostram. -
1SAM|9|9|Olim in Israel sic loquebatur unusquisque vadens consulere Deum: " Venite, et eamus ad videntem "; qui enim propheta dicitur hodie, vocabatur olim videns. -
1SAM|9|10|Et dixit Saul ad puerum suum: " Optimus sermo tuus; veni, eamus ". Et ierunt in civitatem, in qua erat vir Dei.
1SAM|9|11|Cumque ascenderent clivum civitatis, invenerunt puellas egredientes ad hauriendam aquam et dixerunt eis: " Num hic est videns? ".
1SAM|9|12|Quae respondentes dixerunt illis: " Hic est: ecce ante te, festina nunc; hodie enim venit in civitatem, quia sacrificium est hodie populo in excelso.
1SAM|9|13|Ingredientes urbem statim invenietis eum, antequam ascendat excelsum ad vescendum; neque enim comesurus est populus, donec ille veniat, quia ipse benedicit hostiae, et deinceps comedunt, qui vocati sunt. Nunc ergo conscendite, quia statim reperietis eum ".
1SAM|9|14|Et ascenderunt in civitatem. Cumque illi intrarent in urbem, apparuit Samuel egrediens obviam eis, ut ascenderet in excelsum.
1SAM|9|15|Dominus autem revelaverat Samuel, ante unam diem quam veniret Saul, dicens:
1SAM|9|16|" Hac ipsa, quae nunc est hora, cras mittam ad te virum de terra Beniamin, et unges eum ducem super populum meum Israel, et salvabit populum meum de manu Philisthinorum, quia respexi populum meum; venit enim clamor eorum ad me ".
1SAM|9|17|Cumque aspexisset Samuel Saulem, Dominus ait ei: " Ecce vir, quem dixeram tibi; iste dominabitur populo meo ".
1SAM|9|18|Accessit autem Saul ad Samuelem in medio portae et ait: " Indica, oro, mihi: Ubi est domus videntis? ".
1SAM|9|19|Et respondit Samuel Sauli dicens: " Ego sum videns. Ascende ante me in excelsum, ut comedatis mecum hodie. Et dimittam te mane et omnia, quae sunt in corde tuo, indicabo tibi;
1SAM|9|20|et de asinis, quas perdidisti nudiustertius, ne sollicitus sis, quia inventae sunt. Et cuius erunt optima quaeque Israel? Nonne tibi et omni domui patris tui? ".
1SAM|9|21|Respondens autem Saul ait: "Numquid non Beniaminita ego sum de minima tribu Israel, et cognatio mea novissima inter omnes familias de tribu Beniamin? Quare ergo locutus es mihi sermonem istum? ".
1SAM|9|22|Assumens itaque Samuel Saulem et puerum eius introduxit eos in triclinium et dedit eis locum in capite eorum, qui fuerant invitati: erant enim quasi triginta viri.
1SAM|9|23|Dixitque Samuel coco: " Da partem, quam dedi tibi et praecepi, ut reponeres seorsum apud te ".
1SAM|9|24|Levavit autem cocus armum et caudam et posuit ante Saul. Dixitque Samuel: " Ecce quod remansit; pone ante te et comede, quia de industria servatum est tibi, quando populum vocavi ". Et comedit Saul cum Samuel in die illa.
1SAM|9|25|Et descenderunt de excelso in oppidum. Et straverunt pro Saul in solario, et dormivit.
1SAM|9|26|Cumque mane surrexissent, et iam elucesceret, vocavit Samuel Saul in solario dicens: " Surge, ut dimittam te ". Et surrexit Saul. Egressique sunt ambo, ipse videlicet et Samuel.
1SAM|9|27|Cumque descenderent in extrema parte civitatis, Samuel dixit ad Saul: " Dic puero, ut antecedat nos - et ille antecessit C; tu autem subsiste paulisper, ut indicem tibi verbum Domini ".
1SAM|10|1|Tulit autem Samuel lenticulam olei et effudit super caput eius et deosculatus eum ait: " Ecce unxit te Dominus in principem super populum suum, super Israel. Et tu dominaberis populo Domini et tu liberabis eum de manu inimicorum eius, qui in circuitu eius sunt. Et hoc tibi signum quia unxit te Deus in principem super hereditatem suam:
1SAM|10|2|cum abieris hodie a me, invenies duos viros iuxta sepulcrum Rachel in finibus Beniamin, dicentque tibi: "Inventae sunt asinae, ad quas ieras perquirendas; et intermissis pater tuus asinis sollicitus est pro vobis et dicit: Quid faciam de filio meo?".
1SAM|10|3|Cumque abieris inde et ultra transieris et veneris ad quercum Thabor, invenient te ibi tres viri ascendentes ad Deum in Bethel: unus portans tres haedos et alius tres tortas panis et alius portans utrem vini.
1SAM|10|4|Cumque te salutaverint, dabunt tibi duos panes, et accipies de manu eorum.
1SAM|10|5|Post haec venies in Gabaa Dei, ubi est statio Philisthinorum; et, cum ingressus fueris ibi urbem, obviam habebis gregem prophetarum descendentium de excelso et ante eos psalterium et tympanum et tibiam et citharam ipsosque prophetantes.
1SAM|10|6|Et insiliet in te spiritus Domini, et prophetabis cum eis et mutaberis in virum alium.
1SAM|10|7|Quando ergo evenerint signa haec omnia tibi, fac, quaecumque invenerit manus tua, quia Dominus tecum est.
1SAM|10|8|Et descendes ante me in Galgala. Ego quippe descendam ad te, ut offeram oblationem et immolem victimas pacificas. Septem diebus exspectabis, donec veniam ad te et ostendam tibi, quae facias ".
1SAM|10|9|Itaque, cum avertisset umerum suum, ut abiret a Samuele, immutavit ei Deus cor aliud, et venerunt omnia signa haec in die illa.
1SAM|10|10|Veneruntque inde in Gabaa, et ecce grex prophetarum obvius ei; et insiluit super eum spiritus Dei, et prophetavit in medio eorum.
1SAM|10|11|Videntes autem omnes, qui noverant eum heri et nudiustertius, quod esset cum prophetis et prophetaret, dixerunt ad invicem: " Quaenam res accidit filio Cis? Num et Saul inter prophetas? ".
1SAM|10|12|Responditque vir loci illius dicens: " Et quis pater eorum? ". Propterea versum est in proverbium: " Num et Saul inter prophetas? ".
1SAM|10|13|Cessavit autem prophetare et venit in Gabaa;
1SAM|10|14|dixitque patruus Saul ad eum et ad puerum eius: " Quo abistis? ". Qui respondit: " Quaerere asinas; quas cum non repperissemus, venimus ad Samuelem".
1SAM|10|15|Et dixit ei patruus suus: "Indica mihi quid dixerit tibi Samuel".
1SAM|10|16|Et ait Saul ad patruum suum: " Indicavit nobis quia inventae essent asinae ". De sermone autem regni non indicavit ei, quem locutus illi fuerat Samuel.
1SAM|10|17|Et convocavit Samuel populum ad Dominum in Maspha
1SAM|10|18|et ait ad filios Israel: " Haec dicit Dominus, Deus Israel: Ego eduxi Israel de Aegypto et erui vos de manu Aegyptiorum et de manu omnium regnorum, quae affligebant vos.
1SAM|10|19|Vos autem hodie proiecistis Deum vestrum, qui solus salvavit vos de universis malis et tribulationibus vestris, et dixistis: "Nequaquam, sed regem constitue super nos!". Nunc ergo state coram Domino per tribus vestras et per familias ".
1SAM|10|20|Et applicuit Samuel omnes tribus Israel; et cecidit sors in tribum Beniamin.
1SAM|10|21|Et applicuit tribum Beniamin et cognationes eius; et cecidit in cognationem Metri et pervenit usque ad Saul filium Cis. Quaesierunt ergo eum, et non est inventus.
1SAM|10|22|Et consuluerunt post haec Dominum, utrumnam venisset illuc vir. Responditque Dominus: " Ecce absconditus est inter sarcinas ".
1SAM|10|23|Cucurrerunt itaque et tulerunt eum inde; stetitque in medio populi et altior fuit universo populo ab umero et sursum.
1SAM|10|24|Et ait Samuel ad omnem populum: Certe videtis, quem elegit Dominus, quoniam non sit similis ei in omni populo ". Et clamavit cunctus populus et ait: " Vivat rex! ".
1SAM|10|25|Locutus est autem Samuel ad populum legem regni et scripsit in libro et reposuit coram Domino; et dimisit Samuel omnem populum, singulos in domum suam.
1SAM|10|26|Sed et Saul abiit in domum suam in Gabaa; et abierunt cum eo viri fortes, quorum tetigerat Deus corda.
1SAM|10|27|Filii vero Belial dixerunt: " Num salvare nos poterit iste? ". Et despexerunt eum et non attulerunt ei munera; ille vero dissimulabat se audire.
1SAM|11|1|Ascendit autem Naas Am monites et pugnare coepit ad versum Iabes Galaad. Dixeruntque omnes viri Iabes ad Naas: " Habeto nos foederatos, et serviemus tibi ".
1SAM|11|2|Et respondit ad eos Naas Ammonites: " In hoc feriam vobiscum foedus, ut eruam omnium vestrum oculos dextros ponamque vos opprobrium in universo Israel ".
1SAM|11|3|Et dixerunt ad eum seniores Iabes: " Concede nobis septem dies, ut mittamus nuntios in universos terminos Israel; et, si non fuerit qui defendat nos, egrediemur ad te ".
1SAM|11|4|Venerunt ergo nuntii in Gabaa Saulis et locuti sunt verba audiente populo; et levavit omnis populus vocem suam et flevit.
1SAM|11|5|Et ecce Saul veniebat sequens boves de agro et ait: " Quid habet populus quod plorat? ". Et narraverunt ei verba virorum Iabes.
1SAM|11|6|Et insilivit spiritus Domini in Saul, cum audisset verba haec; et iratus est furor eius nimis.
1SAM|11|7|Et assumens par boum concidit in frusta misitque in omnes terminos Israel per manum nuntiorum dicens: " Quicumque non exierit secutusque fuerit Saul et Samuel, sic fiet bobus eius ". Invasit ergo timor Domini populum, et egressi sunt quasi vir unus.
1SAM|11|8|Et recensuit eos in Bezec: fueruntque filiorum Israel trecenta milia; virorum autem Iudae triginta milia.
1SAM|11|9|Et dixit nuntiis, qui venerant: " Sic dicetis viris, qui sunt in Iabes Galaad: Cras erit vobis salus, cum incaluerit sol ". Venerunt ergo nuntii et annuntiaverunt viris Iabes, qui laetati sunt
1SAM|11|10|et dixerunt: "Mane exibimus ad vos, et facietis nobis omne, quod placuerit vobis ".
1SAM|11|11|Et factum est, cum venisset dies crastinus, constituit Saul populum in tres partes; et ingressi sunt media castra in vigilia matutina et percusserunt Ammon, usque dum incalesceret dies. Reliqui autem dispersi sunt, ita ut non relinquerentur in eis duo pariter.
1SAM|11|12|Et ait populus ad Samuel: " Quis est iste qui dixit: "Saul num regnabit super nos?". Date viros, et interficiemus eos ".
1SAM|11|13|Et ait Saul: " Non occidetur quisquam in die hac, quia hodie fecit Dominus salutem in Israel".
1SAM|11|14|Dixit autem Samuel ad populum: " Venite, et eamus in Galgala et innovemus ibi regnum ".
1SAM|11|15|Et perrexit omnis populus in Galgala, et fecerunt ibi regem Saul coram Domino in Galgala; et immolaverunt ibi victimas pacificas coram Domino. Et laetatus est ibi Saul et cuncti viri Israel nimis.
1SAM|12|1|Dixit autem Samuel ad universum Israel: " Ecce audivi vocem vestram iuxta omnia, quae locuti estis ad me, et constitui super vos regem;
1SAM|12|2|et nunc rex graditur ante vos. Ego autem senui et incanui; porro filii mei vobiscum sunt. Itaque conversatus coram vobis ab adulescentia mea usque ad hanc diem;
1SAM|12|3|ecce praesto sum. Loquimini contra me coram Domino et coram christo eius, utrum bovem cuiusquam tulerim an asinum, si quempiam calumniatus sum, si oppressi aliquem, si de manu cuiusquam munus accepi, ut oculos meos clauderem in eius causa. Restituam vobis ".
1SAM|12|4|Et dixerunt: " Non es calumniatus nos neque oppressisti neque tulisti de manu alicuius quippiam ".
1SAM|12|5|Dixitque ad eos: " Testis Dominus adversum vos, et testis christus eius in die hac, quia non inveneritis in manu mea quippiam ". Et dixerunt: " Testis ".
1SAM|12|6|Et ait Samuel ad populum: " Testis est Dominus, qui fecit Moysen et Aaron et eduxit patres nostros de terra Aegypti.
1SAM|12|7|Nunc ergo state, ut iudicio contendam adversum vos coram Domino de omnibus misericordiis Domini, quas fecit vobiscum et cum patribus vestris:
1SAM|12|8|quomodo ingressus est Iacob in Aegyptum, et oppresserunt eos Aegyptii; et clamaverunt patres vestri ad Dominum, et misit Dominus Moysen et Aaron et eduxit patres vestros ex Aegypto et collocavit eos in loco hoc;
1SAM|12|9|qui obliti sunt Domini Dei sui, et tradidit eos in manu Sisarae magistri militiae Asor et in manu Philisthinorum et in manu regis Moab, et pugnaverunt adversum eos.
1SAM|12|10|Postea autem clamaverunt ad Dominum et dixerunt: "Peccavimus, quia dereliquimus Dominum et servivimus Baalim et Astharoth; nunc ergo erue nos de manu inimicorum nostrorum, et serviemus tibi".
1SAM|12|11|Et misit Dominus Ierobbaal et Barac et Iephte et Samuel et eruit vos de manu inimicorum vestrorum per circuitum; et habitastis confidenter.
1SAM|12|12|Videntes autem quod Naas rex filiorum Ammon venisset adversum vos, dixistis mihi: "Nequaquam, sed rex imperabit nobis!", cum Dominus Deus vester regnaret in vobis.
1SAM|12|13|Nunc ergo praesto est rex vester, quem elegistis et petistis; ecce dedit vobis Dominus regem.
1SAM|12|14|Si timueritis Dominum et servieritis ei et audieritis vocem eius et non contempseritis sermonem Domini, eritis et vos et rex, qui imperat vobis, sequentes Dominum Deum vestrum.
1SAM|12|15|Si autem non audieritis vocem Domini, sed contempseritis sermonem Domini, erit manus Domini super vos et super regem vestrum, ut disperdat vos.
1SAM|12|16|Sed et nunc state et videte rem istam grandem, quam facturus est Dominus in conspectu vestro.
1SAM|12|17|Numquid non messis tritici est hodie? Invocabo Dominum, et dabit tonitrua et pluvias; et scietis et videbitis quia grande malum feceritis vobis in conspectu Domini petentes super vos regem ".
1SAM|12|18|Et clamavit Samuel ad Dominum, et dedit Dominus tonitrua et pluviam in die illa.
1SAM|12|19|Et timuit omnis populus nimis Dominum et Samuel; dixitque universus populus ad Samuel: " Ora pro servis tuis ad Dominum Deum tuum, ut non moriamur: addidimus enim universis peccatis nostris malum, ut peteremus nobis regem ".
1SAM|12|20|Dixit autem Samuel ad populum: " Nolite timere. Vos fecistis universum malum hoc; verumtamen nolite recedere a tergo Domini et servite Domino in omni corde vestro;
1SAM|12|21|et nolite declinare post vana, quae non proderunt vobis neque eruent vos, quia vana sunt;
1SAM|12|22|profecto non derelinquet Dominus populum suum propter nomen suum magnum, quia dignatus est Dominus facere vos sibi populum.
1SAM|12|23|Absit autem a me hoc peccatum in Dominum, ut cessem orare pro vobis et docere vos viam bonam et rectam.
1SAM|12|24|Igitur timete Dominum et servite ei in veritate et ex toto corde vestro; vidistis enim magnifica, quae in vobis gesserit.
1SAM|12|25|Quod si perseveraveritis in malitia, et vos et rex vester pariter peribitis ".
1SAM|13|1|Filius annorum Saul, cum regnare coepisset; duobus au tem annis regnavit super Israel.
1SAM|13|2|Et elegit sibi Saul tria milia de Israel: et erant cum Saul duo milia in Machmas et in monte Bethel, mille autem cum Ionathan in Gabaa Beniamin. Porro ceterum populum remisit unumquemque in tabernacula sua.
1SAM|13|3|Et percussit Ionathan stationem Philisthinorum, quae erat in Gabaa. Quod audierunt Philisthim; Saul autem cecinit bucina in omni terra dicens: " Audiant Hebraei! ".
1SAM|13|4|Et universus Israel audivit huiuscemodi famam: " Percussit Saul stationem Philisthinorum; et factus est Israel odiosus Philisthim ". Ergo populus congregatus est post Saul in Galgala.
1SAM|13|5|Et Philisthim congregati sunt ad proeliandum contra Israel: tria milia curruum et sex milia equitum et reliquum vulgus plurimum sicut arena, quae est in litore maris. Et ascendentes castrametati sunt in Machmas ad orientem Bethaven.
1SAM|13|6|Quod cum vidissent viri Israel se in arto sitos - afflictus est enim populus - absconderunt se in speluncis et in abditis, in petris quoque et in antris et in cisternis.
1SAM|13|7|Hebraei autem transierunt Iordanem in terram Gad et Galaad.Cumque adhuc esset Saul in Galgalis, universus populus perterritus est, qui sequebatur eum.
1SAM|13|8|Et exspectavit septem diebus iuxta placitum Samuel, et non venit Samuel in Galgala; dilapsusque est populus ab eo.
1SAM|13|9|Ait ergo Saul: " Afferte mihi holocaustum et pacifica ". Et obtulit holocaustum.
1SAM|13|10|Cumque complesset offerens holocaustum, ecce Samuel veniebat; et egressus est Saul obviam ei, ut salutaret eum.
1SAM|13|11|Locutusque est ad eum Samuel: " Quid fecisti? ". Respondit Saul: " Quia vidi quod dilaberetur populus a me, et tu non veneras iuxta placitos dies, porro Philisthim congregati fuerant in Machmas,
1SAM|13|12|dixi: Nunc descendent Philisthim ad me in Galgala, et faciem Domini non placavi. Necessitate compulsus obtuli holocaustum ".
1SAM|13|13|Dixitque Samuel ad Saul: " Stulte egisti. Utinam custodisses mandata Domini Dei tui, quae praecepit tibi! Profecto nunc confirmasset Dominus regnum tuum super Israel in sempiternum;
1SAM|13|14|sed nequaquam regnum tuum ultra consurget. Quaesivit sibi Dominus virum iuxta cor suum; et constituit eum Dominus ducem super populum suum, eo quod non servaveris, quae praecepit Dominus ".
1SAM|13|15|Surrexit autem Samuel et ascendit de Galgalis et abiit per viam suam. Et reliquus populus ascendit post Saul obviam exercitui bellatorum. Et venerunt de Galgalis in Gabaa Beniamin. Et recensuit Saul populum, qui inventi fuerant cum eo, quasi sescentos viros.
1SAM|13|16|Et Saul et Ionathan filius eius populusque, qui erat cum eis, erat in Gabaa Beniamin; porro Philisthim consederant in Machmas.
1SAM|13|17|Et egressi sunt ad praedandum de castris Philisthinorum tres cunei: unus cuneus pergebat contra viam Ophra ad terram Sual,
1SAM|13|18|porro alius ingrediebatur per viam Bethoron, tertius autem verterat se ad iter termini imminentis valli Seboim contra desertum.
1SAM|13|19|Porro faber ferrarius non inveniebatur in omni terra Israel; caverant enim Philisthim, ne forte facerent Hebraei gladium aut lanceam.
1SAM|13|20|Descendebat ergo omnis Israel ad Philisthim, ut exacueret unusquisque vomerem suum et ligonem et securim et falcem.
1SAM|13|21|Pretium autem exacutionis erat: pro vomeribus et ligonibus duae partes sicli, et tertia pars sicli ad acuendas secures et ad stimulum corrigendum.
1SAM|13|22|Cumque venisset dies proelii Machmas, non est inventus ensis et lancea in manu totius populi, qui erat cum Saul et cum Ionathan, excepto Saul et Ionathan filio eius.
1SAM|13|23|Egressa est autem statio Philisthim ad fauces Machmas.
1SAM|14|1|Et accidit quadam die, ut diceret Ionathan filius Saul ad adulescentem armigerum suum: " Veni, et transeamus ad stationem Philisthim, quae est ibi ex adverso ". Patri autem suo hoc ipsum non indicavit.
1SAM|14|2|Porro Saul morabatur in extrema parte Gabaa sub malogranato, quae erat in Magron; et erat populus cum eo quasi sescentorum virorum.
1SAM|14|3|Et Ahias filius Achitob fratris Ichabod filii Phinees, qui ortus fuerat ex Heli sacerdote Domini in Silo, portabat ephod. Sed et populus ignorabat quod isset Ionathan.
1SAM|14|4|Erant autem inter ascensus, per quos nitebatur Ionathan transire ad stationem Philisthinorum, dens rupis hinc ex una parte et dens rupis illinc ex altera parte: nomen uni Boses et nomen alteri Sene;
1SAM|14|5|unus scopulus prominens ad aquilonem ex adverso Machmas et alter a meridie contra Gabaa.
1SAM|14|6|Dixit autem Ionathan ad adulescentem armigerum suum: " Veni, transeamus ad stationem incircumcisorum horum, si forte faciat Dominus pro nobis; quia non est Domino difficile salvare vel in multitudine vel in paucis ".
1SAM|14|7|Dixitque ei armiger suus: " Fac omnia, quae placent animo tuo. Perge quo cupis; ego ero tecum ubicumque volueris ".
1SAM|14|8|Et ait Ionathan: " Ecce nos transimus ad viros istos. Cumque apparuerimus eis,
1SAM|14|9|si taliter locuti fuerint ad nos: "Manete, donec veniamus ad vos", stemus in loco nostro nec ascendamus ad eos.
1SAM|14|10|Si autem dixerint: "Ascendite ad nos", ascendamus, quia tradidit eos Dominus in manibus nostris; hoc erit nobis signum ".
1SAM|14|11|Apparuit igitur uterque stationi Philisthinorum. Dixeruntque Philisthim: " En Hebraei egrediuntur de cavernis, in quibus absconditi fuerant ".
1SAM|14|12|Et locuti sunt viri de statione ad Ionathan et ad armigerum eius dixeruntque: " Ascendite ad nos, et ostendimus vobis rem ". Et ait Ionathan ad armigerum suum: " Ascendamus; sequere me, tradidit enim eos Dominus in manu Israel ".
1SAM|14|13|Ascendit autem Ionathan reptans manibus et pedibus et armiger eius post eum; Philisthim cadebant ante Ionathan, et eos armiger eius interficiebat sequens eum.
1SAM|14|14|Et facta est plaga prima, qua percussit Ionathan et armiger eius quasi viginti viros in media fere parte iugeri.
1SAM|14|15|Et factus est terror in castris per agros; sed et omnis populus stationis eorum et, qui ierant ad praedandum, obstupuerunt; et conturbata est terra, et factus est terror a Deo.
1SAM|14|16|Et respexerunt speculatores Saul, qui erant in Gabaa Beniamin; et ecce multitudo fluctuabat huc illucque diffugiens.
1SAM|14|17|Et ait Saul populo, qui erat cum eo: " Requirite et videte quis abierit ex nobis ". Cumque requisissent, repertum est non adesse Ionathan et armigerum eius.
1SAM|14|18|Et ait Saul ad Ahiam: " Applica ephod ". Ipse enim portabat ephod in die illa in conspectu filiorum Israel.
1SAM|14|19|Cumque loqueretur Saul ad sacerdotem, tumultus maior fiebat in castris Philisthinorum, crescebatque paulatim et clarius reboabat. Et ait Saul ad sacerdotem: " Contrahe manum tuam ".
1SAM|14|20|Congregati ergo sunt Saul et omnis populus, qui erat cum eo, et venerunt usque ad locum certaminis. Et ecce versus fuerat gladius uniuscuiusque ad proximum suum: perturbatio magna nimis.
1SAM|14|21|Sed et Hebraei, qui fuerant cum Philisthim heri et nudiustertius ascenderantque cum eis in castris, reversi sunt et ipsi, ut essent cum Israel, qui erant cum Saul et Ionathan.
1SAM|14|22|Omnes quoque Israelitae, qui se absconderant in monte Ephraim, audientes quod fugissent Philisthim, sociaverunt se et ipsi cum suis in proelio.
1SAM|14|23|Et salvavit Dominus in die illa Israel; pugna autem pervenit ultra Bethaven.
1SAM|14|24|Et viri Israel comprimebant se in die illa. Adiuravit autem Saul populum dicens: " Maledictus vir, qui comederit panem usque ad vesperam, donec ulciscar de inimicis meis! ". Et non manducavit universus populus panem.
1SAM|14|25|Omneque terrae vulgus venit in saltum, in quo erat mel super faciem agri.
1SAM|14|26|Ingressus est itaque populus saltum, et apparuit fluens mel. Nullusque applicuit manum ad os suum; timebat enim populus iuramentum.
1SAM|14|27|Porro Ionathan non audierat, cum adiuraret pater eius populum; extenditque summitatem virgae, quam habebat in manu, et intinxit in favo mellis et convertit manum suam ad os suum, et illuminati sunt oculi eius.
1SAM|14|28|Respondensque unus de populo ait: " Iureiurando constrinxit pater tuus populum dicens: "Maledictus, qui comederit panem hodie!". Defecit autem populus ".
1SAM|14|29|Dixitque Ionathan: " Turbavit pater meus terram! Videte quia illuminati sunt oculi mei, eo quod gustaverim paululum de melle isto;
1SAM|14|30|quanto magis si comedisset hodie populus de praeda inimicorum suorum, quam repperit? Nonne nunc maior facta fuisset plaga in Philisthim? ".
1SAM|14|31|Percusserunt ergo in die illa Philisthaeos a Machmis usque in Aialon; defatigatus est autem populus nimis.
1SAM|14|32|Et versus ad praedam tulit oves et boves et vitulos; et mactaverunt in terra, comeditque populus cum sanguine.
1SAM|14|33|Nuntiaverunt autem Saul dicentes: " Ecce populus peccat Domino comedens cum sanguine ". Qui ait: " Praevaricati estis! Volvite ad me huc saxum grande ".
1SAM|14|34|Et dixit Saul: " Dispergimini in vulgus et dicite eis, ut adducat ad me unusquisque bovem suum et arietem, et occidite super istud et vescimini; et non peccabitis Domino comedentes cum sanguine ". Adduxit itaque omnis populus, unusquisque quod erat in manu sua illa nocte, et occiderunt ibi.
1SAM|14|35|Aedificavit autem Saul altare Domino. Tuncque primum coepit aedificare altare Domino.
1SAM|14|36|Et dixit Saul: " Irruamus super Philisthim nocte et vastemus eos, usquedum illucescat mane; nec relinquamus de eis virum ". Dixitque populus: " Omne, quod bonum videtur in oculis tuis, fac ". Et ait sacerdos: " Accedamus huc ad Deum ".
1SAM|14|37|Et consuluit Saul Deum: " Num persequar Philisthim? Numquid trades eos in manu Israel? ". Et non respondit ei in die illa.
1SAM|14|38|Dixitque Saul: " Accedite huc, universi duces populi, et scitote et videte per quem acciderit peccatum hoc hodie.
1SAM|14|39|Vivit Dominus, salvator Israel, quia si per Ionathan filium meum factum est, absque retractatione morietur ". Ad quod nullus contradixit ei de omni populo.
1SAM|14|40|Et ait ad universum Israel: " Separamini vos in partem unam, et ego cum Ionathan filio meo ero in parte altera ". Respondit populus ad Saul: " Quod bonum videtur in oculis tuis, fac ".
1SAM|14|41|Et dixit Saul ad Dominum, Deum Israel: " Quid est quod non responderis servo tuo hodie? Si est in me aut in Ionathan filio meo iniquitas ista, Domine, Deus Israel, da Urim; sed, si est haec iniquitas in populo tuo Israel, da Tummim ". Et deprehensus est Ionathan et Saul; populus autem salvus evasit.
1SAM|14|42|Et ait Saul: " Mittite sortem inter me et inter Ionathan filium meum ". Et captus est Ionathan.
1SAM|14|43|Dixit autem Saul ad Ionathan: " Indica mihi quid feceris ". Et indicavit ei Ionathan et ait: " Gustans gustavi in summitate virgae, quae erat in manu mea, paululum mellis et ecce ego morior ".
1SAM|14|44|Et ait Saul: " Haec faciat mihi Deus et haec addat, nisi morte morieris, Ionathan ".
1SAM|14|45|Dixitque populus ad Saul: " Ergone Ionathan morietur, qui fecit salutem hanc magnam in Israel? Hoc nefas est; vivit Dominus, quia non cadet capillus de capite eius in terram, quia cum Deo operatus est hodie ". Liberavit ergo populus Ionathan, ut non moreretur.
1SAM|14|46|Recessitque Saul nec persecutus est Philisthim; porro Philisthim abierunt in loca sua.
1SAM|14|47|At Saul, confirmato regno super Israel, pugnabat per circuitum adversum omnes inimicos eius: contra Moab et filios Ammon et Edom et reges Soba et Philisthaeos; et, quocumque se verterat, superabat.
1SAM|14|48|Fortiter egit et percussit Amalec et eruit Israel de manu vastatorum eius.
1SAM|14|49|Fuerunt autem filii Saul Ionathan et Isui et Melchisua. Nomina duarum filiarum eius: nomen primogenitae Merob et nomen minoris Michol.
1SAM|14|50|Et nomen uxoris Saul Achinoam filia Achimaas, et nomen principis militiae eius Abner filius Ner patrui Saul.
1SAM|14|51|Porro Cis pater Saul et Ner pater Abner fuerunt filii Abiel.
1SAM|14|52|Erat autem bellum potens adversum Philisthaeos omnibus diebus Saul; nam, quemcumque viderat Saul virum fortem et aptum ad proelium, sociabat eum sibi.
1SAM|15|1|Et dixit Samuel ad Saul: " Me misit Dominus, ut unge rem te in regem super populum eius Israel. Nunc ergo audi vocem Domini.
1SAM|15|2|Haec dicit Dominus exercituum: "Recensui, quaecumque fecit Amalec Israeli, quomodo restitit ei in via, cum ascenderet de Aegypto.
1SAM|15|3|Nunc igitur vade et demolire Amalec et percute anathemate universa eius; non parcas ei, sed interfice a viro usque ad mulierem et parvulum atque lactantem, bovem et ovem, camelum et asinum" ".
1SAM|15|4|Convocavit itaque Saul populum et recensuit eos in Telem: ducenta milia peditum et decem milia virorum Iudae.
1SAM|15|5|Cumque venisset Saul usque ad civitatem Amalec, tetendit insidias in torrente
1SAM|15|6|dixitque Saul Cinaeo: " Abite, recedite atque descendite ab Amalec, ne forte perdam te cum eo; tu enim fecisti misericordiam cum omnibus filiis Israel, cum ascenderent de Aegypto ". Et recessit Cinaeus de medio Amalec.
1SAM|15|7|Percussitque Saul Amalec ab Hevila usque ad Sur, quae est e regione Aegypti.
1SAM|15|8|Et apprehendit Agag regem Amalec vivum; omne autem vulgus interfecit in ore gladii.
1SAM|15|9|Et pepercit Saul et populus Agag et optimis gregibus ovium et armentorum, pinguibus scilicet pecoribus et agnis et universis, quae pulchra erant, nec voluerunt disperdere ea; quidquid vero vile fuit et reprobum, hoc demoliti sunt.
1SAM|15|10|Factum est autem verbum Domini ad Samuel dicens:
1SAM|15|11|" Paenitet me quod constituerim Saul regem, quia dereliquit me et verba mea opere non implevit ". Contristatusque est Samuel et clamavit ad Dominum tota nocte.
1SAM|15|12|Cumque de nocte surrexisset Samuel, ut iret ad Saul mane, nuntiatum est Samueli quod venisset Saul in Carmel et erexisset sibi trophaeum et reversus transisset descendissetque in Galgala.
1SAM|15|13|Et cum venisset Samuel ad Saul, dixit ei Saul: " Benedictus tu Domino; implevi verbum Domini ".
1SAM|15|14|Dixitque Samuel: " Et quae est haec vox gregum, quae resonat in auribus meis, et armentorum, quam ego audio? ".
1SAM|15|15|Et ait Saul: " De Amalec adduxerunt ea; pepercit enim populus melioribus ovibus et armentis, ut immolarentur Domino Deo tuo; reliqua vero occidimus ".
1SAM|15|16|Dixit autem Samuel ad Saul: " Sine me, et indicabo tibi, quae locutus sit Dominus ad me nocte ". Dixitque ei: " Loquere ".
1SAM|15|17|Et ait Samuel: " Nonne, cum parvulus esses in oculis tuis, caput in tribubus Israel factus es? Unxitque te Dominus regem super Israel
1SAM|15|18|et misit te Dominus in viam et ait: " Vade et interfice peccatores Amalec et pugnabis contra eos usque ad internecionem eorum ".
1SAM|15|19|Quare ergo non audisti vocem Domini, sed versus ad praedam es et fecisti malum in oculis Domini? ".
1SAM|15|20|Et ait Saul ad Samuelem: " Immo audivi vocem Domini et ambulavi in via, per quam misit me Dominus; et adduxi Agag regem Amalec et Amalec interfeci.
1SAM|15|21|Tulit autem populus de praeda oves et boves, primitias eorum, quae caesa sunt, ut immolet Domino Deo tuo in Galgalis ".
1SAM|15|22|Et ait Samuel: " Numquid vult Dominus holocausta aut victimas et non potius ut oboediatur voci Domini? Melior est enim oboedientia quam victimae, et auscultare magis quam offerre adipem arietum.
1SAM|15|23|Vere peccatum hariolandi est repugnare, et scelus idololatriae nolle acquiescere: pro eo ergo quod abiecisti sermonem Domini, abiecit te, ne sis rex ".
1SAM|15|24|Dixitque Saul ad Samuelem: " Peccavi, quia praevaricatus sum sermonem Domini et verba tua timens populum et oboediens voci eorum;
1SAM|15|25|sed nunc tolle, quaeso, peccatum meum et revertere mecum, ut adorem Dominum ".
1SAM|15|26|Et ait Samuel ad Saul: " Non revertar tecum, quia proiecisti sermonem Domini; et proiecit te Dominus, ne sis rex super Israel ".
1SAM|15|27|Et conversus est Samuel, ut abiret; ille autem apprehendit summitatem pallii eius, quae et scissa est.
1SAM|15|28|Et ait ad eum Samuel: " Scidit Dominus regnum Israel a te hodie et tradidit illud proximo tuo meliori te.
1SAM|15|29|Porro Gloria Israel non mentitur et paenitudine non flectitur; neque enim homo est, ut agat paenitentiam ".
1SAM|15|30|At ille ait: " Peccavi, sed nunc honora me coram senibus populi mei et coram Israel; et revertere mecum, ut adorem Dominum Deum tuum ".
1SAM|15|31|Reversus ergo Samuel secutus est Saulem et adoravit Saul Dominum.
1SAM|15|32|Dixitque Samuel: " Adducite ad me Agag regem Amalec ". Et oblatus est ei Agag tremens. Et dixit Agag: " Certe secessit amaritudo mortis! ".
1SAM|15|33|Et ait Samuel: " Sicut fecit absque liberis mulieres gladius tuus, sic absque liberis erit inter mulieres mater tua ". Et in frusta concidit Samuel Agag coram Domino in Galgalis.
1SAM|15|34|Abiit autem Samuel in Rama; Saul vero ascendit in domum suam in Gabaa Saulis.
1SAM|15|35|Et non vidit Samuel ultra Saul usque ad diem mortis suae; verumtamen lugebat Samuel Saul, quoniam Dominum paenitebat quod constituisset Saul regem super Israel.
1SAM|16|1|Dixitque Dominus ad Samuelem: " Usquequo tu luges Saul, cum ego proiecerim eum, ne regnet super Israel? Imple cornu tuum oleo et veni, ut mittam te ad Isai Bethlehemitem; providi enim in filiis eius mihi regem ".
1SAM|16|2|Et ait Samuel: " Quomodo vadam? Audiet enim Saul et interficiet me ". Et ait Dominus: " Vitulam de armento tolles in manu tua et dices: "Ad immolandum Domino veni".
1SAM|16|3|Et vocabis Isai ad victimam; et ego ostendam tibi quid facias, et unges quemcumque monstravero tibi ".
1SAM|16|4|Fecit ergo Samuel, sicut locutus est ei Dominus, venitque in Bethlehem. Et expaverunt seniores civitatis occurrentes ei dixeruntque: " Pacificusne ingressus tuus? ".
1SAM|16|5|Et ait: " Pacificus; ad immolandum Domino veni. Sanctificamini et venite mecum, ut immolem ". Sanctificavit ergo Isai et filios eius et vocavit eos ad sacrificium.
1SAM|16|6|Cumque ingressi essent, vidit Eliab et ait: " Absque dubio coram Domino est christus eius! ".
1SAM|16|7|Et dixit Dominus ad Samuelem: " Ne respicias vultum eius neque altitudinem staturae eius, quoniam abieci eum; nec iuxta intuitum hominis iudico: homo enim videt ea, quae parent, Dominus autem intuetur cor ".
1SAM|16|8|Et vocavit Isai Abinadab et adduxit eum coram Samuele, qui dixit: " Nec hunc elegit Dominus ".
1SAM|16|9|Adduxit autem Isai Samma, de quo ait: " Etiam hunc non elegit Dominus ".
1SAM|16|10|Adduxit itaque Isai septem filios suos coram Samuele, et ait Samuel ad Isai: " Non elegit Dominus ex istis ".
1SAM|16|11|Dixitque Samuel ad Isai: " Numquid iam completi sunt filii? ". Qui respondit: " Adhuc reliquus est minimus et pascit oves ". Et ait Samuel ad Isai: " Mitte et adduc eum; nec enim discumbemus prius quam huc ille venerit ".
1SAM|16|12|Misit ergo et adduxit eum; erat autem rufus et pulcher aspectu decoraque facie. Et ait Dominus: " Surge, unge eum; ipse est enim ".
1SAM|16|13|Tulit igitur Samuel cornu olei et unxit eum in medio fratrum eius; et directus est spiritus Domini in David a die illa et in reliquum. Surgensque Samuel abiit in Rama.
1SAM|16|14|Spiritus autem Domini recessit a Saul, et exagitabat eum spiritus nequam a Domino.
1SAM|16|15|Dixeruntque servi Saul ad eum: " Ecce spiritus Dei malus exagitat te.
1SAM|16|16|Iubeat dominus noster, et servi tui, qui coram te sunt, quaerant hominem scientem psallere cithara, ut, quando arripuerit te spiritus Dei malus, psallat manu sua, et levius feras ".
1SAM|16|17|Et ait Saul ad servos suos: " Providete mihi aliquem bene psallentem et adducite eum ad me ".
1SAM|16|18|Et respondens unus de pueris ait: " Ecce vidi filium Isai Bethlehemitae scientem psallere et fortissimum robore et virum bellicosum et prudentem in verbis et virum pulchrum; et Dominus est cum eo ".
1SAM|16|19|Misit ergo Saul nuntios ad Isai dicens: " Mitte ad me David filium tuum, qui est in pascuis ".
1SAM|16|20|Tulitque Isai asinum cum pane et utre vini et haedo de capris uno et misit per manum David filii sui Sauli.
1SAM|16|21|Et venit David ad Saul et stetit coram eo; at ille dilexit eum nimis, et factus est eius armiger.
1SAM|16|22|Misitque Saul ad Isai dicens: " Stet David in conspectu meo; invenit enim gratiam in oculis meis ".
1SAM|16|23|Igitur, quandocumque spiritus Dei arripiebat Saul, David tollebat citharam et percutiebat manu sua; et refocillabatur Saul et levius habebat: recedebat enim ab eo spiritus malus.
1SAM|17|1|Congregantes vero Phili sthim agmina sua in proe lium, convenerunt in Socho Iudae et castrametati sunt inter Socho et Azeca in Aphesdommim.
1SAM|17|2|Porro Saul et viri Israel congregati venerunt in vallem Terebinthi et instruxerunt aciem ad pugnandum contra Philisthim.
1SAM|17|3|Et Philisthim stabant super montem ex hac parte, et Israel stabat super montem ex altera parte; vallisque erat inter eos.
1SAM|17|4|Et egressus est vir propugnator de castris Philisthinorum nomine Goliath de Geth altitudinis sex cubitorum et palmi.
1SAM|17|5|Et cassis aerea super caput eius, et lorica squamata induebatur; porro pondus loricae eius quinque milia siclorum aeris.
1SAM|17|6|Et ocreas aereas habebat in cruribus, et acinaces aereus erat inter umeros eius.
1SAM|17|7|Hastile autem hastae eius erat quasi liciatorium texentium, ipsum autem ferrum hastae eius sescentos siclos habebat ferri; et armiger eius antecedebat eum.
1SAM|17|8|Stansque clamabat adversum agmina Israel et dicebat eis: " Quare venitis parati ad proelium? Numquid ego non sum Philisthaeus, et vos servi Saul? Eligite ex vobis virum, et descendat ad singulare certamen!
1SAM|17|9|Si quiverit pugnare mecum et percusserit me, erimus vobis servi; si autem ego praevaluero et percussero eum, vos servi eritis et servietis nobis ".
1SAM|17|10|Et aiebat Philisthaeus: " Ego exprobravi agminibus Israel hodie: Date mihi virum, et ineat mecum singulare certamen! ".
1SAM|17|11|Audiens autem Saul et omnes Israelitae sermones Philisthaei huiuscemodi stupebant et metuebant nimis.
1SAM|17|12|David autem erat filius viri Ephrathaei, de quo supra dictum est, de Bethlehem Iudae, cui erat nomen Isai; qui habebat octo filios et erat vir in diebus Saul senex et grandaevus inter viros.
1SAM|17|13|Abierunt autem tres filii eius maiores post Saul in proelium; et nomina trium filiorum eius, qui perrexerant ad bellum: Eliab primogenitus et secundus Abinadab tertiusque Samma.
1SAM|17|14|David autem erat minimus; tribus ergo maioribus secutis Saulem,
1SAM|17|15|ibat David et revertebatur a Saul, ut pasceret gregem patris sui in Bethlehem.
1SAM|17|16|Procedebat vero Philisthaeus mane et vespere et stabat quadraginta diebus.
1SAM|17|17|Dixit autem Isai ad David filium suum: " Accipe fratribus tuis ephi frumenti tosti et decem panes istos et curre in castra ad fratres tuos.
1SAM|17|18|Et decem formellas casei has deferes ad tribunum, et fratres tuos visitabis, si recte agant; et pignus ab eis referes ".
1SAM|17|19|Saul autem et illi et omnes filii Israel in valle Terebinthi pugnabant adversum Philisthim.
1SAM|17|20|Surrexit itaque David mane et commendavit gregem custodi et onustus abiit, sicut praeceperat ei Isai. Et venit ad carraginem, dum exercitus egrediebatur ad pugnam et vociferabatur in certamine.
1SAM|17|21|Direxerunt ergo Israel et Philisthim aciem adversus aciem.
1SAM|17|22|Derelinquens autem David vasa, quae attulerat, sub manu custodis ad sarcinas, cucurrit ad locum certaminis et interrogabat, si omnia recte agerentur erga fratres suos.
1SAM|17|23|Cumque adhuc ille loqueretur eis, apparuit vir ille propugnator ascendens, Goliath nomine, Philisthaeus de Geth, ex castris Philisthinorum; et loquente eo haec eadem verba, audivit David.
1SAM|17|24|Omnes autem Israelitae, cum vidissent virum, fugerunt a facie eius timentes eum valde.
1SAM|17|25|Et dixit unus quispiam de Israel: " Num vidistis virum hunc, qui ascendit? Ad exprobrandum enim Israeli ascendit. Virum ergo, qui percusserit eum, ditabit rex divitiis magnis et filiam suam dabit ei; et domum patris eius faciet absque tributo in Israel ".
1SAM|17|26|Et ait David ad viros, qui stabant secum, dicens: " Quid dabitur viro, qui percusserit Philisthaeum hunc et tulerit opprobrium de Israel? Quis est enim hic Philisthaeus incircumcisus, qui exprobravit acies Dei viventis? ".
1SAM|17|27|Referebat autem ei populus eundem sermonem dicens: " Haec dabuntur viro, qui percusserit eum ".
1SAM|17|28|Quod cum audisset Eliab frater eius maior, loquente eo cum aliis, iratus est contra David et ait: " Quare venisti et cui dereliquisti pauculas oves illas in deserto? Ego novi superbiam tuam et nequitiam cordis tui, quia ut videres proelium descendisti ".
1SAM|17|29|Et dixit David: " Quid feci? Numquid non verbum est? ".
1SAM|17|30|Et declinavit paululum ab eo ad alium dixitque eundem sermonem; et respondit ei populus verbum sicut prius.
1SAM|17|31|Audita sunt autem verba, quae locutus est David, et annuntiata in conspectu Saul.
1SAM|17|32|Ad quem cum fuisset adductus, locutus est ei: " Non concidat cor cuiusquam in eo; ego servus tuus vadam et pugnabo adversus Philisthaeum istum ".
1SAM|17|33|Et ait Saul ad David: " Non vales resistere Philisthaeo isti nec pugnare adversus eum, quia puer es; hic autem vir bellator ab adulescentia sua ".
1SAM|17|34|Dixitque David ad Saul: " Pascebat servus tuus patris sui gregem, et veniebat leo vel ursus tollebatque arietem de medio gregis.
1SAM|17|35|Et sequebar eos et percutiebam eruebamque de ore eorum; et illi consurgebant adversum me, et apprehendebam mentum eorum et percutiebam interficiebamque eos.
1SAM|17|36|Nam et leonem et ursum interfecit servus tuus; erit igitur et Philisthaeus hic incircumcisus quasi unus ex eis, quia ausus est maledicere exercitum Dei viventis ".
1SAM|17|37|Et ait David: " Dominus, qui eruit me de manu leonis et de manu ursi, ipse liberabit me de manu Philisthaei huius ". Dixit autem Saul ad David: Vade, et Dominus tecum sit ".
1SAM|17|38|Et induit Saul David vestimentis suis et imposuit galeam aeream super caput eius et vestivit eum lorica.
1SAM|17|39|Accinctus ergo David gladio eius super vestem suam coepit tentare, si armatus posset incedere; non enim habebat consuetudinem. Dixitque David ad Saul: " Non possum sic incedere, quia nec usum habeo ". Et deposuit ea
1SAM|17|40|et tulit baculum suum in manu sua; et elegit sibi quinque levissimos lapides de torrente et misit eos in peram pastoralem, qua ut sacculo lapidum utebatur, et fundam manu tulit et processit adversum Philisthaeum.
1SAM|17|41|Ibat autem Philisthaeus incedens et appropinquans adversum David, et armiger eius ante eum.
1SAM|17|42|Cumque inspexisset Philisthaeus et vidisset David, despexit eum; erat enim adulescens rufus et pulcher aspectu.
1SAM|17|43|Et dixit Philisthaeus ad David: " Numquid ego canis sum, quod tu venis ad me cum baculo? ". Et maledixit Philisthaeus David in diis suis;
1SAM|17|44|dixitque ad David: " Veni ad me, et dabo carnes tuas volatilibus caeli et bestiis terrae ".
1SAM|17|45|Dixit autem David ad Philisthaeum: " Tu venis ad me cum gladio et hasta et acinace; ego autem venio ad te in nomine Domini exercituum, Dei agminum Israel, quibus exprobrasti.
1SAM|17|46|Hodie dabit te Dominus in manu mea, et percutiam te et auferam caput tuum a te; et dabo cadaver tuum et cadavera castrorum Philisthim hodie volatilibus caeli et bestiis terrae, ut sciat omnis terra quia est Deus in Israel,
1SAM|17|47|et noverit universa ecclesia haec quia non in gladio nec in hasta salvat Dominus: ipsius enim est bellum, et tradet vos in manus nostras ".
1SAM|17|48|Cum ergo surrexisset Philisthaeus et veniret et appropinquaret contra David, festinavit David et cucurrit ad pugnam adversum Philisthaeum.
1SAM|17|49|Et misit manum suam in peram tulitque unum lapidem et funda iecit; et percussit Philisthaeum in fronte, et infixus est lapis in fronte eius, et cecidit in faciem suam super terram.
1SAM|17|50|Praevaluitque David adversum Philisthaeum in funda et in lapide; percussumque Philisthaeum interfecit. Cumque gladium non haberet in manu, David
1SAM|17|51|cucurrit et stetit super Philisthaeum; et tulit gladium eius et eduxit eum de vagina sua et interfecit eum praeciditque caput eius.Videntes autem Philisthim quod mortuus esset fortissimus eorum fugerunt.
1SAM|17|52|Et consurgentes viri Israel et Iudae vociferati sunt et persecuti Philisthaeos usque dum venirent ad Geth et usque ad portas Accaron. Cecideruntque vulnerati de Philisthim in via a Saarim usque ad Geth et usque ad Accaron.
1SAM|17|53|Et revertentes filii Israel, postquam persecuti fuerant Philisthaeos, praedati sunt castra eorum.
1SAM|17|54|Assumens autem David caput Philisthaei attulit illud in Ierusalem; arma vero eius posuit in tabernaculo.
1SAM|17|55|Eo autem tempore, quo viderat Saul David egredientem contra Philisthaeum, ait ad Abner principem militiae: " De qua stirpe descendit hic adulescens, Abner? ". Dixitque Abner: " Vivit anima tua, rex, quia non novi ".
1SAM|17|56|Et ait rex: " Interroga tu, cuius filius sit iste puer ".
1SAM|17|57|Cumque regressus esset David, percusso Philisthaeo, tulit eum Abner et introduxit coram Saul caput Philisthaei habentem in manu.
1SAM|17|58|Et ait ad eum Saul: " De qua progenie es, o adulescens? ". Dixitque David: " Filius servi tui Isai Bethlehemitae ego sum ".
1SAM|18|1|Et factum est cum complesset loqui ad Saul, anima Ionathan colligata est animae David, et dilexit eum Ionathan quasi animam suam.
1SAM|18|2|Tulitque eum Saul in die illa et non concessit ei, ut reverteretur in domum patris sui.
1SAM|18|3|Inierunt autem Ionathan et David foedus; diligebat enim eum quasi animam suam.
1SAM|18|4|Et exspoliavit se Ionathan tunicam, qua erat vestitus, et dedit eam David et reliqua vestimenta sua usque ad gladium et arcum suum et usque ad balteum.
1SAM|18|5|Egrediebatur quoque David ad omnia, quaecumque misisset eum Saul, et prospere agebat; posuitque eum Saul super viros belli, et acceptus erat in oculis universi populi, etiam in conspectu famulorum Saul.
1SAM|18|6|Porro cum reverterentur, cum rediret David, percusso Philisthaeo, egressae sunt mulieres de universis urbibus Israel cantantes chorosque ducentes in occursum Saul regis in tympanis et in canticis laetitiae et in sistris.
1SAM|18|7|Et praecinebant mulieres ludentes atque dicentes: Percussit Saul milia sua,et David decem milia sua ".
1SAM|18|8|Iratus est autem Saul nimis, et displicuit in oculis eius iste sermo, dixitque: " Dederunt David decem milia et mihi dederunt milia; quid ei superest nisi solum regnum? ".
1SAM|18|9|Non rectis ergo oculis Saul aspiciebat David ex die illa et deinceps.
1SAM|18|10|Post diem autem alteram invasit spiritus Dei malus Saul, et vaticinabatur in medio domus suae; David autem psallebat manu sua sicut per singulos dies, tenebatque Saul lanceam.
1SAM|18|11|Et sustulit eam putans quod configere posset David cum pariete; et declinavit David a facie eius secundo.
1SAM|18|12|Et timuit Saul David, eo quod esset Dominus cum eo et a se recessisset.
1SAM|18|13|Amovit ergo eum Saul a se et fecit eum tribunum super mille viros; et egrediebatur et intrabat in conspectu populi.
1SAM|18|14|In omnibus quoque viis suis David prospere agebat, et Dominus erat cum eo.
1SAM|18|15|Vidit itaque Saul quod prospere ageret nimis et coepit pavere eum;
1SAM|18|16|omnis autem Israel et Iuda diligebat David; ipse enim egrediebatur et ingrediebatur ante eos.
1SAM|18|17|Dixit autem Saul ad David: " Ecce filia mea maior Merob, ipsam dabo tibi uxorem; tantummodo esto mihi vir fortis et proeliare bella Domini ". Saul autem reputabat dicens: " Non sit manus mea in eo, sed sit super illum manus Philisthinorum ".
1SAM|18|18|Ait autem David ad Saul: " Quis ego sum, aut quae est vita mea aut cognatio patris mei in Israel, ut fiam gener regis? ".
1SAM|18|19|Factum est autem tempus, cum deberet dari Merob filia Saul David, data est Hadriel Molathitae uxor.
1SAM|18|20|Dilexit autem Michol filia Saul altera David, et nuntiatum est Saul, et placuit ei;
1SAM|18|21|dixitque Saul: " Dabo eam illi, ut fiat ei in scandalum, et sit super eum manus Philisthinorum ". Dixit ergo Saul ad David altera vice: " Gener meus eris hodie ".
1SAM|18|22|Et mandavit Saul servis suis: " Loquimini ad David secreto dicentes: Ecce places regi, et omnes servi eius diligunt te; nunc ergo esto gener regis" ".
1SAM|18|23|Et locuti sunt servi Saul in auribus David omnia verba haec, et ait David: " Num parum vobis videtur generum esse regis? Ego autem sum vir pauper et tenuis ".
1SAM|18|24|Et renuntiaverunt servi Saul dicentes: " Huiuscemodi verba locutus est David ".
1SAM|18|25|Dixit autem Saul: " Sic loquimini ad David: "Non habet necesse rex sponsalia, nisi tantum centum praeputia Philisthinorum, ut fiat ultio de inimicis regis" ". Porro Saul cogitabat tradere David in manibus Philisthinorum.
1SAM|18|26|Cumque renuntiassent servi eius David verba, quae dixerat Saul, placuit sermo in oculis David, ut fieret gener regis.
1SAM|18|27|Et nondum erant dies impleti, cum David surgens abiit cum viris, qui sub eo erant, et percussit ex Philisthim ducentos viros; et attulit praeputia eorum, et annumeraverunt ea regi, ut esset gener eius.Dedit itaque ei Saul Michol filiam suam uxorem.
1SAM|18|28|Et vidit Saul et intellexit quia Dominus esset cum David; Michol autem filia Saul diligebat eum.
1SAM|18|29|Et Saul magis coepit timere David; factusque est Saul inimicus David cunctis diebus.
1SAM|18|30|Et egressi sunt principes Philisthinorum; et, quotiescumque egrediebantur, prospere agebat David magis quam omnes servi Saul, et celebre factum est nomen eius nimis.
1SAM|19|1|Locutus est autem Saul ad Ionathan filium suum et ad omnes servos suos de occisione David; porro Ionathan filius Saul diligebat David valde.
1SAM|19|2|Et indicavit Ionathan David dicens: " Quaerit Saul pater meus occidere te; quapropter observa te, quaeso, mane; et manebis clam et absconderis.
1SAM|19|3|Ego autem egrediens stabo iuxta patrem meum in agro, ubicumque fueris; et ego loquar de te ad patrem meum et, quodcumque videro, nuntiabo tibi ".
1SAM|19|4|Locutus est ergo Ionathan de David bona ad Saul patrem suum dixitque ad eum: " Ne peccet rex in servum suum David, quia non peccavit tibi, et opera eius bona sunt tibi valde.
1SAM|19|5|Et posuit animam suam in manu sua et percussit Philisthaeum, et fecit Dominus victoriam magnam universo Israeli; vidisti et laetatus es. Quare ergo peccas in sanguine innoxio interficiens David, qui est absque culpa?.
1SAM|19|6|Quod cum audisset Saul, placatus voce Ionathan iuravit: " Vivit Dominus quia non occidetur ".
1SAM|19|7|Vocavit itaque Ionathan David et indicavit ei omnia verba haec; et introduxit lonathan David ad Saul, et fuit ante eum, sicut fuerat heri et nudiustertius.
1SAM|19|8|Motum est autem rursum bellum, et egressus David pugnavit adversum Philisthim percussitque eos plaga magna; et fugerunt a facie eius.
1SAM|19|9|Et factus est spiritus Domini malus in Saul; sedebat autem in domo sua et tenebat lanceam, porro David psallebat in manu sua.
1SAM|19|10|Nisusque est Saul configere lancea David in pariete; et declinavit David a facie Saul, lancea autem, casso vulnere, perlata est in parietem. Et David fugit et salvatus est nocte illa.
1SAM|19|11|Misit ergo Saul satellites suos in domum David, ut custodirent eum, et interficeretur mane.Quod cum annuntiasset David Michol uxor sua dicens: " Nisi salvaveris te nocte hac, cras morieris ",
1SAM|19|12|deposuit eum per fenestram. Porro ille abiit et aufugit atque salvatus est.
1SAM|19|13|Tulit autem Michol theraphim et posuit eum super lectum; et pellem pilosam caprarum posuit ad caput eius et operuit eum vestimentis.
1SAM|19|14|Misit autem Saul nuntios, qui raperent David, et responsum est quod aegrotaret.
1SAM|19|15|Rursumque misit Saul nuntios, ut viderent David, dicens: " Afferte eum ad me in lecto, ut occidatur ".
1SAM|19|16|Cumque venissent nuntii, inventus est theraphim super lectum, et pellis caprarum ad caput eius.
1SAM|19|17|Dixitque Saul ad Michol: " Quare sic illusisti mihi et dimisisti inimicum meum, ut fugeret? ". Et respondit Michol ad Saul: " Quia ipse locutus est mihi: "Dimitte me, alioquin interficiam te" ".
1SAM|19|18|David autem fugiens salvatus est et venit ad Samuel in Rama et nuntiavit ei omnia, quae fecerat sibi Saul. Et abierunt ipse et Samuel et morati sunt in Naioth.
1SAM|19|19|Nuntiatum est autem Sauli a dicentibus: " Ecce David in Naioth in Rama.
1SAM|19|20|Misit ergo Saul nuntios, ut raperent David. Qui cum vidissent cuneum prophetarum vaticinantium et Samuel stantem super eos, factus est in illis spiritus Dei, et vaticinari coeperunt etiam ipsi.
1SAM|19|21|Quod cum nuntiatum esset Sauli, misit alios nuntios; vaticinati sunt autem et illi. Et rursum Saul misit tertios nuntios, qui et ipsi vaticinati sunt.
1SAM|19|22|Abiit autem etiam ipse in Rama et venit usque ad cisternam magnam, quae est in Socho; et interrogavit et dixit: " In quo loco sunt Samuel et David? ". Dictumque est ei: " Ecce in Naioth sunt in Rama ".
1SAM|19|23|Et abiit inde in Naioth in Rama; et factus est etiam super eum spiritus Dei, et ambulabat ingrediens et vaticinans, usquedum veniret in Naioth in Rama.
1SAM|19|24|Et exspoliavit se etiam ipse vestimentis suis et vaticinatus est cum ceteris coram Samuel; et cecidit nudus tota die illa et nocte, unde et exivit proverbium: " Num et Saul inter prophetas? ".
1SAM|20|1|Fugit autem David de Naioth, quae est in Rama, veniensque locutus est coram Ionathan: " Quid feci? Quae est iniquitas mea et quod peccatum meum in patrem tuum, quia quaerit animam meam? ".
1SAM|20|2|Qui dixit ei: " Absit, non morieris; neque enim faciet pater meus quidquam grande vel parvum, nisi prius indicaverit mihi; hoc ergo celavit me pater meus tantummodo? Nequaquam erit istud ".
1SAM|20|3|Et rursum respondit David et ait: " Scit profecto pater tuus quia inveni gratiam in oculis tuis et dixit: "Nesciat hoc Ionathan, ne forte tristetur". Quinimmo vivit Dominus, et vivit anima tua, quia uno tantum gradu ego morsque dividimur ".
1SAM|20|4|Et ait Ionathan ad David: " Quid desiderat anima tua, ut faciam tibi? ".
1SAM|20|5|Dixit autem David ad Ionathan: " Ecce neomenia est crastino, et ego ex more sedere soleo iuxta regem ad vescendum; dimitte ergo me, ut abscondar in agro usque ad vesperam diei tertiae.
1SAM|20|6|Si requisierit me pater tuus, respondebis ei: "Rogavit me David, ut iret celeriter in Bethlehem civitatem suam, quia victimae annuae ibi sunt universis contribulibus eius".
1SAM|20|7|Si dixerit: "Bene", pax erit servo tuo; si autem fuerit iratus, scito quia malum decretum est ab eo.
1SAM|20|8|Fac ergo misericordiam in servum tuum, quia foedus Domini me famulum tuum tecum inire fecisti; si autem est in me aliqua iniquitas, tu me interfice et ad patrem tuum ne introducas me ".
1SAM|20|9|Et ait Ionathan: " Absit hoc a te; neque enim fieri potest ut, si certo cognovero malum decretum esse a patre meo contra te, non annuntiem tibi ".
1SAM|20|10|Responditque David ad Ionathan: " Quis nuntiabit mihi, si quid forte responderit tibi pater tuus dure? ".
1SAM|20|11|Et ait Ionathan ad David: " Veni, egrediamur foras in agrum ". Cumque exissent ambo in agrum,
1SAM|20|12|ait Ionathan ad David: " Vivit Dominus, Deus Israel, investigabo sententiam patris mei hoc fere tempore cras vel perendie; et si aliquid boni fuerit super David, et non statim miserim ad te et notum tibi fecerim,
1SAM|20|13|haec faciat Dominus in Ionathan et haec augeat! Si autem perseveraverit patris mei malitia adversum te, hoc quoque notum faciam tibi et dimittam te, ut vadas in pace. Et sit Dominus tecum, sicut fuit cum patre meo.
1SAM|20|14|Et, si vixero, facies mihi misericordiam Domini; si vero mortuus fuero,
1SAM|20|15|non auferas misericordiam tuam a domo mea usque in sempiternum, quando eradicaverit Dominus inimicos David unumquemque de terra ".
1SAM|20|16|Pepigit ergo foedus Ionathan cum domo David dicens: " Requirat Dominus de manu inimicorum David! ".
1SAM|20|17|Et addidit Ionathan ut faceret David iurare per dilectionem suam erga illum; sicut animam enim suam, ita diligebat eum.
1SAM|20|18|Dixitque ad eum Ionathan: " Cras neomenia est, et requireris;
1SAM|20|19|vacua erit enim sessio tua. Perendie descendes festinus et venies in locum, ubi abscondisti te in die facti illius; et sedebis iuxta acervum illum.
1SAM|20|20|Et ego tres sagittas mittam iuxta eum et iaciam quasi exercens me ad signum.
1SAM|20|21|Mittam quoque et puerum dicens ei: "Vade et affer mihi sagittas".
1SAM|20|22|Si dixero puero: "Ecce sagittae intra te sunt, tolle eas", tu veni ad me, quia pax tibi est, et nihil est mali, vivit Dominus. Si autem sic locutus fuero puero: "Ecce sagittae ultra te sunt", vade, quia dimisit te Dominus.
1SAM|20|23|De verbo autem, quod locuti fuimus, ego et tu, sit Dominus inter me et te usque in sempiternum ".
1SAM|20|24|Absconditus est ergo David in agro; et venit neomenia, et sedit rex ad mensam ad comedendum.
1SAM|20|25|Cumque sedisset rex super cathedram suam secundum consuetudinem, quae erat iuxta parietem, sedit Ionathan ex adverso, et sedit Abner ex latere Saul; vacuusque apparuit locus David.
1SAM|20|26|Et non est locutus Saul quidquam in die illa; cogitabat enim quod forte evenisset ei, ut non esset mundus nec purificatus.
1SAM|20|27|Cumque illuxisset dies secunda post neomeniam, rursum vacuus apparuit locus David; dixitque Saul ad Ionathan filium suum: " Cur non venit filius Isai nec heri nec hodie ad vescendum? ".
1SAM|20|28|Et respondit Ionathan Sauli: " Rogavit me obnixe, ut iret in Bethlehem,
1SAM|20|29|et ait: "Dimitte me, quoniam sacrificium familiae est in civitate, et frater meus ipse accersivit me; nunc ergo, si inveni gratiam in oculis tuis, vadam cito et videbo fratres meos". Ob hanc causam non venit ad mensam regis ".
1SAM|20|30|Iratus autem Saul adversum Ionathan dixit ei: " Fili mulieris perversae, numquid ignoro quia diligis filium Isai in confusionem tuam et in confusionem nuditatis matris tuae?
1SAM|20|31|Omnibus enim diebus, quibus filius Isai vixerit super terram, non stabilieris tu neque regnum tuum; itaque iam nunc mitte et adduc eum ad me, quia filius mortis est ".
1SAM|20|32|Respondens autem Ionathan Sauli patri suo ait: " Quare morietur? Quid fecit? ".
1SAM|20|33|Et arripuit Saul lanceam, ut percuteret eum; et intellexit Ionathan quod definitum esset patri suo, ut interficeret David.
1SAM|20|34|Surrexit ergo Ionathan a mensa in ira furoris et non comedit in die neomeniae secunda panem; contristatus est enim super David, eo quod confudisset eum pater suus.
1SAM|20|35|Cumque illuxisset mane, venit Ionathan in agrum ad locum constitutum a David et puer parvulus cum eo;
1SAM|20|36|et ait ad puerum suum: " Vade et affer mihi sagittas, quas ego iacio ". Cumque puer cucurrisset, iecit sagittam trans puerum.
1SAM|20|37|Venit itaque puer ad locum sagittae, quam miserat Ionathan, et clamavit Ionathan post tergum pueri et ait: " Ecce ibi est sagitta porro ultra te.
1SAM|20|38|Clamavitque Ionathan post tergum pueri: " Festina velociter, ne steteris ". Sustulit autem puer Ionathae sagittam et attulit ad dominum suum
1SAM|20|39|et quid ageretur penitus ignorabat, tantummodo enim Ionathan et David rem noverant.
1SAM|20|40|Dedit igitur Ionathan arma sua puero et dixit ei: " Vade, defer in civitatem ".
1SAM|20|41|Cumque abisset puer, surrexit David de latere acervi et cadens pronus in terram adoravit tertio; et osculantes alterutrum fleverunt pariter, David autem amplius.
1SAM|20|42|Dixit ergo Ionathan ad David: " Vade in pace; iuravimus enim ambo in nomine Domini dicentes: Dominus erit inter me et te et inter semen meum et semen tuum usque in sempiternum ".
1SAM|21|1|Et surrexit David et abiit; sed et Ionathan ingressus est civitatem.
1SAM|21|2|Venit autem David in Nob ad Achimelech sacerdotem, et obstupuit Achimelech eo quod venisset David, et dixit ei: " Quare tu solus et nullus est tecum? ".
1SAM|21|3|Et ait David ad Achimelech sacerdotem: " Rex praecepit mihi negotium et dixit: "Nemo sciat rem, propter quam a me missus es, et cuiusmodi tibi praecepta dederim"; pueris vero condixi in illum et illum locum.
1SAM|21|4|Nunc igitur, si habes ad manum quinque panes, da mihi, aut quidquid inveneris ".
1SAM|21|5|Et respondens sacerdos David ait ei: " Non habeo panes laicos ad manum, sed tantum panem sanctum; si mundi sunt pueri maxime a mulieribus? ".
1SAM|21|6|Et respondit David sacerdoti et dixit ei: " Equidem, si de mulieribus agitur, continuimus nos ab heri et nudiustertius. Quando egrediebar, fuerunt corpora puerorum sancta, quamvis iter esset profanum. Quanto magis hodie sunt sancti quoad corpora ".
1SAM|21|7|Dedit ergo ei sacerdos sanctificatum panem; neque enim erat ibi panis, nisi tantum panes propositionis, qui sublati fuerant a facie Domini, ut ponerentur panes calidi.
1SAM|21|8|Erat autem ibi vir de servis Saul in die illa retentus ante Dominum; et nomen eius Doeg Idumaeus, potentissimus pastorum Saul.
1SAM|21|9|Dixit autem David ad Achimelech: " Si habes hic ad manum hastam aut gladium? Quia gladium meum et arma mea non tuli mecum; negotium enim regis urgebat ".
1SAM|21|10|Et dixit sacerdos: " Ecce hic gladius Goliath Philisthaei, quem percussisti in valle Terebinthi; est involutus pallio post ephod. Si istum vis tollere, tolle, neque enim est alius hic absque eo ". Et ait David: " Non est huic alter similis; da mihi eum ".
1SAM|21|11|Surrexit itaque David et fugit in die illa a facie Saul et venit ad Achis regem Geth.
1SAM|21|12|Dixeruntque ei servi Achis: " Numquid non iste est David rex terrae? Nonne huic cantabant per choros dicentes: "Percussit Saul milia sua, et David decem milia sua"? ".
1SAM|21|13|Posuit autem David sermones istos in corde suo et extimuit valde a facie Achis regis Geth.
1SAM|21|14|Et immutavit os suum coram eis; et insaniebat inter manus eorum et impingebat in ostia portae, defluebantque salivae in barbam.
1SAM|21|15|Et ait Achis ad servos suos: " Vidistis hominem insanum. Quare adduxistis eum ad me?
1SAM|21|16|An desunt nobis furiosi, quod introduxistis istum, ut fureret, me praesente? Hicine ingredietur domum meam? ".
1SAM|22|1|Abiit ergo inde David et fugit in speluncam Odollam; quod cum audissent fratres eius et omnis domus patris eius, descenderunt ad eum illuc.
1SAM|22|2|Et convenerunt ad eum omnes, qui erant in angustia constituti et oppressi aere alieno et amaro animo; et factus est eorum princeps, fueruntque cum eo quasi quadringenti viri.
1SAM|22|3|Et profectus est David inde in Maspha, quae est Moab, et dixit ad regem Moab: " Maneat, oro, pater meus et mater mea vobiscum, donec sciam quid faciat mihi Deus ".
1SAM|22|4|Et reliquit eos ante faciem regis Moab; manseruntque apud eum cunctis diebus, quibus David fuit in praesidio.
1SAM|22|5|Dixitquc Gad propheta ad David: " Noli manere in praesidio. Proficiscere et vade in terram Iudae ". Et profectus David venit in saltum Haret.
1SAM|22|6|Et audivit Saul quod detectus fuisset David et viri, qui erant cum eo. Saul autem, cum maneret in Gabaa et esset sub myrice, quae est in excelso, hastam manu tenens, cunctique servi eius circumstarent eum,
1SAM|22|7|ait ad servos suos, qui assistebant ei: " Audite, Beniaminitae. Etiam omnibus vobis dabit filius Isai agros et vineas et universos vos faciet tribunos et centuriones,
1SAM|22|8|quoniam coniurastis omnes adversum me. Et non est qui mihi renuntiet quod filius meus foedus iunxerit cum filio Isai; non est qui vicem meam doleat ex vobis, nec qui annuntiet mihi quod suscitaverit filius meus servum meum adversum me insidiantem mihi sicut hodie ".
1SAM|22|9|Respondens autem Doeg Idumaeus, qui assistebat cum servis Saul: " Vidi, inquit, filium Isai in Nob apud Achimelech filium Achitob;
1SAM|22|10|qui consuluit pro eo Dominum et cibaria dedit ei, sed et gladium Goliath Philisthaei dedit illi ".
1SAM|22|11|Misit ergo rex ad accersendum Achimelech sacerdotem filium Achitob et omnem domum patris eius, sacerdotum, qui erant in Nob; qui venerunt universi ad regem.
1SAM|22|12|Et ait Saul: " Audi, fili Achitob ". Qui respondit: " Praesto sum, domine ".
1SAM|22|13|Dixitque ad eum Saul: " Quare coniurastis adversum me, tu et filius Isai, et dedisti ei panes et gladium et consuluisti pro eo Deum, ut consurgeret adversum me insidiator, sicut est hodie? ".
1SAM|22|14|Respondensque Achimelech regi ait: " Et quis in omnibus servis tuis sicut David fidelis et gener regis et dux satellitum tuorum et gloriosus in domo tua?
1SAM|22|15|Num hodie coepi consulere pro eo Deum? Absit hoc a me, ne suspicetur rex adversus servum suum rem huiuscemodi, adversus universam domum patris mei; non enim scivit servus tuus quidquam super hoc negotio, vel modicum vel grande ".
1SAM|22|16|Dixitque rex: " Morte morieris, Achimelech, tu et omnis domus patris tui ".
1SAM|22|17|Et ait rex emissariis, qui circumstabant eum: " Convertimini et interficite sacerdotes Domini, nam manus eorum cum David est; scientes quod fugisset, non indicaverunt mihi ". Noluerunt autem servi regis extendere manum suam in sacerdotes Domini.
1SAM|22|18|Et ait rex ad Doeg: " Convertere tu et irrue in sacerdotes ". Conversusque Doeg Idumaeus irruit in sacerdotes; et trucidavit in die illa octoginta quinque viros vestitos ephod lineo.
1SAM|22|19|Nob autem civitatem sacerdotum percussit in ore gladii, viros et mulieres, parvulos et lactantes, bovem et asinum et ovem in ore gladii.
1SAM|22|20|Evadens autem unus filius Achimelech filii Achitob, cuius nomen erat Abiathar, fugit ad David
1SAM|22|21|et annuntiavit ei quod occidisset Saul sacerdotes Domini.
1SAM|22|22|Et ait David ad Abiathar: " Sciebam in die illa quod, cum ibi esset Doeg Idumaeus, procul dubio annuntiaret Saul; ego sum reus omnium animarum domus patris tui.
1SAM|22|23|Mane mecum, ne timeas; qui enim quaerit animam meam, quaerit et animam tuam, mecumque servaberis ".
1SAM|23|1|Et nuntiaverunt David di centes: " Ecce Philisthim op pugnant Ceila et diripiunt areas ".
1SAM|23|2|Consuluit igitur David Dominum dicens: " Num vadam et percutiam Philisthaeos istos? ". Et ait Dominus ad David: " Vade et percuties Philisthaeos et salvabis Ceila ".
1SAM|23|3|Et dixerunt viri, qui erant cum David, ad eum: " Ecce nos hic in Iuda consistentes timemus; quanto magis si ierimus in Ceila adversum agmina Philisthinorum? ".
1SAM|23|4|Rursum ergo David consuluit Dominum, qui respondens ei ait: " Surge et vade in Ceila; ego enim tradam Philisthaeos in manu tua ".
1SAM|23|5|Abiit ergo David et viri eius in Ceila et pugnavit adversum Philisthaeos et abegit iumenta eorum et percussit eos plaga magna: et salvavit David habitatores Ceilae.
1SAM|23|6|Porro cum fugisset Abiathar filius Achimelcch ad David, et ipse cum David in Ceila ephod secum habens descenderat.
1SAM|23|7|Nuntiatum est autem Saul quod venisset David in Ceila, et ait Saul: " Tradidit eum Deus in manus meas; conclususque est introgressus urbem, in qua portae et serae sunt ".
1SAM|23|8|Et convocavit Saul omnem populum, ut ad pugnam descenderet in Ceila et obsideret David et viros eius.
1SAM|23|9|Quod cum rescisset David quia praepararet ei Saul clam malum, dixit ad Abiathar sacerdotem: " Applica ephod ".
1SAM|23|10|Et ait David: " Domine, Deus Israel, audivit famam servus tuus quod disponat Saul venire ad Ceila, ut evertat urbem propter me.
1SAM|23|11|Si tradent me viri Ceilae in manus eius? Et si descendet Saul, sicut audivit servus tuus? Domine, Deus Israel, indica servo tuo ". Et ait Dominus: " Descendet ".
1SAM|23|12|Dixitque David: " Si tradent viri Ceilae me et viros, qui sunt mecum, in manu Saul? ". Et dixit Dominus: " Tradent ".
1SAM|23|13|Surrexit ergo David et viri eius quasi sescenti et egressi de Ceila huc atque illuc vagabantur incerti. Nuntiatumque est Saul quod fugisset David de Ceila, quam ob rem destitit exire.
1SAM|23|14|Morabatur autem David in deserto in locis firmissimis mansitque in monte, in deserto Ziph; et quaerebat eum Saul cunctis diebus, sed non tradidit eum Deus in manus eius.
1SAM|23|15|Et cognovit David quod egressus esset Saul, ut quaereret animam eius; porro David erat in deserto Ziph in Horesa.
1SAM|23|16|Et surrexit Ionathan filius Saul et abiit ad David in Horesa; et confortavit manus eius in Deo dixitque ei:
1SAM|23|17|" Ne timeas, neque enim inveniet te manus Saul patris mei; et tu regnabis super Israel, et ego ero tibi secundus; sed et Saul pater meus scit hoc ".
1SAM|23|18|Percussit igitur uterque foedus coram Domino; mansitque David in Horesa, Ionathan autem reversus est in domum suam.
1SAM|23|19|Ascenderunt autem Ziphaei ad Saul in Gabaa dicentes: " Nonne David latitat apud nos in locis tutissimis in Horesa, in colle Hachila, quae est ad meridiem deserti?
1SAM|23|20|Nunc ergo, si desideravit anima tua, rex, ut descenderes, descende; nostrum autem erit ut tradamus eum in manus regis ".
1SAM|23|21|Dixitque Saul: " Benedicti vos a Domino, quia doluistis vicem meam.
1SAM|23|22|Abite, oro, et diligentius praeparate et curiosius agite; et considerate locum, ubi sit pes eius, vel quis viderit eum ibi; dictum est enim ad me quod callidus sit valde.
1SAM|23|23|Considerate et videte omnia latibula eius, in quibus absconditur, et revertimini ad me ad certum locum, ut vadam vobiscum; quodsi fuerit in regione, perscrutabor eum in cunctis regionibus Iudae ".
1SAM|23|24|At illi surgentes abierunt in Ziph ante Saul.David autem et viri eius erant in deserto Maon, in Araba ad meridiem deserti.
1SAM|23|25|Ivit ergo Saul et socii eius ad quaerendum eum, et nuntiatum est David; descenditque ad petram et versabatur in deserto Maon. Quod cum audisset Saul, persecutus est David in deserto Maon.
1SAM|23|26|Et ibat Saul ad latus montis ex parte una, David autem et viri eius erant in latere montis ex parte altera; porro David praeceps fugiebat a facie Saul. Itaque Saul et viri eius in modum coronae cingebant David et viros eius, ut caperent eos.
1SAM|23|27|Et nuntius venit ad Saul dicens: " Festina et veni, quoniam infuderunt se Philisthim super terram ".
1SAM|23|28|Reversus est ergo Saul desistens persequi David; et perrexit in occursum Philisthinorum. Propter hoc vocaverunt locum illum: " Petram dividentem ".
1SAM|24|1|Ascendit ergo David inde et habitavit in locis tutissimis Engaddi.
1SAM|24|2|Cumque reversus esset Saul, postquam persecutus est Philisthaeos, nuntiaverunt ei dicentes: " Ecce David in deserto est Engaddi ".
1SAM|24|3|Assumens ergo Saul tria milia electorum virorum ex omni Israel perrexit ad investigandum David et viros eius ad rupes ibicum.
1SAM|24|4|Et venit ad caulas ovium, quae se offerebant vianti.Eratque ibi spelunca, quam ingressus est Saul, ut purgaret ventrem; porro David et viri eius in interiore parte speluncae latebant.
1SAM|24|5|Et dixerunt viri David ad eum: " Ecce dies, de qua locutus est Dominus ad te: "Ego trado tibi inimicum tuum, ut facias ei sicut placuerit in oculis tuis" ". Surrexit ergo David et praecidit oram chlamydis Saul silenter.
1SAM|24|6|Post haec cor David percussit eum, eo quod abscidisset oram chlamydis Saul,
1SAM|24|7|dixitque ad viros suos: " Propitius mihi sit Dominus, ne faciam hanc rem domino meo, christo Domini, ut mittam manum meam in eum, quoniam christus Domini est ".
1SAM|24|8|Et cohibuit David viros suos sermonibus et non permisit eos, ut consurgerent in Saul.Porro Saul exsurgens de spelunca pergebat coepto itinere.
1SAM|24|9|Surrexit autem et David post eum et egressus de spelunca clamavit post tergum Saul dicens: " Domine mi rex! ". Et respexit Saul post se, et inclinans se David pronus in terram adoravit
1SAM|24|10|dixitque ad Saul: " Quare audis verba hominum loquentium: "David quaerit malum adversum te?".
1SAM|24|11|Ecce hodie viderunt oculi tui quod tradiderit te Dominus hodie in manu mea in spelunca; et dictum est mihi, ut occiderem te, sed pepercit tibi oculus meus. Dixi enim: Non extendam manum meam in dominum meum, quia christus Domini est
1SAM|24|12|et pater meus. Quin potius vide et cognosce oram chlamydis tuae in manu mea, quoniam, cum praeciderem summitatem chlamydis tuae, nolui occidere te. Animadverte et vide quoniam non est in manu mea malum neque iniquitas, neque peccavi in te; tu autem insidiaris animae meae, ut auferas eam.
1SAM|24|13|Iudicet Dominus inter me et te et ulciscatur me Dominus ex te; manus autem mea non sit in te.
1SAM|24|14|Sicut et in proverbio antiquo dicitur: "Ab impiis egredietur impietas", manus ergo mea non sit in te.
1SAM|24|15|Quem sequitur rex Israel? Quem persequeris? Canem mortuum et pulicem unum.
1SAM|24|16|Sit Dominus iudex et iudicet inter me et te et videat et diiudicet causam meam et eruat me de manu tua ".
1SAM|24|17|Cum autem complesset David loquens sermones huiuscemodi ad Saul, dixit Saul: " Numquid vox haec tua est, fili mi David? ". Et levavit Saul vocem suam et flevit.
1SAM|24|18|Dixitque ad David: " Iustior tu es quam ego; tu enim tribuisti mihi bona, ego autem reddidi tibi mala.
1SAM|24|19|Et tu indicasti hodie, quae feceris mihi bona, quomodo tradiderit me Dominus in manu tua, et non occideris me.
1SAM|24|20|Quis enim, cum invenerit inimicum suum, dimittet eum in via bona? Sed Dominus reddat tibi vicissitudinem hanc, pro eo quod hodie operatus es in me.
1SAM|24|21|Et nunc, quia scio quod certissime regnaturus sis et habiturus in manu tua regnum Israel,
1SAM|24|22|iura mihi in Domino, ne deleas semen meum post me neque auferas nomen meum de domo patris mei ".
1SAM|24|23|Et iuravit David Sauli. Abiit ergo Saul in domum suam, et David et viri eius ascenderunt ad praesidium.
1SAM|25|1|Mortuus est autem Samuel; et congregatus est universus Israel, et planxerunt eum et sepelierunt eum in domo sua in Rama.Consurgensque David descendit in desertum Maon.
1SAM|25|2|Erat autem vir quispiam in solitudine Maon, et possessio eius in Carmel; et homo ille magnus nimis; erantque ei oves tria milia et mille caprae. Et accidit ut tonderet gregem suum in Carmel.
1SAM|25|3|Nomen autem viri illius erat Nabal et nomen uxoris eius Abigail. Eratque mulier illa prudentissima et speciosa; porro vir eius durus et moribus malis; erat autem de genere Chaleb.
1SAM|25|4|Cum ergo audisset David in deserto quod tonderet Nabal gregem suum,
1SAM|25|5|misit decem iuvenes et dixit eis: " Ascendite in Carmel et venietis ad Nabal et salutabitis eum ex nomine meo pacifice
1SAM|25|6|et dicetis fratri meo: "Et tibi pax et domui tuae pax et omnibus, quaecumque habes, sit pax!
1SAM|25|7|Et nunc audivi quod tonsores essent apud te. Pastores autem tui erant nobiscum in deserto; numquam eis molesti fuimus, nec aliquando defuit eis quidquam de grege omni tempore, quo fuerunt nobiscum in Carmel.
1SAM|25|8|Interroga pueros tuos, et indicabunt tibi. Nunc ergo inveniant pueri isti gratiam in oculis tuis, in die enim bona venimus; quodcumque invenerit manus tua, da servis tuis et filio tuo David" ".
1SAM|25|9|Cumque venissent pueri David, locuti sunt ad Nabal omnia verba haec ex nomine David et siluerunt.
1SAM|25|10|Respondens autem Nabal pueris David ait: " Quis est David, et quis est filius Isai? Hodie increverunt servi, qui fugiunt dominos suos.
1SAM|25|11|Tollam ergo panes meos et aquas meas et carnes pecorum, quae occidi, tonsoribus meis et dabo viris, quos nescio unde sint? ".
1SAM|25|12|Regressi sunt itaque pueri David per viam suam et reversi venerunt et nuntiaverunt ei omnia verba haec.
1SAM|25|13|Tunc David ait viris suis: " Accingatur unusquisque gladio suo! ". Et accincti sunt singuli gladio suo, accinctusque est et David ense suo, et secuti sunt David quasi quadringenti viri; porro ducenti remanserunt ad sarcinas.
1SAM|25|14|Abigail autem uxori Nabal nuntiavit unus de pueris suis dicens: " Ecce misit David nuntios de deserto, ut benedicerent domino nostro, sed aversatus est eos.
1SAM|25|15|Homines isti boni satis fuerunt nobis et non molesti; nec quidquam aliquando periit omni tempore, quo sumus conversati cum eis in deserto.
1SAM|25|16|Pro muro erant nobis tam in nocte quam in die omnibus diebus, quibus pavimus apud eos greges.
1SAM|25|17|Quam ob rem considera et recogita quid facias, quoniam malum decretum est adversus dominum nostrum et adversus domum eius universam. Et ipse filius Belial est, ita ut nemo ei possit loqui ".
1SAM|25|18|Festinavit igitur Abigail et tulit ducentos panes et duos utres vini et quinque arietes coctos et quinque sata frumenti tosti et centum ligaturas uvae passae et ducentas massas caricarum et imposuit super asinos.
1SAM|25|19|Dixitque pueris suis: " Praecedite me, ecce ego post tergum sequar vos. Viro autem suo Nabal non indicavit.
1SAM|25|20|Cum ergo ascendisset asinum et descenderet in tegmine montis, David et viri eius descendebant in occursum eius; quibus et illa occurrit.
1SAM|25|21|Et aiebat David: " Vere frustra servavi omnia, quae huius erant in deserto, et non periit quidquam de cunctis, quae ad eum pertinebant; et reddidit mihi malum pro bono.
1SAM|25|22|Haec faciat Deus inimicis David et haec addat, si reliquero de omnibus, quae ad eum pertinent, usque mane quidquid masculini sexus ".
1SAM|25|23|Cum autem vidisset Abigail David, festinavit et descendit de asino et procidit coram David super faciem suam et adoravit super terram.
1SAM|25|24|Et cecidit ad pedes eius et dixit: " In me sit, domine mi, haec iniquitas; loquatur, obsecro, ancilla tua in auribus tuis, et audi verba famulae tuae.
1SAM|25|25|Ne ponat, oro, dominus meus cor suum super virum istum iniquum Nabal, quia secundum nomen suum stultus est, et est stultitia cum eo; ego autem ancilla tua non vidi pueros domini mei, quos misisti.
1SAM|25|26|Nunc ergo, domine mi, vivit Dominus, et vivit anima tua, quia Dominus prohibuit te, ne venires in sanguine et salvares te manu tua; et nunc fiant sicut Nabal inimici tui et qui quaerunt domino meo malum.
1SAM|25|27|Quapropter suscipe benedictionem hanc, quam attulit ancilla tua domino meo, et da pueris, qui sequuntur dominum meum.
1SAM|25|28|Aufer iniquitatem famulae tuae. Faciens enim faciet Dominus domino meo domum fidelem, quia proelia Domini dominus meus proeliatur; malitia ergo non inveniatur in te omnibus diebus vitae tuae.
1SAM|25|29|Si enim surrexerit aliquando homo persequens te et quaerens animam tuam, erit anima domini mei custodita in fasciculo vitae apud Dominum Deum tuum; sed inimicorum tuorum animam ipse iaciat in impetu et circulo fundae.
1SAM|25|30|Cum ergo fecerit Dominus domino meo omnia, quae locutus est, bona de te et constituerit te ducem super Israel,
1SAM|25|31|non erit tibi hoc in singultum et in scrupulum cordis domino meo, quod effuderis sanguinem innoxium et ipse te ultus fueris; et cum benefecerit Dominus domino meo, recordaberis ancillae tuae ".
1SAM|25|32|Et ait David ad Abigail: " Benedictus Dominus, Deus Israel, qui misit te hodie in occursum meum. Et benedicta prudentia tua,
1SAM|25|33|et benedicta tu, quae prohibuisti me hodie, ne irem ad sanguinem et ulciscerer me manu mea.
1SAM|25|34|Alioquin, vivit Dominus, Deus Israel, qui prohibuit me malum facere tibi, nisi cito venisses in occursum mihi, non remansisset Nabal usque ad lucem matutinam quidquid masculini sexus ".
1SAM|25|35|Suscepit ergo David de manu eius omnia, quae attulerat ei, dixitque ei: Vade pacifice in domum tuam. Ecce audivi vocem tuam et honoravi faciem tuam ".
1SAM|25|36|Venit autem Abigail ad Nabal; et ecce erat ei convivium in domo eius quasi convivium regis, et cor Nabal iucundum; erat enim ebrius nimis. Et non indicavit ei verbum pusillum aut grande usque in mane.
1SAM|25|37|Diluculo autem, cum digessisset vinum Nabal, haec indicavit ei uxor sua; et emortuum est cor eius intrinsecus, et factus est quasi lapis.
1SAM|25|38|Cumque pertransissent decem dies, percussit Dominus Nabal, et mortuus est.
1SAM|25|39|Quod cum audisset David mortuum Nabal, ait: " Benedictus Dominus, qui iudicavit causam opprobrii mei de manu Nabal et servum suum custodivit a malo et malitiam Nabal reddidit Dominus in caput eius ".Misit ergo David et locutus est ad Abigail, ut sumeret eam sibi in uxorem.
1SAM|25|40|Et venerunt pueri David ad Abigail in Carmel et locuti sunt ad eam dicentes: " David misit nos ad te, ut accipiat te sibi in uxorem ".
1SAM|25|41|Quae consurgens adoravit prona in terram et ait: " Ecce famula tua sit in ancillam, ut lavet pedes servorum domini mei ".
1SAM|25|42|Et festinavit et surrexit Abigail et ascendit super asinum, et quinque puellae ierunt cum ea pedisequae eius; et secuta est nuntios David et facta est illi uxor.
1SAM|25|43|Sed et Achinoam accepit David de Iezrahel, et fuit utraque uxor eius.
1SAM|25|44|Saul autem dedit Michol filiam suam uxorem David Phalti filio Lais, qui erat de Gallim.
1SAM|26|1|Et venerunt Ziphaei ad Saul in Gabaa dicentes: " Ecce David absconditus est in colle Hachila, quae est ex adverso solitudinis ".
1SAM|26|2|Et surrexit Saul et descendit in desertum Ziph, et cum eo tria milia virorum de electis Israel, ut quaereret David in deserto Ziph.
1SAM|26|3|Et castrametatus est Saul in colle Hachila, quae erat ex adverso solitudinis in via. David autem habitabat in deserto; videns autem quod venisset Saul post se in desertum,
1SAM|26|4|misit exploratores et didicit quod illuc venisset certissime.
1SAM|26|5|Et surrexit David et venit ad locum, ubi erat Saul. Cumque vidisset locum, in quo dormiebat Saul et Abner filius Ner princeps militiae eius, Saulem dormientem in carragine et reliquum vulgus per circuitum eius,
1SAM|26|6|ait David ad Achimelech Hetthaeum et Abisai filium Sarviae fratrem Ioab dicens: " Quis descendet mecum ad Saul in castra? ". Dixitque Abisai: " Ego descendam tecum ".
1SAM|26|7|Venerunt ergo David et Abisai ad populum nocte et invenerunt Saul iacentem et dormientem in carragine et hastam fixam in terra ad caput eius, Abner autem et populum dormientes in circuitu eius.
1SAM|26|8|Dixitque Abisai ad David: " Conclusit Deus hodie inimicum tuum in manus tuas; nunc ergo perfodiam eum lancea in terra semel, et secundo opus non erit ".
1SAM|26|9|Et dixit David ad Abisai: " Ne interficias eum; quis enim extendit manum suam in christum Domini et innocens erit? ".
1SAM|26|10|Et dixit David: " Vivit Dominus quia Dominus percutiet eum, aut dies eius veniet, ut moriatur, aut in proelium descendens peribit.
1SAM|26|11|Propitius mihi sit Dominus, ne extendam manum meam in christum Domini. Nunc igitur tolle hastam, quae est ad caput eius, et scyphum aquae, et abeamus ".
1SAM|26|12|Tulit ergo David hastam et scyphum aquae, qui erat ad caput Saul, et abierunt; et non erat quisquam, qui videret et intellegeret et vigilaret, sed omnes dormiebant, quia sopor Domini irruerat super eos.
1SAM|26|13|Cumque transisset David ex adverso et stetisset in vertice montis de longe, et esset grande intervallum inter eos,
1SAM|26|14|clamavit David ad populum et ad Abner filium Ner dicens: " Nonne respondebis, Abner? ". Et respondens Abner ait: " Quis es tu? Clamasti ad regem! ".
1SAM|26|15|Et ait David ad Abner: " Numquid non vir tu es? Et quis alius similis tui in Israel? Quare ergo non custodisti dominum tuum regem? Ingressus est enim unus de turba, ut interficeret regem dominum tuum.
1SAM|26|16|Non est bonum hoc, quod fecisti. Vivit Dominus quoniam filii mortis estis vos, qui non custodistis dominum vestrum, christum Domini. Nunc ergo vide, ubi sit hasta regis et ubi scyphus aquae, qui erat ad caput eius ".
1SAM|26|17|Cognovit autem Saul vocem David et dixit: " Num vox tua haec est, fili mi David? ". Et ait David: " Vox mea, domine mi rex ".
1SAM|26|18|Et ait: " Quam ob causam dominus meus persequitur servum suum? Quid feci? Aut quod est in manu mea malum?
1SAM|26|19|Nunc ergo audiat, oro, dominus meus rex verba servi sui: Si Dominus incitat te adversum me, odoretur sacrificium; si autem filii hominum, maledicti sint in conspectu Domini, quia eiecerunt me hodie, ut non habitem in hereditate Domini dicentes: "Vade, servi diis alienis".
1SAM|26|20|Et nunc non effundatur sanguis meus in terra longe a facie Domini; quia egressus est rex Israel, ut quaerat pulicem unum, sicut persequitur quis perdicem in montibus ".
1SAM|26|21|Et ait Saul: " Peccavi. Revertere, fili mi David; nequaquam enim ultra malefaciam tibi, eo quod pretiosa fuerit anima mea in oculis tuis hodie; apparet quod stulte egerim et erraverim multum nimis ".
1SAM|26|22|Et respondens David ait: " Ecce hasta regis; transeat unus de pueris et tollat eam.
1SAM|26|23|Dominus autem retribuet unicuique secundum iustitiam suam et fidem; tradidit enim te Dominus hodie in manu mea, et nolui extendere manum meam in christum Domini.
1SAM|26|24|Et sicut magnificata est anima tua hodie in oculis meis, sic magnificetur anima mea in oculis Domini, et liberet me de omni angustia ".
1SAM|26|25|Ait ergo Saul ad David: " Benedictus tu, fili mi David; et quidem faciens facies et potens poteris ". Abiit autem David in viam suam, et Saul reversus est in locum suum.
1SAM|27|1|Et ait David in corde suo: " Aliquando incidam in uno die in manu Saul; nonne melius est ut fugiam et salver in terra Philisthinorum, ut desperet Saul cessetque me quaerere in cunctis finibus Israel? Fugiam ergo manus eius ".
1SAM|27|2|Et surrexit David et abiit ipse et sescenti viri cum eo ad Achis filium Maoch regem Geth.
1SAM|27|3|Et habitavit David cum Achis in Geth ipse et viri eius unusquisque cum domo sua; David et duae uxores eius, Achinoam Iezrahelites et Abigail uxor Nabal de Carmel.
1SAM|27|4|Et nuntiatum est Saul quod fugisset David in Geth, et non addidit ultra ut quaereret eum.
1SAM|27|5|Dixit autem David ad Achis: " Si inveni gratiam in oculis tuis, detur mihi locus in una urbium regionis huius, ut habitem ibi. Cur enim manet servus tuus in civitate regis tecum? ".
1SAM|27|6|Dedit itaque ei Achis in die illa Siceleg; propter quam causam facta est Siceleg regum Iudae usque in diem hanc.
1SAM|27|7|Fuit autem numerus dierum, quibus habitavit David in regione Philisthinorum, annus et quattuor menses.
1SAM|27|8|Et ascendit David et viri eius et agebant praedas de Gesuri et de Gerzi et de Amalecitis; hae enim gentes habitabant terram, quae est a Telem in via Sur et usque ad terram Aegypti.
1SAM|27|9|Et percutiebat David omnem terram nec relinquebat viventem virum et mulierem; tollensque oves et boves et asinos et camelos et vestes revertebatur et veniebat ad Achis.
1SAM|27|10|Dicebat autem ei Achis: " In quem irruistis hodie? ". Respondebatque David: " Contra Nageb Iudae vel contra Nageb Ierameel vel contra Nageb Ceni ".
1SAM|27|11|Viro et mulieri non parcebat David nec adducebat in Geth dicens: " Ne forte loquantur adversum nos: "Haec fecit David" ". Et hoc erat decretum illi omnibus diebus, quibus habitavit in regione Philisthinorum.
1SAM|27|12|Credidit ergo Achis David dicens: " Valde odiosum se fecit populo suo Israel; eritigitur mihi servus sempiternus ".
1SAM|28|1|Factum est autem in diebus illis, congregaverunt Phili sthim agmina sua, ut praepararentur ad bellum contra Israel. Dixitque Achis ad David: " Sciens nunc scito quoniam mecum egredieris in castris tu et viri tui ".
1SAM|28|2|Dixitque David ad Achis: " Ideo tu quoque scies, quae facturus est servus tuus ". Et ait Achis ad David: " Ideo custodem capitis mei ponam te cunctis diebus ".
1SAM|28|3|Samuel autem mortuus erat; planxeratque eum omnis Israel, et sepelierant eum in Rama urbe sua. Et Saul abstulerat magos et hariolos de terra.
1SAM|28|4|Congregatique sunt Philisthim et venerunt et castrametati sunt in Sunam. Congregavit autem et Saul universum Israel, et castrametati sunt in Gelboe.
1SAM|28|5|Et vidit Saul castra Philisthim et timuit, et expavit cor eius nimis.
1SAM|28|6|Consuluitque Dominum, et non respondit ei neque per somnia neque per Urim neque per prophetas.
1SAM|28|7|Dixitque Saul servis suis: " Quaerite mihi mulierem habentem pythonem, et vadam ad eam et sciscitabor per illam ". Et dixerunt servi eius ad eum: Est mulier habens pythonem in Endor ".
1SAM|28|8|Mutavit ergo habitum suum vestitusque est aliis vestimentis et abiit ipse et duo viri cum eo; veneruntque ad mulierem nocte, et ait: " Divina mihi in pythone et suscita mihi, quem dixero tibi ".
1SAM|28|9|Et ait mulier ad eum: " Ecce tu nosti, quanta fecerit Saul et quomodo eraserit magos et hariolos de terra; quare ergo insidiaris animae meae, ut occidar? ".
1SAM|28|10|Et iuravit ei Saul in Domino dicens: " Vivit Dominus quia non veniet tibi quidquam mali propter hanc rem ".
1SAM|28|11|Dixitque ei mulier: " Quem suscitabo tibi? ". Qui ait: " Samuelem suscita mihi ".
1SAM|28|12|Cum autem vidisset mulier Samuelem, exclamavit voce magna et dixit ad Saul: " Quare imposuisti mihi? Tu es enim Saul! ".
1SAM|28|13|Dixitque ei rex: " Noli timere. Quid vidisti? ". Et ait mulier ad Saul: Hominem divinum vidi ascendentem de terra ".
1SAM|28|14|Dixitque ei: " Qualis est forma eius? ". Quae ait: " Vir senex ascendit et ipse amictus est pallio ". Intellexit Saul quod Samuel esset et inclinavit se super faciem suam in terra et adoravit.
1SAM|28|15|Dixit autem Samuel ad Saul: " Quare inquietasti me, ut suscitarer? ". Et ait Saul: " Coartor nimis. Siquidem Philisthim pugnant adversum me, et Deus recessit a me et exaudire me noluit neque in manu prophetarum neque per somnia; vocavi ergo te, ut ostenderes mihi quid faciam ".
1SAM|28|16|Et ait Samuel: " Quid interrogas me, cum Dominus recesserit a te et factus est adversarius tuus?
1SAM|28|17|Fecit enim Dominus, sicut locutus est in manu mea, et scidit regnum de manu tua et dedit illud proximo tuo David,
1SAM|28|18|quia non oboedisti voci Domini neque fecisti iram furoris eius in Amalec. Idcirco quod pateris, fecit tibi Dominus hodie.
1SAM|28|19|Et dabit Dominus etiam Israel tecum in manu Philisthim; cras autem tu et filii tui mecum eritis, sed et castra Israel tradet Dominus in manu Philisthim ".
1SAM|28|20|Statimque Saul cecidit porrectus in terram; extimuerat enim verba Samuel, et robur non erat in eo, quia non comederat panem tota die illa et tota nocte illa.
1SAM|28|21|Accessit itaque mulier ad Saul et vidit quod conturbatus esset valde; dixitque ad eum: " Ecce audivit ancilla tua vocem tuam, et posui animam meam in manu mea et oboedivi sermonibus tuis, quos locutus es ad me.
1SAM|28|22|Nunc igitur audi et tu vocem ancillae tuae, ut ponam coram te buccellam panis, et comedens convalescas, ut possis iter facere ".
1SAM|28|23|Qui renuit et ait: " Non comedam ". Coegerunt autem eum servi sui et mulier; et tandem, audita voce eorum, surrexit de terra et sedit super lectum.
1SAM|28|24|Mulier autem illa habebat vitulum pascualem in domo; et festinavit et occidit eum, tollensque farinam miscuit eam et coxit azyma.
1SAM|28|25|Et posuit ante Saul et ante servos eius. Qui cum comedissent, surrexerunt et abierunt hac eadem nocte.
1SAM|29|1|Congregata sunt ergo Philisthim universa agmina in Aphec; sed et Israel castrametatus est super fontem, qui erat in Iezrahel.
1SAM|29|2|Et principes quidem Philisthim incedebant in centuriis et milibus; David autem et viri eius incedebant in novissimo agmine cum Achis.
1SAM|29|3|Dixeruntque principes Philisthim: " Quid sibi volunt Hebraei isti? ". Et ait Achis ad principes Philisthim: " Nonne iste est David, qui fuit servus Saul regis Israel et est apud me multis diebus vel annis, et non inveni in eo quidquam ex die, qua transfugit ad me, usque ad diem hanc? ".
1SAM|29|4|Irati sunt autem adversus eum principes Philisthim et dixerunt ei: " Revertatur vir iste et sedeat in loco suo, in quo constituisti eum, et non descendat nobiscum in proelium, ne fiat nobis adversarius, cum proeliari coeperimus. Quomodo enim aliter placare poterit dominum suum nisi in capitibus horum virorum?
1SAM|29|5|Nonne iste est David, cui cantabant in choris dicentes: "Percussit Saul milia sua, et David decem milia sua"? ".
1SAM|29|6|Vocavit ergo Achis David et ait ei: " Vivit Dominus quia rectus es tu, et bonus est in conspectu meo exitus tuus et introitus tuus mecum in castris, et non inveni in te quidquam mali ex die, qua venisti ad me, usque ad diem hanc. Sed principibus non places.
1SAM|29|7|Revertere ergo et vade in pace et non offendes oculos principum Philisthim ".
1SAM|29|8|Dixitque David ad Achis: " Quid enim feci, et quid invenisti in me servo tuo a die, qua fui in conspectu tuo, usque in diem hanc, ut non veniam et pugnem contra inimicos domini mei regis? ".
1SAM|29|9|Respondens autem Achis locutus est ad David: " Scio quia bonus es tu in oculis meis sicut angelus Dei; sed principes Philisthim dixerunt: "Non ascendet nobiscum in proelium".
1SAM|29|10|Igitur consurge mane, tu et servi domini tui, qui venerunt tecum, et, cum de nocte surrexeritis et coeperit dilucescere, pergite ".
1SAM|29|11|Surrexit itaque de nocte David ipse et viri eius, ut proficiscerentur mane et reverterentur ad terram Philisthim. Philisthim autem ascenderunt in Iezrahel.
1SAM|30|1|Cumque venissent David et viri eius in Siceleg die tertia, Amalecitae impetum fecerant contra Nageb et contra Siceleg et percusserant Siceleg et succenderant eam igni;
1SAM|30|2|et captivas duxerant mulieres et omnes in ea a minimo usque ad magnum et non interfecerant quemquam, sed secum duxerant et pergebant in itinere suo.
1SAM|30|3|Cum ergo venisset David et viri eius ad civitatem et invenissent eam succensam igni et uxores suas et filios suos et filias ductas esse captivas,
1SAM|30|4|levaverunt David et populus, qui erat cum eo, voces suas et planxerunt, donec deficerent in eis lacrimae.
1SAM|30|5|Siquidem et duae uxores David captivae ductae fuerant, Achinoam Iezrahelites et Abigail uxor Nabal de Carmel.
1SAM|30|6|Et angustiatus est David valde; volebat enim eum populus lapidare, quia amara erat anima uniuscuiusque viri super filiis suis et filiabus. Confortatus est autem David in Domino Deo suo
1SAM|30|7|et ait ad Abiathar sacerdotem filium Achimelech: " Applica ad me ephod. Et applicuit Abiathar ephod ad David.
1SAM|30|8|Et consuluit David Dominum dicens: " Persequar latrunculos hos et comprehendam eos an non? ". Dixitque ei: " Persequere; absque dubio enim comprehendes eos et excuties praedam ".
1SAM|30|9|Abiit ergo David ipse et sescenti viri, qui erant cum eo, et venerunt usque ad torrentem Besor, et lassi quidam substiterunt.
1SAM|30|10|Persecutus est autem David ipse et quadringenti viri; et reliqui substiterunt: ducenti, qui lassi transire non poterant torrentem Besor.
1SAM|30|11|Et invenerunt virum Aegyptium in agro et adduxerunt eum ad David; dederuntque ei panem, et comedit, et dederunt ei aquam bibere,
1SAM|30|12|sed et dederunt ei fragmen massae caricarum et duas ligaturas uvae passae. Quae cum comedisset, reversus est spiritus eius; non enim comederat panem neque biberat aquam tribus diebus et tribus noctibus.
1SAM|30|13|Dixit itaque ei David: " Cuius es tu vel unde? ". Qui ait ei: " Puer Aegyptius ego sum servus viri Amalecitae; dereliquit autem me dominus meus, quia aegrotare coepi nudiustertius.
1SAM|30|14|Siquidem nos erupimus contra Nageb Cherethi et contra Nageb Iudae et Nageb Chaleb et Siceleg succendimus igni ".
1SAM|30|15|Dixitque ei David: " Potes me ducere ad istum cuneum? ". Qui ait: " Iura mihi per Deum quod non occidas me et non tradas me in manu domini mei, et ducam te ad cuneum istum ". Et iuravit ei David.
1SAM|30|16|Qui cum duxisset eum, ecce illi discumbebant super faciem universae terrae comedentes et bibentes et festum celebrantes pro cuncta praeda et spoliis, quae ceperant de terra Philisthim et de terra Iudae.
1SAM|30|17|Et percussit eos David die altera a diluculo usque ad vesperam, et non evasit ex eis quisquam, nisi quadringenti viri adulescentes, qui ascenderant camelos et fugerant.
1SAM|30|18|Eruit ergo David omnia, quae ceperant Amalecitae, et duas uxores suas eruit.
1SAM|30|19|Nec defuit quidquam a parvo usque ad magnum tam de filiis quam de filiabus et de spoliis, et, quaecumque rapuerant, omnia reduxit David.
1SAM|30|20|Cepit ergo David universos greges et armenta, et minaverunt ante faciem eius possessionem hanc dixeruntque: " Haec est praeda David ".
1SAM|30|21|Venit autem David ad ducentos viros, qui lassi substiterant nec sequi potuerant David, et residere eos iusserat in torrente Besor. Qui egressi sunt obviam David et populo, qui erat cum eo. Accedens autem David ad populum salutavit eos pacifice.
1SAM|30|22|Respondensque omnis vir pessimus et iniquus de viris, qui ierant cum David, dixit: " Quia non venerunt nobiscum, non dabimus eis quidquam de praeda, quam eruimus; sed sufficiat unicuique uxor sua et filii; quos cum acceperint, recedant ".
1SAM|30|23|Dixit autem David: " Non sic facietis, fratres mei, de his, quae tradidit Dominus nobis, et custodivit nos et dedit latrunculos, qui eruperant adversum nos, in manu nostra;
1SAM|30|24|nec audiet vos quisquam super sermone hoc; aequa enim pars erit descendentis ad proelium et remanentis ad sarcinas, et similiter divident.
1SAM|30|25|Et factum est hoc ex die illa et deinceps constitutum ut praeceptum et quasi lex in Israel usque ad diem hanc.
1SAM|30|26|Venit ergo David in Siceleg et misit dona de praeda senioribus Iudae proximis suis dicens: " Accipite benedictionem de praeda hostium Domini ";
1SAM|30|27|his, qui erant in Bethul et qui in Ramathnageb et qui in Iether
1SAM|30|28|et qui in Aroer et qui in Sephamoth et qui in Esthemo
1SAM|30|29|et qui in Carmel et qui in urbibus Ierameeli et qui in urbibus Ceni
1SAM|30|30|et qui in Horma et qui in Borasan et qui in Athach
1SAM|30|31|et qui in Hebron et reliquis locis, in quibus commoratus fuerat David ipse et viri eius.
1SAM|31|1|Philisthim autem pugnabant adversum Israel; et fugerunt viri Israel ante faciem Philisthim et ceciderunt interfecti in monte Gelboe.
1SAM|31|2|Irrueruntque Philisthim in Saul et filios eius et percusserunt Ionathan et Abinadab et Melchisua filios Saul.
1SAM|31|3|Totumque pondus proelii versum est in Saul; et consecuti sunt eum viri arcu, et vulneratus est vehementer a sagittariis.
1SAM|31|4|Dixitque Saul ad armigerum suum: " Evagina gladium tuum et percute me, ne forte veniant incircumcisi isti et confodiant me et illudant mihi ". Et noluit armiger eius; erat enim nimio timore perterritus. Arripuit itaque Saul gladium et irruit super eum.
1SAM|31|5|Quod cum vidisset armiger eius, videlicet quod mortuus esset Saul, irruit etiam ipse super gladium suum et mortuus est cum eo.
1SAM|31|6|Mortuus est ergo Saul et tres filii eius et armiger illius et universi viri eius in die illa pariter.
1SAM|31|7|Videntes autem viri Israel, qui erant trans vallem et trans Iordanem, quod fugissent viri Israelitae et quod mortuus esset Saul et filii eius, reliquerunt civitates suas et fugerunt. Veneruntque Philisthim et habitaverunt ibi.
1SAM|31|8|Facta autem die altera, venerunt Philisthim, ut spoliarent interfectos, et invenerunt Saul et tres filios eius iacentes in monte Gelboe.
1SAM|31|9|Et praeciderunt caput Saul et exspoliaverunt eum armis, quae miserunt in terram Philisthinorum per circuitum, ut annuntiaretur in templis idolorum suorum et populo.
1SAM|31|10|Et posuerunt arma eius in templo Astharoth, corpus vero eius suspenderunt in muro Bethsan.
1SAM|31|11|Quod cum audissent habitatores Iabes Galaad, quaecumque fecerant Philisthim Saul,
1SAM|31|12|surrexerunt omnes viri fortissimi et ambulaverunt tota nocte et tulerunt cadaver Saul et cadavera filiorum eius de muro Bethsan; veneruntque Iabes et combusserunt ea ibi.
1SAM|31|13|Et tulerunt ossa eorum et sepelierunt sub myrice in Iabes et ieiunaverunt septem diebus.
