1COR|1|1|Paul, called to be an apostle of Christ Jesus by the will of God, and our brother Sosthenes,
1COR|1|2|To the church of God in Corinth, to those sanctified in Christ Jesus and called to be holy, together with all those everywhere who call on the name of our Lord Jesus Christ--their Lord and ours:
1COR|1|3|Grace and peace to you from God our Father and the Lord Jesus Christ.
1COR|1|4|I always thank God for you because of his grace given you in Christ Jesus.
1COR|1|5|For in him you have been enriched in every way--in all your speaking and in all your knowledge--
1COR|1|6|because our testimony about Christ was confirmed in you.
1COR|1|7|Therefore you do not lack any spiritual gift as you eagerly wait for our Lord Jesus Christ to be revealed.
1COR|1|8|He will keep you strong to the end, so that you will be blameless on the day of our Lord Jesus Christ.
1COR|1|9|God, who has called you into fellowship with his Son Jesus Christ our Lord, is faithful.
1COR|1|10|I appeal to you, brothers, in the name of our Lord Jesus Christ, that all of you agree with one another so that there may be no divisions among you and that you may be perfectly united in mind and thought.
1COR|1|11|My brothers, some from Chloe's household have informed me that there are quarrels among you.
1COR|1|12|What I mean is this: One of you says, "I follow Paul"; another, "I follow Apollos"; another, "I follow Cephas "; still another, "I follow Christ."
1COR|1|13|Is Christ divided? Was Paul crucified for you? Were you baptized into the name of Paul?
1COR|1|14|I am thankful that I did not baptize any of you except Crispus and Gaius,
1COR|1|15|so no one can say that you were baptized into my name.
1COR|1|16|(Yes, I also baptized the household of Stephanas; beyond that, I don't remember if I baptized anyone else.)
1COR|1|17|For Christ did not send me to baptize, but to preach the gospel--not with words of human wisdom, lest the cross of Christ be emptied of its power.
1COR|1|18|For the message of the cross is foolishness to those who are perishing, but to us who are being saved it is the power of God.
1COR|1|19|For it is written: "I will destroy the wisdom of the wise; the intelligence of the intelligent I will frustrate."
1COR|1|20|Where is the wise man? Where is the scholar? Where is the philosopher of this age? Has not God made foolish the wisdom of the world?
1COR|1|21|For since in the wisdom of God the world through its wisdom did not know him, God was pleased through the foolishness of what was preached to save those who believe.
1COR|1|22|Jews demand miraculous signs and Greeks look for wisdom,
1COR|1|23|but we preach Christ crucified: a stumbling block to Jews and foolishness to Gentiles,
1COR|1|24|but to those whom God has called, both Jews and Greeks, Christ the power of God and the wisdom of God.
1COR|1|25|For the foolishness of God is wiser than man's wisdom, and the weakness of God is stronger than man's strength.
1COR|1|26|Brothers, think of what you were when you were called. Not many of you were wise by human standards; not many were influential; not many were of noble birth.
1COR|1|27|But God chose the foolish things of the world to shame the wise; God chose the weak things of the world to shame the strong.
1COR|1|28|He chose the lowly things of this world and the despised things--and the things that are not--to nullify the things that are,
1COR|1|29|so that no one may boast before him.
1COR|1|30|It is because of him that you are in Christ Jesus, who has become for us wisdom from God--that is, our righteousness, holiness and redemption.
1COR|1|31|Therefore, as it is written: "Let him who boasts boast in the Lord."
1COR|2|1|When I came to you, brothers, I did not come with eloquence or superior wisdom as I proclaimed to you the testimony about God.
1COR|2|2|For I resolved to know nothing while I was with you except Jesus Christ and him crucified.
1COR|2|3|I came to you in weakness and fear, and with much trembling.
1COR|2|4|My message and my preaching were not with wise and persuasive words, but with a demonstration of the Spirit's power,
1COR|2|5|so that your faith might not rest on men's wisdom, but on God's power.
1COR|2|6|We do, however, speak a message of wisdom among the mature, but not the wisdom of this age or of the rulers of this age, who are coming to nothing.
1COR|2|7|No, we speak of God's secret wisdom, a wisdom that has been hidden and that God destined for our glory before time began.
1COR|2|8|None of the rulers of this age understood it, for if they had, they would not have crucified the Lord of glory.
1COR|2|9|However, as it is written: "No eye has seen, no ear has heard, no mind has conceived what God has prepared for those who love him"--
1COR|2|10|but God has revealed it to us by his Spirit.
1COR|2|11|The Spirit searches all things, even the deep things of God. For who among men knows the thoughts of a man except the man's spirit within him? In the same way no one knows the thoughts of God except the Spirit of God.
1COR|2|12|We have not received the spirit of the world but the Spirit who is from God, that we may understand what God has freely given us.
1COR|2|13|This is what we speak, not in words taught us by human wisdom but in words taught by the Spirit, expressing spiritual truths in spiritual words.
1COR|2|14|The man without the Spirit does not accept the things that come from the Spirit of God, for they are foolishness to him, and he cannot understand them, because they are spiritually discerned.
1COR|2|15|The spiritual man makes judgments about all things, but he himself is not subject to any man's judgment:
1COR|2|16|"For who has known the mind of the Lord that he may instruct him?" But we have the mind of Christ.
1COR|3|1|Brothers, I could not address you as spiritual but as worldly--mere infants in Christ.
1COR|3|2|I gave you milk, not solid food, for you were not yet ready for it. Indeed, you are still not ready.
1COR|3|3|You are still worldly. For since there is jealousy and quarreling among you, are you not worldly? Are you not acting like mere men?
1COR|3|4|For when one says, "I follow Paul," and another, "I follow Apollos," are you not mere men?
1COR|3|5|What, after all, is Apollos? And what is Paul? Only servants, through whom you came to believe--as the Lord has assigned to each his task.
1COR|3|6|I planted the seed, Apollos watered it, but God made it grow.
1COR|3|7|So neither he who plants nor he who waters is anything, but only God, who makes things grow.
1COR|3|8|The man who plants and the man who waters have one purpose, and each will be rewarded according to his own labor.
1COR|3|9|For we are God's fellow workers; you are God's field, God's building.
1COR|3|10|By the grace God has given me, I laid a foundation as an expert builder, and someone else is building on it. But each one should be careful how he builds.
1COR|3|11|For no one can lay any foundation other than the one already laid, which is Jesus Christ.
1COR|3|12|If any man builds on this foundation using gold, silver, costly stones, wood, hay or straw,
1COR|3|13|his work will be shown for what it is, because the Day will bring it to light. It will be revealed with fire, and the fire will test the quality of each man's work.
1COR|3|14|If what he has built survives, he will receive his reward.
1COR|3|15|If it is burned up, he will suffer loss; he himself will be saved, but only as one escaping through the flames.
1COR|3|16|Don't you know that you yourselves are God's temple and that God's Spirit lives in you?
1COR|3|17|If anyone destroys God's temple, God will destroy him; for God's temple is sacred, and you are that temple.
1COR|3|18|Do not deceive yourselves. If any one of you thinks he is wise by the standards of this age, he should become a "fool" so that he may become wise.
1COR|3|19|For the wisdom of this world is foolishness in God's sight. As it is written: "He catches the wise in their craftiness";
1COR|3|20|and again, "The Lord knows that the thoughts of the wise are futile."
1COR|3|21|So then, no more boasting about men! All things are yours,
1COR|3|22|whether Paul or Apollos or Cephas or the world or life or death or the present or the future--all are yours,
1COR|3|23|and you are of Christ, and Christ is of God.
1COR|4|1|So then, men ought to regard us as servants of Christ and as those entrusted with the secret things of God.
1COR|4|2|Now it is required that those who have been given a trust must prove faithful.
1COR|4|3|I care very little if I am judged by you or by any human court; indeed, I do not even judge myself.
1COR|4|4|My conscience is clear, but that does not make me innocent. It is the Lord who judges me.
1COR|4|5|Therefore judge nothing before the appointed time; wait till the Lord comes. He will bring to light what is hidden in darkness and will expose the motives of men's hearts. At that time each will receive his praise from God.
1COR|4|6|Now, brothers, I have applied these things to myself and Apollos for your benefit, so that you may learn from us the meaning of the saying, "Do not go beyond what is written." Then you will not take pride in one man over against another.
1COR|4|7|For who makes you different from anyone else? What do you have that you did not receive? And if you did receive it, why do you boast as though you did not?
1COR|4|8|Already you have all you want! Already you have become rich! You have become kings--and that without us! How I wish that you really had become kings so that we might be kings with you!
1COR|4|9|For it seems to me that God has put us apostles on display at the end of the procession, like men condemned to die in the arena. We have been made a spectacle to the whole universe, to angels as well as to men.
1COR|4|10|We are fools for Christ, but you are so wise in Christ! We are weak, but you are strong! You are honored, we are dishonored!
1COR|4|11|To this very hour we go hungry and thirsty, we are in rags, we are brutally treated, we are homeless.
1COR|4|12|We work hard with our own hands. When we are cursed, we bless; when we are persecuted, we endure it;
1COR|4|13|when we are slandered, we answer kindly. Up to this moment we have become the scum of the earth, the refuse of the world.
1COR|4|14|I am not writing this to shame you, but to warn you, as my dear children.
1COR|4|15|Even though you have ten thousand guardians in Christ, you do not have many fathers, for in Christ Jesus I became your father through the gospel.
1COR|4|16|Therefore I urge you to imitate me.
1COR|4|17|For this reason I am sending to you Timothy, my son whom I love, who is faithful in the Lord. He will remind you of my way of life in Christ Jesus, which agrees with what I teach everywhere in every church.
1COR|4|18|Some of you have become arrogant, as if I were not coming to you.
1COR|4|19|But I will come to you very soon, if the Lord is willing, and then I will find out not only how these arrogant people are talking, but what power they have.
1COR|4|20|For the kingdom of God is not a matter of talk but of power.
1COR|4|21|What do you prefer? Shall I come to you with a whip, or in love and with a gentle spirit?
1COR|5|1|It is actually reported that there is sexual immorality among you, and of a kind that does not occur even among pagans: A man has his father's wife.
1COR|5|2|And you are proud! Shouldn't you rather have been filled with grief and have put out of your fellowship the man who did this?
1COR|5|3|Even though I am not physically present, I am with you in spirit. And I have already passed judgment on the one who did this, just as if I were present.
1COR|5|4|When you are assembled in the name of our Lord Jesus and I am with you in spirit, and the power of our Lord Jesus is present,
1COR|5|5|hand this man over to Satan, so that the sinful nature may be destroyed and his spirit saved on the day of the Lord.
1COR|5|6|Your boasting is not good. Don't you know that a little yeast works through the whole batch of dough?
1COR|5|7|Get rid of the old yeast that you may be a new batch without yeast--as you really are. For Christ, our Passover lamb, has been sacrificed.
1COR|5|8|Therefore let us keep the Festival, not with the old yeast, the yeast of malice and wickedness, but with bread without yeast, the bread of sincerity and truth.
1COR|5|9|I have written you in my letter not to associate with sexually immoral people--
1COR|5|10|not at all meaning the people of this world who are immoral, or the greedy and swindlers, or idolaters. In that case you would have to leave this world.
1COR|5|11|But now I am writing you that you must not associate with anyone who calls himself a brother but is sexually immoral or greedy, an idolater or a slanderer, a drunkard or a swindler. With such a man do not even eat.
1COR|5|12|What business is it of mine to judge those outside the church? Are you not to judge those inside?
1COR|5|13|God will judge those outside. "Expel the wicked man from among you."
1COR|6|1|If any of you has a dispute with another, dare he take it before the ungodly for judgment instead of before the saints?
1COR|6|2|Do you not know that the saints will judge the world? And if you are to judge the world, are you not competent to judge trivial cases?
1COR|6|3|Do you not know that we will judge angels? How much more the things of this life!
1COR|6|4|Therefore, if you have disputes about such matters, appoint as judges even men of little account in the church!
1COR|6|5|I say this to shame you. Is it possible that there is nobody among you wise enough to judge a dispute between believers?
1COR|6|6|But instead, one brother goes to law against another--and this in front of unbelievers!
1COR|6|7|The very fact that you have lawsuits among you means you have been completely defeated already. Why not rather be wronged? Why not rather be cheated?
1COR|6|8|Instead, you yourselves cheat and do wrong, and you do this to your brothers.
1COR|6|9|Do you not know that the wicked will not inherit the kingdom of God? Do not be deceived: Neither the sexually immoral nor idolaters nor adulterers nor male prostitutes nor homosexual offenders
1COR|6|10|nor thieves nor the greedy nor drunkards nor slanderers nor swindlers will inherit the kingdom of God.
1COR|6|11|And that is what some of you were. But you were washed, you were sanctified, you were justified in the name of the Lord Jesus Christ and by the Spirit of our God.
1COR|6|12|"Everything is permissible for me"--but not everything is beneficial. "Everything is permissible for me"--but I will not be mastered by anything.
1COR|6|13|"Food for the stomach and the stomach for food"--but God will destroy them both. The body is not meant for sexual immorality, but for the Lord, and the Lord for the body.
1COR|6|14|By his power God raised the Lord from the dead, and he will raise us also.
1COR|6|15|Do you not know that your bodies are members of Christ himself? Shall I then take the members of Christ and unite them with a prostitute? Never!
1COR|6|16|Do you not know that he who unites himself with a prostitute is one with her in body? For it is said, "The two will become one flesh."
1COR|6|17|But he who unites himself with the Lord is one with him in spirit.
1COR|6|18|Flee from sexual immorality. All other sins a man commits are outside his body, but he who sins sexually sins against his own body.
1COR|6|19|Do you not know that your body is a temple of the Holy Spirit, who is in you, whom you have received from God? You are not your own;
1COR|6|20|you were bought at a price. Therefore honor God with your body.
1COR|7|1|Now for the matters you wrote about: It is good for a man not to marry.
1COR|7|2|But since there is so much immorality, each man should have his own wife, and each woman her own husband.
1COR|7|3|The husband should fulfill his marital duty to his wife, and likewise the wife to her husband.
1COR|7|4|The wife's body does not belong to her alone but also to her husband. In the same way, the husband's body does not belong to him alone but also to his wife.
1COR|7|5|Do not deprive each other except by mutual consent and for a time, so that you may devote yourselves to prayer. Then come together again so that Satan will not tempt you because of your lack of self-control.
1COR|7|6|I say this as a concession, not as a command.
1COR|7|7|I wish that all men were as I am. But each man has his own gift from God; one has this gift, another has that.
1COR|7|8|Now to the unmarried and the widows I say: It is good for them to stay unmarried, as I am.
1COR|7|9|But if they cannot control themselves, they should marry, for it is better to marry than to burn with passion.
1COR|7|10|To the married I give this command (not I, but the Lord): A wife must not separate from her husband.
1COR|7|11|But if she does, she must remain unmarried or else be reconciled to her husband. And a husband must not divorce his wife.
1COR|7|12|To the rest I say this (I, not the Lord): If any brother has a wife who is not a believer and she is willing to live with him, he must not divorce her.
1COR|7|13|And if a woman has a husband who is not a believer and he is willing to live with her, she must not divorce him.
1COR|7|14|For the unbelieving husband has been sanctified through his wife, and the unbelieving wife has been sanctified through her believing husband. Otherwise your children would be unclean, but as it is, they are holy.
1COR|7|15|But if the unbeliever leaves, let him do so. A believing man or woman is not bound in such circumstances; God has called us to live in peace.
1COR|7|16|How do you know, wife, whether you will save your husband? Or, how do you know, husband, whether you will save your wife?
1COR|7|17|Nevertheless, each one should retain the place in life that the Lord assigned to him and to which God has called him. This is the rule I lay down in all the churches.
1COR|7|18|Was a man already circumcised when he was called? He should not become uncircumcised. Was a man uncircumcised when he was called? He should not be circumcised.
1COR|7|19|Circumcision is nothing and uncircumcision is nothing. Keeping God's commands is what counts.
1COR|7|20|Each one should remain in the situation which he was in when God called him.
1COR|7|21|Were you a slave when you were called? Don't let it trouble you--although if you can gain your freedom, do so.
1COR|7|22|For he who was a slave when he was called by the Lord is the Lord's freedman; similarly, he who was a free man when he was called is Christ's slave.
1COR|7|23|You were bought at a price; do not become slaves of men.
1COR|7|24|Brothers, each man, as responsible to God, should remain in the situation God called him to.
1COR|7|25|Now about virgins: I have no command from the Lord, but I give a judgment as one who by the Lord's mercy is trustworthy.
1COR|7|26|Because of the present crisis, I think that it is good for you to remain as you are.
1COR|7|27|Are you married? Do not seek a divorce. Are you unmarried? Do not look for a wife.
1COR|7|28|But if you do marry, you have not sinned; and if a virgin marries, she has not sinned. But those who marry will face many troubles in this life, and I want to spare you this.
1COR|7|29|What I mean, brothers, is that the time is short. From now on those who have wives should live as if they had none;
1COR|7|30|those who mourn, as if they did not; those who are happy, as if they were not; those who buy something, as if it were not theirs to keep;
1COR|7|31|those who use the things of the world, as if not engrossed in them. For this world in its present form is passing away.
1COR|7|32|I would like you to be free from concern. An unmarried man is concerned about the Lord's affairs--how he can please the Lord.
1COR|7|33|But a married man is concerned about the affairs of this world--how he can please his wife--
1COR|7|34|and his interests are divided. An unmarried woman or virgin is concerned about the Lord's affairs: Her aim is to be devoted to the Lord in both body and spirit. But a married woman is concerned about the affairs of this world--how she can please her husband.
1COR|7|35|I am saying this for your own good, not to restrict you, but that you may live in a right way in undivided devotion to the Lord.
1COR|7|36|If anyone thinks he is acting improperly toward the virgin he is engaged to, and if she is getting along in years and he feels he ought to marry, he should do as he wants. He is not sinning. They should get married.
1COR|7|37|But the man who has settled the matter in his own mind, who is under no compulsion but has control over his own will, and who has made up his mind not to marry the virgin--this man also does the right thing.
1COR|7|38|So then, he who marries the virgin does right, but he who does not marry her does even better.
1COR|7|39|A woman is bound to her husband as long as he lives. But if her husband dies, she is free to marry anyone she wishes, but he must belong to the Lord.
1COR|7|40|In my judgment, she is happier if she stays as she is--and I think that I too have the Spirit of God.
1COR|8|1|Now about food sacrificed to idols: We know that we all possess knowledge. Knowledge puffs up, but love builds up.
1COR|8|2|The man who thinks he knows something does not yet know as he ought to know.
1COR|8|3|But the man who loves God is known by God.
1COR|8|4|So then, about eating food sacrificed to idols: We know that an idol is nothing at all in the world and that there is no God but one.
1COR|8|5|For even if there are so-called gods, whether in heaven or on earth (as indeed there are many "gods" and many "lords"),
1COR|8|6|yet for us there is but one God, the Father, from whom all things came and for whom we live; and there is but one Lord, Jesus Christ, through whom all things came and through whom we live.
1COR|8|7|But not everyone knows this. Some people are still so accustomed to idols that when they eat such food they think of it as having been sacrificed to an idol, and since their conscience is weak, it is defiled.
1COR|8|8|But food does not bring us near to God; we are no worse if we do not eat, and no better if we do.
1COR|8|9|Be careful, however, that the exercise of your freedom does not become a stumbling block to the weak.
1COR|8|10|For if anyone with a weak conscience sees you who have this knowledge eating in an idol's temple, won't he be emboldened to eat what has been sacrificed to idols?
1COR|8|11|So this weak brother, for whom Christ died, is destroyed by your knowledge.
1COR|8|12|When you sin against your brothers in this way and wound their weak conscience, you sin against Christ.
1COR|8|13|Therefore, if what I eat causes my brother to fall into sin, I will never eat meat again, so that I will not cause him to fall.
1COR|9|1|Am I not free? Am I not an apostle? Have I not seen Jesus our Lord? Are you not the result of my work in the Lord?
1COR|9|2|Even though I may not be an apostle to others, surely I am to you! For you are the seal of my apostleship in the Lord.
1COR|9|3|This is my defense to those who sit in judgment on me.
1COR|9|4|Don't we have the right to food and drink?
1COR|9|5|Don't we have the right to take a believing wife along with us, as do the other apostles and the Lord's brothers and Cephas?
1COR|9|6|Or is it only I and Barnabas who must work for a living?
1COR|9|7|Who serves as a soldier at his own expense? Who plants a vineyard and does not eat of its grapes? Who tends a flock and does not drink of the milk?
1COR|9|8|Do I say this merely from a human point of view? Doesn't the Law say the same thing?
1COR|9|9|For it is written in the Law of Moses: "Do not muzzle an ox while it is treading out the grain." Is it about oxen that God is concerned?
1COR|9|10|Surely he says this for us, doesn't he? Yes, this was written for us, because when the plowman plows and the thresher threshes, they ought to do so in the hope of sharing in the harvest.
1COR|9|11|If we have sown spiritual seed among you, is it too much if we reap a material harvest from you?
1COR|9|12|If others have this right of support from you, shouldn't we have it all the more?
1COR|9|13|But we did not use this right. On the contrary, we put up with anything rather than hinder the gospel of Christ. Don't you know that those who work in the temple get their food from the temple, and those who serve at the altar share in what is offered on the altar?
1COR|9|14|In the same way, the Lord has commanded that those who preach the gospel should receive their living from the gospel.
1COR|9|15|But I have not used any of these rights. And I am not writing this in the hope that you will do such things for me. I would rather die than have anyone deprive me of this boast.
1COR|9|16|Yet when I preach the gospel, I cannot boast, for I am compelled to preach. Woe to me if I do not preach the gospel!
1COR|9|17|If I preach voluntarily, I have a reward; if not voluntarily, I am simply discharging the trust committed to me.
1COR|9|18|What then is my reward? Just this: that in preaching the gospel I may offer it free of charge, and so not make use of my rights in preaching it.
1COR|9|19|Though I am free and belong to no man, I make myself a slave to everyone, to win as many as possible.
1COR|9|20|To the Jews I became like a Jew, to win the Jews. To those under the law I became like one under the law (though I myself am not under the law), so as to win those under the law.
1COR|9|21|To those not having the law I became like one not having the law (though I am not free from God's law but am under Christ's law), so as to win those not having the law.
1COR|9|22|To the weak I became weak, to win the weak. I have become all things to all men so that by all possible means I might save some.
1COR|9|23|I do all this for the sake of the gospel, that I may share in its blessings.
1COR|9|24|Do you not know that in a race all the runners run, but only one gets the prize? Run in such a way as to get the prize.
1COR|9|25|Everyone who competes in the games goes into strict training. They do it to get a crown that will not last; but we do it to get a crown that will last forever.
1COR|9|26|Therefore I do not run like a man running aimlessly; I do not fight like a man beating the air.
1COR|9|27|No, I beat my body and make it my slave so that after I have preached to others, I myself will not be disqualified for the prize.
1COR|10|1|For I do not want you to be ignorant of the fact, brothers, that our forefathers were all under the cloud and that they all passed through the sea.
1COR|10|2|They were all baptized into Moses in the cloud and in the sea.
1COR|10|3|They all ate the same spiritual food
1COR|10|4|and drank the same spiritual drink; for they drank from the spiritual rock that accompanied them, and that rock was Christ.
1COR|10|5|Nevertheless, God was not pleased with most of them; their bodies were scattered over the desert.
1COR|10|6|Now these things occurred as examples to keep us from setting our hearts on evil things as they did.
1COR|10|7|Do not be idolaters, as some of them were; as it is written: "The people sat down to eat and drink and got up to indulge in pagan revelry."
1COR|10|8|We should not commit sexual immorality, as some of them did--and in one day twenty-three thousand of them died.
1COR|10|9|We should not test the Lord, as some of them did--and were killed by snakes.
1COR|10|10|And do not grumble, as some of them did--and were killed by the destroying angel.
1COR|10|11|These things happened to them as examples and were written down as warnings for us, on whom the fulfillment of the ages has come.
1COR|10|12|So, if you think you are standing firm, be careful that you don't fall!
1COR|10|13|No temptation has seized you except what is common to man. And God is faithful; he will not let you be tempted beyond what you can bear. But when you are tempted, he will also provide a way out so that you can stand up under it.
1COR|10|14|Therefore, my dear friends, flee from idolatry.
1COR|10|15|I speak to sensible people; judge for yourselves what I say.
1COR|10|16|Is not the cup of thanksgiving for which we give thanks a participation in the blood of Christ? And is not the bread that we break a participation in the body of Christ?
1COR|10|17|Because there is one loaf, we, who are many, are one body, for we all partake of the one loaf.
1COR|10|18|Consider the people of Israel: Do not those who eat the sacrifices participate in the altar?
1COR|10|19|Do I mean then that a sacrifice offered to an idol is anything, or that an idol is anything?
1COR|10|20|No, but the sacrifices of pagans are offered to demons, not to God, and I do not want you to be participants with demons.
1COR|10|21|You cannot drink the cup of the Lord and the cup of demons too; you cannot have a part in both the Lord's table and the table of demons.
1COR|10|22|Are we trying to arouse the Lord's jealousy? Are we stronger than he?
1COR|10|23|"Everything is permissible"--but not everything is beneficial. "Everything is permissible"--but not everything is constructive.
1COR|10|24|Nobody should seek his own good, but the good of others.
1COR|10|25|Eat anything sold in the meat market without raising questions of conscience,
1COR|10|26|for, "The earth is the Lord's, and everything in it."
1COR|10|27|If some unbeliever invites you to a meal and you want to go, eat whatever is put before you without raising questions of conscience.
1COR|10|28|But if anyone says to you, "This has been offered in sacrifice," then do not eat it, both for the sake of the man who told you and for conscience' sake--
1COR|10|29|the other man's conscience, I mean, not yours. For why should my freedom be judged by another's conscience?
1COR|10|30|If I take part in the meal with thankfulness, why am I denounced because of something I thank God for?
1COR|10|31|So whether you eat or drink or whatever you do, do it all for the glory of God.
1COR|10|32|Do not cause anyone to stumble, whether Jews, Greeks or the church of God--
1COR|10|33|even as I try to please everybody in every way. For I am not seeking my own good but the good of many, so that they may be saved.
1COR|11|1|Follow my example, as I follow the example of Christ.
1COR|11|2|I praise you for remembering me in everything and for holding to the teachings, just as I passed them on to you.
1COR|11|3|Now I want you to realize that the head of every man is Christ, and the head of the woman is man, and the head of Christ is God.
1COR|11|4|Every man who prays or prophesies with his head covered dishonors his head.
1COR|11|5|And every woman who prays or prophesies with her head uncovered dishonors her head--it is just as though her head were shaved.
1COR|11|6|If a woman does not cover her head, she should have her hair cut off; and if it is a disgrace for a woman to have her hair cut or shaved off, she should cover her head.
1COR|11|7|A man ought not to cover his head, since he is the image and glory of God; but the woman is the glory of man.
1COR|11|8|For man did not come from woman, but woman from man;
1COR|11|9|neither was man created for woman, but woman for man.
1COR|11|10|For this reason, and because of the angels, the woman ought to have a sign of authority on her head.
1COR|11|11|In the Lord, however, woman is not independent of man, nor is man independent of woman.
1COR|11|12|For as woman came from man, so also man is born of woman. But everything comes from God.
1COR|11|13|Judge for yourselves: Is it proper for a woman to pray to God with her head uncovered?
1COR|11|14|Does not the very nature of things teach you that if a man has long hair, it is a disgrace to him,
1COR|11|15|but that if a woman has long hair, it is her glory? For long hair is given to her as a covering.
1COR|11|16|If anyone wants to be contentious about this, we have no other practice--nor do the churches of God.
1COR|11|17|In the following directives I have no praise for you, for your meetings do more harm than good.
1COR|11|18|In the first place, I hear that when you come together as a church, there are divisions among you, and to some extent I believe it.
1COR|11|19|No doubt there have to be differences among you to show which of you have God's approval.
1COR|11|20|When you come together, it is not the Lord's Supper you eat,
1COR|11|21|for as you eat, each of you goes ahead without waiting for anybody else. One remains hungry, another gets drunk.
1COR|11|22|Don't you have homes to eat and drink in? Or do you despise the church of God and humiliate those who have nothing? What shall I say to you? Shall I praise you for this? Certainly not!
1COR|11|23|For I received from the Lord what I also passed on to you: The Lord Jesus, on the night he was betrayed, took bread,
1COR|11|24|and when he had given thanks, he broke it and said, "This is my body, which is for you; do this in remembrance of me."
1COR|11|25|In the same way, after supper he took the cup, saying, "This cup is the new covenant in my blood; do this, whenever you drink it, in remembrance of me."
1COR|11|26|For whenever you eat this bread and drink this cup, you proclaim the Lord's death until he comes.
1COR|11|27|Therefore, whoever eats the bread or drinks the cup of the Lord in an unworthy manner will be guilty of sinning against the body and blood of the Lord.
1COR|11|28|A man ought to examine himself before he eats of the bread and drinks of the cup.
1COR|11|29|For anyone who eats and drinks without recognizing the body of the Lord eats and drinks judgment on himself.
1COR|11|30|That is why many among you are weak and sick, and a number of you have fallen asleep.
1COR|11|31|But if we judged ourselves, we would not come under judgment.
1COR|11|32|When we are judged by the Lord, we are being disciplined so that we will not be condemned with the world.
1COR|11|33|So then, my brothers, when you come together to eat, wait for each other.
1COR|11|34|If anyone is hungry, he should eat at home, so that when you meet together it may not result in judgment. And when I come I will give further directions.
1COR|12|1|Now about spiritual gifts, brothers, I do not want you to be ignorant.
1COR|12|2|You know that when you were pagans, somehow or other you were influenced and led astray to mute idols.
1COR|12|3|Therefore I tell you that no one who is speaking by the Spirit of God says, "Jesus be cursed," and no one can say, "Jesus is Lord," except by the Holy Spirit.
1COR|12|4|There are different kinds of gifts, but the same Spirit.
1COR|12|5|There are different kinds of service, but the same Lord.
1COR|12|6|There are different kinds of working, but the same God works all of them in all men.
1COR|12|7|Now to each one the manifestation of the Spirit is given for the common good.
1COR|12|8|To one there is given through the Spirit the message of wisdom, to another the message of knowledge by means of the same Spirit,
1COR|12|9|to another faith by the same Spirit, to another gifts of healing by that one Spirit,
1COR|12|10|to another miraculous powers, to another prophecy, to another distinguishing between spirits, to another speaking in different kinds of tongues, and to still another the interpretation of tongues.
1COR|12|11|All these are the work of one and the same Spirit, and he gives them to each one, just as he determines.
1COR|12|12|The body is a unit, though it is made up of many parts; and though all its parts are many, they form one body. So it is with Christ.
1COR|12|13|For we were all baptized by one Spirit into one body--whether Jews or Greeks, slave or free--and we were all given the one Spirit to drink.
1COR|12|14|Now the body is not made up of one part but of many.
1COR|12|15|If the foot should say, "Because I am not a hand, I do not belong to the body," it would not for that reason cease to be part of the body.
1COR|12|16|And if the ear should say, "Because I am not an eye, I do not belong to the body," it would not for that reason cease to be part of the body.
1COR|12|17|If the whole body were an eye, where would the sense of hearing be? If the whole body were an ear, where would the sense of smell be?
1COR|12|18|But in fact God has arranged the parts in the body, every one of them, just as he wanted them to be.
1COR|12|19|If they were all one part, where would the body be?
1COR|12|20|As it is, there are many parts, but one body.
1COR|12|21|The eye cannot say to the hand, "I don't need you!" And the head cannot say to the feet, "I don't need you!"
1COR|12|22|On the contrary, those parts of the body that seem to be weaker are indispensable,
1COR|12|23|and the parts that we think are less honorable we treat with special honor. And the parts that are unpresentable are treated with special modesty,
1COR|12|24|while our presentable parts need no special treatment. But God has combined the members of the body and has given greater honor to the parts that lacked it,
1COR|12|25|so that there should be no division in the body, but that its parts should have equal concern for each other.
1COR|12|26|If one part suffers, every part suffers with it; if one part is honored, every part rejoices with it.
1COR|12|27|Now you are the body of Christ, and each one of you is a part of it.
1COR|12|28|And in the church God has appointed first of all apostles, second prophets, third teachers, then workers of miracles, also those having gifts of healing, those able to help others, those with gifts of administration, and those speaking in different kinds of tongues.
1COR|12|29|Are all apostles? Are all prophets? Are all teachers? Do all work miracles?
1COR|12|30|Do all have gifts of healing? Do all speak in tongues? Do all interpret?
1COR|12|31|But eagerly desire the greater gifts. And now I will show you the most excellent way.
1COR|13|1|If I speak in the tongues of men and of angels, but have not love, I am only a resounding gong or a clanging cymbal.
1COR|13|2|If I have the gift of prophecy and can fathom all mysteries and all knowledge, and if I have a faith that can move mountains, but have not love, I am nothing.
1COR|13|3|If I give all I possess to the poor and surrender my body to the flames, but have not love, I gain nothing.
1COR|13|4|Love is patient, love is kind. It does not envy, it does not boast, it is not proud.
1COR|13|5|It is not rude, it is not self-seeking, it is not easily angered, it keeps no record of wrongs.
1COR|13|6|Love does not delight in evil but rejoices with the truth.
1COR|13|7|It always protects, always trusts, always hopes, always perseveres.
1COR|13|8|Love never fails. But where there are prophecies, they will cease; where there are tongues, they will be stilled; where there is knowledge, it will pass away.
1COR|13|9|For we know in part and we prophesy in part,
1COR|13|10|but when perfection comes, the imperfect disappears.
1COR|13|11|When I was a child, I talked like a child, I thought like a child, I reasoned like a child. When I became a man, I put childish ways behind me.
1COR|13|12|Now we see but a poor reflection as in a mirror; then we shall see face to face. Now I know in part; then I shall know fully, even as I am fully known.
1COR|13|13|And now these three remain: faith, hope and love. But the greatest of these is love.
1COR|14|1|Follow the way of love and eagerly desire spiritual gifts, especially the gift of prophecy.
1COR|14|2|For anyone who speaks in a tongue does not speak to men but to God. Indeed, no one understands him; he utters mysteries with his spirit.
1COR|14|3|But everyone who prophesies speaks to men for their strengthening, encouragement and comfort.
1COR|14|4|He who speaks in a tongue edifies himself, but he who prophesies edifies the church.
1COR|14|5|I would like every one of you to speak in tongues, but I would rather have you prophesy. He who prophesies is greater than one who speaks in tongues, unless he interprets, so that the church may be edified.
1COR|14|6|Now, brothers, if I come to you and speak in tongues, what good will I be to you, unless I bring you some revelation or knowledge or prophecy or word of instruction?
1COR|14|7|Even in the case of lifeless things that make sounds, such as the flute or harp, how will anyone know what tune is being played unless there is a distinction in the notes?
1COR|14|8|Again, if the trumpet does not sound a clear call, who will get ready for battle?
1COR|14|9|So it is with you. Unless you speak intelligible words with your tongue, how will anyone know what you are saying? You will just be speaking into the air.
1COR|14|10|Undoubtedly there are all sorts of languages in the world, yet none of them is without meaning.
1COR|14|11|If then I do not grasp the meaning of what someone is saying, I am a foreigner to the speaker, and he is a foreigner to me.
1COR|14|12|So it is with you. Since you are eager to have spiritual gifts, try to excel in gifts that build up the church.
1COR|14|13|For this reason anyone who speaks in a tongue should pray that he may interpret what he says.
1COR|14|14|For if I pray in a tongue, my spirit prays, but my mind is unfruitful.
1COR|14|15|So what shall I do? I will pray with my spirit, but I will also pray with my mind; I will sing with my spirit, but I will also sing with my mind.
1COR|14|16|If you are praising God with your spirit, how can one who finds himself among those who do not understand say "Amen" to your thanksgiving, since he does not know what you are saying?
1COR|14|17|You may be giving thanks well enough, but the other man is not edified.
1COR|14|18|I thank God that I speak in tongues more than all of you.
1COR|14|19|But in the church I would rather speak five intelligible words to instruct others than ten thousand words in a tongue.
1COR|14|20|Brothers, stop thinking like children. In regard to evil be infants, but in your thinking be adults.
1COR|14|21|In the Law it is written: "Through men of strange tongues and through the lips of foreigners I will speak to this people, but even then they will not listen to me," says the Lord.
1COR|14|22|Tongues, then, are a sign, not for believers but for unbelievers; prophecy, however, is for believers, not for unbelievers.
1COR|14|23|So if the whole church comes together and everyone speaks in tongues, and some who do not understand or some unbelievers come in, will they not say that you are out of your mind?
1COR|14|24|But if an unbeliever or someone who does not understand comes in while everybody is prophesying, he will be convinced by all that he is a sinner and will be judged by all,
1COR|14|25|and the secrets of his heart will be laid bare. So he will fall down and worship God, exclaiming, "God is really among you!"
1COR|14|26|What then shall we say, brothers? When you come together, everyone has a hymn, or a word of instruction, a revelation, a tongue or an interpretation. All of these must be done for the strengthening of the church.
1COR|14|27|If anyone speaks in a tongue, two--or at the most three--should speak, one at a time, and someone must interpret.
1COR|14|28|If there is no interpreter, the speaker should keep quiet in the church and speak to himself and God.
1COR|14|29|Two or three prophets should speak, and the others should weigh carefully what is said.
1COR|14|30|And if a revelation comes to someone who is sitting down, the first speaker should stop.
1COR|14|31|For you can all prophesy in turn so that everyone may be instructed and encouraged.
1COR|14|32|The spirits of prophets are subject to the control of prophets.
1COR|14|33|For God is not a God of disorder but of peace.
1COR|14|34|As in all the congregations of the saints, women should remain silent in the churches. They are not allowed to speak, but must be in submission, as the Law says.
1COR|14|35|If they want to inquire about something, they should ask their own husbands at home; for it is disgraceful for a woman to speak in the church.
1COR|14|36|Did the word of God originate with you? Or are you the only people it has reached?
1COR|14|37|If anybody thinks he is a prophet or spiritually gifted, let him acknowledge that what I am writing to you is the Lord's command.
1COR|14|38|If he ignores this, he himself will be ignored.
1COR|14|39|Therefore, my brothers, be eager to prophesy, and do not forbid speaking in tongues.
1COR|14|40|But everything should be done in a fitting and orderly way.
1COR|15|1|Now, brothers, I want to remind you of the gospel I preached to you, which you received and on which you have taken your stand.
1COR|15|2|By this gospel you are saved, if you hold firmly to the word I preached to you. Otherwise, you have believed in vain.
1COR|15|3|For what I received I passed on to you as of first importance: that Christ died for our sins according to the Scriptures,
1COR|15|4|that he was buried, that he was raised on the third day according to the Scriptures,
1COR|15|5|and that he appeared to Peter, and then to the Twelve.
1COR|15|6|After that, he appeared to more than five hundred of the brothers at the same time, most of whom are still living, though some have fallen asleep.
1COR|15|7|Then he appeared to James, then to all the apostles,
1COR|15|8|and last of all he appeared to me also, as to one abnormally born.
1COR|15|9|For I am the least of the apostles and do not even deserve to be called an apostle, because I persecuted the church of God.
1COR|15|10|But by the grace of God I am what I am, and his grace to me was not without effect. No, I worked harder than all of them--yet not I, but the grace of God that was with me.
1COR|15|11|Whether, then, it was I or they, this is what we preach, and this is what you believed.
1COR|15|12|But if it is preached that Christ has been raised from the dead, how can some of you say that there is no resurrection of the dead?
1COR|15|13|If there is no resurrection of the dead, then not even Christ has been raised.
1COR|15|14|And if Christ has not been raised, our preaching is useless and so is your faith.
1COR|15|15|More than that, we are then found to be false witnesses about God, for we have testified about God that he raised Christ from the dead. But he did not raise him if in fact the dead are not raised.
1COR|15|16|For if the dead are not raised, then Christ has not been raised either.
1COR|15|17|And if Christ has not been raised, your faith is futile; you are still in your sins.
1COR|15|18|Then those also who have fallen asleep in Christ are lost.
1COR|15|19|If only for this life we have hope in Christ, we are to be pitied more than all men.
1COR|15|20|But Christ has indeed been raised from the dead, the firstfruits of those who have fallen asleep.
1COR|15|21|For since death came through a man, the resurrection of the dead comes also through a man.
1COR|15|22|For as in Adam all die, so in Christ all will be made alive.
1COR|15|23|But each in his own turn: Christ, the firstfruits; then, when he comes, those who belong to him.
1COR|15|24|Then the end will come, when he hands over the kingdom to God the Father after he has destroyed all dominion, authority and power.
1COR|15|25|For he must reign until he has put all his enemies under his feet.
1COR|15|26|The last enemy to be destroyed is death.
1COR|15|27|For he "has put everything under his feet." Now when it says that "everything" has been put under him, it is clear that this does not include God himself, who put everything under Christ.
1COR|15|28|When he has done this, then the Son himself will be made subject to him who put everything under him, so that God may be all in all.
1COR|15|29|Now if there is no resurrection, what will those do who are baptized for the dead? If the dead are not raised at all, why are people baptized for them?
1COR|15|30|And as for us, why do we endanger ourselves every hour?
1COR|15|31|I die every day--I mean that, brothers--just as surely as I glory over you in Christ Jesus our Lord.
1COR|15|32|If I fought wild beasts in Ephesus for merely human reasons, what have I gained? If the dead are not raised, "Let us eat and drink, for tomorrow we die."
1COR|15|33|Do not be misled: "Bad company corrupts good character."
1COR|15|34|Come back to your senses as you ought, and stop sinning; for there are some who are ignorant of God--I say this to your shame.
1COR|15|35|But someone may ask, "How are the dead raised? With what kind of body will they come?"
1COR|15|36|How foolish! What you sow does not come to life unless it dies.
1COR|15|37|When you sow, you do not plant the body that will be, but just a seed, perhaps of wheat or of something else.
1COR|15|38|But God gives it a body as he has determined, and to each kind of seed he gives its own body.
1COR|15|39|All flesh is not the same: Men have one kind of flesh, animals have another, birds another and fish another.
1COR|15|40|There are also heavenly bodies and there are earthly bodies; but the splendor of the heavenly bodies is one kind, and the splendor of the earthly bodies is another.
1COR|15|41|The sun has one kind of splendor, the moon another and the stars another; and star differs from star in splendor.
1COR|15|42|So will it be with the resurrection of the dead. The body that is sown is perishable, it is raised imperishable;
1COR|15|43|it is sown in dishonor, it is raised in glory; it is sown in weakness, it is raised in power;
1COR|15|44|it is sown a natural body, it is raised a spiritual body. If there is a natural body, there is also a spiritual body.
1COR|15|45|So it is written: "The first man Adam became a living being"; the last Adam, a lifegiving spirit.
1COR|15|46|The spiritual did not come first, but the natural, and after that the spiritual.
1COR|15|47|The first man was of the dust of the earth, the second man from heaven.
1COR|15|48|As was the earthly man, so are those who are of the earth; and as is the man from heaven, so also are those who are of heaven.
1COR|15|49|And just as we have borne the likeness of the earthly man, so shall we bear the likeness of the man from heaven.
1COR|15|50|I declare to you, brothers, that flesh and blood cannot inherit the kingdom of God, nor does the perishable inherit the imperishable.
1COR|15|51|Listen, I tell you a mystery: We will not all sleep, but we will all be changed--
1COR|15|52|in a flash, in the twinkling of an eye, at the last trumpet. For the trumpet will sound, the dead will be raised imperishable, and we will be changed.
1COR|15|53|For the perishable must clothe itself with the imperishable, and the mortal with immortality.
1COR|15|54|When the perishable has been clothed with the imperishable, and the mortal with immortality, then the saying that is written will come true: "Death has been swallowed up in victory."
1COR|15|55|"Where, O death, is your victory? Where, O death, is your sting?"
1COR|15|56|The sting of death is sin, and the power of sin is the law.
1COR|15|57|But thanks be to God! He gives us the victory through our Lord Jesus Christ.
1COR|15|58|Therefore, my dear brothers, stand firm. Let nothing move you. Always give yourselves fully to the work of the Lord, because you know that your labor in the Lord is not in vain.
1COR|16|1|Now about the collection for God's people: Do what I told the Galatian churches to do.
1COR|16|2|On the first day of every week, each one of you should set aside a sum of money in keeping with his income, saving it up, so that when I come no collections will have to be made.
1COR|16|3|Then, when I arrive, I will give letters of introduction to the men you approve and send them with your gift to Jerusalem.
1COR|16|4|If it seems advisable for me to go also, they will accompany me.
1COR|16|5|After I go through Macedonia, I will come to you--for I will be going through Macedonia.
1COR|16|6|Perhaps I will stay with you awhile, or even spend the winter, so that you can help me on my journey, wherever I go.
1COR|16|7|I do not want to see you now and make only a passing visit; I hope to spend some time with you, if the Lord permits.
1COR|16|8|But I will stay on at Ephesus until Pentecost,
1COR|16|9|because a great door for effective work has opened to me, and there are many who oppose me.
1COR|16|10|If Timothy comes, see to it that he has nothing to fear while he is with you, for he is carrying on the work of the Lord, just as I am.
1COR|16|11|No one, then, should refuse to accept him. Send him on his way in peace so that he may return to me. I am expecting him along with the brothers.
1COR|16|12|Now about our brother Apollos: I strongly urged him to go to you with the brothers. He was quite unwilling to go now, but he will go when he has the opportunity.
1COR|16|13|Be on your guard; stand firm in the faith; be men of courage; be strong.
1COR|16|14|Do everything in love.
1COR|16|15|You know that the household of Stephanas were the first converts in Achaia, and they have devoted themselves to the service of the saints. I urge you, brothers,
1COR|16|16|to submit to such as these and to everyone who joins in the work, and labors at it.
1COR|16|17|I was glad when Stephanas, Fortunatus and Achaicus arrived, because they have supplied what was lacking from you.
1COR|16|18|For they refreshed my spirit and yours also. Such men deserve recognition.
1COR|16|19|The churches in the province of Asia send you greetings. Aquila and Priscilla greet you warmly in the Lord, and so does the church that meets at their house.
1COR|16|20|All the brothers here send you greetings. Greet one another with a holy kiss.
1COR|16|21|I, Paul, write this greeting in my own hand.
1COR|16|22|If anyone does not love the Lord--a curse be on him. Come, O Lord!
1COR|16|23|The grace of the Lord Jesus be with you.
1COR|16|24|My love to all of you in Christ Jesus. Amen.
