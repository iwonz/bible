JAS|1|1|上帝和主耶稣基督的仆人 雅各 问候散居在各处的十二个支派的人。
JAS|1|2|我的弟兄们，你们遭受各种试炼时，都要认为是大喜乐，
JAS|1|3|因为知道你们的信心经过考验，就生忍耐。
JAS|1|4|但要让忍耐发挥完全的功用，使你们能又完全又完整，一无所缺。
JAS|1|5|你们中间若有缺少智慧的，该求那厚赐与众人又不斥责人的上帝，上帝必赐给他。
JAS|1|6|只要凭着信心求，一点也不疑惑；因为那疑惑的人，就像海中的波浪被风吹动翻腾。
JAS|1|7|这样的人不要想从主那里得到什么。
JAS|1|8|三心二意的人，在他一切所行的路上都摇摆不定。
JAS|1|9|卑微的弟兄要因高升而夸耀，
JAS|1|10|富足的却要因被降卑而夸耀，因为富足的人要消逝，如同草上的花一样。
JAS|1|11|太阳出来，热风刮起，草就枯干，花也凋谢，它美丽的样子就消失了；那富足的人在他一生的奔波中也要这样衰残。
JAS|1|12|忍受试炼的人有福了，因为他经过考验以后必得生命的冠冕，这是主应许给爱他之人的。
JAS|1|13|人被诱惑，不可说：“我是被上帝诱惑”；因为上帝是不被恶诱惑的，他也不诱惑人。
JAS|1|14|但每一个人被诱惑是因自己的私欲牵引而被诱惑的。
JAS|1|15|私欲既怀了胎，就生出罪来；罪既长成，就生出死来。
JAS|1|16|我亲爱的弟兄们，不要被欺骗了。
JAS|1|17|各样美善的恩泽和各样完美的赏赐都是从上头来的，从众光之父那里降下来的；在他并没有改变，也没有转动的影儿。
JAS|1|18|他按自己的旨意，用真理的道生了我们，使我们在他所造的万物中成为初熟的果子。
JAS|1|19|我亲爱的弟兄们，你们要明白：你们每一个人要快快地听，慢慢地说，慢慢地动怒，
JAS|1|20|因为人的怒气并不能实现上帝的义。
JAS|1|21|所以，你们要除去一切的污秽和累积的恶毒，要存温柔的心领受所栽种的道，就是能救你们灵魂的道。
JAS|1|22|但是，你们要作行道的人，不要只作听道的人，自己欺骗自己。
JAS|1|23|因为只听道而不行道的，就像人对着镜子观看自己本来的面目，
JAS|1|24|注视后，就离开，立刻忘了自己的相貌如何。
JAS|1|25|惟有查看那完美、使人自由的律法，并且时常遵守的，他不是听了就忘，而是切实行出来，这样的人在所行的事上必然蒙福。
JAS|1|26|若有人自以为虔诚，却不勒住自己的舌头，反欺骗自己的心，这人的虔诚是徒然的。
JAS|1|27|在上帝—我们的父面前，清洁没有玷污的虔诚就是看顾在患难中的孤儿寡妇，并且保守自己不沾染世俗。
JAS|2|1|我的弟兄们，你们信奉我们荣耀的主耶稣基督，就不可按着外貌待人。
JAS|2|2|若有一个人戴着金戒指，穿着华丽的衣服，进入你们的会堂，又有一个穷人穿着肮脏的衣服也进去，
JAS|2|3|而你们只看重那穿华丽衣服的人，说：“请坐在这里”，又对那穷人说：“你站在那里”，或“坐在我脚凳旁”；
JAS|2|4|这岂不是你们偏心待人，用恶意评断人吗？
JAS|2|5|我亲爱的弟兄们，请听，上帝岂不是拣选了世上的贫穷人，使他们在信心上富足，并承受他所应许给那些爱他之人的国吗？
JAS|2|6|你们却羞辱贫穷的人。欺压你们，拉你们到公堂去的，不就是这些富有的人吗？
JAS|2|7|毁谤为你们求告时所奉的尊名的，不就是他们吗？
JAS|2|8|经上记着：“要爱邻 如己”，你们若切实守这至尊的律法，你们就做得很好。
JAS|2|9|但你们若按外貌待人就是犯罪，是被律法定为犯法的。
JAS|2|10|因为凡遵守全部律法的，只违背了一条就是违犯了所有的律法。
JAS|2|11|原来那说“不可奸淫”的，也说“不可杀人”。你就是不奸淫，却杀人，也是成为违犯律法的。
JAS|2|12|既然你们要按使人自由的律法受审判，就要照这律法说话行事。
JAS|2|13|因为对那不怜悯人的，他们要受没有怜悯的审判；怜悯胜过审判。
JAS|2|14|我的弟兄们，若有人说自己有信心，却没有行为，有什么益处呢？这信心能救他吗？
JAS|2|15|若是弟兄或是姊妹没有衣服穿，又缺少日用的饮食；
JAS|2|16|你们中间有人对他们说：“平平安安地去吧！愿你们穿得暖，吃得饱”，却不给他们身体所需要的，这有什么益处呢？
JAS|2|17|信心也是这样，若没有行为是死的。
JAS|2|18|但是有人会说：“你有信心，我有行为。”把你没有行为的信心给我看，我就藉着我的行为把我的信心给你看。
JAS|2|19|你信上帝只有一位，你信得很好；连鬼魔也信，且怕得发抖。
JAS|2|20|你这虚浮的人哪，你愿意知道没有行为的信心是没有用的吗？
JAS|2|21|我们的祖宗 亚伯拉罕 把他儿子 以撒 献在坛上，岂不是因行为得称义吗？
JAS|2|22|可见信心是与他的行为相辅并行，而且信心是因着行为才得以成全的。
JAS|2|23|这正应验了经上所说：“ 亚伯拉罕 信了上帝，这就算他为义”；他又得称为上帝的朋友。
JAS|2|24|这样看来，人称义是因着行为，不是单因着信。
JAS|2|25|同样，妓女 喇合 接待使者，又放他们从另一条路出去，不也是因行为称义吗？
JAS|2|26|所以，就如身体没有灵魂是死的，信心没有行为也是死的。
JAS|3|1|我的弟兄们，不要许多人做教师，因为你们知道，我们做教师的要接受更严厉的审判。
JAS|3|2|原来我们在许多事上都有过失；若有人在言语上没有过失，他就是完全的人，也能勒住自己的全身。
JAS|3|3|我们若把嚼环放在马嘴里使它们驯服，就能控制它们的全身。
JAS|3|4|再看船只，虽然甚大，又被强风猛吹，只用小小的舵就随着掌舵的意思转动。
JAS|3|5|同样，舌头是小肢体，却能说大话。 看哪，最小的火能点燃最大的树林。
JAS|3|6|舌头就是火。在我们百体中，舌头是个不义的世界，能玷污全身，也能烧毁生命的轮子，而且是被地狱的火点燃的。
JAS|3|7|各类的走兽、飞禽、爬虫、水族，本来都可以制伏，也已经被人制伏了；
JAS|3|8|惟独舌头没有人能制伏，是永不静止的邪恶，充满了害死人的毒气。
JAS|3|9|我们用舌头颂赞我们的主—我们的天父，又用舌头诅咒照着上帝形像被造的人。
JAS|3|10|颂赞和诅咒从同一个口出来。我的弟兄们，这是不应该的。
JAS|3|11|泉源能从一个出口发出甜苦两样的水吗？
JAS|3|12|我的弟兄们，无花果树能生橄榄吗？葡萄树能结无花果吗？咸水也不能流出甜水来。
JAS|3|13|你们中间谁是有智慧有见识的呢？他就当在智慧的温柔上显出他的善行来。
JAS|3|14|你们心里若怀着恶毒的嫉妒和自私，就不可自夸，不可说谎话抵挡真理。
JAS|3|15|这样的智慧不是从上头下来的，而是属地上的，属情欲的，属鬼魔的。
JAS|3|16|在何处有嫉妒、自私，在何处就有动乱和各样的坏事。
JAS|3|17|惟独从上头来的智慧，先是清洁，后是和平、温良、柔顺，满有怜悯和美善的果子，没有偏私，没有虚伪。
JAS|3|18|正义的果实是为促进和平的人用和平栽种出来的。
JAS|4|1|你们中间的冲突是哪里来的？争执是哪里来的？不是从你们肢体中交战着的私欲来的吗？
JAS|4|2|你们贪恋，得不着就杀人；你们嫉妒，不能得手就起争执和冲突；你们得不着，是因为你们不求。
JAS|4|3|你们求也得不着，是因为你们妄求，为了要浪费在你们的宴乐中。
JAS|4|4|你们这些淫乱的人哪，岂不知道与世俗为友就是与上帝为敌吗？所以，凡想要与世俗为友的，就是与上帝为敌了。
JAS|4|5|经上说：“上帝爱安置在我们里面的灵，爱到嫉妒的地步。” 你们以为这话是徒然的吗？
JAS|4|6|但是他赐更多的恩典，正如经上说： “上帝抵挡骄傲的人， 但赐恩给谦卑的人。”
JAS|4|7|所以，要顺服上帝。要抵挡魔鬼，魔鬼就必逃避你们；
JAS|4|8|要亲近上帝，上帝就必亲近你们。有罪的人哪，要洁净你们的手！心怀二意的人哪，要清洁你们的心！
JAS|4|9|你们要愁苦，悲哀，哭泣；要将欢笑变为悲哀，欢乐变为愁闷。
JAS|4|10|要在主面前谦卑，他就使你们高升。
JAS|4|11|弟兄们，不可彼此诋毁。诋毁弟兄或评断弟兄的人，就是诋毁律法，评断律法；你若评断律法，就不是遵行律法，而是评断者了。
JAS|4|12|立法者和审判者只有一位；他就是那能拯救人也能毁灭人的。你是谁，竟敢评断你的邻舍！
JAS|4|13|注意！有人说：“今天或明天我们要往某城去，在那里住一年，做买卖赚钱。”
JAS|4|14|其实明天如何，你们还不知道。你们的生命是什么呢？你们 原来是一片云雾，出现片刻就不见了。
JAS|4|15|你们倒应当说：“主若愿意，我们就能活着，也可以做这事或那事。”
JAS|4|16|现今你们竟然狂傲自夸；凡这样的自夸都是邪恶的。
JAS|4|17|所以，人若知道该行善而不去行，这就是他的罪了。
JAS|5|1|注意！你们这些富足人哪，要为将要临到你们身上的灾难哭泣、号啕。
JAS|5|2|你们的财物腐烂了，你们的衣服被虫子蛀了。
JAS|5|3|你们的金银都生锈了；这锈要证明你们的不是，又要像火一样吞吃你们的肉。你们在这末世只知道积蓄钱财。
JAS|5|4|工人给你们收割庄稼，你们克扣他们的工钱；这工钱在喊冤，而且收割工人的冤声已经进入万军之主的耳朵了。
JAS|5|5|你们在地上享奢华宴乐，把自己养肥了，等候宰杀的日子。
JAS|5|6|你们定了义人的罪，把他杀害，他没有抵抗你们。
JAS|5|7|所以弟兄们，你们要忍耐，直到主来。看哪，农夫等候着地里宝贵的出产，耐心地等到它得了秋霖春雨。
JAS|5|8|你们也要忍耐，坚固你们的心，因为主来的日子近了。
JAS|5|9|弟兄们，你们不要彼此埋怨，免得受审判。看哪，审判的主站在门口了。
JAS|5|10|弟兄们，你们要把那先前奉主名说话的众先知作能受苦、能忍耐的榜样。
JAS|5|11|看哪，那些忍耐的人，我们称他们是有福的。你们听见过 约伯 的忍耐，也看见主给他的结局，知道主是充满怜悯和慈悲的。
JAS|5|12|我的弟兄们，最要紧的是不可起誓；不可指着天起誓，也不可指着地起誓，任何誓都不可起。你们说话，是，就说是；不是，就说不是，免得你们落在审判之下。
JAS|5|13|你们中间若有人受苦，他该祷告；有人喜乐，他该歌颂。
JAS|5|14|你们中间若有人病了，他该请教会的长老们来为他祷告，奉主的名为他抹油。
JAS|5|15|出于信心的祈祷必能救那病人，主必叫他起来；他若犯了罪，也必蒙赦免。
JAS|5|16|所以，你们要彼此认罪，互相代求，使你们得医治。义人祈祷所发的力量是大有功效的。
JAS|5|17|以利亚 与我们是同样性情的人，他恳切地祈求不要下雨，地上就三年六个月没有下雨。
JAS|5|18|他又祷告，天就降下雨来，地就有了出产。
JAS|5|19|我的弟兄们，你们中间若有人迷失了真理而有人使他回转，
JAS|5|20|这人该知道，使一个罪人从迷途中回转，会从死亡中把他的灵魂救回来，而且遮盖许多的罪。
