EPH|1|1|Павел, волею Божиею Апостол Иисуса Христа, находящимся в Ефесе святым и верным во Христе Иисусе:
EPH|1|2|благодать вам и мир от Бога Отца нашего и Господа Иисуса Христа.
EPH|1|3|Благословен Бог и Отец Господа нашего Иисуса Христа, благословивший нас во Христе всяким духовным благословением в небесах,
EPH|1|4|так как Он избрал нас в Нем прежде создания мира, чтобы мы были святы и непорочны пред Ним в любви,
EPH|1|5|предопределив усыновить нас Себе чрез Иисуса Христа, по благоволению воли Своей,
EPH|1|6|в похвалу славы благодати Своей, которою Он облагодатствовал нас в Возлюбленном,
EPH|1|7|в Котором мы имеем искупление Кровию Его, прощение грехов, по богатству благодати Его,
EPH|1|8|каковую Он в преизбытке даровал нам во всякой премудрости и разумении,
EPH|1|9|открыв нам тайну Своей воли по Своему благоволению, которое Он прежде положил в Нем,
EPH|1|10|в устроении полноты времен, дабы все небесное и земное соединить под главою Христом.
EPH|1|11|В Нем мы и сделались наследниками, быв предназначены [к тому] по определению Совершающего все по изволению воли Своей,
EPH|1|12|дабы послужить к похвале славы Его нам, которые ранее уповали на Христа.
EPH|1|13|В Нем и вы, услышав слово истины, благовествование вашего спасения, и уверовав в Него, запечатлены обетованным Святым Духом,
EPH|1|14|Который есть залог наследия нашего, для искупления удела [Его], в похвалу славы Его.
EPH|1|15|Посему и я, услышав о вашей вере во Христа Иисуса и о любви ко всем святым,
EPH|1|16|непрестанно благодарю за вас [Бога], вспоминая о вас в молитвах моих,
EPH|1|17|чтобы Бог Господа нашего Иисуса Христа, Отец славы, дал вам Духа премудрости и откровения к познанию Его,
EPH|1|18|и просветил очи сердца вашего, дабы вы познали, в чем состоит надежда призвания Его, и какое богатство славного наследия Его для святых,
EPH|1|19|и как безмерно величие могущества Его в нас, верующих по действию державной силы Его,
EPH|1|20|которою Он воздействовал во Христе, воскресив Его из мертвых и посадив одесную Себя на небесах,
EPH|1|21|превыше всякого Начальства, и Власти, и Силы, и Господства, и всякого имени, именуемого не только в сем веке, но и в будущем,
EPH|1|22|и все покорил под ноги Его, и поставил Его выше всего, главою Церкви,
EPH|1|23|которая есть Тело Его, полнота Наполняющего все во всем.
EPH|2|1|И вас, мертвых по преступлениям и грехам вашим,
EPH|2|2|в которых вы некогда жили, по обычаю мира сего, по [воле] князя, господствующего в воздухе, духа, действующего ныне в сынах противления,
EPH|2|3|между которыми и мы все жили некогда по нашим плотским похотям, исполняя желания плоти и помыслов, и были по природе чадами гнева, как и прочие,
EPH|2|4|Бог, богатый милостью, по Своей великой любви, которою возлюбил нас,
EPH|2|5|и нас, мертвых по преступлениям, оживотворил со Христом, – благодатью вы спасены, –
EPH|2|6|и воскресил с Ним, и посадил на небесах во Христе Иисусе,
EPH|2|7|дабы явить в грядущих веках преизобильное богатство благодати Своей в благости к нам во Христе Иисусе.
EPH|2|8|Ибо благодатью вы спасены через веру, и сие не от вас, Божий дар:
EPH|2|9|не от дел, чтобы никто не хвалился.
EPH|2|10|Ибо мы – Его творение, созданы во Христе Иисусе на добрые дела, которые Бог предназначил нам исполнять.
EPH|2|11|Итак помните, что вы, некогда язычники по плоти, которых называли необрезанными так называемые обрезанные плотским [обрезанием], совершаемым руками,
EPH|2|12|что вы были в то время без Христа, отчуждены от общества Израильского, чужды заветов обетования, не имели надежды и были безбожники в мире.
EPH|2|13|А теперь во Христе Иисусе вы, бывшие некогда далеко, стали близки Кровию Христовою.
EPH|2|14|Ибо Он есть мир наш, соделавший из обоих одно и разрушивший стоявшую посреди преграду,
EPH|2|15|упразднив вражду Плотию Своею, а закон заповедей учением, дабы из двух создать в Себе Самом одного нового человека, устрояя мир,
EPH|2|16|и в одном теле примирить обоих с Богом посредством креста, убив вражду на нем.
EPH|2|17|И, придя, благовествовал мир вам, дальним и близким,
EPH|2|18|потому что через Него и те и другие имеем доступ к Отцу, в одном Духе.
EPH|2|19|Итак вы уже не чужие и не пришельцы, но сограждане святым и свои Богу,
EPH|2|20|быв утверждены на основании Апостолов и пророков, имея Самого Иисуса Христа краеугольным [камнем],
EPH|2|21|на котором все здание, слагаясь стройно, возрастает в святый храм в Господе,
EPH|2|22|на котором и вы устрояетесь в жилище Божие Духом.
EPH|3|1|Для сего–то я, Павел, [сделался] узником Иисуса Христа за вас язычников.
EPH|3|2|Как вы слышали о домостроительстве благодати Божией, данной мне для вас,
EPH|3|3|потому что мне через откровение возвещена тайна (о чем я и выше писал кратко),
EPH|3|4|то вы, читая, можете усмотреть мое разумение тайны Христовой,
EPH|3|5|которая не была возвещена прежним поколениям сынов человеческих, как ныне открыта святым Апостолам Его и пророкам Духом Святым,
EPH|3|6|чтобы и язычникам быть сонаследниками, составляющими одно тело, и сопричастниками обетования Его во Христе Иисусе посредством благовествования,
EPH|3|7|которого служителем сделался я по дару благодати Божией, данной мне действием силы Его.
EPH|3|8|Мне, наименьшему из всех святых, дана благодать сия – благовествовать язычникам неисследимое богатство Христово
EPH|3|9|и открыть всем, в чем состоит домостроительство тайны, сокрывавшейся от вечности в Боге, создавшем все Иисусом Христом,
EPH|3|10|дабы ныне соделалась известною через Церковь начальствам и властям на небесах многоразличная премудрость Божия,
EPH|3|11|по предвечному определению, которое Он исполнил во Христе Иисусе, Господе нашем,
EPH|3|12|в Котором мы имеем дерзновение и надежный доступ через веру в Него.
EPH|3|13|Посему прошу вас не унывать при моих ради вас скорбях, которые суть ваша слава.
EPH|3|14|Для сего преклоняю колени мои пред Отцем Господа нашего Иисуса Христа,
EPH|3|15|от Которого именуется всякое отечество на небесах и на земле,
EPH|3|16|да даст вам, по богатству славы Своей, крепко утвердиться Духом Его во внутреннем человеке,
EPH|3|17|верою вселиться Христу в сердца ваши,
EPH|3|18|чтобы вы, укорененные и утвержденные в любви, могли постигнуть со всеми святыми, что широта и долгота, и глубина и высота,
EPH|3|19|и уразуметь превосходящую разумение любовь Христову, дабы вам исполниться всею полнотою Божиею.
EPH|3|20|А Тому, Кто действующею в нас силою может сделать несравненно больше всего, чего мы просим, или о чем помышляем,
EPH|3|21|Тому слава в Церкви во Христе Иисусе во все роды, от века до века. Аминь.
EPH|4|1|Итак я, узник в Господе, умоляю вас поступать достойно звания, в которое вы призваны,
EPH|4|2|со всяким смиренномудрием и кротостью и долготерпением, снисходя друг ко другу любовью,
EPH|4|3|стараясь сохранять единство духа в союзе мира.
EPH|4|4|Одно тело и один дух, как вы и призваны к одной надежде вашего звания;
EPH|4|5|один Господь, одна вера, одно крещение,
EPH|4|6|один Бог и Отец всех, Который над всеми, и через всех, и во всех нас.
EPH|4|7|Каждому же из нас дана благодать по мере дара Христова.
EPH|4|8|Посему и сказано: восшед на высоту, пленил плен и дал дары человекам.
EPH|4|9|А "восшел" что означает, как не то, что Он и нисходил прежде в преисподние места земли?
EPH|4|10|Нисшедший, Он же есть и восшедший превыше всех небес, дабы наполнить все.
EPH|4|11|И Он поставил одних Апостолами, других пророками, иных Евангелистами, иных пастырями и учителями,
EPH|4|12|к совершению святых, на дело служения, для созидания Тела Христова,
EPH|4|13|доколе все придем в единство веры и познания Сына Божия, в мужа совершенного, в меру полного возраста Христова;
EPH|4|14|дабы мы не были более младенцами, колеблющимися и увлекающимися всяким ветром учения, по лукавству человеков, по хитрому искусству обольщения,
EPH|4|15|но истинною любовью все возращали в Того, Который есть глава Христос,
EPH|4|16|из Которого все тело, составляемое и совокупляемое посредством всяких взаимно скрепляющих связей, при действии в свою меру каждого члена, получает приращение для созидания самого себя в любви.
EPH|4|17|Посему я говорю и заклинаю Господом, чтобы вы более не поступали, как поступают прочие народы, по суетности ума своего,
EPH|4|18|будучи помрачены в разуме, отчуждены от жизни Божией, по причине их невежества и ожесточения сердца их.
EPH|4|19|Они, дойдя до бесчувствия, предались распутству так, что делают всякую нечистоту с ненасытимостью.
EPH|4|20|Но вы не так познали Христа;
EPH|4|21|потому что вы слышали о Нем и в Нем научились, – так как истина во Иисусе, –
EPH|4|22|отложить прежний образ жизни ветхого человека, истлевающего в обольстительных похотях,
EPH|4|23|а обновиться духом ума вашего
EPH|4|24|и облечься в нового человека, созданного по Богу, в праведности и святости истины.
EPH|4|25|Посему, отвергнув ложь, говорите истину каждый ближнему своему, потому что мы члены друг другу.
EPH|4|26|Гневаясь, не согрешайте: солнце да не зайдет во гневе вашем;
EPH|4|27|и не давайте места диаволу.
EPH|4|28|Кто крал, вперед не кради, а лучше трудись, делая своими руками полезное, чтобы было из чего уделять нуждающемуся.
EPH|4|29|Никакое гнилое слово да не исходит из уст ваших, а только доброе для назидания в вере, дабы оно доставляло благодать слушающим.
EPH|4|30|И не оскорбляйте Святаго Духа Божия, Которым вы запечатлены в день искупления.
EPH|4|31|Всякое раздражение и ярость, и гнев, и крик, и злоречие со всякою злобою да будут удалены от вас;
EPH|4|32|но будьте друг ко другу добры, сострадательны, прощайте друг друга, как и Бог во Христе простил вас.
EPH|5|1|Итак, подражайте Богу, как чада возлюбленные,
EPH|5|2|и живите в любви, как и Христос возлюбил нас и предал Себя за нас в приношение и жертву Богу, в благоухание приятное.
EPH|5|3|А блуд и всякая нечистота и любостяжание не должны даже именоваться у вас, как прилично святым.
EPH|5|4|Также сквернословие и пустословие и смехотворство не приличны [вам], а, напротив, благодарение;
EPH|5|5|ибо знайте, что никакой блудник, или нечистый, или любостяжатель, который есть идолослужитель, не имеет наследия в Царстве Христа и Бога.
EPH|5|6|Никто да не обольщает вас пустыми словами, ибо за это приходит гнев Божий на сынов противления;
EPH|5|7|итак, не будьте сообщниками их.
EPH|5|8|Вы были некогда тьма, а теперь – свет в Господе: поступайте, как чада света,
EPH|5|9|потому что плод Духа состоит во всякой благости, праведности и истине.
EPH|5|10|Испытывайте, что благоугодно Богу,
EPH|5|11|и не участвуйте в бесплодных делах тьмы, но и обличайте.
EPH|5|12|Ибо о том, что они делают тайно, стыдно и говорить.
EPH|5|13|Все же обнаруживаемое делается явным от света, ибо все, делающееся явным, свет есть.
EPH|5|14|Посему сказано: "встань, спящий, и воскресни из мертвых, и осветит тебя Христос".
EPH|5|15|Итак, смотрите, поступайте осторожно, не как неразумные, но как мудрые,
EPH|5|16|дорожа временем, потому что дни лукавы.
EPH|5|17|Итак, не будьте нерассудительны, но познавайте, что есть воля Божия.
EPH|5|18|И не упивайтесь вином, от которого бывает распутство; но исполняйтесь Духом,
EPH|5|19|назидая самих себя псалмами и славословиями и песнопениями духовными, поя и воспевая в сердцах ваших Господу,
EPH|5|20|благодаря всегда за все Бога и Отца, во имя Господа нашего Иисуса Христа,
EPH|5|21|повинуясь друг другу в страхе Божием.
EPH|5|22|Жены, повинуйтесь своим мужьям, как Господу,
EPH|5|23|потому что муж есть глава жены, как и Христос глава Церкви, и Он же Спаситель тела.
EPH|5|24|Но как Церковь повинуется Христу, так и жены своим мужьям во всем.
EPH|5|25|Мужья, любите своих жен, как и Христос возлюбил Церковь и предал Себя за нее,
EPH|5|26|чтобы освятить ее, очистив банею водною посредством слова;
EPH|5|27|чтобы представить ее Себе славною Церковью, не имеющею пятна, или порока, или чего–либо подобного, но дабы она была свята и непорочна.
EPH|5|28|Так должны мужья любить своих жен, как свои тела: любящий свою жену любит самого себя.
EPH|5|29|Ибо никто никогда не имел ненависти к своей плоти, но питает и греет ее, как и Господь Церковь,
EPH|5|30|потому что мы члены тела Его, от плоти Его и от костей Его.
EPH|5|31|Посему оставит человек отца своего и мать и прилепится к жене своей, и будут двое одна плоть.
EPH|5|32|Тайна сия велика; я говорю по отношению ко Христу и к Церкви.
EPH|5|33|Так каждый из вас да любит свою жену, как самого себя; а жена да боится своего мужа.
EPH|6|1|Дети, повинуйтесь своим родителям в Господе, ибо сего [требует] справедливость.
EPH|6|2|Почитай отца твоего и мать, это первая заповедь с обетованием:
EPH|6|3|да будет тебе благо, и будешь долголетен на земле.
EPH|6|4|И вы, отцы, не раздражайте детей ваших, но воспитывайте их в учении и наставлении Господнем.
EPH|6|5|Рабы, повинуйтесь господам своим по плоти со страхом и трепетом, в простоте сердца вашего, как Христу,
EPH|6|6|не с видимою только услужливостью, как человекоугодники, но как рабы Христовы, исполняя волю Божию от души,
EPH|6|7|служа с усердием, как Господу, а не как человекам,
EPH|6|8|зная, что каждый получит от Господа по мере добра, которое он сделал, раб ли, или свободный.
EPH|6|9|И вы, господа, поступайте с ними так же, умеряя строгость, зная, что и над вами самими и над ними есть на небесах Господь, у Которого нет лицеприятия.
EPH|6|10|Наконец, братия мои, укрепляйтесь Господом и могуществом силы Его.
EPH|6|11|Облекитесь во всеоружие Божие, чтобы вам можно было стать против козней диавольских,
EPH|6|12|потому что наша брань не против крови и плоти, но против начальств, против властей, против мироправителей тьмы века сего, против духов злобы поднебесной.
EPH|6|13|Для сего приимите всеоружие Божие, дабы вы могли противостать в день злый и, все преодолев, устоять.
EPH|6|14|Итак станьте, препоясав чресла ваши истиною и облекшись в броню праведности,
EPH|6|15|и обув ноги в готовность благовествовать мир;
EPH|6|16|а паче всего возьмите щит веры, которым возможете угасить все раскаленные стрелы лукавого;
EPH|6|17|и шлем спасения возьмите, и меч духовный, который есть Слово Божие.
EPH|6|18|Всякою молитвою и прошением молитесь во всякое время духом, и старайтесь о сем самом со всяким постоянством и молением о всех святых
EPH|6|19|и о мне, дабы мне дано было слово – устами моими открыто с дерзновением возвещать тайну благовествования,
EPH|6|20|для которого я исполняю посольство в узах, дабы я смело проповедывал, как мне должно.
EPH|6|21|А дабы и вы знали о моих обстоятельствах и делах, обо всем известит вас Тихик, возлюбленный брат и верный в Господе служитель,
EPH|6|22|которого я и послал к вам для того самого, чтобы вы узнали о нас и чтобы он утешил сердца ваши.
EPH|6|23|Мир братиям и любовь с верою от Бога Отца и Господа Иисуса Христа.
EPH|6|24|Благодать со всеми, неизменно любящими Господа нашего Иисуса Христа. Аминь.
