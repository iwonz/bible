ACTS|1|1|Primum quidem sermonem feci de omnibus, o Theophile, quae coepit Iesus facere et docere,
ACTS|1|2|usque in diem, qua, cum praecepisset apostolis per Spiritum Sanctum, quos elegit, assumptus est;
ACTS|1|3|quibus et praebuit seipsum vivum post passionem suam in multis argumentis, per dies quadraginta apparens eis et loquens ea, quae sunt de regno Dei.
ACTS|1|4|Et convescens praecepit eis ab Hierosolymis ne discederent, sed exspectarent promissionem Patris: " Quam audistis a me,
ACTS|1|5|quia Ioannes quidem baptizavit aqua, vos autem baptizabimini in Spiritu Sancto non post multos hos dies ".
ACTS|1|6|Igitur qui convenerant, interrogabant eum dicentes: " Domine, si in tempore hoc restitues regnum Israeli? ".
ACTS|1|7|Dixit autem eis: " Non est vestrum nosse tempora vel momenta, quae Pater posuit in sua potestate,
ACTS|1|8|sed accipietis virtutem, superveniente Sancto Spiritu in vos, et eritis mihi testes et in Ierusalem et in omni Iudaea et Samaria et usque ad ultimum terrae ".
ACTS|1|9|Et cum haec dixisset, videntibus illis, elevatus est, et nubes suscepit eum ab oculis eorum.
ACTS|1|10|Cumque intuerentur in caelum, eunte illo, ecce duo viri astiterunt iuxta illos in vestibus albis,
ACTS|1|11|qui et dixerunt: " Viri Galilaei, quid statis aspicientes in caelum? Hic Iesus, qui assumptus est a vobis in caelum, sic veniet quemadmodum vidistis eum euntem in caelum ".
ACTS|1|12|Tunc reversi sunt in Ierusalem a monte, qui vocatur Oliveti, qui est iuxta Ierusalem sabbati habens iter.
ACTS|1|13|Et cum introissent, in cenaculum ascenderunt, ubi manebant et Petrus et Ioannes et Iacobus et Andreas, Philippus et Thomas, Bartholomaeus et Matthaeus, Iacobus Alphaei et Simon Zelotes et Iudas Iacobi.
ACTS|1|14|Hi omnes erant perseverantes unanimiter in oratione cum mulieribus et Maria matre Iesu et fratribus eius.
ACTS|1|15|Et in diebus illis exsurgens Petrus in medio fratrum dixit - erat autem turba hominum simul fere centum viginti C:
ACTS|1|16|" Viri fratres, oportebat impleri Scripturam, quam praedixit Spiritus Sanctus per os David de Iuda, qui fuit dux eorum, qui comprehenderunt Iesum,
ACTS|1|17|quia connumeratus erat in nobis et sortitus est sortem ministerii huius.
ACTS|1|18|Hic quidem possedit agrum de mercede iniquitatis; et pronus factus crepuit medius, et diffusa sunt omnia viscera eius.
ACTS|1|19|Et notum factum est omnibus habitantibus Ierusalem, ita ut appellaretur ager ille lingua eorum Aceldamach, hoc est ager Sanguinis.
ACTS|1|20|Scriptum est enim in libro Psalmorum:Fiat commoratío eius deserta,et non sit qui inhabitet in ea"et: "Episcopatum eius accipiat alius".
ACTS|1|21|Oportet ergo ex his viris, qui nobiscum congregati erant in omni tempore, quo intravit et exivit inter nos Dominus Iesus,
ACTS|1|22|incipiens a baptismate Ioannis usque in diem, qua assumptus est a nobis, testem resurrectionis eius nobiscum fieri unum ex istis ".
ACTS|1|23|Et statuerunt duos, Ioseph, qui vocabatur Barsabbas, qui cognominatus est Iustus, et Matthiam.
ACTS|1|24|Et orantes dixerunt: " Tu, Domine, qui corda nosti omnium, ostende quem elegeris ex his duobus unum
ACTS|1|25|accipere locum ministerii huius et apostolatus, de quo praevaricatus est Iudas, ut abiret in locum suum ".
ACTS|1|26|Et dederunt sortes eis, et cecidit sors super Matthiam, et annumeratus est cum undecim apostolis.
ACTS|2|1|Et cum compleretur dies Pen tecostes, erant omnes pariter in eodem loco.
ACTS|2|2|Et factus est repente de caelo sonus tamquam advenientis spiritus vehementis et replevit totam domum, ubi erant sedentes.
ACTS|2|3|Et apparuerunt illis dispertitae linguae tamquam ignis, seditque supra singulos eorum;
ACTS|2|4|et repleti sunt omnes Spiritu Sancto et coeperunt loqui aliis linguis, prout Spiritus dabat eloqui illis.
ACTS|2|5|Erant autem in Ierusalem habitantes Iudaei, viri religiosi ex omni natione, quae sub caelo est;
ACTS|2|6|facta autem hac voce, convenit multitudo et confusa est, quoniam audiebat unusquisque lingua sua illos loquentes.
ACTS|2|7|Stupebant autem et mirabantur dicentes: " Nonne ecce omnes isti, qui loquuntur, Galilaei sunt?
ACTS|2|8|Et quomodo nos audimus unusquisque propria lingua nostra, in qua nati sumus?
ACTS|2|9|Parthi et Medi et Elamitae et qui habitant Mesopotamiam, Iudaeam quoque et Cappadociam, Pontum et Asiam,
ACTS|2|10|Phrygiam quoque et Pamphyliam, Aegyptum et partes Libyae, quae est circa Cyrenem, et advenae Romani,
ACTS|2|11|Iudaei quoque et proselyti, Cretes et Arabes, audimus loquentes eos nostris linguis magnalia Dei ".
ACTS|2|12|Stupebant autem omnes et haesitabant ad invicem dicentes: " Quidnam hoc vult esse? ";
ACTS|2|13|alii autem irridentes dicebant: " Musto pleni sunt isti ".
ACTS|2|14|Stans autem Petrus cum Undecim levavit vocem suam et locutus est eis: " Viri Iudaei et qui habitatis Ierusalem universi, hoc vobis notum sit, et auribus percipite verba mea.
ACTS|2|15|Non enim, sicut vos aestimatis, hi ebrii sunt, est enim hora diei tertia;
ACTS|2|16|sed hoc est, quod dictum est per prophetam Ioel:
ACTS|2|17|"Et erit: in novissimis diebus, dicit Deus,effundam de Spiritu meo super omnem carnem,et prophetabunt filii vestri et filiae vestrae,et iuvenes vestri visiones videbunt,et seniores vestri somnia somniabunt;
ACTS|2|18|et quidem super servos meos et super ancillas measin diebus illis effundam de Spiritu meo,et prophetabunt.
ACTS|2|19|Et dabo prodigia in caelo sursum et signa in terra deorsum,sanguinem et ignem et vaporem fumi;
ACTS|2|20|sol convertetur in tenebras,et luna in sanguinem,antequam veniat dies Dominimagnus et manifestus.
ACTS|2|21|Et erit:omnis quicumque invocaverit nomen Domini, salvus erit".
ACTS|2|22|Viri Israelitae, audite verba haec: Iesum Nazarenum, virum approbatum a Deo apud vos virtutibus et prodigiis et signis, quae fecit per illum Deus in medio vestri, sicut ipsi scitis,
ACTS|2|23|hunc definito consilio et praescientia Dei traditum per manum iniquorum affigentes interemistis,
ACTS|2|24|quem Deus suscitavit, solutis doloribus mortis, iuxta quod impossibile erat teneri illum ab ea.
ACTS|2|25|David enim dicit circa eum:Providebam Dominum coram me semper, quoniam a dextris meis est, ne commovear.
ACTS|2|26|Propter hoc laetatum est cor meum,et exsultavit lingua mea;insuper et caro mea requiescet in spe.
ACTS|2|27|Quoniam non derelinques animam meam in infernoneque dabis Sanctum tuum videre corruptionem.
ACTS|2|28|Notas fecisti mihi vias vitae,replebis me iucunditate cum facie tua".
ACTS|2|29|Viri fratres, liceat audenter dicere ad vos de patriarcha David, quoniam et defunctus est et sepultus est, et sepulcrum eius est apud nos usque in hodiernum diem;
ACTS|2|30|propheta igitur cum esset et sciret quia iure iurando iurasset illi Deus de fructu lumbi eius sedere super sedem eius,
ACTS|2|31|providens locutus est de resurrectione Christi, quia neque derelictus est in inferno, neque caro eius vidit corruptionem.
ACTS|2|32|Hunc Iesum resuscitavit Deus, cuius omnes nos testes sumus.
ACTS|2|33|Dextera igitur Dei exaltatus, et promissione Spiritus Sancti accepta a Patre, effudit hunc, quem vos videtis et auditis.
ACTS|2|34|Non enim David ascendit in caelos; dicit autem ipse:Dixit Dominus Domino meo: Sede a dextris meis,
ACTS|2|35|donec ponam inimicos tuos scabellum pedum tuorum".
ACTS|2|36|Certissime ergo sciat omnis domus Israel quia et Dominum eum et Christum Deus fecit, hunc Iesum, quem vos crucifixistis ".
ACTS|2|37|His auditis, compuncti sunt corde et dixerunt ad Petrum et reliquos apostolos: " Quid faciemus, viri fratres? ".
ACTS|2|38|Petrus vero ad illos: " Paenitentiam, inquit, agite, et baptizetur unusquisque vestrum in nomine Iesu Christi in remissionem peccatorum vestrorum, et accipietis donum Sancti Spiritus;
ACTS|2|39|vobis enim est repromissio et filiis vestris et omnibus, qui longe sunt, quoscumque advocaverit Dominus Deus noster ".
ACTS|2|40|Aliis etiam verbis pluribus testificatus est et exhortabatur eos dicens: " Salvamini a generatione ista prava ".
ACTS|2|41|Qui ergo, recepto sermone eius, baptizati sunt; et appositae sunt in il la die animae circiter tria milia.
ACTS|2|42|Erant autem perseverantes in doctrina apostolorum et communicatione, in fractione panis et orationibus.
ACTS|2|43|Fiebat autem omni animae timor; multa quoque prodigia et signa per apostolos fiebant.
ACTS|2|44|Omnes autem, qui crediderant, erant pariter et habebant omnia communia;
ACTS|2|45|et possessiones et substantias vendebant et dividebant illas omnibus, prout cuique opus erat;
ACTS|2|46|cotidie quoque perdurantes unanimiter in templo et frangentes circa domos panem, sumebant cibum cum exsultatione et simplicitate cordis,
ACTS|2|47|collaudantes Deum et habentes gratiam ad omnem plebem. Dominus autem augebat, qui salvi fierent cotidie in idipsum.
ACTS|3|1|Petrus autem et Ioannes ascen debant in templum ad horam orationis nonam.
ACTS|3|2|Et quidam vir, qui erat claudus ex utero matris suae, baiulabatur; quem ponebant cotidie ad portam templi, quae dicitur Speciosa, ut peteret eleemosynam ab introeuntibus in templum;
ACTS|3|3|is cum vidisset Petrum et Ioannem incipientes introire in templum, rogabat, ut eleemosynam acciperet.
ACTS|3|4|Intuens autem in eum Petrus cum Ioanne dixit: " Respice in nos ".
ACTS|3|5|At ille intendebat in eos, sperans se aliquid accepturum ab eis.
ACTS|3|6|Petrus autem dixit: " Argentum et aurum non est mihi; quod autem habeo, hoc tibi do: In nomine Iesu Christi Nazareni surge et ambula! ".
ACTS|3|7|Et apprehensa ei manu dextera, allevavit eum; et protinus consolidatae sunt bases eius et tali,
ACTS|3|8|et exsiliens stetit et ambulabat; et intravit cum illis in templum, ambulans et exsiliens et laudans Deum.
ACTS|3|9|Et vidit omnis populus eum ambulantem et laudantem Deum;
ACTS|3|10|cognoscebant autem illum quoniam ipse erat, qui ad eleemosynam sedebat ad Speciosam portam templi, et impleti sunt stupore et exstasi in eo, quod contigerat illi.
ACTS|3|11|Cum teneret autem Petrum et Ioannem, concurrit omnis populus ad eos ad porticum, qui appellatur Salomonis, stupentes.
ACTS|3|12|Videns autem Petrus respondit ad populum: " Viri Israelitae, quid miramini in hoc aut nos quid intuemini, quasi nostra virtute aut pietate fecerimus hunc ambulare?
ACTS|3|13|Deus Abraham et Deus Isaac et Deus Iacob, Deus patrum nostrorum, glorificavit puerum suum Iesum, quem vos quidem tradidistis et negastis ante faciem Pilati, iudicante illo dimitti;
ACTS|3|14|vos autem Sanctum et Iustum negastis et petistis virum homicidam donari vobis,
ACTS|3|15|ducem vero vitae interfecistis, quem Deus suscitavit a mortuis, cuius nos testes sumus.
ACTS|3|16|Et in fide nominis eius hunc, quem videtis et nostis, confirmavit nomen eius; et fides, quae per eum est, dedit huic integritatem istam in conspectu omnium vestrum.
ACTS|3|17|Et nunc, fratres, scio quia per ignorantiam fecistis, sicut et principes vestri;
ACTS|3|18|Deus autem, quae praenuntiavit per os omnium Prophetarum pati Christum suum, implevit sic.
ACTS|3|19|Paenitemini igitur et convertimini, ut deleantur vestra peccata,
ACTS|3|20|ut veniant tempora refrigerii a conspectu Domini, et mittat eum, qui praedestinatus est vobis Christus, Iesum,
ACTS|3|21|quem oportet caelum quidem suscipere usque in tempora restitutionis omnium, quae locutus est Deus per os sanctorum a saeculo suorum prophetarum.
ACTS|3|22|Moyses quidem dixit: "Prophetam vobis suscitabit Dominus Deus vester de fratribus vestris tamquam me; ipsum audietis iuxta omnia, quaecumque locutus fuerit vobis.
ACTS|3|23|Erit autem: omnis anima, quae non audierit prophetam illum, exterminabitur de plebe".
ACTS|3|24|Et omnes prophetae a Samuel et deinceps quotquot locuti sunt, etiam annuntiaverunt dies istos.
ACTS|3|25|Vos estis filii prophetarum et testamenti, quod disposuit Deus ad patres vestros dicens ad Abraham: "Et in semine tuo benedicentur omnes familiae terrae".
ACTS|3|26|Vobis primum Deus suscitans Puerum suum, misit eum benedicentem vobis in avertendo unumquemque a nequitiis vestris ".
ACTS|4|1|Loquentibus autem illis ad populum, supervenerunt eis sa cerdotes et magistratus templi et sadducaei,
ACTS|4|2|dolentes quod docerent populum et annuntiarent in Iesu resurrectionem ex mortuis;
ACTS|4|3|et iniecerunt in eos manus et posuerunt in custodiam in crastinum; erat enim iam vespera.
ACTS|4|4|Multi autem eorum, qui audierant verbum, crediderunt; et factus est numerus virorum quinque milia.
ACTS|4|5|Factum est autem in crastinum, ut congregarentur principes eorum et seniores et scribae in Ierusalem,
ACTS|4|6|et Annas princeps sacerdotum et Caiphas et Ioannes et Alexander et quotquot erant de genere sacerdotali,
ACTS|4|7|et statuentes eos in medio interrogabant: " In qua virtute aut in quo nomine fecistis hoc vos? ".
ACTS|4|8|Tunc Petrus repletus Spiritu Sancto dixit ad eos: " Principes populi et seniores,
ACTS|4|9|si nos hodie diiudicamur in benefacto hominis infirmi, in quo iste salvus factus est,
ACTS|4|10|notum sit omnibus vobis et omni plebi Israel quia in nomine Iesu Christi Nazareni, quem vos crucifixistis, quem Deus suscitavit a mortuis, in hoc iste astat coram vobis sanus.
ACTS|4|11|Hic estlapis, qui reprobatus est a vobis aedificatoribus,qui factus est in caput anguli.
ACTS|4|12|Et non est in alio aliquo salus, nec enim nomen aliud est sub caelo datum in hominibus, in quo oportet nos salvos fieri ".
ACTS|4|13|Videntes autem Petri fiduciam et Ioannis, et comperto quod homines essent sine litteris et idiotae, admirabantur et cognoscebant eos quoniam cum Iesu fuerant;
ACTS|4|14|hominem quoque videntes stantem cum eis, qui curatus fuerat, nihil poterant contradicere.
ACTS|4|15|Iubentes autem eos foras extra concilium secedere, conferebant ad invicem
ACTS|4|16|dicentes: " Quid faciemus hominibus istis? Quoniam quidem notum signum factum est per eos omnibus habitantibus in Ierusalem manifestum, et non possumus negare;
ACTS|4|17|sed ne amplius divulgetur in populum, comminemur eis, ne ultra loquantur in nomine hoc ulli hominum ".
ACTS|4|18|Et vocantes eos denuntiaverunt, ne omnino loquerentur neque docerent in nomine Iesu.
ACTS|4|19|Petrus vero et Ioannes respondentes dixerunt ad eos: " Si iustum est in conspectu Dei vos potius audire quam Deum, iudicate;
ACTS|4|20|non enim possumus nos, quae vidimus et audivimus, non loqui ".
ACTS|4|21|At illi ultra comminantes dimiserunt eos, nequaquam invenientes, quomodo punirent eos, propter populum, quia omnes glorificabant Deum in eo, quod acciderat;
ACTS|4|22|annorum enim erat amplius quadraginta homo, in quo factum erat signum istud sanitatis.
ACTS|4|23|Dimissi autem venerunt ad suos et annuntiaverunt quanta ad eos principes sacerdotum et seniores dixissent.
ACTS|4|24|Qui cum audissent, unanimiter levaverunt vocem ad Deum et dixerunt: " Domine, tu, qui fecisti caelum et terram et mare et omnia, quae in eis sunt,
ACTS|4|25|qui Spiritu Sancto per os patris nostri David pueri tui dixisti:Quare fremuerunt gentes,et populi meditati sunt inania?
ACTS|4|26|Astiterunt reges terrae,et principes convenerunt in unumadversus Dominum et adversus Christum eius".
ACTS|4|27|Convenerunt enim vere in civitate ista adversus sanctum puerum tuum Iesum, quem unxisti, Herodes et Pontius Pilatus cum gentibus et populis Israel
ACTS|4|28|facere, quaecumque manus tua et consilium praedestinavit fieri.
ACTS|4|29|Et nunc, Domine, respice in minas eorum et da servis tuis cum omni fiducia loqui verbum tuum,
ACTS|4|30|in eo quod manum tuam extendas ad sanitatem et signa et prodigia facienda per nomen sancti pueri tui Iesu ".
ACTS|4|31|Et cum orassent, motus est locus, in quo erant congregati, et repleti sunt omnes Sancto Spiritu et loquebantur verbum Dei cum fiducia.
ACTS|4|32|Multitudinis autem credentium erat cor et anima una, nec quisquam eorum, quae possidebant, aliquid suum esse dicebat, sed erant illis omnia communia.
ACTS|4|33|Et virtute magna reddebant apostoli testimonium resurrectionis Domini Iesu, et gratia magna erat super omnibus illis.
ACTS|4|34|Neque enim quisquam egens erat inter illos; quotquot enim possessores agrorum aut domorum erant, vendentes afferebant pretia eorum, quae vendebant,
ACTS|4|35|et ponebant ante pedes apostolorum; dividebatur autem singulis, prout cuique opus erat.
ACTS|4|36|Ioseph autem, qui cognominatus est Barnabas ab apostolis - quod est interpretatum filius Consolationis - Levites, Cyprius genere,
ACTS|4|37|cum haberet agrum, vendidit et attulit pecuniam et posuit ante pedes apostolorum.
ACTS|5|1|Vir autem quidam nomine Ananias cum Sapphira uxore sua vendidit agrum
ACTS|5|2|et subtraxit de pretio, conscia quoque uxore, et afferens partem quandam ad pedes apostolorum posuit.
ACTS|5|3|Dixit autem Petrus: " Anania, cur implevit Satanas cor tuum mentiri te Spiritui Sancto et subtrahere de pretio agri?
ACTS|5|4|Nonne manens tibi manebat et venumdatum in tua erat potestate? Quare posuisti in corde tuo hanc rem? Non es mentitus hominibus sed Deo! ".
ACTS|5|5|Audiens autem Ananias haec verba cecidit et exspiravit; et factus est timor magnus in omnes audientes.
ACTS|5|6|Surgentes autem iuvenes involverunt eum et efferentes sepelierunt.
ACTS|5|7|Factum est autem quasi horarum trium spatium, et uxor ipsius nesciens, quod factum fuerat, introivit.
ACTS|5|8|Respondit autem ei Petrus: " Dic mihi, si tanti agrum vendidistis? ". At illa dixit: " Etiam, tanti ".
ACTS|5|9|Petrus autem ad eam: " Quid est quod convenit vobis tentare Spiritum Domini? Ecce pedes eorum, qui sepelierunt virum tuum, ad ostium, et efferent te ".
ACTS|5|10|Confestim cecidit ante pedes eius et exspiravit; intrantes autem iuvenes invenerunt illam mortuam et efferentes sepelierunt ad virum suum.
ACTS|5|11|Et factus est timor magnus super universam ecclesiam et in omnes, qui audierunt haec.
ACTS|5|12|Per manus autem apostolorum fiebant signa et prodigia multa in plebe; et erant unanimiter omnes in porticu Salomonis.
ACTS|5|13|Ceterorum autem nemo audebat coniungere se illis, sed magnificabat eos populus;
ACTS|5|14|magis autem addebantur credentes Domino multitudines virorum ac mulierum,
ACTS|5|15|ita ut et in plateas efferrent infirmos et ponerent in lectulis et grabatis, ut, veniente Petro, saltem umbra illius obumbraret quemquam eorum.
ACTS|5|16|Concurrebat autem et multitudo vicinarum civitatum Ierusalem, afferentes aegros et vexatos ab spiritibus immundis, qui curabantur omnes.
ACTS|5|17|Exsurgens autem princeps sacerdotum et omnes, qui cum illo erant, quae est haeresis sadducaeorum, repleti sunt zelo
ACTS|5|18|et iniecerunt manus in apostolos et posuerunt illos in custodia publica.
ACTS|5|19|Angelus autem Domini per noctem aperuit ianuas carceris et educens eos dixit:
ACTS|5|20|" Ite et stantes loquimini in templo plebi omnia verba vitae huius ".
ACTS|5|21|Qui cum audissent, intraverunt diluculo in templum et docebant.Adveniens autem princeps sacerdotum et, qui cum eo erant, convocaverunt concilium et omnes seniores filiorum Israel et miserunt in carcerem, ut adducerentur illi.
ACTS|5|22|Cum venissent autem ministri, non invenerunt illos in carcere; reversi autem nuntiaverunt
ACTS|5|23|dicentes: " Carcerem invenimus clausum cum omni diligentia et custodes stantes ad ianuas; aperientes autem intus neminem invenimus! ".
ACTS|5|24|Ut audierunt autem hos sermones, magistratus templi et principes sacerdotum ambigebant de illis quidnam fieret illud.
ACTS|5|25|Adveniens autem quidam nuntiavit eis: " Ecce viri, quos posuistis in carcere, sunt in templo stantes et docentes populum ".
ACTS|5|26|Tunc abiens magistratus cum ministris adducebat illos, non per vim; timebant enim populum, ne lapidarentur.
ACTS|5|27|Et cum adduxissent illos, statuerunt in concilio. Et interrogavit eos princeps sacerdotum
ACTS|5|28|dicens: " Nonne praecipiendo praecepimus vobis, ne doceretis in nomine isto? Et ecce replevistis Ierusalem doctrina vestra et vultis inducere super nos sanguinem hominis istius ".
ACTS|5|29|Respondens autem Petrus et apostoli dixerunt: " Oboedire oportet Deo magis quam hominibus.
ACTS|5|30|Deus patrum nostrorum suscitavit Iesum, quem vos interemistis suspendentes in ligno;
ACTS|5|31|hunc Deus Ducem et Salvatorem exaltavit dextera sua ad dandam paenitentiam Israel et remissionem peccatorum.
ACTS|5|32|Et nos sumus testes horum verborum, et Spiritus Sanctus, quem dedit Deus oboedientibus sibi ".
ACTS|5|33|Haec cum audissent, dissecabantur et volebant interficere illos.
ACTS|5|34|Surgens autem quidam in concilio pharisaeus nomine Gamaliel, legis doctor honorabilis universae plebi, iussit foras ad breve homines fieri
ACTS|5|35|dixitque ad illos: " Viri Israelitae, attendite vobis super hominibus istis quid acturi sitis.
ACTS|5|36|Ante hos enim dies exstitit Theudas dicens esse se aliquem, cui consensit virorum numerus circiter quadringentorum; qui occisus est, et omnes, quicumque credebant ei, dissipati sunt et redacti sunt ad nihilum.
ACTS|5|37|Post hunc exstitit Iudas Galilaeus in diebus census et avertit populum post se; et ipse periit, et omnes, quotquot consentiebant ei, dispersi sunt.
ACTS|5|38|Et nunc dico vobis: Discedite ab hominibus istis et sinite illos. Quoniam si est ex hominibus consilium hoc aut opus hoc, dissolvetur;
ACTS|5|39|si vero ex Deo est, non poteritis dissolvere eos, ne forte et adversus Deum pugnantes inveniamini! ".Consenserunt autem illi
ACTS|5|40|et convocantes apostolos, caesis denuntiaverunt, ne loquerentur in nomine Iesu, et dimiserunt eos.
ACTS|5|41|Et illi quidem ibant gaudentes a conspectu concilii, quoniam digni habiti sunt pro nomine contumeliam pati;
ACTS|5|42|et omni die in templo et circa domos non cessabant docentes et evangelizantes Christum, Iesum.
ACTS|6|1|In diebus autem illis, crescente numero discipulorum, factus est murmur Graecorum adversus Hebraeos, eo quod neglegerentur in ministerio cotidiano viduae eorum.
ACTS|6|2|Convocantes autem Duodecim multitudinem discipulorum, dixerunt: " Non est aequum nos derelinquentes verbum Dei ministrare mensis;
ACTS|6|3|considerate vero, fratres, viros ex vobis boni testimonii septem plenos Spiritu et sapientia, quos constituemus super hoc opus;
ACTS|6|4|nos vero orationi et ministerio verbi instantes erimus ".
ACTS|6|5|Et placuit sermo coram omni multitudine; et elegerunt Stephanum, virum plenum fide et Spiritu Sancto, et Philippum et Prochorum et Nicanorem et Timonem et Parmenam et Nicolaum proselytum Antiochenum,
ACTS|6|6|quos statuerunt ante conspectum apostolorum, et orantes imposuerunt eis manus.
ACTS|6|7|Et verbum Dei crescebat, et multiplicabatur numerus discipulorum in Ierusalem valde; multa etiam turba sacerdotum oboediebat fidei.
ACTS|6|8|Stephanus autem plenus gratia et virtute faciebat prodigia et signa magna in populo.
ACTS|6|9|Surrexerunt autem quidam de synagoga, quae appellatur Libertinorum et Cyrenensium et Alexandrinorum et eorum, qui erant a Cilicia et Asia, disputantes cum Stephano;
ACTS|6|10|et non poterant resistere sapientiae et Spiritui, quo loquebatur.
ACTS|6|11|Tunc submiserunt viros, qui dicerent: " Audivimus eum dicentem verba blasphema in Moysen et Deum ";
ACTS|6|12|et commoverunt plebem et seniores et scribas, et concurrentes rapuerunt eum et adduxerunt in concilium
ACTS|6|13|et statuerunt testes falsos dicentes: " Homo iste non cessat loqui verba adversus locum sanctum et Legem;
ACTS|6|14|audivimus enim eum dicentem quoniam Iesus Nazarenus hic destruet locum istum et mutabit consuetudines, quas tradidit nobis Moyses ".
ACTS|6|15|Et intuentes eum omnes, qui sedebant in concilio, viderunt faciem eius tamquam faciem angeli.
ACTS|7|1|Dixit autem princeps sacerdo tum: " Si haec ita se habent? ".
ACTS|7|2|Qui ait: " Viri fratres et patres, audite. Deus gloriae apparuit patri nostro Abraham, cum esset in Mesopotamia, priusquam moraretur in Charran,
ACTS|7|3|et dixit ad illum: "Exi de terra tua et de cognatione tua et veni in terram, quam tibi monstravero".
ACTS|7|4|Tunc egressus de terra Chaldaeorum habitavit in Charran. Et inde, postquam mortuus est pater eius, transtulit illum in terram istam, in qua nunc vos habitatis;
ACTS|7|5|et non dedit illi hereditatem in ea nec passum pedis et repromisit dare illi eam in possessionem et semini eius post ipsum, cum non haberet filium.
ACTS|7|6|Locutus est autem sic Deus: "Erit semen eius accola in terra aliena, et servituti eos subicient et male tractabunt annis quadringentis;
ACTS|7|7|et gentem, cui servierint, iudicabo ego, dixit Deus; et post haec exibunt et deservient mihi in loco isto".
ACTS|7|8|Et dedit illi testamentum circumcisionis; et sic genuit Isaac et circumcidit eum die octava, et Isaac Iacob, et Iacob duodecim patriarchas.
ACTS|7|9|Et patriarchae aemulantes Ioseph vendiderunt in Aegyptum; et erat Deus cum eo
ACTS|7|10|et eripuit eum ex omnibus tribulationibus eius et dedit ei gratiam et sapientiam in conspectu pharaonis regis Aegypti; et constituit eum praepositum super Aegyptum et super omnem domum suam.
ACTS|7|11|Venit autem fames in universam Aegyptum et Chanaan et tribulatio magna, et non inveniebant cibos patres nostri.
ACTS|7|12|Cum audisset autem Iacob esse frumentum in Aegypto, misit patres nostros primum;
ACTS|7|13|et in secundo cognitus est Ioseph a fratribus suis, et manifestatum est pharaoni genus Ioseph.
ACTS|7|14|Mittens autem Ioseph accersivit Iacob patrem suum et omnem cognationem in animabus septuaginta quinque;
ACTS|7|15|et descendit Iacob in Aegyptum. Et defunctus est ipse et patres nostri;
ACTS|7|16|et translati sunt in Sichem et positi sunt in sepulcro, quod emit Abraham pretio argenti a filiis Hemmor in Sichem.
ACTS|7|17|Cum appropinquaret autem tempus repromissionis, quam confessus erat Deus Abrahae, crevit populus et multiplicatus est in Aegypto,
ACTS|7|18|quoadusque surrexit rex alius super Aegypto, qui non sciebat Ioseph.
ACTS|7|19|Hic circumveniens genus nostrum, afflixit patres, ut exponerent infantes suos, ne vivi servarentur.
ACTS|7|20|Eodem tempore natus est Moyses et erat formosus coram Deo; qui nutritus est tribus mensibus in domo patris.
ACTS|7|21|Exposito autem illo, sustulit eum filia pharaonis et enutrivit eum sibi in filium;
ACTS|7|22|et eruditus est Moyses in omni sapientia Aegyptiorum; et erat potens in verbis et in operibus suis.
ACTS|7|23|Cum autem impleretur ei quadraginta annorum tempus, ascendit in cor eius, ut visitaret fratres suos filios Israel.
ACTS|7|24|Et cum vidisset quendam iniuriam patientem, vindicavit et fecit ultionem ei, qui opprimebatur, percusso Aegyptio.
ACTS|7|25|Existimabat autem intellegere fratres, quoniam Deus per manum ipsius daret salutem illis; at illi non intellexerunt.
ACTS|7|26|Atque sequenti die apparuit illis litigantibus et reconciliabat eos in pacem dicens: "Viri, fratres estis; ut quid nocetis alterutrum?".
ACTS|7|27|Qui autem iniuriam faciebat proximo, reppulit eum dicens: "Quis te constituit principem et iudicem super nos?
ACTS|7|28|Numquid interficere me tu vis, quemadmodum interfecisti heri Aegyptium?".
ACTS|7|29|Fugit autem Moyses propter verbum istud; et factus est advena in terra Madian, ubi generavit filios duos.
ACTS|7|30|Et expletis annis quadraginta, apparuit illi in deserto montis Sinai angelus in ignis flamma rubi.
ACTS|7|31|Moyses autem videns admirabatur visum; accedente autem illo, ut consideraret, facta est vox Domini:
ACTS|7|32|"Ego Deus patrum tuorum, Deus Abraham et Isaac et Iacob". Tremefactus autem Moyses non audebat considerare.
ACTS|7|33|Dixit autem illi Dominus: "Solve calceamentum pedum tuorum; locus enim, in quo stas, terra sancta est.
ACTS|7|34|Videns vidi afflictionem populi mei, qui est in Aegypto, et gemitum eorum audivi et descendi liberare eos; et nunc veni, mittam te in Aegyptum".
ACTS|7|35|Hunc Moysen, quem negaverunt dicentes: "Quis te constituit principem et iudicem?", hunc Deus et principem et redemptorem misit cum manu angeli, qui apparuit illi in rubo.
ACTS|7|36|Hic eduxit illos faciens prodigia et signa in terra Aegypti et in Rubro mari et in deserto annis quadraginta.
ACTS|7|37|Hic est Moyses, qui dixit filiis Israel: "Prophetam vobis suscitabit Deus de fratribus vestris tamquam me".
ACTS|7|38|Hic est qui fuit in ecclesia in solitudine cum angelo, qui loquebatur ei in monte Sinai, et cum patribus nostris; qui accepit verba viva dare nobis;
ACTS|7|39|cui noluerunt oboedire patres nostri, sed reppulerunt et aversi sunt in cordibus suis in Aegyptum
ACTS|7|40|dicentes ad Aaron: "Fac nobis deos, qui praecedant nos; Moyses enim hic, qui eduxit nos de terra Aegypti, nescimus quid factum sit ei".
ACTS|7|41|Et vitulum fecerunt in illis diebus et obtulerunt hostiam simulacro et laetabantur in operibus manuum suarum.
ACTS|7|42|Convertit autem Deus et tradidit eos servire militiae caeli, sicut scriptum est in libro Prophetarum:Numquid victimas et hostias obtulistis mihiannis quadraginta in deserto, domus Israel?
ACTS|7|43|Et suscepistis tabernaculum Molochet sidus dei vestri Rhaephan,figuras, quas fecistis ad adorandum eas.Et transferam vos trans Babylonem".
ACTS|7|44|Tabernaculum testimonii erat patribus nostris in deserto, sicut disposuit, qui loquebatur ad Moysen, ut faceret illud secundum formam, quam viderat;
ACTS|7|45|quod et induxerunt suscipientes patres nostri cum Iesu in possessionem gentium, quas expulit Deus a facie patrum nostrorum, usque in diebus David,
ACTS|7|46|qui invenit gratiam ante Deum et petiit, ut inveniret tabernaculum domui Iacob.
ACTS|7|47|Salomon autem aedificavit illi domum.
ACTS|7|48|Sed non Altissimus in manufactis habitat, sicut propheta dicit:
ACTS|7|49|"Caelum mihi thronus est,terra autem scabellum pedum meorum.Quam domum aedificabitis mihi, dicit Dominus,aut quis locus requietionis meae?
ACTS|7|50|Nonne manus mea fecit haec omnia?".
ACTS|7|51|Duri cervice et incircumcisi cordibus et auribus, vos semper Spiritui Sancto resistitis; sicut patres vestri, et vos.
ACTS|7|52|Quem prophetarum non sunt persecuti patres vestri? Et occiderunt eos, qui praenuntiabant de adventu Iusti, cuius vos nunc proditores et homicidae fuistis,
ACTS|7|53|qui accepistis legem in dispositionibus angelorum et non custodistis ".
ACTS|7|54|Audientes autem haec, dissecabantur cordibus suis et stridebant dentibus in eum.
ACTS|7|55|Cum autem esset plenus Spiritu Sancto, intendens in caelum vidit gloriam Dei et Iesum stantem a dextris Dei
ACTS|7|56|et ait: " Ecce video caelos apertos et Filium hominis a dextris stantem Dei ".
ACTS|7|57|Exclamantes autem voce magna continuerunt aures suas et impetum fecerunt unanimiter in eum
ACTS|7|58|et eicientes extra civitatem lapidabant. Et testes deposuerunt vestimenta sua secus pedes adulescentis, qui vocabatur Saulus.
ACTS|7|59|Et lapidabant Stephanum invocantem et dicentem: " Domine Iesu, suscipe spiritum meum ".
ACTS|7|60|Positis autem genibus clamavit voce magna: " Domine, ne statuas illis hoc peccatum "; et cum hoc dixisset, obdormivit.
ACTS|8|1|Saulus autem erat consentiens neci eius. Facta est autem in illa die persecutio magna in ecclesiam, quae erat Hierosolymis; et omnes dispersi sunt per regiones Iudaeae et Samariae praeter apostolos.
ACTS|8|2|Sepelierunt autem Stephanum viri timorati et fecerunt planctum magnum super illum.
ACTS|8|3|Saulus vero devastabat ecclesiam, per domos intrans et trahens viros ac mulieres tradebat in custodiam.
ACTS|8|4|Igitur qui dispersi erant, pertransierunt evangelizantes verbum.
ACTS|8|5|Philippus autem descendens in civitatem Samariae praedicabat illis Christum.
ACTS|8|6|Intendebant autem turbae his, quae a Philippo dicebantur, unanimiter, audientes et videntes signa, quae faciebat:
ACTS|8|7|ex multis enim eorum, qui habebant spiritus immundos, clamantes voce magna exibant; multi autem paralytici et claudi curati sunt.
ACTS|8|8|Factum est autem magnum gaudium in illa civitate.
ACTS|8|9|Vir autem quidam nomine Simon iampridem erat in civitate magias faciens et dementans gentem Samariae, dicens esse se aliquem magnum;
ACTS|8|10|cui attendebant omnes a minimo usque ad maximum dicentes: " Hic est virtus Dei, quae vocatur Magna ".
ACTS|8|11|Attendebant autem eum, propter quod multo tempore magiis dementasset eos.
ACTS|8|12|Cum vero credidissent Philippo evangelizanti de regno Dei et nomine Iesu Christi, baptizabantur viri ac mulieres.
ACTS|8|13|Tunc Simon et ipse credidit et, cum baptizatus esset, adhaerebat Philippo; videns etiam signa et virtutes magnas fieri stupens admirabatur.
ACTS|8|14|Cum autem audissent apostoli, qui erant Hierosolymis, quia recepit Samaria verbum Dei, miserunt ad illos Petrum et Ioannem;
ACTS|8|15|qui cum descendissent, oraverunt pro ipsis, ut acciperent Spiritum Sanctum:
ACTS|8|16|nondum enim super quemquam illorum venerat, sed baptizati tantum erant in nomine Domini Iesu.
ACTS|8|17|Tunc imposuerunt manus super illos, et accipiebant Spiritum Sanctum.
ACTS|8|18|Cum vidisset autem Simon quia per impositionem manuum apostolorum daretur Spiritus, obtulit eis pecuniam
ACTS|8|19|dicens: " Date et mihi hanc potestatem, ut cuicumque imposuero manus, accipiat Spiritum Sanctum ".
ACTS|8|20|Petrus autem dixit ad eum: " Argentum tuum tecum sit in perditionem, quoniam donum Dei existimasti pecunia possideri!
ACTS|8|21|Non est tibi pars neque sors in verbo isto; cor enim tuum non est rectum coram Deo.
ACTS|8|22|Paenitentiam itaque age ab hac nequitia tua et roga Dominum, si forte remittatur tibi haec cogitatio cordis tui;
ACTS|8|23|in felle enim amaritudinis et obligatione iniquitatis video te esse ".
ACTS|8|24|Respondens autem Simon dixit: " Precamini vos pro me ad Dominum, ut nihil veniat super me horum, quae dixistis ".
ACTS|8|25|Et illi quidem testificati et locuti verbum Domini, redibant Hierosolymam et multis vicis Samaritanorum evangelizabant.
ACTS|8|26|Angelus autem Domini locutus est ad Philippum dicens: " Surge et vade contra meridianum ad viam, quae descendit ab Ierusalem in Gazam; haec est deserta ".
ACTS|8|27|Et surgens abiit; et ecce vir Aethiops eunuchus potens Candacis reginae Aethiopum, qui erat super omnem gazam eius, qui venerat adorare in Ierusalem
ACTS|8|28|et revertebatur sedens super currum suum et legebat prophetam Isaiam.
ACTS|8|29|Dixit autem Spiritus Philippo: " Accede et adiunge te ad currum istum.
ACTS|8|30|Accurrens autem Philippus audivit illum legentem Isaiam prophetam et dixit: " Putasne intellegis, quae legis? ".
ACTS|8|31|Qui ait: " Et quomodo possum, si non aliquis ostenderit mihi? ". Rogavitque Philippum, ut ascenderet et sederet secum.
ACTS|8|32|Locus autem Scripturae, quem legebat, erat hic: Tamquam ovis ad occisionem ductus estet sicut agnus coram tondente se sine voce,sic non aperit os suum.
ACTS|8|33|In humilitate eius iudicium eius sublatum est.Generationem illius quis enarrabit?Quoniam tollitur de terra vita eius ".
ACTS|8|34|Respondens autem eunuchus Philippo dixit: " Obsecro te, de quo propheta dicit hoc? De se an de alio aliquo? ".
ACTS|8|35|Aperiens autem Philippus os suum et incipiens a Scriptura ista, evangelizavit illi Iesum.
ACTS|8|36|Et dum irent per viam, venerunt ad quandam aquam; et ait eunuchus: " Ecce aqua; quid prohibet me baptizari? ".
ACTS|8|37|()
ACTS|8|38|Et iussit stare currum; et descenderunt uterque in aquam Philippus et eunuchus, et baptizavit eum.
ACTS|8|39|Cum autem ascendissent de aqua, Spiritus Domini rapuit Philippum, et amplius non vidit eum eunuchus; ibat autem per viam suam gaudens.
ACTS|8|40|Philippus autem inventus est in Azoto et pertransiens evangelizabat civitatibus cunctis, donec veniret Caesaream.
ACTS|9|1|Saulus autem, adhuc spirans minarum et caedis in discipulos Domini, accessit ad principem sacerdotum
ACTS|9|2|et petiit ab eo epistulas in Damascum ad synagogas, ut, si quos invenisset huius viae viros ac mulieres, vinctos perduceret in Ierusalem.
ACTS|9|3|Et cum iter faceret, contigit ut appropinquaret Damasco; et subito circumfulsit eum lux de caelo,
ACTS|9|4|et cadens in terram audivit vocem dicentem sibi: " Saul, Saul, quid me persequeris? ".
ACTS|9|5|Qui dixit: " Quis es, Domine? ". Et ille: " Ego sum Iesus, quem tu persequeris!
ACTS|9|6|Sed surge et ingredere civitatem, et dicetur tibi quid te oporteat facere ".
ACTS|9|7|Viri autem illi, qui comitabantur cum eo, stabant stupefacti, audientes quidem vocem, neminem autem videntes.
ACTS|9|8|Surrexit autem Saulus de terra; apertisque oculis, nihil videbat; ad manus autem illum trahentes introduxerunt Damascum.
ACTS|9|9|Et erat tribus diebus non videns et non manducavit neque bibit.
ACTS|9|10|Erat autem quidam discipulus Damasci nomine Ananias; et dixit ad illum in visu Dominus: " Anania ". At ille ait: " Ecce ego, Domine ".
ACTS|9|11|Et Dominus ad illum: " Surgens vade in vicum, qui vocatur Rectus, et quaere in domo Iudae Saulum nomine Tarsensem; ecce enim orat
ACTS|9|12|et vidit virum Ananiam nomine introeuntem et imponentem sibi manus, ut visum recipiat ".
ACTS|9|13|Respondit autem Ananias: " Domine, audivi a multis de viro hoc, quanta mala sanctis tuis fecerit in Ierusalem;
ACTS|9|14|et hic habet potestatem a principibus sacerdotum alligandi omnes, qui invocant nomen tuum ".
ACTS|9|15|Dixit autem ad eum Dominus: " Vade, quoniam vas electionis est mihi iste, ut portet nomen meum coram gentibus et regibus et filiis Israel;
ACTS|9|16|ego enim ostendam illi quanta oporteat eum pro nomine meo pati ".
ACTS|9|17|Et abiit Ananias; et introivit in domum et imponens ei manus dixit: " Saul frater, Dominus misit me, Iesus qui apparuit tibi in via, qua veniebas, ut videas et implearis Spiritu Sancto ".
ACTS|9|18|Et confestim ceciderunt ab oculis eius tamquam squamae, et visum recepit. Et surgens baptizatus est
ACTS|9|19|et, cum accepisset cibum, confortatus est.Fuit autem cum discipulis, qui erant Damasci, per dies aliquot;
ACTS|9|20|et continuo in synagogis praedicabat Iesum, quoniam hic est Filius Dei.
ACTS|9|21|Stupebant autem omnes, qui audiebant, et dicebant: " Nonne hic est, qui expugnabat in Ierusalem eos, qui invocabant nomen istud, et huc ad hoc venerat, ut vinctos illos duceret ad principes sacerdotum? ".
ACTS|9|22|Saulus autem magis convalescebat et confundebat Iudaeos, qui habitabant Damasci, affirmans quoniam hic est Christus.
ACTS|9|23|Cum implerentur autem dies multi, consilium fecerunt Iudaei, ut eum interficerent;
ACTS|9|24|notae autem factae sunt Saulo insidiae eorum. Custodiebant autem et portas die ac nocte, ut eum interficerent;
ACTS|9|25|accipientes autem discipuli eius nocte per murum dimiserunt eum submittentes in sporta.
ACTS|9|26|Cum autem venisset in Ierusalem, tentabat iungere se discipulis; et omnes timebant eum, non credentes quia esset discipulus.
ACTS|9|27|Barnabas autem apprehensum illum duxit ad apostolos et narravit illis quomodo in via vidisset Dominum, et quia locutus est ei, et quomodo in Damasco fiducialiter egerit in nomine Iesu.
ACTS|9|28|Et erat cum illis intrans et exiens in Ierusalem, fiducialiter agens in nomine Domini.
ACTS|9|29|Loquebatur quoque et disputabat cum Graecis; illi autem quaerebant occidere eum.
ACTS|9|30|Quod cum cognovissent, fratres deduxerunt eum Caesaream et dimiserunt Tarsum.
ACTS|9|31|Ecclesia quidem per totam Iudaeam et Galilaeam et Samariam habebat pacem; aedificabatur et ambulabat in timore Domini et consolatione Sancti Spiritus crescebat.
ACTS|9|32|Factum est autem Petrum, dum pertransiret universos, devenire et ad sanctos, qui habitabant Lyddae.
ACTS|9|33|Invenit autem ibi hominem quendam nomine Aeneam ab annis octo iacentem in grabato, qui erat paralyticus.
ACTS|9|34|Et ait illi Petrus: " Aenea, sanat te Iesus Christus; surge et sterne tibi ". Et continuo surrexit.
ACTS|9|35|Et viderunt illum omnes, qui inhabitabant Lyddam et Saron, qui conversi sunt ad Dominum.
ACTS|9|36|In Ioppe autem erat quaedam discipula nomine Tabitha, quae interpretata dicitur Dorcas; haec erat plena operibus bonis et eleemosynis, quas faciebat.
ACTS|9|37|Factum est autem in diebus illis ut infirmata moreretur; quam cum lavissent, posuerunt in cenaculo.
ACTS|9|38|Cum autem prope esset Lydda ab Ioppe, discipuli audientes quia Petrus esset in ea, miserunt duos viros ad eum rogantes: " Ne pigriteris venire usque ad nos! ".
ACTS|9|39|Exsurgens autem Petrus venit cum illis; et cum advenisset, duxerunt illum in cenaculum; et circumsteterunt illum omnes viduae flentes et ostendentes tunicas et vestes, quas faciebat Dorcas, cum esset cum illis.
ACTS|9|40|Eiectis autem omnibus foras Petrus, et ponens genua oravit et conversus ad corpus dixit: " Tabitha, surge! ". At illa aperuit oculos suos et, viso Petro, resedit.
ACTS|9|41|Dans autem illi manum erexit eam et, cum vocasset sanctos et viduas, exhibuit eam vivam.
ACTS|9|42|Notum autem factum est per universam Ioppen, et crediderunt multi in Domino.
ACTS|9|43|Factum est autem, ut dies multos moraretur in Ioppe apud quendam Simonem coriarium.
ACTS|10|1|Vir autem quidam in Cae sarea nomine Cornelius, cen turio cohortis, quae dicitur Italica,
ACTS|10|2|religiosus et timens Deum cum omni domo sua, faciens eleemosynas multas plebi et deprecans Deum semper,
ACTS|10|3|vidit in visu manifeste quasi hora nona diei angelum Dei introeuntem ad se et dicentem sibi: " Corneli ".
ACTS|10|4|At ille intuens eum et timore correptus dixit: " Quid est, domine? ". Dixit autem illi: " Orationes tuae et eleemosynae tuae ascenderunt in memoriam in conspectu Dei.
ACTS|10|5|Et nunc mitte viros in Ioppen et accersi Simonem quendam, qui cognominatur Petrus;
ACTS|10|6|hic hospitatur apud Simonem quendam coriarium, cui est domus iuxta mare.
ACTS|10|7|Ut autem discessit angelus, qui loquebatur illi, cum vocasset duos domesticos suos et militem religiosum ex his, qui illi parebant,
ACTS|10|8|et narrasset illis omnia, misit illos in Ioppen.
ACTS|10|9|Postera autem die, iter illis facientibus et appropinquantibus civitati, ascendit Petrus super tectum, ut oraret circa horam sextam.
ACTS|10|10|Et cum esuriret, voluit gustare; parantibus autem eis, cecidit super eum mentis excessus,
ACTS|10|11|et videt caelum apertum et descendens vas quoddam velut linteum magnum quattuor initiis submitti in terram,
ACTS|10|12|in quo erant omnia quadrupedia et serpentia terrae et volatilia caeli.
ACTS|10|13|Et facta est vox ad eum: " Surge, Petre, occide et manduca! ".
ACTS|10|14|Ait autem Petrus: " Nequaquam, Domine, quia numquam manducavi omne commune et immundum ".
ACTS|10|15|Et vox iterum secundo ad eum: " Quae Deus purificavit, ne tu commune dixeris ".
ACTS|10|16|Hoc autem factum est per ter, et statim receptum est vas in caelum.
ACTS|10|17|Et dum intra se haesitaret Petrus quidnam esset visio, quam vidisset, ecce viri, qui missi erant a Cornelio, inquirentes domum Simonis astiterunt ad ianuam
ACTS|10|18|et, cum vocassent, interrogabant si Simon, qui cognominatur Petrus, illic haberet hospitium.
ACTS|10|19|Petro autem cogitante de visione, dixit Spiritus ei: " Ecce viri tres quaerunt te;
ACTS|10|20|surge itaque et descende et vade cum eis nihil dubitans, quia ego misi illos ".
ACTS|10|21|Descendens autem Petrus ad viros dixit: " Ecce ego sum, quem quaeritis; quae causa est, propter quam venistis? ".
ACTS|10|22|Qui dixerunt: " Cornelius centurio, vir iustus et timens Deum et testimonium habens ab universa gente Iudaeorum, responsum accepit ab angelo sancto accersire te in domum suam et audire verba abs te ".
ACTS|10|23|Invitans igitur eos recepit hospitio.Sequenti autem die, surgens profectus est cum eis, et quidam ex fratribus ab Ioppe comitati sunt eum.
ACTS|10|24|Altera autem die introivit Caesaream; Cornelius vero exspectabat illos, convocatis cognatis suis et necessariis amicis.
ACTS|10|25|Et factum est, cum introisset Petrus, obvius ei Cornelius procidens ad pedes adoravit.
ACTS|10|26|Petrus vero levavit eum dicens: " Surge, et ego ipse homo sum ".
ACTS|10|27|Et loquens cum illo intravit et invenit multos, qui convenerant;
ACTS|10|28|dixitque ad illos: " Vos scitis quomodo illicitum sit viro Iudaeo coniungi aut accedere ad alienigenam. Et mihi ostendit Deus neminem communem aut immundum dicere hominem;
ACTS|10|29|propter quod sine dubitatione veni accersitus. Interrogo ergo quam ob causam accersistis me ".
ACTS|10|30|Et Cornelius ait: " A nudius quarta die usque in hanc horam orans eram hora nona in domo mea, et ecce vir stetit ante me in veste candida
ACTS|10|31|et ait: "Corneli, exaudita est oratio tua, et eleemosynae tuae commemoratae sunt in conspectu Dei.
ACTS|10|32|Mitte ergo in Ioppen et accersi Simonem, qui cognominatur Petrus; hic hospitatur in domo Simonis coriarii iuxta mare".
ACTS|10|33|Confestim igitur misi ad te, et tu bene fecisti veniendo. Nunc ergo omnes nos in conspectu Dei adsumus audire omnia, quaecumque tibi praecepta sunt a Domino ".
ACTS|10|34|Aperiens autem Petrus os dixit: " In veritate comperio quoniam non est personarum acceptor Deus,
ACTS|10|35|sed in omni gente, qui timet eum et operatur iustitiam, acceptus est illi.
ACTS|10|36|Verbum misit filiis Israel evangelizans pacem per Iesum Christum; hic est omnium Dominus.
ACTS|10|37|Vos scitis quod factum est verbum per universam Iudaeam incipiens a Galilaea post baptismum, quod praedicavit Ioannes:
ACTS|10|38|Iesum a Nazareth, quomodo unxit eum Deus Spiritu Sancto et virtute, qui pertransivit benefaciendo et sanando omnes oppressos a Diabolo, quoniam Deus erat cum illo.
ACTS|10|39|Et nos testes sumus omnium, quae fecit in regione Iudaeorum et Ierusalem; quem et occiderunt suspendentes in ligno.
ACTS|10|40|Hunc Deus suscitavit tertia die et dedit eum manifestum fieri
ACTS|10|41|non omni populo, sed testibus praeordinatis a Deo, nobis, qui manducavimus et bibimus cum illo postquam resurrexit a mortuis;
ACTS|10|42|et praecepit nobis praedicare populo et testificari quia ipse est, qui constitutus est a Deo iudex vivorum et mortuorum.
ACTS|10|43|Huic omnes Prophetae testimonium perhibent remissionem peccatorum accipere per nomen eius omnes, qui credunt in eum ".
ACTS|10|44|Adhuc loquente Petro verba haec, cecidit Spiritus Sanctus super omnes, qui audiebant verbum.
ACTS|10|45|Et obstupuerunt, qui ex circumcisione fideles, qui venerant cum Petro, quia et in nationes gratia Spiritus Sancti effusa est;
ACTS|10|46|audiebant enim illos loquentes linguis et magnificantes Deum. Tunc respondit Petrus:
ACTS|10|47|" Numquid aquam quis prohibere potest, ut non baptizentur hi, qui Spiritum Sanctum acceperunt sicut et nos? ".
ACTS|10|48|Et iussit eos in nomine Iesu Christi baptizari. Tunc rogaverunt eum, ut maneret aliquot diebus.
ACTS|11|1|Audierunt autem apostoli et fratres, qui erant in Iudaea, quoniam et gentes receperunt verbum Dei.
ACTS|11|2|Cum ascendisset autem Petrus in Ierusalem, disceptabant adversus illum, qui erant ex circumcisione,
ACTS|11|3|dicentes: " Introisti ad viros praeputium habentes et manducasti cum illis! ".
ACTS|11|4|Incipiens autem Petrus exponebat illis ex ordine dicens:
ACTS|11|5|" Ego eram in civitate Ioppe orans et vidi in excessu mentis visionem, descendens vas quoddam velut linteum magnum quattuor initiis submitti de caelo et venit usque ad me;
ACTS|11|6|in quod intuens considerabam et vidi quadrupedia terrae et bestias et reptilia et volatilia caeli.
ACTS|11|7|Audivi autem et vocem dicentem mihi: "Surgens, Petre, occide et manduca!".
ACTS|11|8|Dixi autem: Nequaquam, Domine, quia commune aut immundum numquam introivit in os meum.
ACTS|11|9|Respondit autem vox secundo de caelo: "Quae Deus mundavit, tu ne commune dixeris".
ACTS|11|10|Hoc autem factum est per ter, et retracta sunt rursum omnia in caelum.
ACTS|11|11|Et ecce confestim tres viri astiterunt in domo, in qua eramus, missi a Caesarea ad me.
ACTS|11|12|Dixit autem Spiritus mihi, ut irem cum illis nihil haesitans. Venerunt autem mecum et sex fratres isti, et ingressi sumus in domum viri.
ACTS|11|13|Narravit autem nobis quomodo vidisset angelum ad domum suam stantem et dicentem: "Mitte in Ioppen et accersi Simonem, qui cognominatur Petrus,
ACTS|11|14|qui loquetur tibi verba, in quibus salvus eris tu et universa domus tua".
ACTS|11|15|Cum autem coepissem loqui, decidit Spiritus Sanctus super eos, sicut et super nos in initio.
ACTS|11|16|Recordatus sum autem verbi Domini, sicut dicebat: "Ioannes quidem baptizavit aqua, vos autem baptizabimini in Spiritu Sancto".
ACTS|11|17|Si ergo aequale donum dedit illis Deus sicut et nobis, qui credidimus in Dominum Iesum Christum, ego quis eram qui possem prohibere Deum? ".
ACTS|11|18|His autem auditis, acquieverunt et glorificaverunt Deum dicentes: " Ergo et gentibus Deus paenitentiam ad vitam dedit ".
ACTS|11|19|Et illi quidem, qui dispersi fuerant a tribulatione, quae facta fuerat sub Stephano, perambulaverunt usque Phoenicen et Cyprum et Antiochiam, nemini loquentes verbum; nisi solis Iudaeis.
ACTS|11|20|Erant autem quidam ex eis viri Cyprii et Cyrenaei, qui, cum introissent Antiochiam, loquebantur et ad Graecos evangelizantes Dominum Iesum.
ACTS|11|21|Et erat manus Domini cum eis; multusque numerus credentium conversus est ad Dominum.
ACTS|11|22|Auditus est autem sermo in auribus ecclesiae, quae erat in Ierusalem, super istis, et miserunt Barnabam usque Antiochiam;
ACTS|11|23|qui cum pervenisset et vidisset gratiam Dei, gavisus est et hortabatur omnes proposito cordis permanere in Domino,
ACTS|11|24|quia erat vir bonus et plenus Spiritu Sancto et fide. Et apposita est turba multa Domino.
ACTS|11|25|Profectus est autem Tarsum, ut quaereret Saulum;
ACTS|11|26|quem cum invenisset, perduxit Antiochiam. Factum est autem eis, ut annum totum conversarentur in ecclesia et docerent turbam multam, et cognominarentur primum Antiochiae discipuli Christiani.
ACTS|11|27|In his autem diebus supervenerunt ab Hierosolymis prophetae Antiochiam;
ACTS|11|28|et surgens unus ex eis nomine Agabus significavit per Spiritum famem magnam futuram in universo orbe terrarum; quae facta est sub Claudio.
ACTS|11|29|Discipuli autem, prout quis habebat, proposuerunt singuli eorum in ministerium mittere habitantibus in Iudaea fratribus;
ACTS|11|30|quod et fecerunt, mittentes ad presbyteros per manum Barnabae et Sauli.
ACTS|12|1|Illo autem tempore, misit Herodes rex manus, ut affli geret quosdam de ecclesia.
ACTS|12|2|Occidit autem Iacobum fratrem Ioannis gladio.
ACTS|12|3|Videns autem quia placeret Iudaeis, apposuit apprehendere et Petrum - erant autem dies Azymorum -
ACTS|12|4|quem cum apprehendisset, misit in carcerem tradens quattuor quaternionibus militum custodire eum, volens post Pascha producere eum populo.
ACTS|12|5|Et Petrus quidem servabatur in carcere; oratio autem fiebat sine intermissione ab ecclesia ad Deum pro eo.
ACTS|12|6|Cum autem producturus eum esset Herodes, in ipsa nocte erat Petrus dormiens inter duos milites vinctus catenis duabus, et custodes ante ostium custodiebant carcerem.
ACTS|12|7|Et ecce angelus Domini astitit, et lumen refulsit in habitaculo; percusso autem latere Petri, suscitavit eum dicens: " Surge velociter! ". Et ceciderunt catenae de manibus eius.
ACTS|12|8|Dixit autem angelus ad eum: " Praecingere et calcea te sandalia tua! ". Et fecit sic. Et dicit illi: " Circumda tibi vestimentum tuum et sequere me! ".
ACTS|12|9|Et exiens sequebatur et nesciebat quia verum est, quod fiebat per angelum; aestimabat autem se visum videre.
ACTS|12|10|Transeuntes autem primam custodiam et secundam venerunt ad portam ferream, quae ducit ad civitatem, quae ultro aperta est eis, et exeuntes processerunt vicum unum, et continuo discessit angelus ab eo.
ACTS|12|11|Et Petrus ad se reversus dixit: " Nunc scio vere quia misit Dominus angelum suum et eripuit me de manu Herodis et de omni exspectatione plebis Iudaeorum ".
ACTS|12|12|Consideransque venit ad domum Mariae matris Ioannis, qui cognominatur Marcus, ubi erant multi congregati et orantes.
ACTS|12|13|Pulsante autem eo ostium ianuae, processit puella ad audiendum, nomine Rhode;
ACTS|12|14|et ut cognovit vocem Petri, prae gaudio non aperuit ianuam, sed intro currens nuntiavit stare Petrum ante ianuam.
ACTS|12|15|At illi dixerunt ad eam: " Insanis! ". Illa autem affirmabat sic se habere. Illi autem dicebant: " Angelus eius est ".
ACTS|12|16|Petrus autem perseverabat pulsans; cum autem aperuissent, viderunt eum et obstupuerunt.
ACTS|12|17|Annuens autem eis manu, ut tacerent, enarravit quomodo Dominus eduxisset eum de carcere dixitque: " Nuntiate Iacobo ct fratribus haec ". Et egressus abiit in alium locum.
ACTS|12|18|Facta autem die, erat non parva turbatio inter milites, quidnam de Petro factum esset.
ACTS|12|19|Herodes autem, cum requisisset eum et non invenisset, interrogatis custodibus, iussit eos abduci; descendensque a Iudaea in Caesaream ibi commorabatur.
ACTS|12|20|Erat autem iratus Tyriis et Sidoniis; at illi unanimes venerunt ad eum et, persuaso Blasto, qui erat super cubiculum regis, postulabant pacem, eo quod aleretur regio eorum ab annona regis.
ACTS|12|21|Statuto autem die, Herodes, vestitus veste regia, sedens pro tribunalicontionabatur ad eos;
ACTS|12|22|populus autem acclamabat: " Dei vox et non hominis! ".
ACTS|12|23|Confestim autem percussit eum angelus Domini, eo quod non dedisset gloriam Deo; et consumptus a vermibus exspiravit.
ACTS|12|24|Verbum autem Dei crescebat et multiplicabatur.
ACTS|12|25|Barnabas autem et Saulus reversi sunt in Ierusalem expleto ministerio, assumpto Ioanne, qui cognominatus est Marcus.
ACTS|13|1|Erant autem in ecclesia, quae erat Antiochiae, pro phetae et doctores: Barnabas et Simeon, qui vocabatur Niger, et Lucius Cyrenensis et Manaen, qui erat Herodis tetrarchae collactaneus, et Saulus.
ACTS|13|2|Ministrantibus autem illis Domino et ieiunantibus, dixit Spiritus Sanctus: " Separate mihi Barnabam et Saulum in opus, ad quod vocavi eos ".
ACTS|13|3|Tunc ieiunantes et orantes imponentesque eis manus dimiserunt illos.
ACTS|13|4|Et ipsi quidem missi ab Spiritu Sancto devenerunt Seleuciam et inde navigaverunt Cyprum
ACTS|13|5|et, cum venissent Salamina, praedicabant verbum Dei in synagogis Iudaeorum; habebant autem et Ioannem ministrum.
ACTS|13|6|Et cum perambulassent universam insulam usque Paphum, invenerunt quendam virum magum pseudoprophetam Iudaeum, cui nomen Bariesu,
ACTS|13|7|qui erat cum proconsule Sergio Paulo, viro prudente. Hic, accitis Barnaba et Saulo, quaesivit audire verbum Dei;
ACTS|13|8|resistebat autem illis Elymas, magus, sic enim interpretatur nomen eius, quaerens avertere proconsulem a fide.
ACTS|13|9|Saulus autem, qui et Paulus, repletus Spiritu Sancto, intuens in eum
ACTS|13|10|dixit: " O plene omni dolo et omni fallacia, fili Diaboli, inimice omnis iustitiae, non desines subvertere vias Domini rectas?
ACTS|13|11|Et nunc, ecce manus Domini super te; et eris caecus, non videns solem usque ad tempus ". Et confestim cecidit in eum caligo et tenebrae, et circumiens quaerebat, qui eum manum darent.
ACTS|13|12|Tunc proconsul, cum vidisset factum, credidit admirans super doctrinam Domini.
ACTS|13|13|Et cum a Papho navigassent, qui erant cum Paulo, venerunt Pergen Pamphyliae; Ioannes autem discedens ab eis reversus est Hierosolymam.
ACTS|13|14|Illi vero pertranseuntes, a Perge venerunt Antiochiam Pisidiae, et ingressi synagogam die sabbatorum sederunt.
ACTS|13|15|Post lectionem autem Legis et Prophetarum, miserunt principes synagogae ad eos dicentes: " Viri fratres, si quis est in vobis sermo exhortationis ad plebem, dicite! ".
ACTS|13|16|Surgens autem Paulus et manu silentium indicens ait: " Viri Israelitae et qui timetis Deum, audite.
ACTS|13|17|Deus plebis huius Israel elegit patres nostros et plebem exaltavit, cum essent incolae in terra Aegypti, et in brachio excelso eduxit eos ex ea;
ACTS|13|18|et per quadraginta fere annorum tempus mores eorum sustinuit in deserto;
ACTS|13|19|et destruens gentes septem in terra Chanaan sorte distribuit terram eorum,
ACTS|13|20|quasi quadringentos et quinquaginta annos. Et post haec dedit iudices usque ad Samuel prophetam.
ACTS|13|21|Et exinde postulaverunt regem, et dedit illis Deus Saul filium Cis, virum de tribu Beniamin, annis quadraginta.
ACTS|13|22|Et amoto illo, suscitavit illis David in regem, cui et testimonium perhibens dixit: "Inveni David filium Iesse, virum secundum cor meum, qui faciet omnes voluntates meas".
ACTS|13|23|Huius Deus ex semine secundum promissionem eduxit Israel salvatorem Iesum,
ACTS|13|24|praedicante Ioanne ante adventum eius baptismum paenitentiae omni populo Israel.
ACTS|13|25|Cum impleret autem Ioannes cursum suum, dicebat: "Quid me arbitramini esse? Non sum ego; sed ecce venit post me, cuius non sum dignus calceamenta pedum solvere".
ACTS|13|26|Viri fratres, filii generis Abraham et qui in vobis timent Deum, nobis verbum salutis huius missum est.
ACTS|13|27|Qui enim habitabant Ierusalem et principes eorum, hunc ignorantes et voces Prophetarum, quae per omne sabbatum leguntur, iudicantes impleverunt;
ACTS|13|28|et nullam causam mortis invenientes petierunt a Pilato, ut interficeretur;
ACTS|13|29|cumque consummassent omnia, quae de eo scripta erant, deponentes eum de ligno posuerunt in monumento.
ACTS|13|30|Deus vero suscitavit eum a mortuis;
ACTS|13|31|qui visus est per dies multos his, qui simul ascenderant cum eo de Galilaea in Ierusalem, qui nunc sunt testes eius ad plebem.
ACTS|13|32|Et nos vobis evangelizamus eam, quae ad patres promissio facta est,
ACTS|13|33|quoniam hanc Deus adimplevit filiis eorum, nobis resuscitans Iesum, sicut et in Psalmo secundo scriptum est:Filius meus es tu; ego hodie genui te".
ACTS|13|34|Quod autem suscitaverit eum a mortuis, amplius iam non reversurum in corruptionem, ita dixit: "Dabo vobis sancta David fidelia".
ACTS|13|35|Ideoque et in alio dicit:Non dabis Sanctum tuum videre corruptionem".
ACTS|13|36|David enim sua generatione cum administrasset voluntati Dei, dormivit et appositus est ad patres suos et vidit corruptionem;
ACTS|13|37|quem vero Deus suscitavit, non vidit corruptionem.
ACTS|13|38|Notum igitur sit vobis, viri fratres, quia per hunc vobis remissio peccatorum annuntiatur; ab omnibus, quibus non potuistis in lege Moysi iustificari,
ACTS|13|39|in hoc omnis, qui credit, iustificatur.
ACTS|13|40|Videte ergo, ne superveniat, quod dictum est in Prophetis:
ACTS|13|41|"Videte, contemptores,et admiramini et disperdimini,quia opus operor ego in diebus vestris,opus, quod non credetis, si quis enarraverit vobis!" ".
ACTS|13|42|Exeuntibus autem illis, rogabant, ut sequenti sabbato loquerentur sibi verba haec.
ACTS|13|43|Cumque dimissa esset synagoga, secuti sunt multi Iudaeorum et colentium proselytorum Paulum et Barnabam, qui loquentes suadebant eis, ut permanerent in gratia Dei.
ACTS|13|44|Sequenti vero sabbato paene universa civitas convenit audire verbum Domini.
ACTS|13|45|Videntes autem turbas Iudaei, repleti sunt zelo; et contradicebant his, quae a Paulo dicebantur, blasphemantes.
ACTS|13|46|Tunc audenter Paulus et Barnabas dixerunt: " Vobis oportebat primum loqui verbum Dei; sed quoniam repellitis illud et indignos vos iudicatis aeternae vitae, ecce convertimur ad gentes.
ACTS|13|47|Sic enim praecepit nobis Dominus:Posui te in lumen gentium,ut sis in salutem usque ad extremum terrae" ".
ACTS|13|48|Audientes autem gentes gaudebant et glorificabant verbum Domini, et crediderunt, quotquot erant praeordinati ad vitam aeternam;
ACTS|13|49|ferebatur autem verbum Domini per universam regionem.
ACTS|13|50|Iudaei autem concitaverunt honestas inter colentes mulieres et primos civitatis et excitaverunt persecutionem in Paulum et Barnabam et eiecerunt eos de finibus suis.
ACTS|13|51|At illi, excusso pulvere pedum in eos, venerunt Iconium;
ACTS|13|52|discipuli quoque replebantur gaudio et Spiritu Sancto.
ACTS|14|1|Factum est autem Iconii, ut eodem modo introirent syna gogam Iudaeorum et ita loquerentur, ut crederet Iudaeorum et Graecorum copiosa multitudo.
ACTS|14|2|Qui vero increduli fuerunt Iudaei, suscitaverunt et exacerbaverunt animas gentium adversus fratres.
ACTS|14|3|Multo igitur tempore demorati sunt, fiducialiter agentes in Domino, testimonium perhibente verbo gratiae suae, dante signa et prodigia fieri per manus eorum.
ACTS|14|4|Divisa est autem multitudo civitatis: et quidam quidem erant cum Iudaeis, quidam vero cum apostolis.
ACTS|14|5|Cum autem factus esset impetus gentilium et Iudaeorum cum principibus suis, ut contumeliis afficerent et lapidarent eos,
ACTS|14|6|intellegentes confugerunt ad civitates Lycaoniae, Lystram et Derben et ad regionem in circuitu
ACTS|14|7|et ibi evangelizantes erant.
ACTS|14|8|Et quidam vir in Lystris infirmus pedibus sedebat, claudus ex utero matris suae, qui numquam ambulaverat.
ACTS|14|9|Hic audivit Paulum loquentem; qui intuitus eum et videns quia haberet fidem, ut salvus fieret,
ACTS|14|10|dixit magna voce: " Surge super pedes tuos rectus! ". Et exsilivit et ambulabat.
ACTS|14|11|Turbae autem cum vidissent, quod fecerat Paulus, levaverunt vocem suam Lycaonice dicentes: " Dii similes facti hominibus descenderunt ad nos! ";
ACTS|14|12|et vocabant Barnabam Iovem, Paulum vero Mercurium, quoniam ipse erat dux verbi.
ACTS|14|13|Sacerdos quoque templi Iovis, quod erat ante civitatem, tauros et coronas ad ianuas afferens cum populis, volebat sacrificare.
ACTS|14|14|Quod ubi audierunt apostoli Barnabas et Paulus, conscissis tunicis suis, exsilierunt in turbam clamantes
ACTS|14|15|et dicentes: " Viri, quid haec facitis? Et nos mortales sumus similes vobis homines, evangelizantes vobis ab his vanis converti ad Deum vivum, qui fecit caelum et terram et mare et omnia, quae in eis sunt.
ACTS|14|16|Qui in praeteritis generationibus permisit omnes gentes ambulare in viis suis;
ACTS|14|17|et quidem non sine testimonio semetipsum reliquit benefaciens, de caelo dans vobis pluvias et tempora fructifera, implens cibo et laetitia corda vestra ".
ACTS|14|18|Et haec dicentes vix sedaverunt turbas, ne sibi immolarent.
ACTS|14|19|Supervenerunt autem ab Antiochia et Iconio Iudaei et persuasis turbis lapidantesque Paulum trahebant extra civitatem aestimantes eum mortuum esse.
ACTS|14|20|Circumdantibus autem eum discipulis, surgens intravit civitatem. Et postera die profectus est cum Barnaba in Derben.
ACTS|14|21|Cumque evangelizassent civitati illi et docuissent multos, reversi sunt Lystram et Iconium et Antiochiam
ACTS|14|22|confirmantes animas discipulorum, exhortantes, ut permanerent in fide, et quoniam per multas tribulationes oportet nos intrare in regnum Dei.
ACTS|14|23|Et cum ordinassent illis per singulas ecclesias presbyteros et orassent cum ieiunationibus, commendaverunt eos Domino, in quem crediderant.
ACTS|14|24|Transeuntesque Pisidiam venerunt Pamphyliam;
ACTS|14|25|et loquentes in Perge verbum descenderunt in Attaliam.
ACTS|14|26|Et inde navigaverunt Antiochiam, unde erant traditi gratiae Dei in opus, quod compleverunt.
ACTS|14|27|Cum autem venissent et congregassent ecclesiam, rettulerunt quanta fecisset Deus cum illis et quia aperuisset gentibus ostium fidei.
ACTS|14|28|Morati sunt autem tempus non modicum cum discipulis.
ACTS|15|1|Et quidam descendentes de Iudaea docebant fratres: " Nisi circumcidamini secundum morem Moysis, non potestis salvi fieri ".
ACTS|15|2|Facta autem seditione et conquisitione non minima Paulo et Barnabae adversum illos, statuerunt, ut ascenderent Paulus et Barnabas et quidam alii ex illis ad apostolos et presbyteros in Ierusalem super hac quaestione.
ACTS|15|3|Illi igitur deducti ab ecclesia pertransiebant Phoenicen et Samariam narrantes conversionem gentium et faciebant gaudium magnum omnibus fratribus.
ACTS|15|4|Cum autem venissent Hierosolymam, suscepti sunt ab ecclesia et apostolis et presbyteris et annuntiaverunt quanta Deus fecisset cum illis.
ACTS|15|5|Surrexerunt autem quidam de haeresi pharisaeorum, qui crediderant, dicentes: " Oportet circumcidere eos, praecipere quoque servare legem Moysis! ".
ACTS|15|6|Conveneruntque apostoli et presbyteri videre de verbo hoc.
ACTS|15|7|Cum autem magna conquisitio fieret, surgens Petrus dixit ad eos: " Viri fratres, vos scitis quoniam ab antiquis diebus in vobis elegit Deus per os meum audire gentes verbum evangelii et credere;
ACTS|15|8|et qui novit corda, Deus, testimonium perhibuit illis dans Spiritum Sanctum sicut et nobis;
ACTS|15|9|et nihil discrevit inter nos et illos fide purificans corda eorum.
ACTS|15|10|Nunc ergo quid tentatis Deum imponere iugum super cervicem discipulorum, quod neque patres nostri neque nos portare potuimus?
ACTS|15|11|Sed per gratiam Domini Iesu credimus salvari quemadmodum et illi ".
ACTS|15|12|Tacuit autem omnis multitudo, et audiebant Barnabam et Paulum narrantes quanta fecisset Deus signa et prodigia in gentibus per eos.
ACTS|15|13|Et postquam tacuerunt, respondit Iacobus dicens: " Viri fratres, audite me.
ACTS|15|14|Simeon narravit quemadmodum primum Deus visitavit sumere ex gentibus populum nomini suo;
ACTS|15|15|et huic concordant verba Prophetarum, sicut scriptum est:
ACTS|15|16|"Post haec revertaret reaedificabo tabernaculum David, quod decidit,et diruta eius reaedificabo et erigam illud.
ACTS|15|17|ut requirant reliqui hominum Dominumet omnes gentes, super quas invocatum est nomen meum,dicit Dominus faciens haec
ACTS|15|18|nota a saeculo".
ACTS|15|19|Propter quod ego iudico non inquietari eos, qui ex gentibus convertuntur ad Deum,
ACTS|15|20|sed scribere ad eos, ut abstineant se a contaminationibus simulacrorum et fornicatione et suffocato et sanguine.
ACTS|15|21|Moyses enim a generationibus antiquis habet in singulis civitatibus, qui eum praedicent in synagogis, ubi per omne sabbatum legitur ".
ACTS|15|22|Tunc placuit apostolis et presbyteris cum omni ecclesia electos viros ex eis mittere Antiochiam cum Paulo et Barnaba: Iudam, qui cognominatur Barsabbas, et Silam, viros primos in fratribus,
ACTS|15|23|scribentes per manum eorum: " Apostoli et presbyteri fratres his, qui sunt Antiochiae et Syriae et Ciliciae, fratribus ex gentibus, salutem!
ACTS|15|24|Quoniam audivimus quia quidam ex nobis, quibus non mandavimus, exeuntes turbaverunt vos verbis evertentes animas vestras,
ACTS|15|25|placuit nobis collectis in unum eligere viros et mittere ad vos cum carissimis nobis Barnaba et Paulo,
ACTS|15|26|hominibus, qui tradiderunt animas suas pro nomine Domini nostri Iesu Christi.
ACTS|15|27|Misimus ergo Iudam et Silam, qui et ipsi verbis referent eadem.
ACTS|15|28|Visum est enim Spiritui Sancto et nobis nihil ultra imponere vobis oneris quam haec necessario:
ACTS|15|29|abstinere ab idolothytis et sanguine et suffocatis et fornicatione; a quibus custodientes vos bene agetis. Valete ".
ACTS|15|30|Illi igitur dimissi descenderunt Antiochiam et, congregata multitudine, tradiderunt epistulam;
ACTS|15|31|quam cum legissent, gavisi sunt super consolatione.
ACTS|15|32|Iudas quoque et Silas, cum et ipsi essent prophetae, verbo plurimo consolati sunt fratres et confirmaverunt.
ACTS|15|33|Facto autem tempore, dimissi sunt cum pace a fratribus ad eos, qui miserant illos.
ACTS|15|34|()
ACTS|15|35|Paulus autem et Barnabas demorabantur Antiochiae docentes et evangelizantes cum aliis pluribus verbum Domini.
ACTS|15|36|Post aliquot autem dies dixit ad Barnabam Paulus: " Revertentes visitemus fratres per universas civitates, in quibus praedicavimus verbum Domini, quomodo se habeant ".
ACTS|15|37|Barnabas autem volebat secum assumere et Ioannem, qui cognominatur Marcus;
ACTS|15|38|Paulus autem iudicabat eum, qui discessisset ab eis a Pamphylia et non isset cum eis in opus, non debere recipi eum.
ACTS|15|39|Facta est autem exacerbatio, ita ut discederent ab invicem, et Barnabas, assumpto Marco, navigaret Cyprum.
ACTS|15|40|Paulus vero, electo Sila, profectus est, traditus gratiae Domini a fratribus;
ACTS|15|41|perambulabat autem Syriam et Ciliciam confirmans ecclesias.
ACTS|16|1|Pervenit autem in Derben et Lystram. Et ecce discipulus quidam erat ibi nomine Timotheus, filius mulieris Iudaeae fidelis, patre autem Graeco;
ACTS|16|2|huic testimonium reddebant, qui in Lystris erant et Iconii fratres.
ACTS|16|3|Hunc voluit Paulus secum proficisci et assumens circumcidit eum propter Iudaeos, qui erant in illis locis; sciebant enim omnes quod pater eius Graecus esset.
ACTS|16|4|Cum autem pertransirent civitates, tradebant eis custodire dogmata, quae erant decreta ab apostolis et presbyteris, qui essent Hierosolymis.
ACTS|16|5|Ecclesiae quidem confirmabantur fide et abundabant numero cotidie.
ACTS|16|6|Transierunt autem Phrygiam et Galatiae regionem, vetati a Sancto Spiritu loqui verbum in Asia;
ACTS|16|7|cum venissent autem circa Mysiam, tentabant ire Bithyniam, et non permisit eos Spiritus Iesu;
ACTS|16|8|cum autem praeterissent Mysiam, descenderunt Troadem.
ACTS|16|9|Et visio per noctem Paulo ostensa est: vir Macedo quidam erat stans et deprecans eum et dicens: " Transiens in Macedoniam, adiuva nos! ".
ACTS|16|10|Ut autem visum vidit, statim quaesivimus proficisci in Macedoniam, certi facti quia vocasset nos Deus evangelizare eis.
ACTS|16|11|Navigantes autem a Troade recto cursu venimus Samothraciam et sequenti die Neapolim
ACTS|16|12|et inde Philippos, quae est prima partis Macedoniae civitas, colonia. Eramus autem in hac urbe diebus aliquot commorantes.
ACTS|16|13|Die autem sabbatorum egressi sumus foras portam iuxta flumen, ubi putabamus orationem esse, et sedentes loquebamur mulieribus, quae convenerant.
ACTS|16|14|Et quaedam mulier nomine Lydia, purpuraria civitatis Thyatirenorum colens Deum, audiebat, cuius Dominus aperuit cor intendere his, quae dicebantur a Paulo.
ACTS|16|15|Cum autem baptizata esset et domus eius, deprecata est dicens: " Si iudicastis me fidelem Domino esse, introite in domum meam et manete "; et coegit nos.
ACTS|16|16|Factum est autem, euntibus nobis ad orationem, puellam quandam habentem spiritum pythonem obviare nobis, quae quaestum magnum praestabat dominis suis divinando.
ACTS|16|17|Haec subsecuta Paulum et nos clamabat dicens: " Isti homines servi Dei Altissimi sunt, qui annuntiant vobis viam salutis ".
ACTS|16|18|Hoc autem faciebat multis diebus. Dolens autem Paulus et conversus spiritui dixit: " Praecipio tibi in nomine Iesu Christi exire ab ea "; et exiit eadem hora.
ACTS|16|19|Videntes autem domini eius quia exivit spes quaestus eorum, apprehendentes Paulum et Silam traxerunt in forum ad principes;
ACTS|16|20|et producentes eos magistratibus dixerunt: " Hi homines conturbant civitatem nostram, cum sint Iudaei,
ACTS|16|21|et annuntiant mores, quos non licet nobis suscipere neque facere, cum simus Romani ".
ACTS|16|22|Et concurrit plebs adversus eos; et magistratus, scissis tunicis eorum, iusserunt virgis caedi
ACTS|16|23|et, cum multas plagas eis imposuissent, miserunt eos in carcerem, praecipientes custodi, ut caute custodiret eos;
ACTS|16|24|qui cum tale praeceptum accepisset, misit eos in interiorem carcerem et pedes eorum strinxit in ligno.
ACTS|16|25|Media autem nocte, Paulus et Silas orantes laudabant Deum, et audiebant eos, qui in custodia erant;
ACTS|16|26|subito vero terraemotus factus est magnus, ita ut moverentur fundamenta carceris, et aperta sunt statim ostia omnia, et universorum vincula soluta sunt.
ACTS|16|27|Expergefactus autem custos carceris et videns apertas ianuas carceris, evaginato gladio volebat se interficere, aestimans fugisse vinctos.
ACTS|16|28|Clamavit autem Paulus magna voce dicens: " Nihil feceris tibi mali; universi enim hic sumus ".
ACTS|16|29|Petitoque lumine, intro cucurrit et tremefactus procidit Paulo et Silae;
ACTS|16|30|et producens eos foras ait: " Domini, quid me oportet facere, ut salvus fiam? ".
ACTS|16|31|At illi dixerunt: " Crede in Domino Iesu et salvus eris tu et domus tua.
ACTS|16|32|Et locuti sunt ei verbum Domini cum omnibus, qui erant in domo eius.
ACTS|16|33|Et tollens eos in illa hora noctis lavit eos a plagis, et baptizatus est ipse et omnes eius continuo;
ACTS|16|34|cumque perduxisset eos in domum, apposuit mensam et laetatus est cum omni domo sua credens Deo.
ACTS|16|35|Et cum dies factus esset, miserunt magistratus lictores dicentes: " Dimitte homines illos! ".
ACTS|16|36|Nuntiavit autem custos carceris verba haec Paulo: " Miserunt magistratus, ut dimittamini; nunc igitur exeuntes ite in pace ".
ACTS|16|37|Paulus autem dixit eis: " Caesos nos publice, indemnatos, cum homines Romani essemus, miserunt in carcerem; et nunc occulte nos eiciunt? Non ita, sed veniant et ipsi nos educant ".
ACTS|16|38|Nuntiaverunt autem magistratibus lictores verba haec. Timueruntque audito quod Romani essent;
ACTS|16|39|et venientes deprecati sunt eos et educentes rogabant, ut egrederentur urbem.
ACTS|16|40|Exeuntes autem de carcere introierunt ad Lydiam et, visis fratribus, consolati sunt eos et profecti sunt.
ACTS|17|1|Cum autem perambulassent Amphipolim et Apolloniam, venerunt Thessalonicam, ubi erat synagoga Iudaeorum.
ACTS|17|2|Secundum consuetudinem autem suam Paulus introivit ad eos et per sabbata tria disserebat eis de Scripturis
ACTS|17|3|adaperiens et comprobans quia Christum oportebat pati et resurgere a mortuis, et: " Hic est Christus, Iesus, quem ego annuntio vobis ".
ACTS|17|4|Et quidam ex eis crediderunt et adiuncti sunt Paulo et Silae et de colentibus Graecis multitudo magna et mulieres nobiles non paucae.
ACTS|17|5|Zelantes autem Iudaei assumentesque de foro viros quosdam malos et turba facta concitaverunt civitatem; et assistentes domui Iasonis quaerebant eos producere in populum.
ACTS|17|6|Et cum non invenissent eos, trahebant Iasonem et quosdam fratres ad politarchas clamantes: " Qui orbem concitaverunt, isti et huc venerunt,
ACTS|17|7|quos suscepit Iason; et hi omnes contra decreta Caesaris faciunt, regem alium dicentes esse, Iesum ".
ACTS|17|8|Concitaverunt autem plebem et politarchas audientes haec;
ACTS|17|9|et accepto satis ab Iasone et a ceteris, dimiserunt eos.
ACTS|17|10|Fratres vero confestim per noctem dimiserunt Paulum et Silam in Beroeam; qui cum advenissent, in synagogam Iudaeorum introierunt.
ACTS|17|11|Hi autem erant nobiliores eorum, qui sunt Thessalonicae, qui susceperunt verbum cum omni aviditate, cotidie scrutantes Scripturas, si haec ita se haberent.
ACTS|17|12|Et multi quidem crediderunt ex eis et Graecarum mulierum honestarum et virorum non pauci.
ACTS|17|13|Cum autem cognovissent in Thessalonica Iudaei quia et Beroeae annuntiatum est a Paulo verbum Dei, venerunt et illuc commoventes et turbantes multitudinem.
ACTS|17|14|Statimque tunc Paulum dimiserunt fratres, ut iret usque ad mare; Silas autem et Timotheus remanserunt ibi.
ACTS|17|15|Qui autem deducebant Paulum, perduxerunt usque Athenas; et accepto mandato ad Silam et Timotheum, ut quam celerrime venirent ad illum, profecti sunt.
ACTS|17|16|Paulus autem cum Athenis eos exspectaret, irritabatur spiritus eius in ipso videns idololatriae deditam civitatem.
ACTS|17|17|Disputabat igitur in synagoga cum Iudaeis et colentibus et in foro per omnes dies ad eos, qui aderant.
ACTS|17|18|Quidam autem ex Epicureis et Stoicis philosophi disserebant cum eo. Et quidam dicebant: " Quid vult seminiverbius hic dicere? "; alii vero: " Novorum daemoniorum videtur annuntiator esse ", quia Iesum et resurrectionem evangelizabat.
ACTS|17|19|Et apprehensum eum ad Areopagum duxerunt dicentes: " Possumus scire quae est haec nova, quae a te dicitur, doctrina?
ACTS|17|20|Mira enim quaedam infers auribus nostris; volumus ergo scire quidnam velint haec esse ".
ACTS|17|21|Athenienses autem omnes et advenae hospites ad nihil aliud vacabant nisi aut dicere aut audire aliquid novi.
ACTS|17|22|Stans autem Paulus in medio Areopagi ait: " Viri Athenienses, per omnia quasi superstitiosiores vos video;
ACTS|17|23|praeteriens enim et videns simulacra vestra inveni et aram, in qua scriptum erat: "Ignoto deo". Quod ergo ignorantes colitis, hoc ego annuntio vobis.
ACTS|17|24|Deus, qui fecit mundum et omnia, quae in eo sunt, hic, caeli et terrae cum sit Dominus, non in manufactis templis inhabitat
ACTS|17|25|nec manibus humanis colitur indigens aliquo, cum ipse det omnibus vitam et inspirationem et omnia;
ACTS|17|26|fecitque ex uno omne genus hominum inhabitare super universam faciem terrae, definiens statuta tempora et terminos habitationis eorum,
ACTS|17|27|quaerere Deum, si forte attrectent eum et inveniant, quamvis non longe sit ab unoquoque nostrum.
ACTS|17|28|In ipso enim vivimus et movemur et sumus, sicut et quidam vestrum poetarum dixerunt:Ipsius enim et genus sumus".
ACTS|17|29|Genus ergo cum simus Dei, non debemus aestimare auro aut argento aut lapidi, sculpturae artis et cogitationis hominis, divinum esse simile.
ACTS|17|30|Et tempora quidem ignorantiae despiciens Deus, nunc annuntiat hominibus, ut omnes ubique paenitentiam agant,
ACTS|17|31|eo quod statuit diem, in qua iudicaturus est orbem in iustitia in viro, quem constituit, fidem praebens omnibus suscitans eum a mortuis ".
ACTS|17|32|Cum audissent autem resurrectionem mortuorum, quidam quidem irridebant, quidam vero dixerunt: " Audiemus te de hoc iterum ".
ACTS|17|33|Sic Paulus exivit de medio eorum.
ACTS|17|34|Quidam vero viri adhaerentes ei crediderunt; in quibus et Dionysius Areopagita et mulier nomine Damaris et alii cum eis.
ACTS|18|1|Post haec discedens ab Athe nis venit Corinthum.
ACTS|18|2|Et in veniens quendam Iudaeum nomine Aquilam, Ponticum genere, qui nuper venerat ab Italia, et Priscillam uxorem eius, eo quod praecepisset Claudius discedere omnes Iudaeos a Roma, accessit ad eos
ACTS|18|3|et, quia eiusdem erat artis, manebat apud eos et operabatur; erant autem scenofactoriae artis.
ACTS|18|4|Disputabat autem in synagoga per omne sabbatum suadebatque Iudaeis et Graecis.
ACTS|18|5|Cum venissent autem de Macedonia Silas et Timotheus, instabat verbo Paulus testificans Iudaeis esse Christum Iesum.
ACTS|18|6|Contradicentibus autem eis et blasphemantibus, excutiens vestimenta dixit ad eos: " Sanguis vester super caput vestrum! Mundus ego. Ex hoc nunc ad gentes vadam ".
ACTS|18|7|Et migrans inde intravit in domum cuiusdam nomine Titi Iusti, colentis Deum, cuius domus erat coniuncta synagogae.
ACTS|18|8|Crispus autem archisynagogus credidit Domino cum omni domo sua, et multi Corinthiorum audientes credebant et baptizabantur.
ACTS|18|9|Dixit autem Dominus nocte per visionem Paulo: " Noli timere, sed loquere et ne taceas,
ACTS|18|10|quia ego sum tecum, et nemo apponetur tibi, ut noceat te, quoniam populus est mihi multus in hac civitate ".
ACTS|18|11|Sedit autem annum et sex menses docens apud eos verbum Dei.
ACTS|18|12|Gallione autem proconsule Achaiae, insurrexerunt uno animo Iudaei in Paulum et adduxerunt eum ad tribunal
ACTS|18|13|dicentes: " Contra legem hic persuadet hominibus colere Deum ".
ACTS|18|14|Incipiente autem Paulo aperire os, dixit Gallio ad Iudaeos: " Si quidem esset iniquum aliquid aut facinus pessimum, o Iudaei, merito vos sustinerem;
ACTS|18|15|si vero quaestiones sunt de verbo et nominibus et lege vestra, vos ipsi videritis; iudex ego horum nolo esse ".
ACTS|18|16|Et minavit eos a tribunali.
ACTS|18|17|Apprehendentes autem omnes Sosthenen, principem synagogae, percutiebant ante tribunal; et nihil horum Gallioni curae erat.
ACTS|18|18|Paulus vero, cum adhuc sustinuisset dies multos, fratribus valefaciens navigabat Syriam, et cum eo Priscilla et Aquila, qui sibi totonderat in Cenchreis caput; habebat enim votum.
ACTS|18|19|Deveneruntque Ephesum, et illos ibi reliquit; ipse vero ingressus synagogam disputabat cum Iudaeis.
ACTS|18|20|Rogantibus autem eis, ut ampliore tempore maneret, non consensit,
ACTS|18|21|sed valefaciens et dicens: " Iterum revertar ad vos Deo volente ", navigavit ab Epheso;
ACTS|18|22|et descendens Caesaream ascendit et salutavit ecclesiam et descendit Antiochiam.
ACTS|18|23|Et facto ibi aliquanto tempore, profectus est perambulans ex ordine Galaticam regionem et Phrygiam, confirmans omnes discipulos.
ACTS|18|24|Iudaeus autem quidam Apollo nomine, Alexandrinus natione, vir eloquens, devenit Ephesum, potens in Scripturis.
ACTS|18|25|Hic erat catechizatus viam Domini; et fervens spiritu loquebatur et docebat diligenter ea, quae sunt de Iesu, sciens tantum baptisma Ioannis.
ACTS|18|26|Hic ergo coepit fiducialiter agere in synagoga; quem cum audissent Priscilla et Aquila, assumpserunt eum et diligentius exposuerunt ei viam Dei.
ACTS|18|27|Cum autem vellet transire in Achaiam, exhortati fratres scripserunt discipulis, ut susciperent eum; qui cum venisset, contulit multum his, qui crediderant per gratiam;
ACTS|18|28|vehementer enim Iudaeos revincebat publice, ostendens per Scripturas esse Christum Iesum.
ACTS|19|1|Factum est autem, cum Apollo esset Corinthi, ut Paulus, peragratis superioribus partibus, veniret Ephesum et inveniret quosdam discipulos;
ACTS|19|2|dixitque ad eos: " Si Spiritum Sanctum accepistis credentes? ". At illi ad eum: " Sed neque, si Spiritus Sanctus est, audivimus ".
ACTS|19|3|Ille vero ait: " In quo ergo baptizati estis? ". Qui dixerunt: " In Ioannis baptismate ".
ACTS|19|4|Dixit autem Paulus: " Ioannes baptizavit baptisma paenitentiae, populo dicens in eum, qui venturus esset post ipsum ut crederent, hoc est in Iesum ".
ACTS|19|5|His auditis, baptizati sunt in nomine Domini Iesu;
ACTS|19|6|et cum imposuisset illis manus Paulus, venit Spiritus Sanctus super eos, et loquebantur linguis et prophetabant.
ACTS|19|7|Erant autem omnes viri fere duodecim.
ACTS|19|8|Introgressus autem synagogam cum fiducia loquebatur per tres menses disputans et suadens de regno Dei.
ACTS|19|9|Cum autem quidam indurarentur et non crederent maledicentes viam coram multitudine, discedens ab eis segregavit discipulos, cotidie disputans in schola Tyranni.
ACTS|19|10|Hoc autem factum est per biennium, ita ut omnes, qui habitabant in Asia, audirent verbum Domini, Iudaei atque Graeci.
ACTS|19|11|Virtutesque non quaslibet Deus faciebat per manus Pauli,
ACTS|19|12|ita ut etiam super languidos deferrentur a corpore eius sudaria vel semicinctia, et recederent ab eis languores, et spiritus nequam egrederentur.
ACTS|19|13|Tentaverunt autem quidam et de circumeuntibus Iudaeis exorcistis invocare super eos, qui habebant spiritus malos, nomen Domini Iesu dicentes: " Adiuro vos per Iesum, quem Paulus praedicat ".
ACTS|19|14|Erant autem cuiusdam Scevae Iudaei principis sacerdotum septem filii, qui hoc faciebant.
ACTS|19|15|Respondens autem spiritus nequam dixit eis: " Iesum novi et Paulum scio; vos autem qui estis? ".
ACTS|19|16|Et insiliens homo in eos, in quo erat spiritus malus, dominatus amborum invaluit contra eos, ita ut nudi et vulnerati effugerent de domo illa.
ACTS|19|17|Hoc autem notum factum est omnibus Iudaeis atque Graecis, qui habitabant Ephesi, et cecidit timor super omnes illos, et magnificabatur nomen Domini Iesu.
ACTS|19|18|Multique credentium veniebant confitentes et annuntiantes actus suos.
ACTS|19|19|Multi autem ex his, qui fuerant curiosa sectati, conferentes libros combusserunt coram omnibus; et computaverunt pretia illorum et invenerunt argenti quinquaginta milia.
ACTS|19|20|Ita fortiter verbum Domini crescebat et convalescebat.
ACTS|19|21|His autem expletis, proposuit Paulus in Spiritu, transita Macedonia et Achaia, ire Hierosolymam, dicens: " Postquam fuero ibi, oportet me et Romam videre ".
ACTS|19|22|Mittens autem in Macedoniam duos ex ministrantibus sibi, Timotheum et Erastum, ipse remansit ad tempus in Asia.
ACTS|19|23|Facta est autem in illo tempore turbatio non minima de via.
ACTS|19|24|Demetrius enim quidam nomine, argentarius, faciens aedes argenteas Dianae praestabat artificibus non modicum quaestum;
ACTS|19|25|quos congregans et eos, qui eiusmodi erant opifices, dixit: " Viri, scitis quia de hoc artificio acquisitio est nobis;
ACTS|19|26|et videtis et auditis quia non solum Ephesi, sed paene totius Asiae Paulus hic suadens avertit multam turbam dicens quoniam non sunt dii, qui manibus fiunt.
ACTS|19|27|Non solum autem haec periclitatur nobis pars in redargutionem venire, sed et magnae deae Dianae templum in nihilum reputari, et destrui incipiet maiestas eius, quam tota Asia et orbis colit ".
ACTS|19|28|His auditis, repleti sunt ira et clamabant dicentes: " Magna Diana Ephesiorum! ";
ACTS|19|29|et impleta est civitas confusione, et impetum fecerunt uno animo in theatrum, rapto Gaio et Aristarcho Macedonibus, comitibus Pauli.
ACTS|19|30|Paulo autem volente intrare in populum, non permiserunt discipuli;
ACTS|19|31|quidam autem de Asiarchis, qui erant amici eius, miserunt ad eum rogantes, ne se daret in theatrum.
ACTS|19|32|Alii autem aliud clamabant; erat enim ecclesia confusa, et plures nesciebant qua ex causa convenissent.
ACTS|19|33|De turba autem instruxerunt Alexandrum, propellentibus eum Iudaeis; Alexander ergo, manu silentio postulato, volebat rationem reddere populo.
ACTS|19|34|Quem ut cognoverunt Iudaeum esse, vox facta est una omnium quasi per horas duas clamantium: " Magna Diana Ephesiorum ".
ACTS|19|35|Et cum sedasset scriba turbam, dixit: " Viri Ephesii, quis enim est hominum, qui nesciat Ephesiorum civitatem cultricem esse magnae Dianae et simulacri a Iove delapsi?
ACTS|19|36|Cum ergo his contradici non possit, oportet vos sedatos esse et nihil temere agere.
ACTS|19|37|Adduxistis enim homines istos neque sacrilegos neque blasphemantes deam nostram.
ACTS|19|38|Quod si Demetrius et, qui cum eo sunt, artifices habent adversus aliquem causam, conventus forenses aguntur, et proconsules sunt: accusent invicem.
ACTS|19|39|Si quid autem ulterius quaeritis, in legitima ecclesia poterit absolvi.
ACTS|19|40|Nam et periclitamur argui seditionis hodiernae, cum nullus obnoxius sit, de quo non possimus reddere rationem concursus istius ". Et cum haec dixisset, dimisit ecclesiam.
ACTS|20|1|Postquam autem cessavit tumultus, accersitis Paulus discipulis et exhortatus eos, valedixit et profectus est, ut iret in Macedoniam.
ACTS|20|2|Cum autem perambulasset partes illas et exhortatus eos fuisset multo sermone, venit ad Graeciam;
ACTS|20|3|cumque fecisset menses tres, factae sunt illi insidiae a Iudaeis navigaturo in Syriam, habuitque consilium, ut reverteretur per Macedoniam.
ACTS|20|4|Comitabatur autem eum Sopater Pyrrhi Beroeensis, Thessalonicensium vero Aristarchus et Secundus et Gaius Derbeus et Timotheus, Asiani vero Tychicus et Trophimus.
ACTS|20|5|Hi cum praecessissent, sustinebant nos Troade;
ACTS|20|6|nos vero navigavimus post dies Azymorum a Philippis et venimus ad eos Troadem in diebus quinque, ubi demorati sumus diebus septem.
ACTS|20|7|In una autem sabbatorum, cum convenissemus ad frangendum panem, Paulus disputabat eis, profecturus in crastinum, protraxitque sermonem usque in mediam noctem.
ACTS|20|8|Erant autem lampades copiosae in cenaculo, ubi eramus congregati;
ACTS|20|9|sedens autem quidam adulescens nomine Eutychus super fenestram, cum mergeretur somno gravi, disputante diutius Paulo, eductus somno cecidit de tertio cenaculo deorsum et sublatus est mortuus.
ACTS|20|10|Cum descendisset autem Paulus, incubuit super eum et complexus dixit: " Nolite turbari, anima enim ipsius in eo est! ".
ACTS|20|11|Ascendens autem frangensque panem et gustans satisque allocutus usque in lucem, sic profectus est.
ACTS|20|12|Adduxerunt autem puerum viventem et consolati sunt non minime.
ACTS|20|13|Nos autem praecedentes navi enavigavimus in Asson, inde suscepturi Paulum; sic enim disposuerat volens ipse per terram iter facere.
ACTS|20|14|Cum autem convenisset nos in Asson, assumpto eo, venimus Mitylenen
ACTS|20|15|et inde navigantes sequenti die pervenimus contra Chium et alia applicuimus Samum et sequenti venimus Miletum.
ACTS|20|16|Proposuerat enim Paulus transnavigare Ephesum, ne qua mora illi fieret in Asia; festinabat enim, si possibile sibi esset, ut diem Pentecosten faceret Hierosolymis.
ACTS|20|17|A Mileto autem mittens Ephesum convocavit presbyteros ecclesiae.
ACTS|20|18|Qui cum venissent ad eum, dixit eis: " Vos scitis a prima die, qua ingressus sum in Asiam, qualiter vobiscum per omne tempus fuerim,
ACTS|20|19|serviens Domino cum omni humilitate et lacrimis et tentationibus, quae mihi acciderunt in insidiis Iudaeorum;
ACTS|20|20|quomodo nihil subtraxerim utilium, quominus annuntiarem vobis et docerem vos publice et per domos,
ACTS|20|21|testificans Iudaeis atque Graecis in Deum paenitentiam et fidem in Dominum nostrum Iesum.
ACTS|20|22|Et nunc ecce alligatus ego Spiritu vado in Ierusalem, quae in ea eventura sint mihi ignorans,
ACTS|20|23|nisi quod Spiritus Sanctus per omnes civitates protestatur mihi dicens quoniam vincula et tribulationes me manent.
ACTS|20|24|Sed nihili facio animam meam pretiosam mihi, dummodo consummem cursum meum et ministerium, quod accepi a Domino Iesu, testificari evangelium gratiae Dei.
ACTS|20|25|Et nunc ecce ego scio quia amplius non videbitis faciem meam vos omnes, per quos transivi praedicans regnum;
ACTS|20|26|quapropter contestor vos hodierna die, quia mundus sum a sanguine omnium;
ACTS|20|27|non enim subterfugi, quominus annuntiarem omne consilium Dei vobis.
ACTS|20|28|Attendite vobis et universo gregi, in quo vos Spiritus Sanctus posuit episcopos, pascere ecclesiam Dei, quam acquisivit sanguine suo.
ACTS|20|29|Ego scio quoniam intrabunt post discessionem meam lupi graves in vos non parcentes gregi;
ACTS|20|30|et ex vobis ipsis exsurgent viri loquentes perversa, ut abstrahant discipulos post se.
ACTS|20|31|Propter quod vigilate, memoria retinentes quoniam per triennium nocte et die non cessavi cum lacrimis monens unumquemque vestrum.
ACTS|20|32|Et nunc commendo vos Deo et verbo gratiae ipsius, qui potens est aedificare et dare hereditatem in sanctificatis omnibus.
ACTS|20|33|Argentum aut aurum aut vestem nullius concupivi;
ACTS|20|34|ipsi scitis quoniam ad ea, quae mihi opus erant et his, qui mecum sunt, ministraverunt manus istae.
ACTS|20|35|Omnia ostendi vobis quoniam sic laborantes oportet suscipere infirmos, ac meminisse verborum Domini Iesu, quoniam ipse dixit: "Beatius est magis dare quam accipere!" ".
ACTS|20|36|Et cum haec dixisset, positis genibus suis, cum omnibus illis oravit.
ACTS|20|37|Magnus autem fletus factus est omnium; et procumbentes super collum Pauli osculabantur eum
ACTS|20|38|dolentes maxime in verbo, quod dixerat, quoniam amplius faciem eius non essent visuri. Et deducebant eum ad navem.
ACTS|21|1|Cum autem factum esset, ut navigaremus abstracti ab eis, recto cursu venimus Cho et sequenti die Rhodum et inde Patara;
ACTS|21|2|et cum invenissemus navem transfretantem in Phoenicen, ascendentes navigavimus.
ACTS|21|3|Cum paruissemus autem Cypro, et relinquentes eam ad sinistram navigabamus in Syriam et venimus Tyrum, ibi enim navis erat expositura onus.
ACTS|21|4|Inventis autem discipulis, mansimus ibi diebus septem; qui Paulo dicebant per Spiritum, ne iret Hierosolymam.
ACTS|21|5|Et explicitis diebus, profecti ibamus, deducentibus nos omnibus cum uxoribus et filiis usque foras civitatem; et positis genibus in litore orantes,
ACTS|21|6|valefecimus invicem et ascendimus in navem; illi autem redierunt in sua.
ACTS|21|7|Nos vero, navigatione explicita, a Tyro devenimus Ptolemaida et, salutatis fratribus, mansimus die una apud illos.
ACTS|21|8|Alia autem die profecti venimus Caesaream et intrantes in domum Philippi evangelistae, qui erat de septem, mansimus apud eum.
ACTS|21|9|Huic autem erant filiae quattuor virgines prophetantes.
ACTS|21|10|Et cum moraremur plures dies, supervenit quidam a Iudaea propheta nomine Agabus;
ACTS|21|11|is cum venisset ad nos et tulisset zonam Pauli, alligans sibi pedes et manus dixit: " Haec dicit Spiritus Sanctus: Virum, cuius est zona haec, sic alligabunt in Ierusalem Iudaei et tradent in manus gentium ".
ACTS|21|12|Quod cum audissemus, rogabamus nos et, qui loci illius erant, ne ipse ascenderet Ierusalem.
ACTS|21|13|Tunc respondit Paulus: " Quid facitis flentes et affligentes cor meum? Ego enim non solum alligari sed et mori in Ierusalem paratus sum propter nomen Domini Iesu ".
ACTS|21|14|Et cum ei suadere non possemus, quievimus dicentes: " Domini voluntas fiat! ".
ACTS|21|15|Post dies autem istos praeparati ascendebamus Hierosolymam;
ACTS|21|16|venerunt autem et ex discipulis a Caesarea nobiscum adducentes apud quem hospitaremur, Mnasonem quendam Cyprium, antiquum discipulum.
ACTS|21|17|Et cum venissemus Hierosolymam, libenter exceperunt nos fratres.
ACTS|21|18|Sequenti autem die introibat Paulus nobiscum ad Iacobum, omnesque collecti sunt presbyteri.
ACTS|21|19|Quos cum salutasset, narrabat per singula, quae fecisset Deus in gentibus per ministerium ipsius.
ACTS|21|20|At illi cum audissent, glorificabant Deum dixeruntque ei: " Vides, frater, quot milia sint in Iudaeis, qui crediderunt, et omnes aemulatores sunt legis;
ACTS|21|21|audierunt autem de te quia discessionem doceas a Moyse omnes, qui per gentes sunt, Iudaeos, dicens non debere circumcidere eos filios suos neque secundum consuetudines ambulare.
ACTS|21|22|Quid ergo est? Utique audient te supervenisse.
ACTS|21|23|Hoc ergo fac, quod tibi dicimus. Sunt nobis viri quattuor votum habentes super se;
ACTS|21|24|his assumptis, sanctifica te cum illis et impende pro illis, ut radant capita, et scient omnes quia, quae de te audierunt, nihil sunt, sed ambulas et ipse custodiens legem.
ACTS|21|25|De his autem, qui crediderunt, gentibus nos scripsimus iudicantes, ut abstineant ab idolothyto et sanguine et suffocato et fornicatione ".
ACTS|21|26|Tunc Paulus, assumptis viris, postera die purificatus cum illis intravit in templum annuntians expletionem dierum purificationis, donec offerretur pro unoquoque eorum oblatio.
ACTS|21|27|Dum autem septem dies consummarentur, hi, qui de Asia erant, Iudaei cum vidissent eum in templo, concitaverunt omnem turbam et iniecerunt ei manus
ACTS|21|28|clamantes: " Viri Israelitae, adiuvate! Hic est homo, qui adversus populum et legem et locum hunc omnes ubique docens, insuper et Graecos induxit in templum et polluit sanctum locum istum ".
ACTS|21|29|Viderant enim Trophimum Ephesium in civitate cum ipso, quem aestimabant quoniam in templum induxisset Paulus.
ACTS|21|30|Commotaque est civitas tota, et facta est concursio populi, et apprehendentes Paulum trahebant eum extra templum, et statim clausae sunt ianuae.
ACTS|21|31|Quaerentibus autem eum occidere, nuntiatum est tribuno cohortis quia tota confunditur Ierusalem,
ACTS|21|32|qui statim, assumptis militibus et centurionibus, decucurrit ad illos; qui cum vidissent tribunum et milites, cessaverunt percutere Paulum.
ACTS|21|33|Tunc accedens tribunus apprehendit eum et iussit alligari catenis duabus et interrogabat quis esset et quid fecisset.
ACTS|21|34|Alii autem aliud clamabant in turba; et cum non posset certum cognoscere prae tumultu, iussit duci eum in castra.
ACTS|21|35|Et cum venisset ad gradus, contigit ut portaretur a militibus propter vim turbae;
ACTS|21|36|sequebatur enim multitudo populi clamantes: " Tolle eum! ".
ACTS|21|37|Et cum coepisset induci in castra, Paulus dicit tribuno: " Si licet mihi loqui aliquid ad te? ". Qui dixit: " Graece nosti?
ACTS|21|38|Nonne tu es Aegyptius, qui ante hos dies tumultum concitasti et eduxisti in desertum quattuor milia virorum sicariorum? ".
ACTS|21|39|Et dixit Paulus: " Ego homo sum quidem Iudaeus a Tarso Ciliciae, non ignotae civitatis municeps; rogo autem te, permitte mihi loqui ad populum.
ACTS|21|40|Et cum ille permisisset, Paulus stans in gradibus annuit manu ad plebem et, magno silentio facto, allocutus est Hebraea lingua dicens:
ACTS|22|1|" Viri fratres et patres, audi te a me, quam ad vos nunc reddo, rationem.
ACTS|22|2|Cum audissent autem quia Hebraea lingua loquebatur ad illos, magis praestiterunt silentium. Et dixit:
ACTS|22|3|" Ego sum vir Iudaeus, natus Tarso Ciliciae, enutritus autem in ista civitate, secus pedes Gamaliel eruditus iuxta veritatem paternae legis, aemulator Dei, sicut et vos omnes estis hodie.
ACTS|22|4|Qui hanc viam persecutus sum usque ad mortem, alligans et tradens in custodias viros ac mulieres,
ACTS|22|5|sicut et princeps sacerdotum testimonium mihi reddit et omne concilium; a quibus et epistulas accipiens ad fratres, Damascum pergebam, ut adducerem et eos, qui ibi essent, vinctos in Ierusalem, uti punirentur.
ACTS|22|6|Factum est autem, eunte me et appropinquante Damasco, circa mediam diem subito de caelo circumfulsit me lux copiosa;
ACTS|22|7|et decidi in terram et audivi vocem dicentem mihi: "Saul, Saul, quid me persequeris?".
ACTS|22|8|Ego autem respondi: "Quis es, Domine?". Dixitque ad me: "Ego sum Iesus Nazarenus, quem tu persequeris".
ACTS|22|9|Et, qui mecum erant, lumen quidem viderunt, vocem autem non audierunt eius, qui loquebatur mecum.
ACTS|22|10|Et dixi: "Quid faciam, Domine?". Dominus autem dixit ad me: "Surgens vade Damascum, et ibi tibi dicetur de omnibus, quae statutum est tibi, ut faceres".
ACTS|22|11|Et cum non viderem prae claritate luminis illius, ad manum deductus a comitibus veni Damascum.
ACTS|22|12|Ananias autem quidam vir religiosus secundum legem, testimonium habens ab omnibus habitantibus Iudaeis,
ACTS|22|13|veniens ad me et astans dixit mihi: "Saul frater, respice!". Et ego eadem hora respexi in eum.
ACTS|22|14|At ille dixit: "Deus patrum nostrorum praeordinavit te, ut cognosceres voluntatem eius et videres Iustum et audires vocem ex ore eius,
ACTS|22|15|quia eris testis illi ad omnes homines eorum, quae vidisti et audisti.
ACTS|22|16|Et nunc quid moraris? Exsurgens baptizare et ablue peccata tua, invocato nomine ipsius".
ACTS|22|17|Factum est autem, revertenti mihi in Ierusalem et oranti in templo fieri me in stupore mentis
ACTS|22|18|et videre illum dicentem mihi: "Festina et exi velociter ex Ierusalem, quoniam non recipient testimonium tuum de me".
ACTS|22|19|Et ego dixi: "Domine, ipsi sciunt quia ego eram concludens in carcerem et caedens per synagogas eos, qui credebant in te;
ACTS|22|20|et cum funderetur sanguis Stephani testis tui, et ipse astabam et consentiebam et custodiebam vestimenta interficientium illum".
ACTS|22|21|Et dixit ad me: "Vade, quoniam ego in nationes longe mittam te" ".
ACTS|22|22|Audiebant autem eum usque ad hoc verbum et levaverunt vocem suam dicentes: " Tolle de terra eiusmodi, non enim fas est eum vivere! ".
ACTS|22|23|Vociferantibus autem eis et proicientibus vestimenta sua et pulverem iactantibus in aerem,
ACTS|22|24|iussit tribunus induci eum in castra dicens flagellis eum interrogari, ut sciret propter quam causam sic acclamarent ei.
ACTS|22|25|Et cum astrinxissent eum loris, dixit astanti centurioni Paulus: " Si hominem Romanum et indemnatum licet vobis flagellare? ".
ACTS|22|26|Quo audito, centurio accedens ad tribunum nuntiavit dicens: " Quid acturus es? Hic enim homo Romanus est ".
ACTS|22|27|Accedens autem tribunus dixit illi: " Dic mihi, tu Romanus es? ". At ille dixit: " Etiam ".
ACTS|22|28|Et respondit tribunus: " Ego multa summa civitatem hanc consecutus sum. Et Paulus ait: " Ego autem et natus sum ".
ACTS|22|29|Protinus ergo discesserunt ab illo, qui eum interrogaturi erant; tribunus quoque timuit, postquam rescivit quia Romanus esset, et quia alligasset eum.
ACTS|22|30|Postera autem die, volens scire diligenter qua ex causa accusaretur a Iudaeis, solvit eum et iussit principes sacerdotum convenire et omne concilium et producens Paulum statuit coram illis.
ACTS|23|1|Intendens autem concilium Paulus ait: " Viri fratres, ego omni conscientia bona conversatus sum ante Deum usque in hodiernum diem ".
ACTS|23|2|Princeps autem sacerdotum Ananias praecepit astantibus sibi percutere os eius.
ACTS|23|3|Tunc Paulus ad eum dixit: " Percutiet te Deus, paries dealbate! Et tu sedes iudicans me secundum legem et contra legem iubes me percuti? ".
ACTS|23|4|Et, qui astabant, dixerunt: " Summum sacerdotem Dei maledicis?".
ACTS|23|5|Dixit autem Paulus: " Nesciebam, fratres, quia princeps est sacerdotum; scriptum est enim: "Principem populi tui non maledices" ".
ACTS|23|6|Sciens autem Paulus quia una pars esset sadducaeorum, et altera pharisaeorum, exclamabat in concilio: " Viri fratres, ego pharisaeus sum, filius pharisaeorum; de spe et resurrectione mortuorum ego iudicor ".
ACTS|23|7|Et cum haec diceret, facta est dissensio inter pharisaeos et sadducaeos; et divisa est multitudo.
ACTS|23|8|Sadducaei enim dicunt non esse resurrectionem neque angelum neque spiritum; pharisaei autem utrumque confitentur.
ACTS|23|9|Factus est autem clamor magnus; et surgentes scribae quidam partis pharisaeorum pugnabant dicentes: " Nihil mali invenimus in homine isto: quod si spiritus locutus est ei aut angelus ";
ACTS|23|10|et cum magna dissensio facta esset, timens tribunus ne discerperetur Paulus ab ipsis, iussit milites descendere, ut raperent eum de medio eorum ac deducerent in castra.
ACTS|23|11|Sequenti autem nocte, assistens ei Dominus ait: " Constans esto! Sicut enim testificatus es, quae sunt de me, in Ierusalem, sic te oportet et Romae testificari ".
ACTS|23|12|Facta autem die, faciebant concursum Iudaei et devoverunt se dicentes neque manducaturos neque bibituros, donec occiderent Paulum.
ACTS|23|13|Erant autem plus quam quadraginta, qui hanc coniurationem fecerant;
ACTS|23|14|qui accedentes ad principes sacerdotum et seniores dixerunt: " Devotione devovimus nos nihil gustaturos, donec occidamus Paulum.
ACTS|23|15|Nunc ergo vos notum facite tribuno cum concilio, ut producat illum ad vos, tamquam aliquid certius cognituri de eo; nos vero, priusquam appropiet, parati sumus interficere illum ".
ACTS|23|16|Quod cum audisset filius sororis Pauli insidias, venit et intravit in castra nuntiavitque Paulo.
ACTS|23|17|Vocans autem Paulus ad se unum ex centurionibus ait: " Adulescentem hunc perduc ad tribunum, habet enim aliquid indicare illi ".
ACTS|23|18|Et ille quidem assumens eum duxit ad tribunum et ait: " Vinctus Paulus vocans rogavit me hunc adulescentem perducere ad te, habentem aliquid loqui tibi ".
ACTS|23|19|Apprehendens autem tribunus manum illius, secessit cum eo seorsum et interrogabat: " Quid est, quod habes indicare mihi? ".
ACTS|23|20|Ille autem dixit: " Iudaei constituerunt rogare te, ut crastina die Paulum producas in concilium, quasi aliquid certius inquisiturum sit de illo.
ACTS|23|21|Tu ergo ne credideris illis; insidiantur enim ei ex eis viri amplius quadraginta, qui se devoverunt non manducare neque bibere, donec interficiant eum; et nunc parati sunt exspectantes promissum tuum ".
ACTS|23|22|Tribunus igitur dimisit adulescentem praecipiens, ne cui eloqueretur quoniam " haec nota mihi fecisti ".
ACTS|23|23|Et vocatis duobus centurionibus, dixit: " Parate milites ducentos, ut eant usque Caesaream, et equites septuaginta et lancearios ducentos, a tertia hora noctis,
ACTS|23|24|et iumenta praeparate ", ut imponentes Paulum salvum perducerent ad Felicem praesidem,
ACTS|23|25|scribens epistulam habentem formam hanc:
ACTS|23|26|" Claudius Lysias optimo praesidi Felici salutem.
ACTS|23|27|Virum hunc comprehensum a Iudaeis et incipientem interfici ab eis, superveniens cum exercitu eripui, cognito quia Romanus est.
ACTS|23|28|Volensque scire causam, propter quam accusabant illum, deduxi in concilium eorum;
ACTS|23|29|quem inveni accusari de quaestionibus legis ipsorum, nihil vero dignum morte aut vinculis habentem crimen.
ACTS|23|30|Et cum mihi perlatum esset de insidiis, quae in virum pararentur, confestim misi ad te denuntians et accusatoribus, ut dicant adversum eum apud te ".
ACTS|23|31|Milites ergo, secundum praeceptum sibi assumentes Paulum, duxerunt per noctem in Antipatridem;
ACTS|23|32|et postera die, dimissis equitibus, ut abirent cum eo, reversi sunt ad castra.
ACTS|23|33|Qui cum venissent Caesaream et tradidissent epistulam praesidi, statuerunt ante illum et Paulum.
ACTS|23|34|Cum legisset autem et interrogasset de qua provincia esset, et cognoscens quia de Cilicia:
ACTS|23|35|" Audiam te, inquit, cum et accusatores tui venerint "; iussitque in praetorio Herodis custodiri eum.
ACTS|24|1|Post quinque autem dies, descendit princeps sacerdo tum Ananias cum senioribus quibusdam et Tertullo quodam oratore, qui adierunt praesidem adversus Paulum.
ACTS|24|2|Et citato eo, coepit accusare Tertullus dicens: " Cum in multa pace agamus per te, et multa corrigantur genti huic per tuam providentiam,
ACTS|24|3|semper et ubique suscipimus, optime Felix, cum omni gratiarum actione.
ACTS|24|4|Ne diutius autem te protraham, oro, breviter audias nos pro tua clementia.
ACTS|24|5|Invenimus enim hunc hominem pestiferum et concitantem seditiones omnibus Iudaeis, qui sunt in universo orbe, et auctorem seditionis sectae Nazarenorum,
ACTS|24|6|qui etiam templum violare conatus est, quem et apprehendimus,
ACTS|24|7|()
ACTS|24|8|a quo poteris ipse diiudicans de omnibus istis cognoscere, de quibus nos accusamus eum ".
ACTS|24|9|Adiecerunt autem et Iudaei dicentes haec ita se habere.
ACTS|24|10|Respondit autem Paulus, annuente sibi praeside dicere: " Ex multis annis esse te iudicem genti huic sciens bono animo de causa mea rationem reddam,
ACTS|24|11|cum possis cognoscere quia non plus sunt dies mihi quam duodecim, ex quo ascendi adorare in Ierusalem,
ACTS|24|12|et neque in templo invenerunt me cum aliquo disputantem aut concursum facientem turbae neque in synagogis neque in civitate,
ACTS|24|13|neque probare possunt tibi, de quibus nunc accusant me.
ACTS|24|14|Confiteor autem hoc tibi, quod secundum viam, quam dicunt haeresim, sic deservio patrio Deo credens omnibus, quae secundum Legem sunt et in Prophetis scripta,
ACTS|24|15|spem habens in Deum, quam et hi ipsi exspectant, resurrectionem futuram iustorum et iniquorum.
ACTS|24|16|In hoc et ipse studeo sine offendiculo conscientiam habere ad Deum et ad homines semper.
ACTS|24|17|Post annos autem plures, eleemosynas facturus in gentem meam veni et oblationes;
ACTS|24|18|in quibus invenerunt me purificatum in templo, non cum turba neque cum tumultu;
ACTS|24|19|quidam autem ex Asia Iudaei, quos oportebat apud te praesto esse et accusare, si quid haberent adversum me;
ACTS|24|20|aut hi ipsi dicant quid invenerint iniquitatis, cum starem in concilio,
ACTS|24|21|nisi de una hac voce, qua clamavi inter eos stans: De resurrectione mortuorum ego iudicor hodie apud vos! ".
ACTS|24|22|Distulit autem illos Felix certissime sciens ea, quae de hac via sunt, dicens: " Cum tribunus Lysias descenderit, cognoscam causam vestram ",
ACTS|24|23|iubens centurioni custodiri eum et habere mitigationem, nec quemquam prohibere de suis ministrare ei.
ACTS|24|24|Post aliquot autem dies, adveniens Felix cum Drusilla uxore sua, quae erat Iudaea, vocavit Paulum et audivit ab eo de fide, quae est in Christum Iesum.
ACTS|24|25|Disputante autem illo de iustitia et continentia et de iudicio futuro, timefactus Felix respondit: " Quod nunc attinet, vade; tempore autem opportuno accersiam te ",
ACTS|24|26|simul et sperans quia pecunia daretur sibi a Paulo; propter quod et frequenter accersiens eum loquebatur cum eo.
ACTS|24|27|Biennio autem expleto, accepit successorem Felix Porcium Festum; volensque gratiam praestare Iudaeis, Felix reliquit Paulum vinctum.
ACTS|25|1|Festus ergo cum venisset in provinciam, post triduum ascendit Hierosolymam a Caesarea;
ACTS|25|2|adieruntque eum principes sacerdotum et primi Iudaeorum adversus Paulum, et rogabant eum
ACTS|25|3|postulantes gratiam adversum eum, ut iuberet perduci eum in Ierusalem, insidias tendentes, ut eum interficerent in via.
ACTS|25|4|Festus igitur respondit servari Paulum in Caesarea, se autem maturius profecturum:
ACTS|25|5|" Qui ergo in vobis, ait, potentes sunt, descendentes simul, si quod est in viro crimen, accusent eum ".
ACTS|25|6|Demoratus autem inter eos dies non amplius quam octo aut decem, descendit Caesaream; et altera die sedit pro tribunali et iussit Paulum adduci.
ACTS|25|7|Qui cum perductus esset, circumsteterunt eum, qui ab Hierosolyma descenderant, Iudaei, multas et graves causas obicientes, quas non poterant probare,
ACTS|25|8|Paulo rationem reddente: " Neque in legem Iudaeorum neque in templum neque in Caesarem quidquam peccavi ".
ACTS|25|9|Festus autem volens Iudaeis gratiam praestare, respondens Paulo dixit: " Vis Hierosolymam ascendere et ibi de his iudicari apud me? ".
ACTS|25|10|Dixit autem Paulus: " Ad tribunal Caesaris sto, ubi me oportet iudicari. Iudaeis nihil nocui, sicut et tu melius nosti.
ACTS|25|11|Si ergo iniuste egi et dignum morte aliquid feci, non recuso mori; si vero nihil est eorum, quae hi accusant me, nemo potest me illis donare. Caesarem appello! ".
ACTS|25|12|Tunc Festus cum consilio locutus respondit: " Caesarem appellasti; ad Caesarem ibis ".
ACTS|25|13|Et cum dies aliquot transacti essent, Agrippa rex et Berenice descenderunt Caesaream et salutaverunt Festum.
ACTS|25|14|Et cum dies plures ibi demorarentur, Festus regi indicavit de Paulo dicens: " Vir quidam est derelictus a Felice vinctus,
ACTS|25|15|de quo, cum essem Hierosolymis, adierunt me principes sacerdotum et seniores Iudaeorum postulantes adversus illum damnationem;
ACTS|25|16|ad quos respondi, quia non est consuetudo Romanis donare aliquem hominem, priusquam is, qui accusatur, praesentes habeat accusatores locumque defendendi se ab accusatione accipiat.
ACTS|25|17|Cum ergo huc convenissent, sine ulla dilatione sequenti die sedens pro tribunali iussi adduci virum;
ACTS|25|18|de quo, cum stetissent accusatores, nullam causam deferebant, de quibus ego suspicabar malis;
ACTS|25|19|quaestiones vero quasdam de sua superstitione habebant adversus eum et de quodam Iesu defuncto, quem affirmabat Paulus vivere.
ACTS|25|20|Haesitans autem ego de huiusmodi quaestione, dicebam si vellet ire Hierosolymam et ibi iudicari de istis.
ACTS|25|21|Paulo autem appellante, ut servaretur ad Augusti cognitionem, iussi servari eum, donec mittam eum ad Caesarem ".
ACTS|25|22|Agrippa autem ad Festum: " Volebam et ipse hominem audire! ". " Cras, inquit, audies eum ".
ACTS|25|23|Altera autem die, cum venisset Agrippa et Berenice cum multa ambitione, et introissent in auditorium cum tribunis et viris principalibus civitatis, et iubente Festo, adductus est Paulus.
ACTS|25|24|Et dicit Festus: " Agrippa rex et omnes, qui simul adestis nobiscum viri, videtis hunc, de quo omnis multitudo Iudaeorum interpellavit me Hierosolymis et hic, clamantes non oportere eum vivere amplius.
ACTS|25|25|Ego vero comperi nihil dignum eum morte fecisse, ipso autem hoc appellante Augustum, iudicavi mittere.
ACTS|25|26|De quo quid certum scribam domino, non habeo; propter quod produxi eum ad vos et maxime ad te, rex Agrippa, ut, interrogatione facta, habeam quid scribam;
ACTS|25|27|sine ratione enim mihi videtur mittere vinctum et causas eius non significare ".
ACTS|26|1|Agrippa vero ad Paulum ait: " Permittitur tibi loqui pro temetipso ". Tunc Paulus, extenta manu, coepit rationem reddere:
ACTS|26|2|" De omnibus, quibus accusor a Iudaeis, rex Agrippa, aestimo me beatum, apud te cum sim defensurus me hodie,
ACTS|26|3|maxime te sciente omnia, quae apud Iudaeos sunt consuetudines et quaestiones; propter quod, obsecro, patienter me audias.
ACTS|26|4|Et quidem vitam meam a iuventute, quae ab initio fuit in gente mea et in Hierosolymis, noverunt omnes Iudaei;
ACTS|26|5|praescientes me ab initio, si velint testimonium perhibere, quoniam secundum diligentissimam sectam nostrae religionis vixi pharisaeus.
ACTS|26|6|Et nunc propter spem eius, quae ad patres nostros repromissionis facta est a Deo, sto iudicio subiectus,
ACTS|26|7|in quam duodecim tribus nostrae cum perseverantia nocte ac die deservientes sperant devenire; de qua spe accusor a Iudaeis, rex!
ACTS|26|8|Quid incredibile iudicatur apud vos, si Deus mortuos suscitat?
ACTS|26|9|Et ego quidem existimaveram me adversus nomen Iesu Nazareni debere multa contraria agere;
ACTS|26|10|quod et feci Hierosolymis, et multos sanctorum ego in carceribus inclusi, a principibus sacerdotum potestate accepta, et cum occiderentur, detuli sententiam;
ACTS|26|11|et per omnes synagogas frequenter puniens eos compellebam blasphemare, et abundantius insaniens in eos persequebar usque in exteras civitates.
ACTS|26|12|In quibus, dum irem Damascum cum potestate et permissu principum sacerdotum,
ACTS|26|13|die media in via vidi, rex, de caelo supra splendorem solis circumfulgens me lumen et eos, qui mecum simul ibant;
ACTS|26|14|omnesque nos cum decidissemus in terram, audivi vocem loquentem mihi Hebraica lingua: "Saul, Saul, quid me persequeris? Durum est tibi contra stimulum calcitrare".
ACTS|26|15|Ego autem dixi: "Quis es, Domine?". Dominus autem dixit: "Ego sum Iesus, quem tu persequeris.
ACTS|26|16|Sed exsurge et sta super pedes tuos; ad hoc enim apparui tibi, ut constituam te ministrum et testem eorum, quae vidisti, et eorum, quibus apparebo tibi,
ACTS|26|17|eripiens te de populo et de gentibus, in quas ego mitto te
ACTS|26|18|aperire oculos eorum, ut convertantur a tenebris ad lucem et de potestate Satanae ad Deum, ut accipiant remissionem peccatorum et sortem inter sanctificatos per fidem, quae est in me".
ACTS|26|19|Unde, rex Agrippa, non fui incredulus caelestis visionis,
ACTS|26|20|sed his, qui sunt Damasci primum et Hierosolymis, et in omnem regionem Iudaeae et gentibus annuntiabam, ut paenitentiam agerent et converterentur ad Deum digna paenitentiae opera facientes.
ACTS|26|21|Hac ex causa me Iudaei, cum essem in templo comprehensum, tentabant interficere.
ACTS|26|22|Auxilium igitur assecutus a Deo usque in hodiernum diem sto testificans minori atque maiori, nihil extra dicens quam ea, quae Prophetae sunt locuti futura esse et Moyses:
ACTS|26|23|si passibilis Christus, si primus ex resurrectione mortuorum lumen annuntiaturus est populo et gentibus ".
ACTS|26|24|Sic autem eo rationem reddente, Festus magna voce dixit: " Insanis, Paule; multae te litterae ad insaniam convertunt! ".
ACTS|26|25|At Paulus: " Non insanio, inquit, optime Feste, sed veritatis et sobrietatis verba eloquor.
ACTS|26|26|Scit enim de his rex, ad quem et audenter loquor; latere enim eum nihil horum arbitror, neque enim in angulo hoc gestum est.
ACTS|26|27|Credis, rex Agrippa, Prophetis? Scio quia credis ".
ACTS|26|28|Agrippa autem ad Paulum: " In modico suades me Christianum fieri! ".
ACTS|26|29|Et Paulus: " Optarem apud Deum et in modico et in magno non tantum te sed et omnes hos, qui audiunt me hodie, fieri tales, qualis et ego sum, exceptis vinculis his! ".
ACTS|26|30|Et exsurrexit rex et praeses et Berenice et qui assidebant eis;
ACTS|26|31|et cum secessissent, loquebantur ad invicem dicentes: " Nihil morte aut vinculis dignum quid facit homo iste ".
ACTS|26|32|Agrippa autem Festo dixit: " Dimitti poterat homo hic, si non appellasset Caesarem ".
ACTS|27|1|Ut autem iudicatum est na vigare nos in Italiam, tradiderunt et Paulum et quosdam alios vinctos centurioni nomine Iulio, cohortis Augustae.
ACTS|27|2|Ascendentes autem navem Hadramyttenam, incipientem navigare circa Asiae loca, sustulimus, perseverante nobiscum Aristarcho Macedone Thessalonicensi;
ACTS|27|3|sequenti autem die, devenimus Sidonem, et humane tractans Iulius Paulum permisit ad amicos ire et curam sui agere.
ACTS|27|4|Et inde cum sustulissemus, subnavigavimus Cypro, propterea quod essent venti contrarii;
ACTS|27|5|et pelagus Ciliciae et Pamphyliae navigantes venimus Myram, quae est Lyciae.
ACTS|27|6|Et ibi inveniens centurio navem Alexandrinam navigantem in Italiam transposuit nos in eam.
ACTS|27|7|Et cum multis diebus tarde navigaremus et vix devenissemus contra Cnidum, prohibente nos vento, subnavigavimus Cretae secundum Salmonem;
ACTS|27|8|et vix iuxta eam navigantes venimus in locum quendam, qui vocatur Boni Portus, cui iuxta erat civitas Lasaea.
ACTS|27|9|Multo autem tempore peracto, et cum iam non esset tuta navigatio, eo quod et ieiunium iam praeterisset, monebat Paulus
ACTS|27|10|dicens eis: " Viri, video quoniam cum iniuria et multo damno non solum oneris et navis sed etiam animarum nostrarum incipit esse navigatio ".
ACTS|27|11|Centurio autem gubernatori et nauclero magis credebat quam his, quae a Paulo dicebantur.
ACTS|27|12|Et cum aptus portus non esset ad hiemandum, plurimi statuerunt consilium enavigare inde, si quo modo possent devenientes Phoenicen hiemare, portum Cretae respicientem ad africum et ad caurum.
ACTS|27|13|Aspirante autem austro, aestimantes propositum se tenere, cum sustulissent, propius legebant Cretam.
ACTS|27|14|Non post multum autem misit se contra ipsam ventus typhonicus, qui vocatur euroaquilo;
ACTS|27|15|cumque arrepta esset navis et non posset conari in ventum, data nave flatibus, ferebamur.
ACTS|27|16|Insulam autem quandam decurrentes, quae vocatur Cauda, potuimus vix obtinere scapham,
ACTS|27|17|qua sublata, adiutoriis utebantur accingentes navem; et timentes, ne in Syrtim inciderent, submisso vase, sic ferebantur.
ACTS|27|18|Valide autem nobis tempestate iactatis, sequenti die iactum fecerunt
ACTS|27|19|et tertia die suis manibus armamenta navis proiecerunt.
ACTS|27|20|Neque sole autem neque sideribus apparentibus per plures dies, et tempestate non exigua imminente, iam auferebatur spes omnis salutis nostrae.
ACTS|27|21|Et cum multa ieiunatio fuisset, tunc stans Paulus in medio eorum dixit: Oportebat quidem, o viri, audito me, non tollere a Creta lucrique facere iniuriam hanc et iacturam.
ACTS|27|22|Et nunc suadeo vobis bono animo esse, nulla enim amissio animae erit ex vobis praeterquam navis;
ACTS|27|23|astitit enim mihi hac nocte angelus Dei, cuius sum ego, cui et deservio,
ACTS|27|24|dicens: "Ne timeas, Paule; Caesari te oportet assistere, et ecce donavit tibi Deus omnes, qui navigant tecum".
ACTS|27|25|Propter quod bono animo estote, viri; credo enim Deo, quia sic erit, quemadmodum dictum est mihi.
ACTS|27|26|In insulam autem quandam oportet nos incidere ".
ACTS|27|27|Sed posteaquam quarta decima nox supervenit, cum ferremur in Hadria, circa mediam noctem suspicabantur nautae apparere sibi aliquam regionem.
ACTS|27|28|Qui submittentes bolidem invenerunt passus viginti; et pusillum inde separati et rursum submittentes invenerunt passus quindecim;
ACTS|27|29|timentes autem, ne in aspera loca incideremus, de puppi mittentes ancoras quattuor optabant diem fieri.
ACTS|27|30|Nautis vero quaerentibus fugere de navi, cum demisissent scapham in mare sub obtentu, quasi a prora inciperent ancoras extendere,
ACTS|27|31|dixit Paulus centurioni et militibus: " Nisi hi in navi manserint, vos salvi fieri non potestis ".
ACTS|27|32|Tunc absciderunt milites funes scaphae et passi sunt eam excidere.
ACTS|27|33|Donec autem lux inciperet fieri, rogabat Paulus omnes sumere cibum dicens: " Quarta decima hodie die exspectantes ieiuni permanetis nihil accipientes;
ACTS|27|34|propter quod rogo vos accipere cibum, hoc enim pro salute vestra est, quia nullius vestrum capillus de capite peribit ".
ACTS|27|35|Et cum haec dixisset et sumpsisset panem, gratias egit Deo in conspectu omnium et, cum fregisset, coepit manducare.
ACTS|27|36|Animaequiores autem facti omnes et ipsi assumpserunt cibum.
ACTS|27|37|Eramus vero universae animae in navi ducentae septuaginta sex.
ACTS|27|38|Et satiati cibo alleviabant navem iactantes triticum in mare.
ACTS|27|39|Cum autem dies factus esset, terram non agnoscebant; sinum vero quendam considerabant habentem litus, in quem cogitabant, si possent, eicere navem.
ACTS|27|40|Et cum ancoras abstulissent, committebant mari simul laxantes iuncturas gubernaculorum et, levato artemone, secundum flatum aurae tendebant ad litus.
ACTS|27|41|Et cum incidissent in locum dithalassum, impegerunt navem; et prora quidem fixa manebat immobilis, puppis vero solvebatur a vi fluctuum.
ACTS|27|42|Militum autem consilium fuit, ut custodias occiderent, ne quis, cum enatasset, effugeret;
ACTS|27|43|centurio autem volens servare Paulum prohibuit eos a consilio iussitque eos, qui possent natare, mittere se primos et ad terram exire
ACTS|27|44|et ceteros, quosdam in tabulis, quosdam vero super ea, quae de navi essent; et sic factum est ut omnes evaderent ad terram.
ACTS|28|1|Et cum evasissemus, tunc cognovimus quia Melita in sula vocatur.
ACTS|28|2|Barbari vero praestabant non modicam humanitatem nobis; accensa enim pyra, suscipiebant nos omnes propter imbrem, qui imminebat, et frigus.
ACTS|28|3|Cum congregasset autem Paulus sarmentorum aliquantam multitudinem et imposuisset super ignem, vipera, a calore cum processisset, invasit manum eius.
ACTS|28|4|Ut vero viderunt barbari pendentem bestiam de manu eius, ad invicem dicebant: " Utique homicida est homo hic, qui cum evaserit de mari, Ultio non permisit vivere ".
ACTS|28|5|Et ille quidem excutiens bestiam in ignem, nihil mali passus est;
ACTS|28|6|at illi exspectabant eum in tumorem convertendum aut subito casurum et mori. Diu autem illis exspectantibus et videntibus nihil mali in eo fieri, convertentes se dicebant eum esse deum.
ACTS|28|7|In locis autem illis erant praedia principis insulae nomine Publii, qui nos suscipiens triduo benigne hospitio recepit.
ACTS|28|8|Contigit autem patrem Publii febribus et dysenteria vexatum iacere, ad quem Paulus intravit et, cum orasset et imposuisset ei manus, sanavit eum.
ACTS|28|9|Quo facto, et ceteri, qui in insula habebant infirmitates, accedebant et curabantur;
ACTS|28|10|qui etiam multis honoribus nos honoraverunt et navigantibus imposuerunt, quae necessaria erant.
ACTS|28|11|Post menses autem tres, navigavimus in navi Alexandrina, quae in insula hiemaverat, cui erat insigne Castorum.
ACTS|28|12|Et cum venissemus Syracusam, mansimus ibi triduo;
ACTS|28|13|inde solventes devenimus Rhegium. Et post unum diem, superveniente austro, secunda die venimus Puteolos,
ACTS|28|14|ubi, inventis fratribus, rogati sumus manere apud eos dies septem; et sic venimus Romam.
ACTS|28|15|Et inde cum audissent de nobis fratres, occurrerunt nobis usque ad Appii Forum et Tres Tabernas; quos cum vidisset Paulus, gratias agens Deo, accepit fiduciam.
ACTS|28|16|Cum introissemus autem Romam, permissum est Paulo manere sibimet cum custodiente se milite.
ACTS|28|17|Factum est autem, ut post tertium diem convocaret primos Iudaeorum; cumque convenissent dicebat eis: " Ego, viri fratres, nihil adversus plebem faciens aut mores paternos, vinctus ab Hierosolymis traditus sum in manus Romanorum,
ACTS|28|18|qui cum interrogationem de me habuissent, volebant dimittere, eo quod nulla causa esset mortis in me;
ACTS|28|19|contradicentibus autem Iudaeis, coactus sum appellare Caesarem, non quasi gentem meam habens aliquid accusare.
ACTS|28|20|Propter hanc igitur causam rogavi vos videre et alloqui; propter spem enim Israel catena hac circumdatus sum ".
ACTS|28|21|At illi dixerunt ad eum: " Nos neque litteras accepimus de te a Iudaea, neque adveniens aliquis fratrum nuntiavit aut locutus est quid de te malum.
ACTS|28|22|Rogamus autem a te audire quae sentis; nam de secta hac notum est nobis quia ubique ei contradicitur ".
ACTS|28|23|Cum constituissent autem illi diem, venerunt ad eum in hospitium plures, quibus exponebat testificans regnum Dei suadensque eos de Iesu ex Lege Moysis et Prophetis a mane usque ad vesperam.
ACTS|28|24|Et quidam credebant his, quae dicebantur, quidam vero non credebant;
ACTS|28|25|cumque invicem non essent consentientes, discedebant, dicente Paulo unum verbum: " Bene Spiritus Sanctus locutus est per Isaiam prophetam ad patres vestros
ACTS|28|26|dicens:Vade ad populum istum et dic:Auditu audietis et non intellegetis,et videntes videbitis et non perspicietis.
ACTS|28|27|Incrassatum est enim cor populi huius,et auribus graviter audieruntet oculos suos compresserunt,ne forte videant oculiset auribus audiantet corde intellegant et convertantur,et sanabo illos".
ACTS|28|28|Notum ergo sit vobis quoniam gentibus missum est hoc salutare Dei; ipsi et audient! ".
ACTS|28|29|()
ACTS|28|30|Mansit autem biennio toto in suo conducto; et suscipiebat omnes, qui ingrediebantur ad eum,
ACTS|28|31|praedicans regnum Dei et docens quae sunt de Domino Iesu Christo cum omni fiducia sine prohibitione.
