ZECH|1|1|In the eighth month, in the second year of Darius, came the word of the LORD unto Zechariah, the son of Berechiah, the son of Iddo the prophet, saying,
ZECH|1|2|The LORD hath been sore displeased with your fathers.
ZECH|1|3|Therefore say thou unto them, Thus saith the LORD of hosts; Turn ye unto me, saith the LORD of hosts, and I will turn unto you, saith the LORD of hosts.
ZECH|1|4|Be ye not as your fathers, unto whom the former prophets have cried, saying, Thus saith the LORD of hosts; Turn ye now from your evil ways, and from your evil doings: but they did not hear, nor hearken unto me, saith the LORD.
ZECH|1|5|Your fathers, where are they? and the prophets, do they live for ever?
ZECH|1|6|But my words and my statutes, which I commanded my servants the prophets, did they not take hold of your fathers? and they returned and said, Like as the LORD of hosts thought to do unto us, according to our ways, and according to our doings, so hath he dealt with us.
ZECH|1|7|Upon the four and twentieth day of the eleventh month, which is the month Sebat, in the second year of Darius, came the word of the LORD unto Zechariah, the son of Berechiah, the son of Iddo the prophet, saying,
ZECH|1|8|I saw by night, and behold a man riding upon a red horse, and he stood among the myrtle trees that were in the bottom; and behind him were there red horses, speckled, and white.
ZECH|1|9|Then said I, O my lord, what are these? And the angel that talked with me said unto me, I will shew thee what these be.
ZECH|1|10|And the man that stood among the myrtle trees answered and said, These are they whom the LORD hath sent to walk to and fro through the earth.
ZECH|1|11|And they answered the angel of the LORD that stood among the myrtle trees, and said, We have walked to and fro through the earth, and, behold, all the earth sitteth still, and is at rest.
ZECH|1|12|Then the angel of the LORD answered and said, O LORD of hosts, how long wilt thou not have mercy on Jerusalem and on the cities of Judah, against which thou hast had indignation these threescore and ten years?
ZECH|1|13|And the LORD answered the angel that talked with me with good words and comfortable words.
ZECH|1|14|So the angel that communed with me said unto me, Cry thou, saying, Thus saith the LORD of hosts; I am jealous for Jerusalem and for Zion with a great jealousy.
ZECH|1|15|And I am very sore displeased with the heathen that are at ease: for I was but a little displeased, and they helped forward the affliction.
ZECH|1|16|Therefore thus saith the LORD; I am returned to Jerusalem with mercies: my house shall be built in it, saith the LORD of hosts, and a line shall be stretched forth upon Jerusalem.
ZECH|1|17|Cry yet, saying, Thus saith the LORD of hosts; My cities through prosperity shall yet be spread abroad; and the LORD shall yet comfort Zion, and shall yet choose Jerusalem.
ZECH|1|18|Then lifted I up mine eyes, and saw, and behold four horns.
ZECH|1|19|And I said unto the angel that talked with me, What be these? And he answered me, These are the horns which have scattered Judah, Israel, and Jerusalem.
ZECH|1|20|And the LORD shewed me four carpenters.
ZECH|1|21|Then said I, What come these to do? And he spake, saying, These are the horns which have scattered Judah, so that no man did lift up his head: but these are come to fray them, to cast out the horns of the Gentiles, which lifted up their horn over the land of Judah to scatter it.
ZECH|2|1|I lifted up mine eyes again, and looked, and behold a man with a measuring line in his hand.
ZECH|2|2|Then said I, Whither goest thou? And he said unto me, To measure Jerusalem, to see what is the breadth thereof, and what is the length thereof.
ZECH|2|3|And, behold, the angel that talked with me went forth, and another angel went out to meet him,
ZECH|2|4|And said unto him, Run, speak to this young man, saying, Jerusalem shall be inhabited as towns without walls for the multitude of men and cattle therein:
ZECH|2|5|For I, saith the LORD, will be unto her a wall of fire round about, and will be the glory in the midst of her.
ZECH|2|6|Ho, ho, come forth, and flee from the land of the north, saith the LORD: for I have spread you abroad as the four winds of the heaven, saith the LORD.
ZECH|2|7|Deliver thyself, O Zion, that dwellest with the daughter of Babylon.
ZECH|2|8|For thus saith the LORD of hosts; After the glory hath he sent me unto the nations which spoiled you: for he that toucheth you toucheth the apple of his eye.
ZECH|2|9|For, behold, I will shake mine hand upon them, and they shall be a spoil to their servants: and ye shall know that the LORD of hosts hath sent me.
ZECH|2|10|Sing and rejoice, O daughter of Zion: for, lo, I come, and I will dwell in the midst of thee, saith the LORD.
ZECH|2|11|And many nations shall be joined to the LORD in that day, and shall be my people: and I will dwell in the midst of thee, and thou shalt know that the LORD of hosts hath sent me unto thee.
ZECH|2|12|And the LORD shall inherit Judah his portion in the holy land, and shall choose Jerusalem again.
ZECH|2|13|Be silent, O all flesh, before the LORD: for he is raised up out of his holy habitation.
ZECH|3|1|And he shewed me Joshua the high priest standing before the angel of the LORD, and Satan standing at his right hand to resist him.
ZECH|3|2|And the LORD said unto Satan, The LORD rebuke thee, O Satan; even the LORD that hath chosen Jerusalem rebuke thee: is not this a brand plucked out of the fire?
ZECH|3|3|Now Joshua was clothed with filthy garments, and stood before the angel.
ZECH|3|4|And he answered and spake unto those that stood before him, saying, Take away the filthy garments from him. And unto him he said, Behold, I have caused thine iniquity to pass from thee, and I will clothe thee with change of raiment.
ZECH|3|5|And I said, Let them set a fair mitre upon his head. So they set a fair mitre upon his head, and clothed him with garments. And the angel of the LORD stood by.
ZECH|3|6|And the angel of the LORD protested unto Joshua, saying,
ZECH|3|7|Thus saith the LORD of hosts; If thou wilt walk in my ways, and if thou wilt keep my charge, then thou shalt also judge my house, and shalt also keep my courts, and I will give thee places to walk among these that stand by.
ZECH|3|8|Hear now, O Joshua the high priest, thou, and thy fellows that sit before thee: for they are men wondered at: for, behold, I will bring forth my servant the BRANCH.
ZECH|3|9|For behold the stone that I have laid before Joshua; upon one stone shall be seven eyes: behold, I will engrave the graving thereof, saith the LORD of hosts, and I will remove the iniquity of that land in one day.
ZECH|3|10|In that day, saith the LORD of hosts, shall ye call every man his neighbour under the vine and under the fig tree.
ZECH|4|1|And the angel that talked with me came again, and waked me, as a man that is wakened out of his sleep.
ZECH|4|2|And said unto me, What seest thou? And I said, I have looked, and behold a candlestick all of gold, with a bowl upon the top of it, and his seven lamps thereon, and seven pipes to the seven lamps, which are upon the top thereof:
ZECH|4|3|And two olive trees by it, one upon the right side of the bowl, and the other upon the left side thereof.
ZECH|4|4|So I answered and spake to the angel that talked with me, saying, What are these, my lord?
ZECH|4|5|Then the angel that talked with me answered and said unto me, Knowest thou not what these be? And I said, No, my lord.
ZECH|4|6|Then he answered and spake unto me, saying, This is the word of the LORD unto Zerubbabel, saying, Not by might, nor by power, but by my spirit, saith the LORD of hosts.
ZECH|4|7|Who art thou, O great mountain? before Zerubbabel thou shalt become a plain: and he shall bring forth the headstone thereof with shoutings, crying, Grace, grace unto it.
ZECH|4|8|Moreover the word of the LORD came unto me, saying,
ZECH|4|9|The hands of Zerubbabel have laid the foundation of this house; his hands shall also finish it; and thou shalt know that the LORD of hosts hath sent me unto you.
ZECH|4|10|For who hath despised the day of small things? for they shall rejoice, and shall see the plummet in the hand of Zerubbabel with those seven; they are the eyes of the LORD, which run to and fro through the whole earth.
ZECH|4|11|Then answered I, and said unto him, What are these two olive trees upon the right side of the candlestick and upon the left side thereof?
ZECH|4|12|And I answered again, and said unto him, What be these two olive branches which through the two golden pipes empty the golden oil out of themselves?
ZECH|4|13|And he answered me and said, Knowest thou not what these be? And I said, No, my lord.
ZECH|4|14|Then said he, These are the two anointed ones, that stand by the LORD of the whole earth.
ZECH|5|1|Then I turned, and lifted up mine eyes, and looked, and behold a flying roll.
ZECH|5|2|And he said unto me, What seest thou? And I answered, I see a flying roll; the length thereof is twenty cubits, and the breadth thereof ten cubits.
ZECH|5|3|Then said he unto me, This is the curse that goeth forth over the face of the whole earth: for every one that stealeth shall be cut off as on this side according to it; and every one that sweareth shall be cut off as on that side according to it.
ZECH|5|4|I will bring it forth, saith the LORD of hosts, and it shall enter into the house of the thief, and into the house of him that sweareth falsely by my name: and it shall remain in the midst of his house, and shall consume it with the timber thereof and the stones thereof.
ZECH|5|5|Then the angel that talked with me went forth, and said unto me, Lift up now thine eyes, and see what is this that goeth forth.
ZECH|5|6|And I said, What is it? And he said, This is an ephah that goeth forth. He said moreover, This is their resemblance through all the earth.
ZECH|5|7|And, behold, there was lifted up a talent of lead: and this is a woman that sitteth in the midst of the ephah.
ZECH|5|8|And he said, This is wickedness. And he cast it into the midst of the ephah; and he cast the weight of lead upon the mouth thereof.
ZECH|5|9|Then lifted I up mine eyes, and looked, and, behold, there came out two women, and the wind was in their wings; for they had wings like the wings of a stork: and they lifted up the ephah between the earth and the heaven.
ZECH|5|10|Then said I to the angel that talked with me, Whither do these bear the ephah?
ZECH|5|11|And he said unto me, To build it an house in the land of Shinar: and it shall be established, and set there upon her own base.
ZECH|6|1|And I turned, and lifted up mine eyes, and looked, and, behold, there came four chariots out from between two mountains; and the mountains were mountains of brass.
ZECH|6|2|In the first chariot were red horses; and in the second chariot black horses;
ZECH|6|3|And in the third chariot white horses; and in the fourth chariot grisled and bay horses.
ZECH|6|4|Then I answered and said unto the angel that talked with me, What are these, my lord?
ZECH|6|5|And the angel answered and said unto me, These are the four spirits of the heavens, which go forth from standing before the LORD of all the earth.
ZECH|6|6|The black horses which are therein go forth into the north country; and the white go forth after them; and the grisled go forth toward the south country.
ZECH|6|7|And the bay went forth, and sought to go that they might walk to and fro through the earth: and he said, Get you hence, walk to and fro through the earth. So they walked to and fro through the earth.
ZECH|6|8|Then cried he upon me, and spake unto me, saying, Behold, these that go toward the north country have quieted my spirit in the north country.
ZECH|6|9|And the word of the LORD came unto me, saying,
ZECH|6|10|Take of them of the captivity, even of Heldai, of Tobijah, and of Jedaiah, which are come from Babylon, and come thou the same day, and go into the house of Josiah the son of Zephaniah;
ZECH|6|11|Then take silver and gold, and make crowns, and set them upon the head of Joshua the son of Josedech, the high priest;
ZECH|6|12|And speak unto him, saying, Thus speaketh the LORD of hosts, saying, Behold the man whose name is The BRANCH; and he shall grow up out of his place, and he shall build the temple of the LORD:
ZECH|6|13|Even he shall build the temple of the LORD; and he shall bear the glory, and shall sit and rule upon his throne; and he shall be a priest upon his throne: and the counsel of peace shall be between them both.
ZECH|6|14|And the crowns shall be to Helem, and to Tobijah, and to Jedaiah, and to Hen the son of Zephaniah, for a memorial in the temple of the LORD.
ZECH|6|15|And they that are far off shall come and build in the temple of the LORD, and ye shall know that the LORD of hosts hath sent me unto you. And this shall come to pass, if ye will diligently obey the voice of the LORD your God.
ZECH|7|1|And it came to pass in the fourth year of king Darius, that the word of the LORD came unto Zechariah in the fourth day of the ninth month, even in Chisleu;
ZECH|7|2|When they had sent unto the house of God Sherezer and Regemmelech, and their men, to pray before the LORD,
ZECH|7|3|And to speak unto the priests which were in the house of the LORD of hosts, and to the prophets, saying, Should I weep in the fifth month, separating myself, as I have done these so many years?
ZECH|7|4|Then came the word of the LORD of hosts unto me, saying,
ZECH|7|5|Speak unto all the people of the land, and to the priests, saying, When ye fasted and mourned in the fifth and seventh month, even those seventy years, did ye at all fast unto me, even to me?
ZECH|7|6|And when ye did eat, and when ye did drink, did not ye eat for yourselves, and drink for yourselves?
ZECH|7|7|Should ye not hear the words which the LORD hath cried by the former prophets, when Jerusalem was inhabited and in prosperity, and the cities thereof round about her, when men inhabited the south and the plain?
ZECH|7|8|And the word of the LORD came unto Zechariah, saying,
ZECH|7|9|Thus speaketh the LORD of hosts, saying, Execute true judgment, and shew mercy and compassions every man to his brother:
ZECH|7|10|And oppress not the widow, nor the fatherless, the stranger, nor the poor; and let none of you imagine evil against his brother in your heart.
ZECH|7|11|But they refused to hearken, and pulled away the shoulder, and stopped their ears, that they should not hear.
ZECH|7|12|Yea, they made their hearts as an adamant stone, lest they should hear the law, and the words which the LORD of hosts hath sent in his spirit by the former prophets: therefore came a great wrath from the LORD of hosts.
ZECH|7|13|Therefore it is come to pass, that as he cried, and they would not hear; so they cried, and I would not hear, saith the LORD of hosts:
ZECH|7|14|But I scattered them with a whirlwind among all the nations whom they knew not. Thus the land was desolate after them, that no man passed through nor returned: for they laid the pleasant land desolate.
ZECH|8|1|Again the word of the LORD of hosts came to me, saying,
ZECH|8|2|Thus saith the LORD of hosts; I was jealous for Zion with great jealousy, and I was jealous for her with great fury.
ZECH|8|3|Thus saith the LORD; I am returned unto Zion, and will dwell in the midst of Jerusalem: and Jerusalem shall be called a city of truth; and the mountain of the LORD of hosts the holy mountain.
ZECH|8|4|Thus saith the LORD of hosts; There shall yet old men and old women dwell in the streets of Jerusalem, and every man with his staff in his hand for very age.
ZECH|8|5|And the streets of the city shall be full of boys and girls playing in the streets thereof.
ZECH|8|6|Thus saith the LORD of hosts; If it be marvellous in the eyes of the remnant of this people in these days, should it also be marvellous in mine eyes? saith the LORD of hosts.
ZECH|8|7|Thus saith the LORD of hosts; Behold, I will save my people from the east country, and from the west country;
ZECH|8|8|And I will bring them, and they shall dwell in the midst of Jerusalem: and they shall be my people, and I will be their God, in truth and in righteousness.
ZECH|8|9|Thus saith the LORD of hosts; Let your hands be strong, ye that hear in these days these words by the mouth of the prophets, which were in the day that the foundation of the house of the LORD of hosts was laid, that the temple might be built.
ZECH|8|10|For before these days there was no hire for man, nor any hire for beast; neither was there any peace to him that went out or came in because of the affliction: for I set all men every one against his neighbour.
ZECH|8|11|But now I will not be unto the residue of this people as in the former days, saith the LORD of hosts.
ZECH|8|12|For the seed shall be prosperous; the vine shall give her fruit, and the ground shall give her increase, and the heavens shall give their dew; and I will cause the remnant of this people to possess all these things.
ZECH|8|13|And it shall come to pass, that as ye were a curse among the heathen, O house of Judah, and house of Israel; so will I save you, and ye shall be a blessing: fear not, but let your hands be strong.
ZECH|8|14|For thus saith the LORD of hosts; As I thought to punish you, when your fathers provoked me to wrath, saith the LORD of hosts, and I repented not:
ZECH|8|15|So again have I thought in these days to do well unto Jerusalem and to the house of Judah: fear ye not.
ZECH|8|16|These are the things that ye shall do; Speak ye every man the truth to his neighbour; execute the judgment of truth and peace in your gates:
ZECH|8|17|And let none of you imagine evil in your hearts against his neighbour; and love no false oath: for all these are things that I hate, saith the LORD.
ZECH|8|18|And the word of the LORD of hosts came unto me, saying,
ZECH|8|19|Thus saith the LORD of hosts; The fast of the fourth month, and the fast of the fifth, and the fast of the seventh, and the fast of the tenth, shall be to the house of Judah joy and gladness, and cheerful feasts; therefore love the truth and peace.
ZECH|8|20|Thus saith the LORD of hosts; It shall yet come to pass, that there shall come people, and the inhabitants of many cities:
ZECH|8|21|And the inhabitants of one city shall go to another, saying, Let us go speedily to pray before the LORD, and to seek the LORD of hosts: I will go also.
ZECH|8|22|Yea, many people and strong nations shall come to seek the LORD of hosts in Jerusalem, and to pray before the LORD.
ZECH|8|23|Thus saith the LORD of hosts; In those days it shall come to pass, that ten men shall take hold out of all languages of the nations, even shall take hold of the skirt of him that is a Jew, saying, We will go with you: for we have heard that God is with you.
ZECH|9|1|The burden of the word of the LORD in the land of Hadrach, and Damascus shall be the rest thereof: when the eyes of man, as of all the tribes of Israel, shall be toward the LORD.
ZECH|9|2|And Hamath also shall border thereby; Tyrus, and Zidon, though it be very wise.
ZECH|9|3|And Tyrus did build herself a strong hold, and heaped up silver as the dust, and fine gold as the mire of the streets.
ZECH|9|4|Behold, the LORD will cast her out, and he will smite her power in the sea; and she shall be devoured with fire.
ZECH|9|5|Ashkelon shall see it, and fear; Gaza also shall see it, and be very sorrowful, and Ekron; for her expectation shall be ashamed; and the king shall perish from Gaza, and Ashkelon shall not be inhabited.
ZECH|9|6|And a bastard shall dwell in Ashdod, and I will cut off the pride of the Philistines.
ZECH|9|7|And I will take away his blood out of his mouth, and his abominations from between his teeth: but he that remaineth, even he, shall be for our God, and he shall be as a governor in Judah, and Ekron as a Jebusite.
ZECH|9|8|And I will encamp about mine house because of the army, because of him that passeth by, and because of him that returneth: and no oppressor shall pass through them any more: for now have I seen with mine eyes.
ZECH|9|9|Rejoice greatly, O daughter of Zion; shout, O daughter of Jerusalem: behold, thy King cometh unto thee: he is just, and having salvation; lowly, and riding upon an ass, and upon a colt the foal of an ass.
ZECH|9|10|And I will cut off the chariot from Ephraim, and the horse from Jerusalem, and the battle bow shall be cut off: and he shall speak peace unto the heathen: and his dominion shall be from sea even to sea, and from the river even to the ends of the earth.
ZECH|9|11|As for thee also, by the blood of thy covenant I have sent forth thy prisoners out of the pit wherein is no water.
ZECH|9|12|Turn you to the strong hold, ye prisoners of hope: even to day do I declare that I will render double unto thee;
ZECH|9|13|When I have bent Judah for me, filled the bow with Ephraim, and raised up thy sons, O Zion, against thy sons, O Greece, and made thee as the sword of a mighty man.
ZECH|9|14|And the LORD shall be seen over them, and his arrow shall go forth as the lightning: and the LORD God shall blow the trumpet, and shall go with whirlwinds of the south.
ZECH|9|15|The LORD of hosts shall defend them; and they shall devour, and subdue with sling stones; and they shall drink, and make a noise as through wine; and they shall be filled like bowls, and as the corners of the altar.
ZECH|9|16|And the LORD their God shall save them in that day as the flock of his people: for they shall be as the stones of a crown, lifted up as an ensign upon his land.
ZECH|9|17|For how great is his goodness, and how great is his beauty! corn shall make the young men cheerful, and new wine the maids.
ZECH|10|1|Ask ye of the LORD rain in the time of the latter rain; so the LORD shall make bright clouds, and give them showers of rain, to every one grass in the field.
ZECH|10|2|For the idols have spoken vanity, and the diviners have seen a lie, and have told false dreams; they comfort in vain: therefore they went their way as a flock, they were troubled, because there was no shepherd.
ZECH|10|3|Mine anger was kindled against the shepherds, and I punished the goats: for the LORD of hosts hath visited his flock the house of Judah, and hath made them as his goodly horse in the battle.
ZECH|10|4|Out of him came forth the corner, out of him the nail, out of him the battle bow, out of him every oppressor together.
ZECH|10|5|And they shall be as mighty men, which tread down their enemies in the mire of the streets in the battle: and they shall fight, because the LORD is with them, and the riders on horses shall be confounded.
ZECH|10|6|And I will strengthen the house of Judah, and I will save the house of Joseph, and I will bring them again to place them; for I have mercy upon them: and they shall be as though I had not cast them off: for I am the LORD their God, and will hear them.
ZECH|10|7|And they of Ephraim shall be like a mighty man, and their heart shall rejoice as through wine: yea, their children shall see it, and be glad; their heart shall rejoice in the LORD.
ZECH|10|8|I will hiss for them, and gather them; for I have redeemed them: and they shall increase as they have increased.
ZECH|10|9|And I will sow them among the people: and they shall remember me in far countries; and they shall live with their children, and turn again.
ZECH|10|10|I will bring them again also out of the land of Egypt, and gather them out of Assyria; and I will bring them into the land of Gilead and Lebanon; and place shall not be found for them.
ZECH|10|11|And he shall pass through the sea with affliction, and shall smite the waves in the sea, and all the deeps of the river shall dry up: and the pride of Assyria shall be brought down, and the sceptre of Egypt shall depart away.
ZECH|10|12|And I will strengthen them in the LORD; and they shall walk up and down in his name, saith the LORD.
ZECH|11|1|Open thy doors, O Lebanon, that the fire may devour thy cedars.
ZECH|11|2|Howl, fir tree; for the cedar is fallen; because the mighty are spoiled: howl, O ye oaks of Bashan; for the forest of the vintage is come down.
ZECH|11|3|There is a voice of the howling of the shepherds; for their glory is spoiled: a voice of the roaring of young lions; for the pride of Jordan is spoiled.
ZECH|11|4|Thus saith the LORD my God; Feed the flock of the slaughter;
ZECH|11|5|Whose possessors slay them, and hold themselves not guilty: and they that sell them say, Blessed be the LORD; for I am rich: and their own shepherds pity them not.
ZECH|11|6|For I will no more pity the inhabitants of the land, saith the LORD: but, lo, I will deliver the men every one into his neighbour's hand, and into the hand of his king: and they shall smite the land, and out of their hand I will not deliver them.
ZECH|11|7|And I will feed the flock of slaughter, even you, O poor of the flock. And I took unto me two staves; the one I called Beauty, and the other I called Bands; and I fed the flock.
ZECH|11|8|Three shepherds also I cut off in one month; and my soul lothed them, and their soul also abhorred me.
ZECH|11|9|Then said I, I will not feed you: that that dieth, let it die; and that that is to be cut off, let it be cut off; and let the rest eat every one the flesh of another.
ZECH|11|10|And I took my staff, even Beauty, and cut it asunder, that I might break my covenant which I had made with all the people.
ZECH|11|11|And it was broken in that day: and so the poor of the flock that waited upon me knew that it was the word of the LORD.
ZECH|11|12|And I said unto them, If ye think good, give me my price; and if not, forbear. So they weighed for my price thirty pieces of silver.
ZECH|11|13|And the LORD said unto me, Cast it unto the potter: a goodly price that I was prised at of them. And I took the thirty pieces of silver, and cast them to the potter in the house of the LORD.
ZECH|11|14|Then I cut asunder mine other staff, even Bands, that I might break the brotherhood between Judah and Israel.
ZECH|11|15|And the LORD said unto me, Take unto thee yet the instruments of a foolish shepherd.
ZECH|11|16|For, lo, I will raise up a shepherd in the land, which shall not visit those that be cut off, neither shall seek the young one, nor heal that that is broken, nor feed that that standeth still: but he shall eat the flesh of the fat, and tear their claws in pieces.
ZECH|11|17|Woe to the idol shepherd that leaveth the flock! the sword shall be upon his arm, and upon his right eye: his arm shall be clean dried up, and his right eye shall be utterly darkened.
ZECH|12|1|The burden of the word of the LORD for Israel, saith the LORD, which stretcheth forth the heavens, and layeth the foundation of the earth, and formeth the spirit of man within him.
ZECH|12|2|Behold, I will make Jerusalem a cup of trembling unto all the people round about, when they shall be in the siege both against Judah and against Jerusalem.
ZECH|12|3|And in that day will I make Jerusalem a burdensome stone for all people: all that burden themselves with it shall be cut in pieces, though all the people of the earth be gathered together against it.
ZECH|12|4|In that day, saith the LORD, I will smite every horse with astonishment, and his rider with madness: and I will open mine eyes upon the house of Judah, and will smite every horse of the people with blindness.
ZECH|12|5|And the governors of Judah shall say in their heart, The inhabitants of Jerusalem shall be my strength in the LORD of hosts their God.
ZECH|12|6|In that day will I make the governors of Judah like an hearth of fire among the wood, and like a torch of fire in a sheaf; and they shall devour all the people round about, on the right hand and on the left: and Jerusalem shall be inhabited again in her own place, even in Jerusalem.
ZECH|12|7|The LORD also shall save the tents of Judah first, that the glory of the house of David and the glory of the inhabitants of Jerusalem do not magnify themselves against Judah.
ZECH|12|8|In that day shall the LORD defend the inhabitants of Jerusalem; and he that is feeble among them at that day shall be as David; and the house of David shall be as God, as the angel of the LORD before them.
ZECH|12|9|And it shall come to pass in that day, that I will seek to destroy all the nations that come against Jerusalem.
ZECH|12|10|And I will pour upon the house of David, and upon the inhabitants of Jerusalem, the spirit of grace and of supplications: and they shall look upon me whom they have pierced, and they shall mourn for him, as one mourneth for his only son, and shall be in bitterness for him, as one that is in bitterness for his firstborn.
ZECH|12|11|In that day shall there be a great mourning in Jerusalem, as the mourning of Hadadrimmon in the valley of Megiddon.
ZECH|12|12|And the land shall mourn, every family apart; the family of the house of David apart, and their wives apart; the family of the house of Nathan apart, and their wives apart;
ZECH|12|13|The family of the house of Levi apart, and their wives apart; the family of Shimei apart, and their wives apart;
ZECH|12|14|All the families that remain, every family apart, and their wives apart.
ZECH|13|1|In that day there shall be a fountain opened to the house of David and to the inhabitants of Jerusalem for sin and for uncleanness.
ZECH|13|2|And it shall come to pass in that day, saith the LORD of hosts, that I will cut off the names of the idols out of the land, and they shall no more be remembered: and also I will cause the prophets and the unclean spirit to pass out of the land.
ZECH|13|3|And it shall come to pass, that when any shall yet prophesy, then his father and his mother that begat him shall say unto him, Thou shalt not live; for thou speakest lies in the name of the LORD: and his father and his mother that begat him shall thrust him through when he prophesieth.
ZECH|13|4|And it shall come to pass in that day, that the prophets shall be ashamed every one of his vision, when he hath prophesied; neither shall they wear a rough garment to deceive:
ZECH|13|5|But he shall say, I am no prophet, I am an husbandman; for man taught me to keep cattle from my youth.
ZECH|13|6|And one shall say unto him, What are these wounds in thine hands? Then he shall answer, Those with which I was wounded in the house of my friends.
ZECH|13|7|Awake, O sword, against my shepherd, and against the man that is my fellow, saith the LORD of hosts: smite the shepherd, and the sheep shall be scattered: and I will turn mine hand upon the little ones.
ZECH|13|8|And it shall come to pass, that in all the land, saith the LORD, two parts therein shall be cut off and die; but the third shall be left therein.
ZECH|13|9|And I will bring the third part through the fire, and will refine them as silver is refined, and will try them as gold is tried: they shall call on my name, and I will hear them: I will say, It is my people: and they shall say, The LORD is my God.
ZECH|14|1|Behold, the day of the LORD cometh, and thy spoil shall be divided in the midst of thee.
ZECH|14|2|For I will gather all nations against Jerusalem to battle; and the city shall be taken, and the houses rifled, and the women ravished; and half of the city shall go forth into captivity, and the residue of the people shall not be cut off from the city.
ZECH|14|3|Then shall the LORD go forth, and fight against those nations, as when he fought in the day of battle.
ZECH|14|4|And his feet shall stand in that day upon the mount of Olives, which is before Jerusalem on the east, and the mount of Olives shall cleave in the midst thereof toward the east and toward the west, and there shall be a very great valley; and half of the mountain shall remove toward the north, and half of it toward the south.
ZECH|14|5|And ye shall flee to the valley of the mountains; for the valley of the mountains shall reach unto Azal: yea, ye shall flee, like as ye fled from before the earthquake in the days of Uzziah king of Judah: and the LORD my God shall come, and all the saints with thee.
ZECH|14|6|And it shall come to pass in that day, that the light shall not be clear, nor dark:
ZECH|14|7|But it shall be one day which shall be known to the LORD, not day, nor night: but it shall come to pass, that at evening time it shall be light.
ZECH|14|8|And it shall be in that day, that living waters shall go out from Jerusalem; half of them toward the former sea, and half of them toward the hinder sea: in summer and in winter shall it be.
ZECH|14|9|And the LORD shall be king over all the earth: in that day shall there be one LORD, and his name one.
ZECH|14|10|All the land shall be turned as a plain from Geba to Rimmon south of Jerusalem: and it shall be lifted up, and inhabited in her place, from Benjamin's gate unto the place of the first gate, unto the corner gate, and from the tower of Hananeel unto the king's winepresses.
ZECH|14|11|And men shall dwell in it, and there shall be no more utter destruction; but Jerusalem shall be safely inhabited.
ZECH|14|12|And this shall be the plague wherewith the LORD will smite all the people that have fought against Jerusalem; Their flesh shall consume away while they stand upon their feet, and their eyes shall consume away in their holes, and their tongue shall consume away in their mouth.
ZECH|14|13|And it shall come to pass in that day, that a great tumult from the LORD shall be among them; and they shall lay hold every one on the hand of his neighbour, and his hand shall rise up against the hand of his neighbour.
ZECH|14|14|And Judah also shall fight at Jerusalem; and the wealth of all the heathen round about shall be gathered together, gold, and silver, and apparel, in great abundance.
ZECH|14|15|And so shall be the plague of the horse, of the mule, of the camel, and of the ass, and of all the beasts that shall be in these tents, as this plague.
ZECH|14|16|And it shall come to pass, that every one that is left of all the nations which came against Jerusalem shall even go up from year to year to worship the King, the LORD of hosts, and to keep the feast of tabernacles.
ZECH|14|17|And it shall be, that whoso will not come up of all the families of the earth unto Jerusalem to worship the King, the LORD of hosts, even upon them shall be no rain.
ZECH|14|18|And if the family of Egypt go not up, and come not, that have no rain; there shall be the plague, wherewith the LORD will smite the heathen that come not up to keep the feast of tabernacles.
ZECH|14|19|This shall be the punishment of Egypt, and the punishment of all nations that come not up to keep the feast of tabernacles.
ZECH|14|20|In that day shall there be upon the bells of the horses, HOLINESS UNTO THE LORD; and the pots in the LORD's house shall be like the bowls before the altar.
ZECH|14|21|Yea, every pot in Jerusalem and in Judah shall be holiness unto the LORD of hosts: and all they that sacrifice shall come and take of them, and seethe therein: and in that day there shall be no more the Canaanite in the house of the LORD of hosts.
