1THESS|1|1|Павел и Силуан и Тимофей – церкви Фессалоникской в Боге Отце и Господе Иисусе Христе: благодать вам и мир от Бога Отца нашего и Господа Иисуса Христа.
1THESS|1|2|Всегда благодарим Бога за всех вас, вспоминая о вас в молитвах наших,
1THESS|1|3|непрестанно памятуя ваше дело веры и труд любви и терпение упования на Господа нашего Иисуса Христа пред Богом и Отцем нашим,
1THESS|1|4|зная избрание ваше, возлюбленные Богом братия;
1THESS|1|5|потому что наше благовествование у вас было не в слове только, но и в силе и во Святом Духе, и со многим удостоверением, как вы [сами] знаете, каковы были мы для вас между вами.
1THESS|1|6|И вы сделались подражателями нам и Господу, приняв слово при многих скорбях с радостью Духа Святаго,
1THESS|1|7|так что вы стали образцом для всех верующих в Македонии и Ахаии.
1THESS|1|8|Ибо от вас пронеслось слово Господне не только в Македонии и Ахаии, но и во всяком месте прошла [слава] о вере вашей в Бога, так что нам ни о чем не нужно рассказывать.
1THESS|1|9|Ибо сами они сказывают о нас, какой вход имели мы к вам, и как вы обратились к Богу от идолов, [чтобы] служить Богу живому и истинному
1THESS|1|10|и ожидать с небес Сына Его, Которого Он воскресил из мертвых, Иисуса, избавляющего нас от грядущего гнева.
1THESS|2|1|Вы сами знаете, братия, о нашем входе к вам, что он был не бездейственный;
1THESS|2|2|но, прежде пострадав и быв поруганы в Филиппах, как вы знаете, мы дерзнули в Боге нашем проповедать вам благовестие Божие с великим подвигом.
1THESS|2|3|Ибо в учении нашем нет ни заблуждения, ни нечистых [побуждений], ни лукавства;
1THESS|2|4|но, как Бог удостоил нас того, чтобы вверить [нам] благовестие, так мы и говорим, угождая не человекам, но Богу, испытующему сердца наши.
1THESS|2|5|Ибо никогда не было у нас перед вами ни слов ласкательства, как вы знаете, ни видов корысти: Бог свидетель!
1THESS|2|6|Не ищем славы человеческой ни от вас, ни от других:
1THESS|2|7|мы могли явиться с важностью, как Апостолы Христовы, но были тихи среди вас, подобно как кормилица нежно обходится с детьми своими.
1THESS|2|8|Так мы, из усердия к вам, восхотели передать вам не только благовестие Божие, но и души наши, потому что вы стали нам любезны.
1THESS|2|9|Ибо вы помните, братия, труд наш и изнурение: ночью и днем работая, чтобы не отяготить кого из вас, мы проповедывали у вас благовестие Божие.
1THESS|2|10|Свидетели вы и Бог, как свято и праведно и безукоризненно поступали мы перед вами, верующими,
1THESS|2|11|потому что вы знаете, как каждого из вас, как отец детей своих,
1THESS|2|12|мы просили и убеждали и умоляли поступать достойно Бога, призвавшего вас в Свое Царство и славу.
1THESS|2|13|Посему и мы непрестанно благодарим Бога, что, приняв от нас слышанное слово Божие, вы приняли не [как] слово человеческое, но [как] слово Божие, – каково оно есть по истине, – которое и действует в вас, верующих.
1THESS|2|14|Ибо вы, братия, сделались подражателями церквам Божиим во Христе Иисусе, находящимся в Иудее, потому что и вы то же претерпели от своих единоплеменников, что и те от Иудеев,
1THESS|2|15|которые убили и Господа Иисуса и Его пророков, и нас изгнали, и Богу не угождают, и всем человекам противятся,
1THESS|2|16|которые препятствуют нам говорить язычникам, чтобы спаслись, и через это всегда наполняют меру грехов своих; но приближается на них гнев до конца.
1THESS|2|17|Мы же, братия, быв разлучены с вами на короткое время лицем, а не сердцем, тем с большим желанием старались увидеть лице ваше.
1THESS|2|18|И потому мы, я Павел, и раз и два хотели прийти к вам, но воспрепятствовал нам сатана.
1THESS|2|19|Ибо кто наша надежда, или радость, или венец похвалы? Не и вы ли пред Господом нашим Иисусом Христом в пришествие Его?
1THESS|2|20|Ибо вы – слава наша и радость.
1THESS|3|1|И потому, не терпя более, мы восхотели остаться в Афинах одни,
1THESS|3|2|и послали Тимофея, брата нашего и служителя Божия и сотрудника нашего в благовествовании Христовом, чтобы утвердить вас и утешить в вере вашей,
1THESS|3|3|чтобы никто не поколебался в скорбях сих: ибо вы сами знаете, что так нам суждено.
1THESS|3|4|Ибо мы и тогда, как были у вас, предсказывали вам, что будем страдать, как и случилось, и вы знаете.
1THESS|3|5|Посему и я, не терпя более, послал узнать о вере вашей, чтобы как не искусил вас искуситель и не сделался тщетным труд наш.
1THESS|3|6|Теперь же, когда пришел к нам от вас Тимофей и принес нам добрую весть о вере и любви вашей, и что вы всегда имеете добрую память о нас, желая нас видеть, как и мы вас,
1THESS|3|7|то мы, при всей скорби и нужде нашей, утешились вами, братия, ради вашей веры;
1THESS|3|8|ибо теперь мы живы, когда вы стоите в Господе.
1THESS|3|9|Какую благодарность можем мы воздать Богу за вас, за всю радость, которою радуемся о вас пред Богом нашим,
1THESS|3|10|ночь и день всеусердно молясь о том, чтобы видеть лице ваше и дополнить, чего недоставало вере вашей?
1THESS|3|11|Сам же Бог и Отец наш и Господь наш Иисус Христос да управит путь наш к вам.
1THESS|3|12|А вас Господь да исполнит и преисполнит любовью друг к другу и ко всем, какою мы исполнены к вам,
1THESS|3|13|чтобы утвердить сердца ваши непорочными во святыне пред Богом и Отцем нашим в пришествие Господа нашего Иисуса Христа со всеми святыми Его. Аминь.
1THESS|4|1|За сим, братия, просим и умоляем вас Христом Иисусом, чтобы вы, приняв от нас, как должно вам поступать и угождать Богу, более в том преуспевали,
1THESS|4|2|ибо вы знаете, какие мы дали вам заповеди от Господа Иисуса.
1THESS|4|3|Ибо воля Божия есть освящение ваше, чтобы вы воздерживались от блуда;
1THESS|4|4|чтобы каждый из вас умел соблюдать свой сосуд в святости и чести,
1THESS|4|5|а не в страсти похотения, как и язычники, не знающие Бога;
1THESS|4|6|чтобы вы ни в чем не поступали с братом своим противозаконно и корыстолюбиво: потому что Господь – мститель за все это, как и прежде мы говорили вам и свидетельствовали.
1THESS|4|7|Ибо призвал нас Бог не к нечистоте, но к святости.
1THESS|4|8|Итак непокорный непокорен не человеку, но Богу, Который и дал нам Духа Своего Святаго.
1THESS|4|9|О братолюбии же нет нужды писать к вам; ибо вы сами научены Богом любить друг друга,
1THESS|4|10|ибо вы так и поступаете со всеми братиями по всей Македонии. Умоляем же вас, братия, более преуспевать
1THESS|4|11|и усердно стараться о том, чтобы жить тихо, делать свое [дело] и работать своими собственными руками, как мы заповедывали вам;
1THESS|4|12|чтобы вы поступали благоприлично перед внешними и ни в чем не нуждались.
1THESS|4|13|Не хочу же оставить вас, братия, в неведении об умерших, дабы вы не скорбели, как прочие, не имеющие надежды.
1THESS|4|14|Ибо, если мы веруем, что Иисус умер и воскрес, то и умерших в Иисусе Бог приведет с Ним.
1THESS|4|15|Ибо сие говорим вам словом Господним, что мы живущие, оставшиеся до пришествия Господня, не предупредим умерших,
1THESS|4|16|потому что Сам Господь при возвещении, при гласе Архангела и трубе Божией, сойдет с неба, и мертвые во Христе воскреснут прежде;
1THESS|4|17|потом мы, оставшиеся в живых, вместе с ними восхищены будем на облаках в сретение Господу на воздухе, и так всегда с Господом будем.
1THESS|4|18|Итак утешайте друг друга сими словами.
1THESS|5|1|О временах же и сроках нет нужды писать к вам, братия,
1THESS|5|2|ибо сами вы достоверно знаете, что день Господень так придет, как тать ночью.
1THESS|5|3|Ибо, когда будут говорить: "мир и безопасность", тогда внезапно постигнет их пагуба, подобно как мука родами [постигает] имеющую во чреве, и не избегнут.
1THESS|5|4|Но вы, братия, не во тьме, чтобы день застал вас, как тать.
1THESS|5|5|Ибо все вы – сыны света и сыны дня: мы – не [сыны] ночи, ни тьмы.
1THESS|5|6|Итак, не будем спать, как и прочие, но будем бодрствовать и трезвиться.
1THESS|5|7|Ибо спящие спят ночью, и упивающиеся упиваются ночью.
1THESS|5|8|Мы же, будучи [сынами] дня, да трезвимся, облекшись в броню веры и любви и в шлем надежды спасения,
1THESS|5|9|потому что Бог определил нас не на гнев, но к получению спасения через Господа нашего Иисуса Христа,
1THESS|5|10|умершего за нас, чтобы мы, бодрствуем ли, или спим, жили вместе с Ним.
1THESS|5|11|Посему увещавайте друг друга и назидайте один другого, как вы и делаете.
1THESS|5|12|Просим же вас, братия, уважать трудящихся у вас, и предстоятелей ваших в Господе, и вразумляющих вас,
1THESS|5|13|и почитать их преимущественно с любовью за дело их; будьте в мире между собою.
1THESS|5|14|Умоляем также вас, братия, вразумляйте бесчинных, утешайте малодушных, поддерживайте слабых, будьте долготерпеливы ко всем.
1THESS|5|15|Смотрите, чтобы кто кому не воздавал злом за зло; но всегда ищите добра и друг другу и всем.
1THESS|5|16|Всегда радуйтесь.
1THESS|5|17|Непрестанно молитесь.
1THESS|5|18|За все благодарите: ибо такова о вас воля Божия во Христе Иисусе.
1THESS|5|19|Духа не угашайте.
1THESS|5|20|Пророчества не уничижайте.
1THESS|5|21|Все испытывайте, хорошего держитесь.
1THESS|5|22|Удерживайтесь от всякого рода зла.
1THESS|5|23|Сам же Бог мира да освятит вас во всей полноте, и ваш дух и душа и тело во всей целости да сохранится без порока в пришествие Господа нашего Иисуса Христа.
1THESS|5|24|Верен Призывающий вас, Который и сотворит [сие].
1THESS|5|25|Братия! молитесь о нас.
1THESS|5|26|Приветствуйте всех братьев лобзанием святым.
1THESS|5|27|Заклинаю вас Господом прочитать сие послание всем святым братиям.
1THESS|5|28|Благодать Господа нашего Иисуса Христа с вами. Аминь.
