1SAM|1|1|fuit vir unus de Ramathaimsophim de monte Ephraim et nomen eius Helcana filius Hieroam filii Heliu filii Thau filii Suph Ephratheus
1SAM|1|2|et habuit duas uxores nomen uni Anna et nomen secundae Fenenna fueruntque Fenennae filii Annae autem non erant liberi
1SAM|1|3|et ascendebat vir ille de civitate sua statutis diebus ut adoraret et sacrificaret Domino exercituum in Silo erant autem ibi duo filii Heli Ofni et Finees sacerdotes Domini
1SAM|1|4|venit ergo dies et immolavit Helcana deditque Fenennae uxori suae et cunctis filiis eius et filiabus partes
1SAM|1|5|Annae autem dedit partem unam tristis quia Annam diligebat Dominus autem concluserat vulvam eius
1SAM|1|6|adfligebat quoque eam aemula eius et vehementer angebat in tantum ut exprobraret quod conclusisset Dominus vulvam eius
1SAM|1|7|sicque faciebat per singulos annos cum redeunte tempore ascenderent templum Domini et sic provocabat eam porro illa flebat et non capiebat cibum
1SAM|1|8|dixit ergo ei Helcana vir suus Anna cur fles et quare non comedis et quam ob rem adfligitur cor tuum numquid non ego melior sum tibi quam decem filii
1SAM|1|9|surrexit autem Anna postquam comederat in Silo et biberat et Heli sacerdote sedente super sellam ante postes templi Domini
1SAM|1|10|cum esset amaro animo oravit Dominum flens largiter
1SAM|1|11|et votum vovit dicens Domine exercituum si respiciens videris adflictionem famulae tuae et recordatus mei fueris nec oblitus ancillae tuae dederisque servae tuae sexum virilem dabo eum Domino omnes dies vitae eius et novacula non ascendet super caput eius
1SAM|1|12|factum est ergo cum illa multiplicaret preces coram Domino ut Heli observaret os eius
1SAM|1|13|porro Anna loquebatur in corde suo tantumque labia illius movebantur et vox penitus non audiebatur aestimavit igitur eam Heli temulentam
1SAM|1|14|dixitque ei usquequo ebria eris digere paulisper vinum quo mades
1SAM|1|15|respondens Anna nequaquam inquit domine mi nam mulier infelix nimis ego sum vinumque et omne quod inebriare potest non bibi sed effudi animam meam in conspectu Domini
1SAM|1|16|ne reputes ancillam tuam quasi unam de filiabus Belial quia ex multitudine doloris et maeroris mei locuta sum usque in praesens
1SAM|1|17|tunc Heli ait ei vade in pace et Deus Israhel det tibi petitionem quam rogasti eum
1SAM|1|18|et illa dixit utinam inveniat ancilla tua gratiam in oculis tuis et abiit mulier in viam suam et comedit vultusque eius non sunt amplius in diversa mutati
1SAM|1|19|et surrexerunt mane et adoraverunt coram Domino reversique sunt et venerunt in domum suam Ramatha cognovit autem Helcana Annam uxorem suam et recordatus est eius Dominus
1SAM|1|20|et factum est post circulum dierum concepit Anna et peperit filium vocavitque nomen eius Samuhel eo quod a Domino postulasset eum
1SAM|1|21|ascendit autem vir Helcana et omnis domus eius ut immolaret Domino hostiam sollemnem et votum suum
1SAM|1|22|et Anna non ascendit dixit enim viro suo non vadam donec ablactetur infans et ducam eum et appareat ante conspectum Domini et maneat ibi iugiter
1SAM|1|23|et ait ei Helcana vir suus fac quod bonum tibi videtur et mane donec ablactes eum precorque ut impleat Dominus verbum suum mansit ergo mulier et lactavit filium suum donec amoveret eum a lacte
1SAM|1|24|et adduxit eum secum postquam ablactaverat in vitulis tribus et tribus modiis farinae et amphora vini et adduxit eum ad domum Domini in Silo puer autem erat adhuc infantulus
1SAM|1|25|et immolaverunt vitulum et obtulerunt puerum Heli
1SAM|1|26|et ait obsecro mi domine vivit anima tua domine ego sum illa mulier quae steti coram te hic orans Dominum
1SAM|1|27|pro puero isto oravi et dedit Dominus mihi petitionem meam quam postulavi eum
1SAM|1|28|idcirco et ego commodavi eum Domino cunctis diebus quibus fuerit accommodatus Domino et adoraverunt ibi Dominum et oravit Anna et ait
1SAM|2|1|exultavit cor meum in Domino exaltatum est cornu meum in Domino dilatatum est os meum super inimicos meos quia laetata sum in salutari tuo
1SAM|2|2|non est sanctus ut est Dominus neque enim est alius extra te et non est fortis sicut Deus noster
1SAM|2|3|nolite multiplicare loqui sublimia gloriantes recedant vetera de ore vestro quoniam Deus scientiarum Dominus est et ipsi praeparantur cogitationes
1SAM|2|4|arcus fortium superatus est et infirmi accincti sunt robore
1SAM|2|5|saturati prius pro pane se locaverunt et famelici saturati sunt donec sterilis peperit plurimos et quae multos habebat filios infirmata est
1SAM|2|6|Dominus mortificat et vivificat deducit ad infernum et reducit
1SAM|2|7|Dominus pauperem facit et ditat humiliat et sublevat
1SAM|2|8|suscitat de pulvere egenum et de stercore elevat pauperem ut sedeat cum principibus et solium gloriae teneat Domini enim sunt cardines terrae et posuit super eos orbem
1SAM|2|9|pedes sanctorum suorum servabit et impii in tenebris conticescent quia non in fortitudine roborabitur vir
1SAM|2|10|Dominum formidabunt adversarii eius super ipsos in caelis tonabit Dominus iudicabit fines terrae et dabit imperium regi suo et sublimabit cornu christi sui
1SAM|2|11|et abiit Helcana Ramatha in domum suam puer autem erat minister in conspectu Domini ante faciem Heli sacerdotis
1SAM|2|12|porro filii Heli filii Belial nescientes Dominum
1SAM|2|13|neque officium sacerdotum ad populum sed quicumque immolasset victimam veniebat puer sacerdotis dum coquerentur carnes et habebat fuscinulam tridentem in manu sua
1SAM|2|14|et mittebat eam in lebetem vel in caldariam aut in ollam sive in caccabum et omne quod levabat fuscinula tollebat sacerdos sibi sic faciebant universo Israheli venientium in Silo
1SAM|2|15|etiam antequam adolerent adipem veniebat puer sacerdotis et dicebat immolanti da mihi carnem ut coquam sacerdoti non enim accipiam a te carnem coctam sed crudam
1SAM|2|16|dicebatque illi immolans incendatur primum iuxta morem hodie adeps et tolle tibi quantumcumque desiderat anima tua qui respondens aiebat ei nequaquam nunc enim dabis alioquin tollam vi
1SAM|2|17|erat ergo peccatum puerorum grande nimis coram Domino quia detrahebant homines sacrificio Domini
1SAM|2|18|Samuhel autem ministrabat ante faciem Domini puer accinctus ephod lineo
1SAM|2|19|et tunicam parvam faciebat ei mater sua quam adferebat statutis diebus ascendens cum viro suo ut immolaret hostiam sollemnem
1SAM|2|20|et benedixit Heli Helcanae et uxori eius dixitque reddat Dominus tibi semen de muliere hac pro fenore quod commodasti Domino et abierunt in locum suum
1SAM|2|21|visitavit ergo Dominus Annam et concepit et peperit tres filios et duas filias et magnificatus est puer Samuhel apud Dominum
1SAM|2|22|Heli autem erat senex valde et audivit omnia quae faciebant filii sui universo Israheli et quomodo dormiebant cum mulieribus quae observabant ad ostium tabernaculi
1SAM|2|23|et dixit eis quare facitis res huiuscemodi quas ego audio res pessimas ab omni populo
1SAM|2|24|nolite filii mi non enim est bona fama quam ego audio ut transgredi faciatis populum Domini
1SAM|2|25|si peccaverit vir in virum placari ei potest Deus si autem in Domino peccaverit vir quis orabit pro eo et non audierunt vocem patris sui quia voluit Dominus occidere eos
1SAM|2|26|puer autem Samuhel proficiebat atque crescebat et placebat tam Deo quam hominibus
1SAM|2|27|venit autem vir Dei ad Heli et ait ad eum haec dicit Dominus numquid non aperte revelatus sum domui patris tui cum essent in Aegypto in domo Pharaonis
1SAM|2|28|et elegi eum ex omnibus tribubus Israhel mihi in sacerdotem ut ascenderet altare meum et adoleret mihi incensum et portaret ephod coram me et dedi domui patris tui omnia de sacrificiis filiorum Israhel
1SAM|2|29|quare calce abicitis victimam meam et munera mea quae praecepi ut offerrentur in templo et magis honorasti filios tuos quam me ut comederetis primitias omnis sacrificii Israhel populi mei
1SAM|2|30|propterea ait Dominus Deus Israhel loquens locutus sum ut domus tua et domus patris tui ministraret in conspectu meo usque in sempiternum nunc autem dicit Dominus absit hoc a me sed quicumque glorificaverit me glorificabo eum qui autem contemnunt me erunt ignobiles
1SAM|2|31|ecce dies veniunt et praecidam brachium tuum et brachium domus patris tui ut non sit senex in domo tua
1SAM|2|32|et videbis aemulum tuum in templo in universis prosperis Israhel et non erit senex in domo tua omnibus diebus
1SAM|2|33|verumtamen non auferam penitus virum ex te ab altari meo sed ut deficiant oculi tui et tabescat anima tua et pars magna domus tuae morietur cum ad virilem aetatem venerit
1SAM|2|34|hoc autem erit tibi signum quod venturum est duobus filiis tuis Ofni et Finees in die uno morientur ambo
1SAM|2|35|et suscitabo mihi sacerdotem fidelem qui iuxta cor meum et animam meam faciat et aedificabo ei domum fidelem et ambulabit coram christo meo cunctis diebus
1SAM|2|36|futurum est autem ut quicumque remanserit in domo tua veniat ut oretur pro eo et offerat nummum argenteum et tortam panis dicatque dimitte me obsecro ad unam partem sacerdotalem ut comedam buccellam panis
1SAM|3|1|puer autem Samuhel ministrabat Domino coram Heli et sermo Domini erat pretiosus in diebus illis non erat visio manifesta
1SAM|3|2|factum est ergo in die quadam Heli iacebat in loco suo et oculi eius caligaverant nec poterat videre
1SAM|3|3|lucerna Dei antequam extingueretur Samuhel autem dormiebat in templo Domini ubi erat arca Dei
1SAM|3|4|et vocavit Dominus Samuhel qui respondens ait ecce ego
1SAM|3|5|et cucurrit ad Heli et dixit ecce ego vocasti enim me qui dixit non vocavi revertere dormi et abiit et dormivit
1SAM|3|6|et adiecit Dominus vocare rursum Samuhel consurgensque Samuhel abiit ad Heli et dixit ecce ego quia vocasti me qui respondit non vocavi te fili mi revertere et dormi
1SAM|3|7|porro Samuhel necdum sciebat Dominum neque revelatus fuerat ei sermo Domini
1SAM|3|8|et adiecit Dominus et vocavit adhuc Samuhel tertio qui consurgens abiit ad Heli
1SAM|3|9|et ait ecce ego quia vocasti me intellexit igitur Heli quia Dominus vocaret puerum et ait ad Samuhel vade et dormi et si deinceps vocaverit te dices loquere Domine quia audit servus tuus abiit ergo Samuhel et dormivit in loco suo
1SAM|3|10|et venit Dominus et stetit et vocavit sicut vocaverat secundo Samuhel Samuhel et ait Samuhel loquere quia audit servus tuus
1SAM|3|11|et dixit Dominus ad Samuhel ecce ego facio verbum in Israhel quod quicumque audierit tinnient ambae aures eius
1SAM|3|12|in die illo suscitabo adversum Heli omnia quae locutus sum super domum eius incipiam et conplebo
1SAM|3|13|praedixi enim ei quod iudicaturus essem domum eius in aeternum propter iniquitatem eo quod noverat indigne agere filios suos et non corripuit eos
1SAM|3|14|idcirco iuravi domui Heli quod non expietur iniquitas domus eius victimis et muneribus usque in aeternum
1SAM|3|15|dormivit autem Samuhel usque mane aperuitque ostia domus Domini et Samuhel timebat indicare visionem Heli
1SAM|3|16|vocavit ergo Heli Samuhelem et dixit Samuhel fili mi qui respondens ait praesto sum
1SAM|3|17|et interrogavit eum quis est sermo quem locutus est ad te oro te ne celaveris me haec faciat tibi Deus et haec addat si absconderis a me sermonem ex omnibus verbis quae dicta sunt tibi
1SAM|3|18|indicavit itaque ei Samuhel universos sermones et non abscondit ab eo et ille respondit Dominus est quod bonum est in oculis suis faciat
1SAM|3|19|crevit autem Samuhel et Dominus erat cum eo et non cecidit ex omnibus verbis eius in terram
1SAM|3|20|et cognovit universus Israhel a Dan usque Bersabee quod fidelis Samuhel propheta esset Domini
1SAM|3|21|et addidit Dominus ut appareret in Silo quoniam revelatus fuerat Dominus Samuheli in Silo iuxta verbum Domini et evenit sermo Samuhelis universo Israheli
1SAM|4|1|egressus est namque Israhel obviam Philisthim in proelium et castrametatus est iuxta lapidem Adiutorii porro Philisthim venerunt in Afec
1SAM|4|2|et instruxerunt aciem contra Israhel inito autem certamine terga vertit Israhel Philistheis et caesa sunt in illo certamine passim per agros quasi quattuor milia virorum
1SAM|4|3|et reversus est populus ad castra dixeruntque maiores natu de Israhel quare percussit nos Dominus hodie coram Philisthim adferamus ad nos de Silo arcam foederis Domini et veniat in medium nostri ut salvet nos de manu inimicorum nostrorum
1SAM|4|4|misit ergo populus in Silo et tulerunt inde arcam foederis Domini exercituum sedentis super cherubin erantque duo filii Heli cum arca foederis Domini Ofni et Finees
1SAM|4|5|cumque venisset arca foederis Domini in castra vociferatus est omnis Israhel clamore grandi et personuit terra
1SAM|4|6|et audierunt Philisthim vocem clamoris dixeruntque quaenam haec est vox clamoris magni in castris Hebraeorum et cognoverunt quod arca Domini venisset in castra
1SAM|4|7|timueruntque Philisthim dicentes venit Deus in castra et ingemuerunt
1SAM|4|8|vae nobis non enim fuit tanta exultatio heri et nudius tertius vae nobis quis nos servabit de manu deorum sublimium istorum hii sunt dii qui percusserunt Aegyptum omni plaga in deserto
1SAM|4|9|confortamini et estote viri Philisthim ne serviatis Hebraeis sicut illi servierunt vobis confortamini et bellate
1SAM|4|10|pugnaverunt ergo Philisthim et caesus est Israhel et fugit unusquisque in tabernaculum suum et facta est plaga magna nimis et ceciderunt de Israhel triginta milia peditum
1SAM|4|11|et arca Dei capta est duoque filii Heli mortui sunt Ofni et Finees
1SAM|4|12|currens autem vir de Beniamin ex acie venit in Silo in die illo scissa veste et conspersus pulvere caput
1SAM|4|13|cumque ille venisset Heli sedebat super sellam contra viam aspectans erat enim cor eius pavens pro arca Domini vir autem ille postquam ingressus est nuntiavit urbi et ululavit omnis civitas
1SAM|4|14|et audivit Heli sonitum clamoris dixitque quis est hic sonitus tumultus huius at ille festinavit et venit et adnuntiavit Heli
1SAM|4|15|Heli autem erat nonaginta et octo annorum et oculi eius caligaverant et videre non poterat
1SAM|4|16|et dixit ad Heli ego sum qui veni de proelio et ego qui de acie fugi hodie cui ille ait quid actum est fili mi
1SAM|4|17|respondens autem qui nuntiabat fugit inquit Israhel coram Philisthim et ruina magna facta est in populo insuper et duo filii tui mortui sunt Ofni et Finees et arca Dei capta est
1SAM|4|18|cumque ille nominasset arcam Dei cecidit de sella retrorsum iuxta ostium et fractis cervicibus mortuus est senex enim erat vir et grandevus et ipse iudicavit Israhel quadraginta annis
1SAM|4|19|nurus autem eius uxor Finees praegnans erat vicinaque partui et audito nuntio quod capta esset arca Dei et mortuus socer suus et vir suus incurvavit se et peperit inruerant enim in eam dolores subiti
1SAM|4|20|in ipso autem momento mortis eius dixerunt ei quae stabant circa eam ne timeas quia filium peperisti quae non respondit eis neque animadvertit
1SAM|4|21|et vocavit puerum Hicabod dicens translata est gloria de Israhel quia capta est arca Dei et pro socero suo et pro viro suo
1SAM|4|22|et ait translata est gloria ab Israhel eo quod capta esset arca Dei
1SAM|5|1|Philisthim autem tulerunt arcam Dei et asportaverunt eam a lapide Adiutorii in Azotum
1SAM|5|2|tulerunt Philisthim arcam Dei et intulerunt eam in templum Dagon et statuerunt eam iuxta Dagon
1SAM|5|3|cumque surrexissent diluculo Azotii altera die ecce Dagon iacebat pronus in terram ante arcam Domini et tulerunt Dagon et restituerunt eum in loco suo
1SAM|5|4|rursumque mane die alio consurgentes invenerunt Dagon iacentem super faciem suam in terram coram arca Domini caput autem Dagon et duae palmae manuum eius abscisae erant super limen
1SAM|5|5|porro Dagon truncus solus remanserat in loco suo propter hanc causam non calcant sacerdotes Dagon et omnes qui ingrediuntur templum eius super limen Dagon in Azoto usque in hodiernum diem
1SAM|5|6|adgravata autem est manus Domini super Azotios et demolitus est eos et percussit in secretiori parte natium Azotum et fines eius
1SAM|5|7|videntes autem viri azotii huiuscemodi plagam dixerunt non maneat arca Dei Israhel apud nos quoniam dura est manus eius super nos et super Dagon deum nostrum
1SAM|5|8|et mittentes congregaverunt omnes satrapas Philisthinorum ad se et dixerunt quid faciemus de arca Dei Israhel responderuntque Getthei circumducatur arca Dei Israhel et circumduxerunt arcam Dei Israhel
1SAM|5|9|illis autem circumducentibus eam fiebat manus Dei per singulas civitates interfectionis magnae nimis et percutiebat viros uniuscuiusque urbis a parvo usque ad maiorem et conputrescebant prominentes extales eorum
1SAM|5|10|miserunt ergo arcam Dei in Accaron cumque venisset arca Dei in Accaron exclamaverunt Accaronitae dicentes adduxerunt ad nos arcam Dei Israhel ut interficiat nos et populum nostrum
1SAM|5|11|miserunt itaque et congregaverunt omnes satrapas Philisthinorum qui dixerunt dimittite arcam Dei Israhel et revertatur in locum suum et non interficiat nos cum populo nostro
1SAM|5|12|fiebat enim pavor mortis in singulis urbibus et gravissima valde manus Dei viri quoque qui mortui non fuerant percutiebantur in secretiori parte natium et ascendebat ululatus uniuscuiusque civitatis in caelum
1SAM|6|1|fuit ergo arca Domini in regione Philisthinorum septem mensibus
1SAM|6|2|et vocaverunt Philisthim sacerdotes et divinos dicentes quid faciemus de arca Dei indicate nobis quomodo remittemus eam in locum suum qui dixerunt
1SAM|6|3|si remittitis arcam Dei Israhel nolite dimittere eam vacuam sed quod debetis reddite ei pro peccato et tunc curabimini et scietis quare non recedat manus eius a vobis
1SAM|6|4|qui dixerunt quid est quod pro delicto reddere debeamus ei responderuntque illi
1SAM|6|5|iuxta numerum provinciarum Philisthim quinque anos aureos facietis et quinque mures aureos quia plaga una fuit omnibus vobis et satrapis vestris facietisque similitudines anorum vestrorum et similitudines murium qui demoliti sunt terram et dabitis Deo Israhel gloriam si forte relevet manum suam a vobis et a diis vestris et a terra vestra
1SAM|6|6|quare gravatis corda vestra sicut adgravavit Aegyptus et Pharao cor suum nonne postquam percussus est tunc dimisit eos et abierunt
1SAM|6|7|nunc ergo arripite et facite plaustrum novum unum et duas vaccas fetas quibus non est inpositum iugum iungite in plaustro et recludite vitulos earum domi
1SAM|6|8|tolletisque arcam Domini et ponetis in plaustro et vasa aurea quae exsolvistis ei pro delicto ponetis in capsella ad latus eius et dimittite eam ut vadat
1SAM|6|9|et aspicietis et si quidem per viam finium suorum ascenderit contra Bethsames ipse fecit nobis malum hoc grande sin autem minime sciemus quia nequaquam manus eius tetigit nos sed casu accidit
1SAM|6|10|fecerunt ergo illi hoc modo et tollentes duas vaccas quae lactabant vitulos iunxerunt ad plaustrum vitulosque earum concluserunt domi
1SAM|6|11|et posuerunt arcam Dei super plaustrum et capsellam quae habebat mures aureos et similitudinem anorum
1SAM|6|12|ibant autem in directum vaccae per viam quae ducit Bethsames et itinere uno gradiebantur pergentes et mugientes et non declinabant neque ad dextram neque ad sinistram sed et satrapae Philisthinorum sequebantur usque ad terminos Bethsames
1SAM|6|13|porro Bethsamitae metebant triticum in valle et elevantes oculos viderunt arcam et gavisi sunt cum vidissent
1SAM|6|14|et plaustrum venit in agrum Iosue Bethsamitae et stetit ibi erat autem ibi lapis magnus et conciderunt ligna plaustri vaccasque inposuerunt super ea holocaustum Domino
1SAM|6|15|Levitae autem deposuerunt arcam Dei et capsellam quae erat iuxta eam in qua erant vasa aurea et posuerunt super lapidem grandem viri autem bethsamitae obtulerunt holocausta et immolaverunt victimas in die illa Domino
1SAM|6|16|et quinque satrapae Philisthinorum viderunt et reversi sunt in Accaron in die illa
1SAM|6|17|hii sunt autem ani aurei quos reddiderunt Philisthim pro delicto Domino Azotus unum Gaza unum Ascalon unum Geth unum Accaron unum
1SAM|6|18|et mures aureos secundum numerum urbium Philisthim quinque provinciarum ab urbe murata usque ad villam quae erat absque muro et usque ad Abel magnum super quem posuerunt arcam Domini quae erat usque in illa die in agro Iosue Bethsamitis
1SAM|6|19|percussit autem de viris bethsamitibus eo quod vidissent arcam Domini et percussit de populo septuaginta viros et quinquaginta milia plebis luxitque populus quod percussisset Dominus plebem plaga magna
1SAM|6|20|et dixerunt viri bethsamitae quis poterit stare in conspectu Domini Dei sancti huius et ad quem ascendet a nobis
1SAM|6|21|miseruntque nuntios ad habitatores Cariathiarim dicentes reduxerunt Philisthim arcam Domini descendite et ducite eam ad vos
1SAM|7|1|venerunt ergo viri Cariathiarim et duxerunt arcam Domini et intulerunt eam in domum Abinadab in Gabaa Eleazarum autem filium eius sanctificaverunt ut custodiret arcam Domini
1SAM|7|2|et factum est ex qua die mansit arca in Cariathiarim multiplicati sunt dies erat quippe iam annus vicesimus et requievit omnis domus Israhel post Dominum
1SAM|7|3|ait autem Samuhel ad universam domum Israhel dicens si in toto corde vestro revertimini ad Dominum auferte deos alienos de medio vestrum et Astharoth et praeparate corda vestra Domino et servite ei soli et eruet vos de manu Philisthim
1SAM|7|4|abstulerunt ergo filii Israhel Baalim et Astharoth et servierunt Domino soli
1SAM|7|5|dixit autem Samuhel congregate universum Israhel in Masphat ut orem pro vobis Dominum
1SAM|7|6|et convenerunt in Masphat hauseruntque aquam et effuderunt in conspectu Domini et ieiunaverunt in die illa et dixerunt ibi peccavimus Domino iudicavitque Samuhel filios Israhel in Masphat
1SAM|7|7|et audierunt Philisthim quod congregati essent filii Israhel in Masphat et ascenderunt satrapae Philisthinorum ad Israhel quod cum audissent filii Israhel timuerunt a facie Philisthinorum
1SAM|7|8|dixeruntque ad Samuhel ne cesses pro nobis clamare ad Dominum Deum nostrum ut salvet nos de manu Philisthinorum
1SAM|7|9|tulit autem Samuhel agnum lactantem unum et obtulit illum holocaustum integrum Domino et clamavit Samuhel ad Dominum pro Israhel et exaudivit eum Dominus
1SAM|7|10|factum est ergo cum Samuhel offerret holocaustum Philistheos inire proelium contra Israhel intonuit autem Dominus fragore magno in die illa super Philisthim et exterruit eos et caesi sunt a filiis Israhel
1SAM|7|11|egressique viri Israhel de Masphat persecuti sunt Philistheos et percusserunt eos usque ad locum qui erat subter Bethchar
1SAM|7|12|tulit autem Samuhel lapidem unum et posuit eum inter Masphat et inter Sen et vocavit nomen eius lapis Adiutorii dixitque hucusque auxiliatus est nobis Dominus
1SAM|7|13|et humiliati sunt Philisthim nec adposuerunt ultra ut venirent in terminos Israhel facta est itaque manus Domini super Philistheos cunctis diebus Samuhel
1SAM|7|14|et redditae sunt urbes quas tulerant Philisthim ab Israhel Israheli ab Accaron usque Geth et terminos suos liberavit Israhel de manu Philisthinorum eratque pax inter Israhel et Amorreum
1SAM|7|15|iudicabat quoque Samuhel Israhel cunctis diebus vitae suae
1SAM|7|16|et ibat per singulos annos circumiens Bethel et Galgal et Masphat et iudicabat Israhelem in supradictis locis
1SAM|7|17|revertebaturque in Ramatha ibi enim erat domus eius et ibi iudicabat Israhelem aedificavit etiam ibi altare Domino
1SAM|8|1|factum est autem cum senuisset Samuhel posuit filios suos iudices Israhel
1SAM|8|2|fuitque nomen filii eius primogeniti Iohel et nomen secundi Abia iudicum in Bersabee
1SAM|8|3|et non ambulaverunt filii illius in viis eius sed declinaverunt post avaritiam acceperuntque munera et perverterunt iudicium
1SAM|8|4|congregati ergo universi maiores natu Israhel venerunt ad Samuhel in Ramatha
1SAM|8|5|dixeruntque ei ecce tu senuisti et filii tui non ambulant in viis tuis constitue nobis regem ut iudicet nos sicut universae habent nationes
1SAM|8|6|displicuitque sermo in oculis Samuhelis eo quod dixissent da nobis regem ut iudicet nos et oravit Samuhel Dominum
1SAM|8|7|dixit autem Dominus ad Samuhel audi vocem populi in omnibus quae loquuntur tibi non enim te abiecerunt sed me ne regnem super eos
1SAM|8|8|iuxta omnia opera sua quae fecerunt a die qua eduxi eos de Aegypto usque ad diem hanc sicut dereliquerunt me et servierunt diis alienis sic faciunt etiam tibi
1SAM|8|9|nunc ergo audi vocem eorum verumtamen contestare eos et praedic eis ius regis qui regnaturus est super eos
1SAM|8|10|dixit itaque Samuhel omnia verba Domini ad populum qui petierat a se regem
1SAM|8|11|et ait hoc erit ius regis qui imperaturus est vobis filios vestros tollet et ponet in curribus suis facietque sibi equites et praecursores quadrigarum suarum
1SAM|8|12|et constituet sibi tribunos et centuriones et aratores agrorum suorum et messores segetum et fabros armorum et curruum suorum
1SAM|8|13|filias quoque vestras faciet sibi unguentarias et focarias et panificas
1SAM|8|14|agros quoque vestros et vineas et oliveta optima tollet et dabit servis suis
1SAM|8|15|sed et segetes vestras et vinearum reditus addecimabit ut det eunuchis et famulis suis
1SAM|8|16|servos etiam vestros et ancillas et iuvenes optimos et asinos auferet et ponet in opere suo
1SAM|8|17|greges vestros addecimabit vosque eritis ei servi
1SAM|8|18|et clamabitis in die illa a facie regis vestri quem elegistis vobis et non exaudiet vos Dominus in die illa
1SAM|8|19|noluit autem populus audire vocem Samuhel sed dixerunt nequaquam rex enim erit super nos
1SAM|8|20|et erimus nos quoque sicut omnes gentes et iudicabit nos rex noster et egredietur ante nos et pugnabit bella nostra pro nobis
1SAM|8|21|et audivit Samuhel omnia verba populi et locutus est ea in auribus Domini
1SAM|8|22|dixit autem Dominus ad Samuhel audi vocem eorum et constitue super eos regem et ait Samuhel ad viros Israhel vadat unusquisque in civitatem suam
1SAM|9|1|et erat vir de Beniamin nomine Cis filius Abihel filii Seror filii Bechoreth filii Afia filii viri Iemini fortis robore
1SAM|9|2|et erat ei filius vocabulo Saul electus et bonus et non erat vir de filiis Israhel melior illo ab umero et sursum eminebat super omnem populum
1SAM|9|3|perierant autem asinae Cis patris Saul et dixit Cis ad Saul filium suum tolle tecum unum de pueris et consurgens vade et quaere asinas qui cum transissent per montem Ephraim
1SAM|9|4|et per terram Salisa et non invenissent transierunt etiam per terram Salim et non erant sed et per terram Iemini et minime reppererunt
1SAM|9|5|cum autem venissent in terram Suph dixit Saul ad puerum suum qui erat cum eo veni et revertamur ne forte dimiserit pater meus asinas et sollicitus sit pro nobis
1SAM|9|6|qui ait ei ecce est vir Dei in civitate hac vir nobilis omne quod loquitur absque ambiguitate venit nunc ergo eamus illuc si forte indicet nobis de via nostra propter quam venimus
1SAM|9|7|dixitque Saul ad puerum suum ecce ibimus quid feremus ad virum panis defecit in sitarciis nostris et sportulam non habemus ut demus homini Dei nec quicquam aliud
1SAM|9|8|rursum puer respondit Sauli et ait ecce inventa est in manu mea quarta pars stateris argenti demus homini Dei ut indicet nobis viam nostram
1SAM|9|9|olim in Israhel sic loquebatur unusquisque vadens consulere Deum venite et eamus ad videntem qui enim propheta dicitur hodie vocabatur olim videns
1SAM|9|10|et dixit Saul ad puerum suum optimus sermo tuus veni eamus et ierunt in civitatem in qua erat vir Dei
1SAM|9|11|cumque ascenderent clivum civitatis invenerunt puellas egredientes ad hauriendam aquam et dixerunt eis num hic est videns
1SAM|9|12|quae respondentes dixerunt illis hic est ecce ante te festina nunc hodie enim venit in civitate quia sacrificium est hodie populo in excelso
1SAM|9|13|ingredientes urbem statim invenietis eum antequam ascendat excelsum ad vescendum neque enim comesurus est populus donec ille veniat quia ipse benedicit hostiae et deinceps comedunt qui vocati sunt nunc ergo conscendite quia hodie repperietis eum
1SAM|9|14|et ascenderunt in civitatem cumque illi ambularent in medio urbis apparuit Samuhel egrediens obviam eis ut ascenderet in excelsum
1SAM|9|15|Dominus autem revelaverat auriculam Samuhel ante unam diem quam veniret Saul dicens
1SAM|9|16|hac ipsa quae nunc est hora cras mittam ad te virum de terra Beniamin et ungues eum ducem super populum meum Israhel et salvabit populum meum de manu Philisthinorum quia respexi populum meum venit enim clamor eorum ad me
1SAM|9|17|cumque aspexisset Samuhel Saulem Dominus ait ei ecce vir quem dixeram tibi iste dominabitur populo meo
1SAM|9|18|accessit autem Saul ad Samuhelem in medio portae et ait indica oro mihi ubi est domus videntis
1SAM|9|19|et respondit Samuhel Sauli dicens ego sum videns ascende ante me in excelsum ut comedatis mecum hodie et dimittam te mane et omnia quae sunt in corde tuo indicabo tibi
1SAM|9|20|et de asinis quas perdidisti nudius tertius ne sollicitus sis quia inventae sunt et cuius erunt optima quaeque Israhel nonne tibi et omni domui patris tui
1SAM|9|21|respondens autem Saul ait numquid non filius Iemini ego sum de minima tribu Israhel et cognatio mea novissima inter omnes familias de tribu Beniamin quare ergo locutus es mihi sermonem istum
1SAM|9|22|adsumens itaque Samuhel Saulem et puerum eius introduxit eos in triclinium et dedit eis locum in capite eorum qui fuerant invitati erant enim quasi triginta viri
1SAM|9|23|dixitque Samuhel coco da partem quam dedi tibi et praecepi ut reponeres seorsum apud te
1SAM|9|24|levavit autem cocus armum et posuit ante Saul dixitque Samuhel ecce quod remansit pone ante te et comede quia de industria servatum est tibi quando populum vocavi et comedit Saul cum Samuhel in die illa
1SAM|9|25|et descenderunt de excelso in oppidum et locutus est cum Saul in solario
1SAM|9|26|cumque mane surrexissent et iam dilucesceret vocavit Samuhel Saul in solarium dicens surge ut dimittam te et surrexit Saul egressique sunt ambo ipse videlicet et Samuhel
1SAM|9|27|cumque descenderent in extrema parte civitatis Samuhel dixit ad Saul dic puero ut antecedat nos et transeat tu autem subsiste paulisper ut indicem tibi verbum Domini
1SAM|10|1|tulit autem Samuhel lenticulam olei et effudit super caput eius et deosculatus eum ait ecce unxit te Dominus super hereditatem suam in principem
1SAM|10|2|cum abieris hodie a me invenies duos viros iuxta sepulchrum Rachel in finibus Beniamin in meridie dicentque tibi inventae sunt asinae ad quas ieras perquirendas et intermissis pater tuus asinis sollicitus est pro vobis et dicit quid faciam de filio meo
1SAM|10|3|cumque abieris inde et ultra transieris et veneris ad quercum Thabor invenient te ibi tres viri ascendentes ad Deum in Bethel unus portans tres hedos et alius tres tortas panis et alius portans lagoenam vini
1SAM|10|4|cumque te salutaverint dabunt tibi duos panes et accipies de manu eorum
1SAM|10|5|post haec venies in collem Domini ubi est statio Philisthinorum et cum ingressus fueris ibi urbem obviam habebis gregem prophetarum descendentium de excelso et ante eos psalterium et tympanum et tibiam et citharam ipsosque prophetantes
1SAM|10|6|et insiliet in te spiritus Domini et prophetabis cum eis et mutaberis in virum alium
1SAM|10|7|quando ergo evenerint signa haec omnia tibi fac quaecumque invenerit manus tua quia Dominus tecum est
1SAM|10|8|et descendes ante me in Galgala ego quippe descendam ad te ut offeras oblationem et immoles victimas pacificas septem diebus expectabis donec veniam ad te et ostendam tibi quae facias
1SAM|10|9|itaque cum avertisset umerum suum ut abiret a Samuhele inmutavit ei Deus cor aliud et venerunt omnia signa haec in die illa
1SAM|10|10|veneruntque ad praedictum collem et ecce cuneus prophetarum obvius ei et insilivit super eum spiritus Dei et prophetavit in medio eorum
1SAM|10|11|videntes autem omnes qui noverant eum heri et nudius tertius quod esset cum prophetis et prophetaret dixerunt ad invicem quaenam res accidit filio Cis num et Saul in prophetis
1SAM|10|12|responditque alius ad alterum dicens et quis pater eorum propterea versum est in proverbium num et Saul inter prophetas
1SAM|10|13|cessavit autem prophetare et venit ad excelsum
1SAM|10|14|dixitque patruus Saul ad eum et ad puerum eius quo abistis qui responderunt quaerere asinas quas cum non repperissemus venimus ad Samuhelem
1SAM|10|15|et dixit ei patruus suus indica mihi quid dixerit tibi Samuhel
1SAM|10|16|et ait Saul ad patruum suum indicavit nobis quia inventae essent asinae de sermone autem regni non indicavit ei quem locutus illi fuerat Samuhel
1SAM|10|17|et convocavit Samuhel populum ad Dominum in Maspha
1SAM|10|18|et ait ad filios Israhel haec dicit Dominus Deus Israhel ego eduxi Israhel de Aegypto et erui vos de manu Aegyptiorum et de manu omnium regum qui adfligebant vos
1SAM|10|19|vos autem hodie proiecistis Deum vestrum qui solus salvavit vos de universis malis et tribulationibus vestris et dixistis nequaquam sed regem constitue super nos nunc ergo state coram Domino per tribus vestras et per familias
1SAM|10|20|et adplicuit Samuhel omnes tribus Israhel et cecidit sors tribus Beniamin
1SAM|10|21|et adplicuit tribum Beniamin et cognationes eius et cecidit cognatio Metri et pervenit usque ad Saul filium Cis quaesierunt ergo eum et non est inventus
1SAM|10|22|et consuluerunt post haec Dominum utrumnam venturus esset illuc responditque Dominus ecce absconditus est domi
1SAM|10|23|cucurrerunt itaque et tulerunt eum inde stetitque in medio populi et altior fuit universo populo ab umero et sursum
1SAM|10|24|et ait Samuhel ad omnem populum certe videtis quem elegit Dominus quoniam non sit similis ei in omni populo et clamavit cunctus populus et ait vivat rex
1SAM|10|25|locutus est autem Samuhel ad populum legem regni et scripsit in libro et reposuit coram Domino et dimisit Samuhel omnem populum singulos in domum suam
1SAM|10|26|sed et Saul abiit in domum suam in Gabaath et abiit cum eo pars exercitus quorum tetigerat Deus corda
1SAM|10|27|filii vero Belial dixerunt num salvare nos poterit iste et despexerunt eum et non adtulerunt ei munera ille vero dissimulabat se audire
1SAM|11|1|ascendit autem Naas Ammonites et pugnare coepit adversus Iabesgalaad dixeruntque omnes viri Iabes ad Naas habeto nos foederatos et serviemus tibi
1SAM|11|2|et respondit ad eos Naas Ammonites in hoc feriam vobiscum foedus ut eruam omnium vestrum oculos dextros ponamque vos obprobrium in universo Israhel
1SAM|11|3|et dixerunt ad eum seniores Iabes concede nobis septem dies ut mittamus nuntios in universos terminos Israhel et si non fuerit qui defendat nos egrediemur ad te
1SAM|11|4|venerunt ergo nuntii in Gabaath Saulis et locuti sunt verba audiente populo et levavit omnis populus vocem suam et flevit
1SAM|11|5|et ecce Saul veniebat sequens boves de agro et ait quid habet populus quod plorat et narraverunt ei verba virorum Iabes
1SAM|11|6|et insilivit spiritus Domini in Saul cum audisset verba haec et iratus est furor eius nimis
1SAM|11|7|et adsumens utrumque bovem concidit in frusta misitque in omnes terminos Israhel per manum nuntiorum dicens quicumque non exierit secutusque fuerit Saul et Samuhelem sic fiet bubus eius invasit ergo timor Domini populum et egressi sunt quasi vir unus
1SAM|11|8|et recensuit eos in Bezec fueruntque filiorum Israhel trecenta milia virorum autem Iuda triginta milia
1SAM|11|9|et dixerunt nuntiis qui venerant sic dicetis viris qui sunt in Iabesgalaad cras erit vobis salus cum incaluerit sol venerunt ergo nuntii et adnuntiaverunt viris Iabes qui laetati sunt
1SAM|11|10|et dixerunt mane exibimus ad vos et facietis nobis omne quod placuerit vobis
1SAM|11|11|et factum est cum venisset dies crastinus constituit Saul populum in tres partes et ingressus est media castra in vigilia matutina et percussit Ammon usque dum incalesceret dies reliqui autem dispersi sunt ita ut non relinquerentur in eis duo pariter
1SAM|11|12|et ait populus ad Samuhel quis est iste qui dixit Saul non regnabit super nos date viros et interficiemus eos
1SAM|11|13|et ait Saul non occidetur quisquam in die hac quia hodie fecit Dominus salutem in Israhel
1SAM|11|14|dixit autem Samuhel ad populum venite et eamus in Galgala et innovemus ibi regnum
1SAM|11|15|et perrexit omnis populus in Galgala et fecerunt ibi regem Saul coram Domino in Galgala et immolaverunt ibi victimas pacificas coram Domino et laetatus est ibi Saul et cuncti viri Israhel nimis
1SAM|12|1|dixit autem Samuhel ad universum Israhel ecce audivi vocem vestram iuxta omnia quae locuti estis ad me et constitui super vos regem
1SAM|12|2|et nunc rex graditur ante vos ego autem senui et incanui porro filii mei vobiscum sunt itaque conversatus coram vobis ab adulescentia mea usque ad diem hanc ecce praesto sum
1SAM|12|3|loquimini de me coram Domino et coram christo eius utrum bovem cuiusquam tulerim an asinum si quempiam calumniatus sum si oppressi aliquem si de manu cuiusquam munus accepi et contemnam illud hodie restituamque vobis
1SAM|12|4|et dixerunt non es calumniatus nos neque oppressisti neque tulisti de manu alicuius quippiam
1SAM|12|5|dixitque ad eos testis Dominus adversus vos et testis christus eius in die hac quia non inveneritis in manu mea quippiam et dixerunt testis
1SAM|12|6|et ait Samuhel ad populum Dominus qui fecit Mosen et Aaron et eduxit patres nostros de terra Aegypti
1SAM|12|7|nunc ergo state ut iudicio contendam adversum vos coram Domino de omnibus misericordiis Domini quas fecit vobiscum et cum patribus vestris
1SAM|12|8|quomodo ingressus est Iacob in Aegyptum et clamaverunt patres vestri ad Dominum et misit Dominus Mosen et Aaron et eduxit patres vestros ex Aegypto et conlocavit eos in loco hoc
1SAM|12|9|qui obliti sunt Domini Dei sui et tradidit eos in manu Sisarae magistri militiae Asor et in manu Philisthinorum et in manu regis Moab et pugnaverunt adversum eos
1SAM|12|10|postea autem clamaverunt ad Dominum et dixerunt peccavimus quia dereliquimus Dominum et servivimus Baalim et Astharoth nunc ergo erue nos de manu inimicorum nostrorum et serviemus tibi
1SAM|12|11|et misit Dominus Hierobaal et Bedan et Ieptha et Samuhel et eruit vos de manu inimicorum vestrorum per circuitum et habitastis confidenter
1SAM|12|12|videntes autem quod Naas rex filiorum Ammon venisset adversum vos dixistis mihi nequaquam sed rex imperabit nobis cum Dominus Deus vester regnaret in vobis
1SAM|12|13|nunc ergo praesto est rex vester quem elegistis et petistis ecce dedit vobis Dominus regem
1SAM|12|14|si timueritis Dominum et servieritis ei et audieritis vocem eius et non exasperaveritis os Domini eritis et vos et rex qui imperat vobis sequentes Dominum Deum vestrum
1SAM|12|15|si autem non audieritis vocem Domini sed exasperaveritis sermonem Domini erit manus Domini super vos et super patres vestros
1SAM|12|16|sed et nunc state et videte rem istam grandem quam facturus est Dominus in conspectu vestro
1SAM|12|17|numquid non messis tritici est hodie invocabo Dominum et dabit voces et pluvias et scietis et videbitis quia grande malum feceritis vobis in conspectu Domini petentes super vos regem
1SAM|12|18|et clamavit Samuhel ad Dominum et dedit Dominus voces et pluviam in die illa
1SAM|12|19|et timuit omnis populus nimis Dominum et Samuhelem dixitque universus populus ad Samuhel ora pro servis tuis ad Dominum Deum tuum ut non moriamur addidimus enim universis peccatis nostris malum ut peteremus nobis regem
1SAM|12|20|dixit autem Samuhel ad populum nolite timere vos fecistis universum malum hoc verumtamen nolite recedere a tergo Domini et servite Domino in omni corde vestro
1SAM|12|21|et nolite declinare post vana quae non proderunt vobis neque eruent vos quia vana sunt
1SAM|12|22|et non derelinquet Dominus populum suum propter nomen suum magnum quia iuravit Dominus facere vos sibi populum
1SAM|12|23|absit autem a me hoc peccatum in Domino ut cessem orare pro vobis et docebo vos viam bonam et rectam
1SAM|12|24|igitur timete Dominum et servite ei in veritate et ex toto corde vestro vidistis enim magnifica quae in vobis gesserit
1SAM|12|25|quod si perseveraveritis in malitia et vos et rex vester pariter peribitis
1SAM|13|1|filius unius anni Saul cum regnare coepisset duobus autem annis regnavit super Israhel
1SAM|13|2|et elegit sibi Saul tria milia de Israhel et erant cum Saul duo milia in Machmas et in monte Bethel mille autem cum Ionathan in Gabaath Beniamin porro ceterum populum remisit unumquemque in tabernacula sua
1SAM|13|3|et percussit Ionathan stationem Philisthim quae erat in Gabaa quod cum audissent Philisthim Saul cecinit bucina in omni terra dicens audiant Hebraei
1SAM|13|4|et universus Israhel audivit huiuscemodi famam percussit Saul stationem Philisthinorum et erexit se Israhel adversum Philisthim clamavit ergo populus post Saul in Galgala
1SAM|13|5|et Philisthim congregati sunt ad proeliandum contra Israhel triginta milia curruum et sex milia equitum et reliquum vulgus sicut harena quae est in litore maris plurima et ascendentes castrametati sunt in Machmas ad orientem Bethaven
1SAM|13|6|quod cum vidissent viri Israhel se in arto sitos adflictus est enim populus absconderunt se in speluncis et in abditis in petris quoque et in antris et in cisternis
1SAM|13|7|Hebraei autem transierunt Iordanem terram Gad et Galaad cumque adhuc esset Saul in Galgal universus populus perterritus est qui sequebatur eum
1SAM|13|8|et expectavit septem diebus iuxta placitum Samuhel et non venit Samuhel in Galgala dilapsusque est populus ab eo
1SAM|13|9|ait ergo Saul adferte mihi holocaustum et pacifica et obtulit holocaustum
1SAM|13|10|cumque conplesset offerens holocaustum ecce Samuhel veniebat et egressus est Saul obviam ei ut salutaret eum
1SAM|13|11|locutusque est ad eum Samuhel quid fecisti respondit Saul quia vidi quod dilaberetur populus a me et tu non veneras iuxta placitos dies porro Philisthim congregati fuerant in Machmas
1SAM|13|12|dixi nunc descendent Philisthim ad me in Galgala et faciem Domini non placavi necessitate conpulsus obtuli holocaustum
1SAM|13|13|dixitque Samuhel ad Saul stulte egisti nec custodisti mandata Domini Dei tui quae praecepit tibi quod si non fecisses iam nunc praeparasset Dominus regnum tuum super Israhel in sempiternum
1SAM|13|14|sed nequaquam regnum tuum ultra consurget quaesivit sibi Dominus virum iuxta cor suum et praecepit ei Dominus ut esset dux super populum suum eo quod non servaveris quae praecepit Dominus
1SAM|13|15|surrexit autem Samuhel et ascendit de Galgalis in Gabaa Beniamin et recensuit Saul populum qui inventi fuerant cum eo quasi sescentos viros
1SAM|13|16|et Saul et Ionathan filius eius populusque qui inventus fuerat cum eis erat in Gabaa Beniamin porro Philisthim consederant in Machmas
1SAM|13|17|et egressi sunt ad praedandum de castris Philisthim tres cunei unus cuneus pergebat contra viam Ephra ad terram Saul
1SAM|13|18|porro alius ingrediebatur per viam Bethoron tertius autem verterat se ad iter termini inminentis valli Seboim contra desertum
1SAM|13|19|porro faber ferrarius non inveniebatur in omni terra Israhel caverant enim Philisthim ne forte facerent Hebraei gladium aut lanceam
1SAM|13|20|descendebat ergo omnis Israhel ad Philisthim ut exacueret unusquisque vomerem suum et ligonem et securim et sarculum
1SAM|13|21|retunsae itaque erant acies vomerum et ligonum et tridentum et securium usque ad stimulum corrigendum
1SAM|13|22|cumque venisset dies proelii non est inventus ensis et lancea in manu totius populi qui erat cum Saul et cum Ionathan excepto Saul et Ionathan filio eius
1SAM|13|23|egressa est autem statio Philisthim ut transcenderet in Machmas
1SAM|14|1|et accidit quadam die ut diceret Ionathan filius Saul ad adulescentem armigerum suum veni et transeamus ad stationem Philisthim quae est trans locum illum patri autem suo hoc ipsum non indicavit
1SAM|14|2|porro Saul morabatur in extrema parte Gabaa sub malogranato quae erat in Magron et erat populus cum eo quasi sescentorum virorum
1SAM|14|3|et Ahias filius Achitob fratris Ichabod filii Finees qui ortus fuerat ex Heli sacerdote Domini in Silo portabat ephod sed et populus ignorabat quod isset Ionathan
1SAM|14|4|erant autem inter ascensus per quos nitebatur Ionathan transire ad stationem Philisthinorum eminentes petrae ex utraque parte et quasi in modum dentium scopuli hinc inde praerupti nomen uni Boses et nomen alteri Sene
1SAM|14|5|unus scopulus prominens ad aquilonem ex adverso Machmas et alter a meridie contra Gabaa
1SAM|14|6|dixit autem Ionathan ad adulescentem armigerum suum veni transeamus ad stationem incircumcisorum horum si forte faciat Dominus pro nobis quia non est Domino difficile salvare vel in multitudine vel in paucis
1SAM|14|7|dixitque ei armiger suus fac omnia quae placent animo tuo perge quo cupis ero tecum ubicumque volueris
1SAM|14|8|et ait Ionathan ecce nos transimus ad viros istos cumque apparuerimus eis
1SAM|14|9|si taliter locuti fuerint ad nos manete donec veniamus ad vos stemus in loco nostro nec ascendamus ad eos
1SAM|14|10|si autem dixerint ascendite ad nos ascendamus quia tradidit eos Dominus in manibus nostris hoc erit nobis signum
1SAM|14|11|apparuit igitur uterque stationi Philisthinorum dixeruntque Philisthim en Hebraei egrediuntur de cavernis in quibus absconditi fuerant
1SAM|14|12|et locuti sunt viri de statione ad Ionathan et ad armigerum eius dixeruntque ascendite ad nos et ostendimus vobis rem et ait Ionathan ad armigerum suum ascendamus sequere me tradidit enim eos Dominus in manu Israhel
1SAM|14|13|ascendit autem Ionathan reptans manibus et pedibus et armiger eius post eum itaque alii cadebant ante Ionathan alios armiger eius interficiebat sequens eum
1SAM|14|14|et facta est plaga prima quam percussit Ionathan et armiger eius quasi viginti virorum in media parte iugeri quam par boum in die arare consuevit
1SAM|14|15|et factum est miraculum in castris per agros sed et omnis populus stationis eorum qui ierant ad praedandum obstipuit et conturbata est terra et accidit quasi miraculum a Deo
1SAM|14|16|et respexerunt speculatores Saul qui erant in Gabaa Beniamin et ecce multitudo prostrata et huc illucque diffugiens
1SAM|14|17|et ait Saul populo qui erat cum eo requirite et videte quis abierit ex nobis cumque requisissent reppertum est non adesse Ionathan et armigerum eius
1SAM|14|18|et ait Saul ad Ahiam adplica arcam Dei erat enim ibi arca Dei in die illa cum filiis Israhel
1SAM|14|19|cumque loqueretur Saul ad sacerdotem tumultus magnus exortus est in castris Philisthinorum crescebatque paulatim et clarius reboabat et ait Saul ad sacerdotem contrahe manum tuam
1SAM|14|20|conclamavit ergo Saul et omnis populus qui erat cum eo et venerunt usque ad locum certaminis et ecce versus fuerat gladius uniuscuiusque ad proximum suum et caedes magna nimis
1SAM|14|21|sed et Hebraei qui fuerant cum Philisthim heri et nudius tertius ascenderantque cum eis in castris reversi sunt ut essent cum Israhele qui erant cum Saul et Ionathan
1SAM|14|22|omnes quoque Israhelitae qui se absconderant in monte Ephraim audientes quod fugissent Philisthim sociaverunt se cum suis in proelio
1SAM|14|23|et salvavit Dominus in die illa Israhel pugna autem pervenit usque Bethaven
1SAM|14|24|et vir Israhel sociatus sibi est in die illa adiuravit autem Saul populum dicens maledictus vir qui comederit panem usque ad vesperam donec ulciscar de inimicis meis et non manducavit universus populus panem
1SAM|14|25|omneque terrae vulgus venit in saltum in quo erat mel super faciem agri
1SAM|14|26|ingressus est itaque populus saltum et apparuit fluens mel nullusque adplicuit manum ad os suum timebat enim populus iuramentum
1SAM|14|27|porro Ionathan non audierat cum adiuraret pater eius populum extenditque summitatem virgae quam habebat in manu et intinxit in favo mellis et convertit manum suam ad os suum et inluminati sunt oculi eius
1SAM|14|28|respondensque unus de populo ait iureiurando constrinxit pater tuus populum dicens maledictus qui comederit panem hodie defecerat autem populus
1SAM|14|29|dixitque Ionathan turbavit pater meus terram vidistis ipsi quia inluminati sunt oculi mei eo quod gustaverim paululum de melle isto
1SAM|14|30|quanto magis si comedisset populus de praeda inimicorum suorum quam repperit nonne maior facta fuisset plaga in Philisthim
1SAM|14|31|percusserunt ergo in die illa Philistheos a Machmis usque in Ahialon defatigatus est autem populus nimis
1SAM|14|32|et versus ad praedam tulit oves et boves et vitulos et mactaverunt in terra comeditque populus cum sanguine
1SAM|14|33|nuntiaverunt autem Saul dicentes quod populus peccasset Domino comedens cum sanguine qui ait praevaricati estis volvite ad me iam nunc saxum grande
1SAM|14|34|et dixit Saul dispergimini in vulgus et dicite eis ut adducat ad me unusquisque bovem suum et arietem et occidite super istud et vescimini et non peccabitis Domino comedentes cum sanguine adduxit itaque omnis populus unusquisque bovem in manu sua usque ad noctem et occiderunt ibi
1SAM|14|35|aedificavit autem Saul altare Domini tuncque primum coepit aedificare altare Domini
1SAM|14|36|et dixit Saul inruamus super Philisthim nocte et vastemus eos usque dum inlucescat mane nec relinquamus de eis virum dixitque populus omne quod bonum videtur in oculis tuis fac et ait sacerdos accedamus huc ad Deum
1SAM|14|37|et consuluit Saul Deum num persequar Philisthim si trades eos in manu Israhel et non respondit ei in die illa
1SAM|14|38|dixitque Saul adplicate huc universos angulos populi et scitote et videte per quem acciderit peccatum hoc hodie
1SAM|14|39|vivit Dominus salvator Israhel quia si per Ionathan filium meum factum est absque retractatione morietur ad quod nullus contradixit ei de omni populo
1SAM|14|40|et ait ad universum Israhel separamini vos in partem unam et ego cum Ionathan filio meo ero in parte una respondit populus ad Saul quod bonum videtur in oculis tuis fac
1SAM|14|41|et dixit Saul ad Dominum Deum Israhel da indicium et deprehensus est Ionathan et Saul populus autem exivit
1SAM|14|42|et ait Saul mittite sortem inter me et inter Ionathan filium meum et captus est Ionathan
1SAM|14|43|dixit autem Saul ad Ionathan indica mihi quid feceris et indicavit ei Ionathan et ait gustans gustavi in summitate virgae quae erat in manu mea paululum mellis et ecce ego morior
1SAM|14|44|et ait Saul haec faciat mihi Deus et haec addat quia morte morieris Ionathan
1SAM|14|45|dixitque populus ad Saul ergone Ionathan morietur qui fecit salutem hanc magnam in Israhel hoc nefas est vivit Dominus si ceciderit capillus de capite eius in terram quia cum Deo operatus est hodie liberavit ergo populus Ionathan ut non moreretur
1SAM|14|46|recessitque Saul nec persecutus est Philisthim porro Philisthim abierunt in loca sua
1SAM|14|47|at Saul confirmato regno super Israhel pugnabat per circuitum adversum omnes inimicos eius contra Moab et filios Ammon et Edom et reges Suba et Philistheos et quocumque se verterat superabat
1SAM|14|48|congregatoque exercitu percussit Amalech et eruit Israhel de manu vastatorum eius
1SAM|14|49|fuerunt autem filii Saul Ionathan et Iesui et Melchisua nomina duarum filiarum eius nomen primogenitae Merob et nomen minoris Michol
1SAM|14|50|et nomen uxoris Saul Ahinoem filia Ahimaas et nomina principum militiae eius Abner filius Ner patruelis Saul
1SAM|14|51|Cis fuerat pater Saul et Ner pater Abner filius Abihel
1SAM|14|52|erat autem bellum potens adversum Philistheos omnibus diebus Saul nam quemcumque viderat Saul virum fortem et aptum ad proelium sociabat eum sibi
1SAM|15|1|et dixit Samuhel ad Saul me misit Dominus ut unguerem te in regem super populum eius Israhel nunc ergo audi vocem Domini
1SAM|15|2|haec dicit Dominus exercituum recensui quaecumque fecit Amalech Israheli quomodo restitit ei in via cum ascenderet de Aegypto
1SAM|15|3|nunc igitur vade et percute Amalech et demolire universa eius non parcas ei sed interfice a viro usque ad mulierem et parvulum atque lactantem bovem et ovem camelum et asinum
1SAM|15|4|praecepit itaque Saul populo et recensuit eos quasi agnos ducenta milia peditum et decem milia virorum Iuda
1SAM|15|5|cumque venisset Saul usque ad civitatem Amalech tetendit insidias in torrente
1SAM|15|6|dixitque Saul Cineo abite recedite atque descendite ab Amalech ne forte involvam te cum eo tu enim fecisti misericordiam cum omnibus filiis Israhel cum ascenderent de Aegypto et recessit Cineus de medio Amalech
1SAM|15|7|percussitque Saul Amalech ab Evila donec venias Sur quae est e regione Aegypti
1SAM|15|8|et adprehendit Agag regem Amalech vivum omne autem vulgus interfecit in ore gladii
1SAM|15|9|et pepercit Saul et populus Agag et optimis gregibus ovium et armentorum et vestibus et arietibus et universis quae pulchra erant nec voluerunt disperdere ea quicquid vero vile fuit et reprobum hoc demoliti sunt
1SAM|15|10|factum est autem verbum Domini ad Samuhel dicens
1SAM|15|11|paenitet me quod constituerim Saul regem quia dereliquit me et verba mea opere non implevit contristatusque est Samuhel et clamavit ad Dominum tota nocte
1SAM|15|12|cumque de nocte surrexisset Samuhel ut iret ad Saul mane nuntiatum est Samuheli eo quod venisset Saul in Carmelum et erexisset sibi fornicem triumphalem et reversus transisset descendissetque in Galgala venit ergo Samuhel ad Saul et
1SAM|15|13|dixit ei Saul benedictus tu Domino implevi verbum Domini
1SAM|15|14|dixitque Samuhel et quae est haec vox gregum quae resonat in auribus meis et armentorum quam ego audio
1SAM|15|15|et ait Saul de Amalech adduxerunt ea pepercit enim populus melioribus ovibus et armentis ut immolarentur Domino Deo tuo reliqua vero occidimus
1SAM|15|16|dixit autem Samuhel ad Saul sine me et indicabo tibi quae locutus sit Dominus ad me nocte dixitque ei loquere
1SAM|15|17|et ait Samuhel nonne cum parvulus esses in oculis tuis caput in tribubus Israhel factus es unxitque te Dominus regem super Israhel
1SAM|15|18|et misit te Dominus in via et ait vade et interfice peccatores Amalech et pugnabis contra eos usque ad internicionem eorum
1SAM|15|19|quare ergo non audisti vocem Domini sed versus ad praedam es et fecisti malum in oculis Domini
1SAM|15|20|et ait Saul ad Samuhelem immo audivi vocem Domini et ambulavi in via per quam misit me Dominus et adduxi Agag regem Amalech et Amalech interfeci
1SAM|15|21|tulit autem populus de praeda oves et boves primitias eorum quae caesa sunt ut immolet Domino Deo suo in Galgalis
1SAM|15|22|et ait Samuhel numquid vult Dominus holocausta aut victimas et non potius ut oboediatur voci Domini melior est enim oboedientia quam victimae et auscultare magis quam offerre adipem arietum
1SAM|15|23|quoniam quasi peccatum ariolandi est repugnare et quasi scelus idolatriae nolle adquiescere pro eo ergo quod abiecisti sermonem Domini abiecit te ne sis rex
1SAM|15|24|dixitque Saul ad Samuhel peccavi quia praevaricatus sum sermonem Domini et verba tua timens populum et oboediens voci eorum
1SAM|15|25|sed nunc porta quaeso peccatum meum et revertere mecum ut adorem Dominum
1SAM|15|26|et ait Samuhel ad Saul non revertar tecum quia proiecisti sermonem Domini et proiecit te Dominus ne sis rex super Israhel
1SAM|15|27|et conversus est Samuhel ut abiret ille autem adprehendit summitatem pallii eius quae et scissa est
1SAM|15|28|et ait ad eum Samuhel scidit Dominus regnum Israhel a te hodie et tradidit illud proximo tuo meliori te
1SAM|15|29|porro Triumphator in Israhel non parcet et paenitudine non flectetur neque enim homo est ut agat paenitentiam
1SAM|15|30|at ille ait peccavi sed nunc honora me coram senibus populi mei et coram Israhel et revertere mecum ut adorem Dominum Deum tuum
1SAM|15|31|reversus ergo Samuhel secutus est Saulem et adoravit Saul Dominum
1SAM|15|32|dixitque Samuhel adducite ad me Agag regem Amalech et oblatus est ei Agag pinguissimus et dixit Agag sicine separat amara mors
1SAM|15|33|et ait Samuhel sicut fecit absque liberis mulieres gladius tuus sic absque liberis erit inter mulieres mater tua et in frusta concidit Samuhel Agag coram Domino in Galgalis
1SAM|15|34|abiit autem Samuhel in Ramatha Saul vero ascendit in domum suam in Gabaath
1SAM|15|35|et non vidit Samuhel ultra Saul usque ad diem mortis suae verumtamen lugebat Samuhel Saul quoniam Dominum paenitebat quod constituisset regem Saul super Israhel
1SAM|16|1|dixitque Dominus ad Samuhel usquequo tu luges Saul cum ego proiecerim eum ne regnet super Israhel imple cornu tuum oleo et veni ut mittam te ad Isai Bethleemitem providi enim in filiis eius mihi regem
1SAM|16|2|et ait Samuhel quomodo vadam audiet enim Saul et interficiet me et ait Dominus vitulum de armento tolles in manu tua et dices ad immolandum Domino veni
1SAM|16|3|et vocabis Isai ad victimam et ego ostendam tibi quid facias et ungues quemcumque monstravero tibi
1SAM|16|4|fecit ergo Samuhel sicut locutus est ei Dominus venitque in Bethleem et admirati sunt seniores civitatis occurrentes ei dixeruntque pacificus ingressus tuus
1SAM|16|5|et ait pacificus ad immolandum Domino veni sanctificamini et venite mecum ut immolem sanctificavit ergo Isai et filios eius et vocavit eos ad sacrificium
1SAM|16|6|cumque ingressi essent vidit Heliab et ait num coram Domino est christus eius
1SAM|16|7|et dixit Dominus ad Samuhel ne respicias vultum eius neque altitudinem staturae eius quoniam abieci eum nec iuxta intuitum hominis iudico homo enim videt ea quae parent Dominus autem intuetur cor
1SAM|16|8|et vocavit Isai Abinadab et adduxit eum coram Samuhel qui dixit nec hunc elegit Dominus
1SAM|16|9|adduxit autem Isai Samma de quo ait etiam hunc non elegit Dominus
1SAM|16|10|adduxit itaque Isai septem filios suos coram Samuhel et ait Samuhel ad Isai non elegit Dominus ex istis
1SAM|16|11|dixitque Samuhel ad Isai numquid iam conpleti sunt filii qui respondit adhuc reliquus est parvulus et pascit oves et ait Samuhel ad Isai mitte et adduc eum nec enim discumbemus priusquam ille huc venerit
1SAM|16|12|misit ergo et adduxit eum erat autem rufus et pulcher aspectu decoraque facie et ait Dominus surge ungue eum ipse est enim
1SAM|16|13|tulit igitur Samuhel cornu olei et unxit eum in medio fratrum eius et directus est spiritus Domini in David a die illa et in reliquum surgensque Samuhel abiit in Ramatha
1SAM|16|14|spiritus autem Domini recessit a Saul et exagitabat eum spiritus nequam a Domino
1SAM|16|15|dixeruntque servi Saul ad eum ecce spiritus Dei malus exagitat te
1SAM|16|16|iubeat dominus noster et servi tui qui coram te sunt quaerant hominem scientem psallere cithara ut quando arripuerit te spiritus Dei malus psallat manu sua et levius feras
1SAM|16|17|et ait Saul ad servos suos providete mihi aliquem bene psallentem et adducite eum ad me
1SAM|16|18|et respondens unus de pueris ait ecce vidi filium Isai Bethleemitem scientem psallere et fortissimum robore et virum bellicosum et prudentem in verbis et virum pulchrum et Dominus est cum eo
1SAM|16|19|misit ergo Saul nuntios ad Isai dicens mitte ad me David filium tuum qui est in pascuis
1SAM|16|20|tulitque Isai asinum plenum panibus et lagoenam vini et hedum de capris unum et misit per manum David filii sui Saul
1SAM|16|21|et venit David ad Saul et stetit coram eo at ille dilexit eum nimis et factus est eius armiger
1SAM|16|22|misitque Saul ad Isai dicens stet David in conspectu meo invenit enim gratiam in oculis meis
1SAM|16|23|igitur quandocumque spiritus Dei arripiebat Saul tollebat David citharam et percutiebat manu sua et refocilabatur Saul et levius habebat recedebat enim ab eo spiritus malus
1SAM|17|1|congregantes vero Philisthim agmina sua in proelium convenerunt in Soccho Iudae et castrametati sunt inter Soccho et Azeca in finibus Dommim
1SAM|17|2|porro Saul et viri Israhel congregati venerunt in valle Terebinthi et direxerunt aciem ad pugnandum contra Philisthim
1SAM|17|3|et Philisthim stabant super montem ex hac parte et Israhel stabat super montem ex altera parte vallisque erat inter eos
1SAM|17|4|et egressus est vir spurius de castris Philisthinorum nomine Goliath de Geth altitudinis sex cubitorum et palmo
1SAM|17|5|et cassis aerea super caput eius et lorica hamata induebatur porro pondus loricae eius quinque milia siclorum aeris
1SAM|17|6|et ocreas aereas habebat in cruribus et clypeus aereus tegebat umeros eius
1SAM|17|7|hastile autem hastae eius erat quasi liciatorium texentium ipsum autem ferrum hastae eius sescentos siclos habebat ferri et armiger eius antecedebat eum
1SAM|17|8|stansque clamabat adversum falangas Israhel et dicebat eis quare venitis parati ad proelium numquid ego non sum Philistheus et vos servi Saul eligite ex vobis virum et descendat ad singulare certamen
1SAM|17|9|si quiverit pugnare mecum et percusserit me erimus vobis servi si autem ego praevaluero et percussero eum vos servi eritis et servietis nobis
1SAM|17|10|et aiebat Philistheus ego exprobravi agminibus Israhelis hodie date mihi virum et ineat mecum singulare certamen
1SAM|17|11|audiens autem Saul et omnes viri israhelitae sermones Philisthei huiuscemodi stupebant et metuebant nimis
1SAM|17|12|David autem erat filius viri ephrathei de quo supra dictum est de Bethleem Iuda cui erat nomen Isai qui habebat octo filios et erat vir in diebus Saul senex et grandevus inter viros
1SAM|17|13|abierunt autem tres filii eius maiores post Saul in proelium et nomina trium filiorum eius qui perrexerant ad bellum Heliab primogenitus et secundus Abinadab tertiusque Samma
1SAM|17|14|David autem erat minimus tribus ergo maioribus secutis Saulem
1SAM|17|15|abiit David et reversus est a Saul ut pasceret gregem patris sui in Bethleem
1SAM|17|16|procedebat vero Philistheus mane et vespere et stabat quadraginta diebus
1SAM|17|17|dixit autem Isai ad David filium suum accipe fratribus tuis oephi pulentae et decem panes istos et curre in castra ad fratres tuos
1SAM|17|18|et decem formellas casei has deferes ad tribunum et fratres tuos visitabis si recte agant et cum quibus ordinati sint disce
1SAM|17|19|Saul autem et illi et omnes filii Israhel in valle Terebinthi pugnabant adversum Philisthim
1SAM|17|20|surrexit itaque David mane et commendavit gregem custodi et onustus abiit sicut praeceperat ei Isai et venit ad locum Magala et ad exercitum qui egressus ad pugnam vociferatus erat in certamine
1SAM|17|21|direxerat enim aciem Israhel sed et Philisthim ex adverso fuerant praeparati
1SAM|17|22|derelinquens ergo David vasa quae adtulerat sub manu custodis ad sarcinas cucurrit ad locum certaminis et interrogabat si omnia recte agerentur erga fratres suos
1SAM|17|23|cumque adhuc ille loqueretur eis apparuit vir ille spurius ascendens Goliath nomine Philistheus de Geth ex castris Philisthinorum et loquente eo haec eadem verba audivit David
1SAM|17|24|omnes autem Israhelitae cum vidissent virum fugerunt a facie eius timentes eum valde
1SAM|17|25|et dixit unus quispiam de Israhel num vidisti virum hunc qui ascendit ad exprobrandum enim Israheli ascendit virum ergo qui percusserit eum ditabit rex divitiis magnis et filiam suam dabit ei et domum patris eius faciet absque tributo in Israhel
1SAM|17|26|et ait David ad viros qui stabant secum dicens quid dabitur viro qui percusserit Philistheum hunc et tulerit obprobrium de Israhel quis est enim hic Philistheus incircumcisus qui exprobravit acies Dei viventis
1SAM|17|27|referebat autem ei populus eundem sermonem dicens haec dabuntur viro qui percusserit eum
1SAM|17|28|quod cum audisset Heliab frater eius maior loquente eo cum aliis iratus est contra David et ait quare venisti et quare dereliquisti pauculas oves illas in deserto ego novi superbiam tuam et nequitiam cordis tui quia ut videres proelium descendisti
1SAM|17|29|et dixit David quid feci numquid non verbum est
1SAM|17|30|et declinavit paululum ab eo ad alium dixitque eundem sermonem et respondit ei populus verbum sicut et prius
1SAM|17|31|audita sunt autem verba quae locutus est David et adnuntiata in conspectu Saul
1SAM|17|32|ad quem cum fuisset adductus locutus est ei non concidat cor cuiusquam in eo ego servus tuus vadam et pugnabo adversus Philistheum
1SAM|17|33|et ait Saul ad David non vales resistere Philistheo isti nec pugnare adversum eum quia puer es hic autem vir bellator ab adulescentia sua
1SAM|17|34|dixitque David ad Saul pascebat servus tuus patris sui gregem et veniebat leo vel ursus tollebatque arietem de medio gregis
1SAM|17|35|et sequebar eos et percutiebam eruebamque de ore eorum et illi consurgebant adversum me et adprehendebam mentum eorum et suffocabam interficiebamque eos
1SAM|17|36|nam et leonem et ursum interfeci ego servus tuus erit igitur et Philistheus hic incircumcisus quasi unus ex eis quia ausus est maledicere exercitum Dei viventis
1SAM|17|37|et ait David Dominus qui eruit me de manu leonis et de manu ursi ipse liberabit me de manu Philisthei huius dixit autem Saul ad David vade et Dominus tecum sit
1SAM|17|38|et induit Saul David vestimentis suis et inposuit galeam aeream super caput eius et vestivit eum lorica
1SAM|17|39|accinctus ergo David gladio eius super veste sua coepit temptare si armatus posset incedere non enim habebat consuetudinem dixitque David ad Saul non possum sic incedere quia nec usum habeo et deposuit ea
1SAM|17|40|et tulit baculum suum quem semper habebat in manibus et elegit sibi quinque limpidissimos lapides de torrente et misit eos in peram pastoralem quam habebat secum et fundam manu tulit et processit adversum Philistheum
1SAM|17|41|ibat autem Philistheus incedens et adpropinquans adversum David et armiger eius ante eum
1SAM|17|42|cumque inspexisset Philistheus et vidisset David despexit eum erat enim adulescens rufus et pulcher aspectu
1SAM|17|43|et dixit Philistheus ad David numquid ego canis sum quod tu venis ad me cum baculo et maledixit Philistheus David in diis suis
1SAM|17|44|dixitque ad David veni ad me et dabo carnes tuas volatilibus caeli et bestiis terrae
1SAM|17|45|dixit autem David ad Philistheum tu venis ad me cum gladio et hasta et clypeo ego autem venio ad te in nomine Domini exercituum Dei agminum Israhel quibus exprobrasti
1SAM|17|46|hodie et dabit te Dominus in manu mea et percutiam te et auferam caput tuum a te et dabo cadaver castrorum Philisthim hodie volatilibus caeli et bestiis terrae ut sciat omnis terra quia est Deus in Israhel
1SAM|17|47|et noverit universa ecclesia haec quia non in gladio nec in hasta salvat Dominus ipsius est enim bellum et tradet vos in manus nostras
1SAM|17|48|cum ergo surrexisset Philistheus et veniret et adpropinquaret contra David festinavit David et cucurrit ad pugnam ex adverso Philisthei
1SAM|17|49|et misit manum suam in peram tulitque unum lapidem et funda iecit et percussit Philistheum in fronte et infixus est lapis in fronte eius et cecidit in faciem suam super terram
1SAM|17|50|praevaluitque David adversus Philistheum in funda et in lapide percussumque Philistheum interfecit cumque gladium non haberet in manu David
1SAM|17|51|cucurrit et stetit super Philistheum et tulit gladium eius et eduxit de vagina sua et interfecit eum praeciditque caput eius videntes autem Philisthim quod mortuus esset fortissimus eorum fugerunt
1SAM|17|52|et consurgentes viri Israhel et Iuda vociferati sunt et persecuti Philistheos usque dum venirent in vallem et usque ad portas Accaron cecideruntque vulnerati de Philisthim in via Sarim usque ad Geth et usque Accaron
1SAM|17|53|et revertentes filii Israhel postquam persecuti fuerant Philistheos invaserunt castra eorum
1SAM|17|54|adsumens autem David caput Philisthei adtulit illud in Hierusalem arma vero eius posuit in tabernaculo suo
1SAM|17|55|eo autem tempore quo viderat Saul David egredientem contra Philistheum ait ad Abner principem militiae de qua stirpe descendit hic adulescens Abner dixitque Abner vivit anima tua rex si novi
1SAM|17|56|et ait rex interroga tu cuius filius sit iste puer
1SAM|17|57|cumque regressus esset David percusso Philistheo tulit eum Abner et introduxit coram Saul caput Philisthei habentem in manu
1SAM|17|58|et ait ad eum Saul de qua progenie es o adulescens dixitque David filius servi tui Isai Bethleemitae ego sum
1SAM|18|1|et factum est cum conplesset loqui ad Saul anima Ionathan conligata est animae David et dilexit eum Ionathan quasi animam suam
1SAM|18|2|tulitque eum Saul in die illa et non concessit ei ut reverteretur in domum patris sui
1SAM|18|3|inierunt autem Ionathan et David foedus diligebat enim eum quasi animam suam
1SAM|18|4|nam expoliavit se Ionathan tunicam qua erat vestitus et dedit eam David et reliqua vestimenta sua usque ad gladium et arcum suum et usque ad balteum
1SAM|18|5|egrediebatur quoque David ad omnia quaecumque misisset eum Saul et prudenter se agebat posuitque eum Saul super viros belli et acceptus erat in oculis universi populi maximeque in conspectu famulorum Saul
1SAM|18|6|porro cum reverteretur percusso Philistheo David egressae sunt mulieres de universis urbibus Israhel cantantes chorosque ducentes in occursum Saul regis in tympanis laetitiae et in sistris
1SAM|18|7|et praecinebant mulieres ludentes atque dicentes percussit Saul mille et David decem milia
1SAM|18|8|iratus est autem Saul nimis et displicuit in oculis eius iste sermo dixitque dederunt David decem milia et mihi dederunt mille quid ei superest nisi solum regnum
1SAM|18|9|non rectis ergo oculis Saul aspiciebat David ex die illa et deinceps
1SAM|18|10|post diem autem alteram invasit spiritus Dei malus Saul et prophetabat in medio domus suae David autem psallebat manu sua sicut per singulos dies tenebatque Saul lanceam
1SAM|18|11|et misit eam putans quod configere posset David cum pariete et declinavit David a facie eius secundo
1SAM|18|12|et timuit Saul David eo quod esset Dominus cum eo et a se recessisset
1SAM|18|13|amovit ergo eum Saul a se et fecit eum tribunum super mille viros et egrediebatur et intrabat in conspectu populi
1SAM|18|14|in omnibus quoque viis suis David prudenter agebat et Dominus erat cum eo
1SAM|18|15|vidit itaque Saul quod prudens esset nimis et coepit cavere eum
1SAM|18|16|omnis autem Israhel et Iuda diligebat David ipse enim egrediebatur et ingrediebatur ante eos
1SAM|18|17|dixit autem Saul ad David ecce filia mea maior Merob ipsam dabo tibi uxorem tantummodo esto vir fortis et proeliare bella Domini Saul autem reputabat dicens non sit manus mea in eo sed sit super illum manus Philisthinorum
1SAM|18|18|ait autem David ad Saul quis ego sum aut quae est vita mea aut cognatio patris mei in Israhel ut fiam gener regis
1SAM|18|19|factum est autem tempus cum deberet dari Merob filia Saul David data est Hadrihel Molathitae uxor
1SAM|18|20|dilexit autem Michol filia Saul altera David et nuntiatum est Saul et placuit ei
1SAM|18|21|dixitque Saul dabo eam illi ut fiat ei in scandalum et sit super eum manus Philisthinorum dixit ergo Saul ad David in duabus rebus gener meus eris hodie
1SAM|18|22|et mandavit Saul servis suis loquimini ad David clam me dicentes ecce places regi et omnes servi eius diligunt te nunc ergo esto gener regis
1SAM|18|23|et locuti sunt servi Saul in auribus David omnia verba haec et ait David num parum vobis videtur generum esse regis ego autem sum vir pauper et tenuis
1SAM|18|24|et renuntiaverunt servi Saul dicentes huiuscemodi verba locutus est David
1SAM|18|25|dixit autem Saul sic loquimini ad David non habet necesse rex sponsalia nisi tantum centum praeputia Philisthinorum ut fiat ultio de inimicis regis porro Saul cogitabat tradere David in manibus Philisthinorum
1SAM|18|26|cumque renuntiassent servi eius David verba quae diximus placuit sermo in oculis David ut fieret gener regis
1SAM|18|27|et post dies paucos surgens David abiit cum viris qui sub eo erant et percussis Philisthim ducentis viris adtulit praeputia eorum et adnumeravit ea regi ut esset gener eius dedit itaque ei Saul Michol filiam suam uxorem
1SAM|18|28|et vidit Saul et intellexit quia Dominus esset cum David Michol autem filia Saul diligebat eum
1SAM|18|29|et Saul magis coepit timere David factusque est Saul inimicus David cunctis diebus
1SAM|18|30|et egressi sunt principes Philisthinorum a principio autem egressionis eorum prudentius se gerebat David quam omnes servi Saul et celebre factum est nomen eius nimis
1SAM|19|1|locutus est autem Saul ad Ionathan filium suum et ad omnes servos suos ut occiderent David porro Ionathan filius Saul diligebat David valde
1SAM|19|2|et indicavit Ionathan David dicens quaerit Saul pater meus occidere te quapropter observa te quaeso mane et manebis clam et absconderis
1SAM|19|3|ego autem egrediens stabo iuxta patrem meum in agro ubicumque fueris et ego loquar de te ad patrem meum et quodcumque videro nuntiabo tibi
1SAM|19|4|locutus est ergo Ionathan de David bona ad Saul patrem suum dixitque ad eum ne pecces rex in servum tuum David quia non peccavit tibi et opera eius bona sunt tibi valde
1SAM|19|5|et posuit animam suam in manu sua et percussit Philistheum et fecit Dominus salutem magnam universo Israhel vidisti et laetatus es quare ergo peccas in sanguine innoxio interficiens David qui est absque culpa
1SAM|19|6|quod cum audisset Saul placatus voce Ionathae iuravit vivit Dominus quia non occidetur
1SAM|19|7|vocavit itaque Ionathan David et indicavit ei omnia verba haec et introduxit Ionathan David ad Saul et fuit ante eum sicut fuerat heri et nudius tertius
1SAM|19|8|motum est autem rursus bellum et egressus David pugnavit adversus Philisthim percussitque eos plaga magna et fugerunt a facie eius
1SAM|19|9|et factus est spiritus Domini malus in Saul sedebat autem in domo sua et tenebat lanceam porro David psallebat in manu sua
1SAM|19|10|nisusque est Saul configere lancea David in pariete et declinavit David a facie Saul lancea autem casso vulnere perlata est in parietem et David fugit et salvatus est nocte illa
1SAM|19|11|misit ergo Saul satellites suos in domum David ut custodirent eum et interficeretur mane quod cum adnuntiasset David Michol uxor sua dicens nisi salvaveris te nocte hac cras morieris
1SAM|19|12|deposuit eum per fenestram porro ille abiit et aufugit atque salvatus est
1SAM|19|13|tulit autem Michol statuam et posuit eam super lectum et pellem pilosam caprarum posuit ad caput eius et operuit eam vestimentis
1SAM|19|14|misit autem Saul apparitores qui raperent David et responsum est quod aegrotaret
1SAM|19|15|rursumque misit Saul nuntios ut viderent David dicens adferte eum ad me in lecto ut occidatur
1SAM|19|16|cumque venissent nuntii inventum est simulacrum super lectum et pellis caprarum ad caput eius
1SAM|19|17|dixitque Saul ad Michol quare sic inlusisti mihi et dimisisti inimicum meum ut fugeret et respondit Michol ad Saul quia ipse locutus est mihi dimitte me alioquin interficiam te
1SAM|19|18|David autem fugiens salvatus est et venit ad Samuhel in Ramatha et nuntiavit ei omnia quae fecerat sibi Saul et abierunt ipse et Samuhel et morati sunt in Nahioth
1SAM|19|19|nuntiatum est autem Sauli a dicentibus ecce David in Nahioth in Rama
1SAM|19|20|misit ergo Saul lictores ut raperent David qui cum vidissent cuneum prophetarum vaticinantium et Samuhel stantem super eos factus est etiam in illis spiritus Domini et prophetare coeperunt etiam ipsi
1SAM|19|21|quod cum nuntiatum esset Sauli misit alios nuntios prophetaverunt autem et illi et rursum Saul misit tertios nuntios qui et ipsi prophetaverunt
1SAM|19|22|abiit autem etiam ipse in Ramatha et venit usque ad cisternam magnam quae est in Soccho et interrogavit et dixit in quo loco sunt Samuhel et David dictumque est ei ecce in Nahioth sunt in Rama
1SAM|19|23|et abiit in Nahioth in Rama et factus est etiam super eum spiritus Dei et ambulabat ingrediens et prophetabat usque dum veniret in Nahioth in Rama
1SAM|19|24|et expoliavit se etiam ipse vestimentis suis et prophetavit cum ceteris coram Samuhel et cecidit nudus tota die illa et nocte unde et exivit proverbium num et Saul inter prophetas
1SAM|20|1|fugit autem David de Nahioth quae erat in Rama veniensque locutus est coram Ionathan quid feci quae est iniquitas mea et quod peccatum meum in patrem tuum quia quaerit animam meam
1SAM|20|2|qui dixit ei absit non morieris neque enim faciet pater meus quicquam grande vel parvum nisi prius indicaverit mihi hunc ergo celavit me pater meus sermonem tantummodo nequaquam erit istud
1SAM|20|3|et iuravit rursum David et ille ait scit profecto pater tuus quia inveni gratiam in oculis tuis et dicet nesciat hoc Ionathan ne forte tristetur quinimmo vivit Dominus et vivit anima tua quia uno tantum ut ita dicam gradu ego morsque dividimur
1SAM|20|4|et ait Ionathan ad David quodcumque dixerit mihi anima tua faciam tibi
1SAM|20|5|dixit autem David ad Ionathan ecce kalendae sunt crastino et ego ex more sedere soleo iuxta regem ad vescendum dimitte ergo me ut abscondar in agro usque ad vesperam diei tertiae
1SAM|20|6|si requisierit me pater tuus respondebis ei rogavit me David ut iret celeriter in Bethleem civitatem suam quia victimae sollemnes ibi sunt universis contribulibus eius
1SAM|20|7|si dixerit bene pax erit servo tuo si autem fuerit iratus scito quia conpleta est malitia eius
1SAM|20|8|fac ergo misericordiam in servum tuum quia foedus Domini me famulum tuum tecum inire fecisti si autem est in me aliqua iniquitas tu me interfice et ad patrem tuum ne introducas me
1SAM|20|9|et ait Ionathan absit hoc a te neque enim fieri potest ut si certo cognovero conpletam patris mei esse malitiam contra te non adnuntiem tibi
1SAM|20|10|responditque David ad Ionathan quis nuntiabit mihi si quid forte responderit tibi pater tuus dure
1SAM|20|11|et ait Ionathan ad David veni egrediamur in agrum cumque exissent ambo in agrum
1SAM|20|12|ait Ionathan ad David Domine Deus Israhel si investigavero sententiam patris mei crastino vel perendie et aliquid boni fuerit super David et non statim misero ad te et notum tibi fecero
1SAM|20|13|haec faciat Dominus Ionathan et haec augeat si autem perseveraverit patris mei malitia adversum te revelabo aurem tuam et dimittam te ut vadas in pace et sit Dominus tecum sicut fuit cum patre meo
1SAM|20|14|et si vixero facies mihi misericordiam Domini si vero mortuus fuero
1SAM|20|15|non auferas misericordiam tuam a domo mea usque in sempiternum quando eradicaverit Dominus inimicos David unumquemque de terra
1SAM|20|16|pepigit ergo foedus Ionathan cum domo David et requisivit Dominus de manu inimicorum David
1SAM|20|17|et addidit Ionathan deierare David eo quod diligeret illum sicut animam enim suam ita diligebat eum
1SAM|20|18|dixitque ad eum Ionathan cras kalendae sunt et requireris
1SAM|20|19|requiretur enim sessio tua usque perendie descendes ergo festinus et venies in locum ubi celandus es in die qua operari licet et sedebis iuxta lapidem cui est nomen Ezel
1SAM|20|20|et ego tres sagittas mittam iuxta eum et iaciam quasi exercens me ad signum
1SAM|20|21|mittam quoque et puerum dicens ei vade et adfer mihi sagittas
1SAM|20|22|si dixero puero ecce sagittae intra te sunt tolle eas tu veni ad me quia pax tibi est et nihil est mali vivit Dominus si autem sic locutus fuero puero ecce sagittae ultra te sunt vade quia dimisit te Dominus
1SAM|20|23|de verbo autem quod locuti fuimus ego et tu sit Dominus inter me et te usque in sempiternum
1SAM|20|24|absconditus est ergo David in agro et venerunt kalendae et sedit rex ad comedendum panem
1SAM|20|25|cumque sedisset rex super cathedram suam secundum consuetudinem quae erat iuxta parietem surrexit Ionathan et sedit Abner ex latere Saul vacuusque apparuit locus David
1SAM|20|26|et non est locutus Saul quicquam in die illa cogitabat enim quod forte evenisset ei ut non esset mundus nec purificatus
1SAM|20|27|cumque inluxisset dies secunda post kalendas rursum vacuus apparuit locus David dixitque Saul ad Ionathan filium suum cur non venit filius Isai nec heri nec hodie ad vescendum
1SAM|20|28|et respondit Ionathan Sauli rogavit me obnixe ut iret in Bethleem
1SAM|20|29|et ait dimitte me quoniam sacrificium sollemne est in civitate unus de fratribus meis accersivit me nunc ergo si inveni gratiam in oculis tuis vadam cito et videbo fratres meos ob hanc causam non venit ad mensam regis
1SAM|20|30|iratus autem Saul adversus Ionathan dixit ei fili mulieris virum ultro rapientis numquid ignoro quia diligis filium Isai in confusionem tuam et in confusionem ignominiosae matris tuae
1SAM|20|31|omnibus enim diebus quibus filius Isai vixerit super terram non stabilieris tu neque regnum tuum itaque iam nunc mitte et adduc eum ad me quia filius mortis est
1SAM|20|32|respondens autem Ionathan Sauli patri suo ait quare moritur quid fecit
1SAM|20|33|et arripuit Saul lanceam ut percuteret eum et intellexit Ionathan quod definitum esset patri suo ut interficeret David
1SAM|20|34|surrexit ergo Ionathan a mensa in ira furoris et non comedit in die kalendarum secunda panem contristatus est enim super David eo quod confudisset eum pater suus
1SAM|20|35|cumque inluxisset mane venit Ionathan in agrum iuxta placitum David et puer parvulus cum eo
1SAM|20|36|et ait ad puerum suum vade et adfer mihi sagittas quas ego iacio cumque puer cucurrisset iecit aliam sagittam trans puerum
1SAM|20|37|venit itaque puer ad locum iaculi quod miserat Ionathan et clamavit Ionathan post tergum pueri et ait ecce ibi est sagitta porro ultra te
1SAM|20|38|clamavitque Ionathan post tergum pueri festina velociter ne steteris collegit autem puer Ionathae sagittas et adtulit ad dominum suum
1SAM|20|39|et quid ageretur penitus ignorabat tantummodo enim Ionathan et David rem noverant
1SAM|20|40|dedit igitur Ionathan arma sua puero et dixit ei vade defer in civitatem
1SAM|20|41|cumque abisset puer surrexit David de loco qui vergebat ad austrum et cadens pronus in terram adoravit tertio et osculantes alterutrum fleverunt pariter David autem amplius
1SAM|20|42|dixit ergo Ionathan ad David vade in pace quaecumque iuravimus ambo in nomine Domini dicentes Dominus sit inter me et te et inter semen meum et semen tuum usque in sempiternum
1SAM|20|43|et surrexit et abiit sed et Ionathan ingressus est civitatem
1SAM|21|1|venit autem David in Nobe ad Ahimelech sacerdotem et obstipuit Ahimelech eo quod venisset David et dixit ei quare tu solus et nullus est tecum
1SAM|21|2|et ait David ad Ahimelech sacerdotem rex praecepit mihi sermonem et dixit nemo sciat rem propter quam a me missus es et cuiusmodi tibi praecepta dederim nam et pueris condixi in illum et illum locum
1SAM|21|3|nunc igitur si quid habes ad manum vel quinque panes da mihi aut quicquid inveneris
1SAM|21|4|et respondens sacerdos David ait ei non habeo panes laicos ad manum sed tantum panem sanctum si mundi sunt pueri maxime a mulieribus
1SAM|21|5|et respondit David sacerdoti et dixit ei equidem si de mulieribus agitur continuimus nos ab heri et nudius tertius quando egrediebamur et fuerunt vasa puerorum sancta porro via haec polluta est sed et ipsa hodie sanctificabitur in vasis
1SAM|21|6|dedit ergo ei sacerdos sanctificatum panem neque enim erat ibi panis nisi tantum panes propositionis qui sublati fuerant a facie Domini ut ponerentur panes calidi
1SAM|21|7|erat autem ibi vir de servis Saul in die illa intus in tabernaculo Domini et nomen eius Doec Idumeus potentissimus pastorum Saul
1SAM|21|8|dixit autem David ad Ahimelech si habes hic ad manum hastam aut gladium quia gladium meum et arma mea non tuli mecum sermo enim regis urguebat
1SAM|21|9|et dixit sacerdos gladius Goliath Philisthei quem percussisti in valle Terebinthi est involutus pallio post ephod si istum vis tollere tolle neque enim est alius hic absque eo et ait David non est huic alter similis da mihi eum
1SAM|21|10|surrexit itaque David et fugit in die illa a facie Saul et venit ad Achis regem Geth
1SAM|21|11|dixeruntque ei servi Achis numquid non iste est David rex terrae nonne huic cantabant per choros dicentes percussit Saul mille et David decem milia
1SAM|21|12|posuit autem David sermones istos in corde suo et extimuit valde a facie Achis regis Geth
1SAM|21|13|et inmutavit os suum coram eis et conlabebatur inter manus eorum et inpingebat in ostia portae defluebantque salivae eius in barbam
1SAM|21|14|et ait Achis ad servos suos vidistis hominem insanum quare adduxistis eum ad me
1SAM|21|15|an desunt nobis furiosi quod introduxistis istum ut fureret me praesente hicine ingredietur domum meam
1SAM|22|1|abiit ergo inde David et fugit in speluncam Odollam quod cum audissent fratres eius et omnis domus patris eius descenderunt ad eum illuc
1SAM|22|2|et convenerunt ad eum omnes qui erant in angustia constituti et oppressi aere alieno et amaro animo et factus est eorum princeps fueruntque cum eo quasi quadringenti viri
1SAM|22|3|et profectus est David inde in Maspha quae est Moab et dixit ad regem Moab maneat oro pater meus et mater mea vobiscum donec sciam quid faciat mihi Deus
1SAM|22|4|et reliquit eos ante faciem regis Moab manseruntque apud eum cunctis diebus quibus David fuit in praesidio
1SAM|22|5|dixitque Gad propheta ad David noli manere in praesidio proficiscere et vade in terram Iuda et profectus David venit in saltum Hareth
1SAM|22|6|et audivit Saul quod apparuisset David et viri qui erant cum eo Saul autem cum maneret in Gabaa et esset in nemore quod est in Rama hastam manu tenens cunctique socii eius circumstarent eum
1SAM|22|7|ait ad servos suos qui adsistebant ei audite filii Iemini numquid omnibus vobis dabit filius Isai agros et vineas et universos vos faciet tribunos et centuriones
1SAM|22|8|quoniam coniurastis omnes adversum me et non est qui mihi renuntiet maxime cum et filius meus foedus iunxerit cum filio Isai non est qui vicem meam doleat ex vobis nec qui adnuntiet mihi eo quod suscitaverit filius meus servum meum adversum me insidiantem mihi usque hodie
1SAM|22|9|respondens autem Doec Idumeus qui adsistebat et erat primus inter servos Saul vidi inquit filium Isai in Nobe apud Ahimelech filium Achitob
1SAM|22|10|qui consuluit pro eo Dominum et cibaria dedit ei sed et gladium Goliath Philisthei dedit illi
1SAM|22|11|misit ergo rex ad accersiendum Ahimelech filium Achitob sacerdotem et omnem domum patris eius sacerdotum qui erant in Nobe qui venerunt universi ad regem
1SAM|22|12|et ait Saul audi fili Achitob qui respondit praesto sum domine
1SAM|22|13|dixitque ad eum Saul quare coniurastis adversum me tu et filius Isai et dedisti ei panes et gladium et consuluisti pro eo Deum ut consurgeret adversum me insidiator usque hodie permanens
1SAM|22|14|respondensque Ahimelech regi ait et quis in omnibus servis tuis sicut David fidelis et gener regis et pergens ad imperium tuum et gloriosus in domo tua
1SAM|22|15|num hodie coepi consulere pro eo Deum absit hoc a me ne suspicetur rex adversus servum suum rem huiuscemodi in universa domo patris mei non enim scivit servus tuus quicquam super hoc negotio vel modicum vel grande
1SAM|22|16|dixitque rex morte morieris Ahimelech tu et omnis domus patris tui
1SAM|22|17|et ait rex emissariis qui circumstabant eum convertimini et interficite sacerdotes Domini nam manus eorum cum David est scientes quod fugisset non indicaverunt mihi noluerunt autem servi regis extendere manum suam in sacerdotes Domini
1SAM|22|18|et ait rex Doec convertere tu et inrue in sacerdotes conversusque Doec Idumeus inruit in sacerdotes et trucidavit in die illa octoginta quinque viros vestitos ephod lineo
1SAM|22|19|Nobe autem civitatem sacerdotum percussit in ore gladii viros et mulieres parvulos et lactantes bovem et asinum et ovem in ore gladii
1SAM|22|20|evadens autem unus filius Ahimelech filii Achitob cuius nomen erat Abiathar fugit ad David
1SAM|22|21|et adnuntiavit ei quod occidisset Saul sacerdotes Domini
1SAM|22|22|et ait David ad Abiathar sciebam in die illa quod cum ibi esset Doec Idumeus procul dubio adnuntiaret Saul ego sum reus omnium animarum patris tui
1SAM|22|23|mane mecum ne timeas si quis quaesierit animam meam quaeret et animam tuam mecumque servaberis
1SAM|23|1|et nuntiaverunt David dicentes ecce Philisthim obpugnant Ceila et diripiunt areas
1SAM|23|2|consuluit igitur David Dominum dicens num vadam et percutiam Philistheos istos et ait Dominus ad David vade et percuties Philistheos et salvabis Ceila
1SAM|23|3|et dixerunt viri qui erant cum David ad eum ecce nos hic in Iudaea consistentes timemus quanto magis si ierimus in Ceila adversum agmina Philisthinorum
1SAM|23|4|rursum ergo David consuluit Dominum qui respondens ei ait surge et vade in Ceila ego enim tradam Philistheos in manu tua
1SAM|23|5|abiit David et viri eius in Ceila et pugnavit adversum Philistheos et abegit iumenta eorum et percussit eos plaga magna et salvavit David habitatores Ceilae
1SAM|23|6|porro eo tempore quo fugiebat Abiathar filius Ahimelech ad David in Ceila ephod secum habens descenderat
1SAM|23|7|nuntiatum est autem Saul quod venisset David in Ceila et ait Saul tradidit eum Deus in manus meas conclususque est introgressus urbem in qua portae et serae
1SAM|23|8|et praecepit Saul omni populo ut ad pugnam descenderet in Ceila et obsideret David et viros eius
1SAM|23|9|quod cum rescisset David quia praepararet ei Saul clam malum dixit ad Abiathar sacerdotem adplica ephod
1SAM|23|10|et ait David Domine Deus Israhel audivit famam servus tuus quod disponat Saul venire ad Ceila ut evertat urbem propter me
1SAM|23|11|si tradent me viri Ceila in manus eius et si descendet Saul sicut audivit servus tuus Domine Deus Israhel indica servo tuo et ait Dominus descendet
1SAM|23|12|dixitque David si tradent viri Ceilae me et viros qui sunt mecum in manu Saul et dixit Dominus tradent
1SAM|23|13|surrexit ergo David et viri eius quasi sescenti et egressi de Ceila huc atque illuc vagabantur incerti nuntiatumque est Saul quod fugisset David de Ceila quam ob rem dissimulavit exire
1SAM|23|14|morabatur autem David in deserto in locis firmissimis mansitque in monte solitudinis Ziph quaerebat tamen eum Saul cunctis diebus et non tradidit eum Deus in manus eius
1SAM|23|15|et vidit David quod egressus esset Saul ut quaereret animam eius porro David erat in deserto Ziph in silva
1SAM|23|16|et surrexit Ionathan filius Saul et abiit ad David in silva et confortavit manus eius in Deo dixitque ei
1SAM|23|17|ne timeas neque enim inveniet te manus Saul patris mei et tu regnabis super Israhel et ego ero tibi secundus sed et Saul pater meus scit hoc
1SAM|23|18|percussit igitur uterque foedus coram Domino mansitque David in silva Ionathas autem reversus est in domum suam
1SAM|23|19|ascenderunt autem Ziphei ad Saul in Gabaa dicentes nonne David latitat apud nos in locis tutissimis silvae in colle Achilae quae est ad dexteram deserti
1SAM|23|20|nunc ergo sicut desideravit anima tua ut descenderes descende nostrum autem erit ut tradamus eum in manus regis
1SAM|23|21|dixitque Saul benedicti vos a Domino quia doluistis vicem meam
1SAM|23|22|abite oro et diligentius praeparate et curiosius agite et considerate locum ubi sit pes eius vel quis viderit eum ibi recogitat enim de me quod callide insidier ei
1SAM|23|23|considerate et videte omnia latibula eius in quibus absconditur et revertimini ad me ad rem certam ut vadam vobiscum quod si etiam in terra se abstruserit perscrutabor eum in cunctis milibus Iuda
1SAM|23|24|at illi surgentes abierunt in Ziph ante Saul David autem et viri eius erant in deserto Maon in campestribus ad dextram Iesimuth
1SAM|23|25|ivit ergo Saul et socii eius ad quaerendum et nuntiatum est David statimque descendit ad petram et versabatur in deserto Maon quod cum audisset Saul persecutus est David in deserto Maon
1SAM|23|26|et ibat Saul ad latus montis ex parte una David autem et viri eius erant in latere montis ex parte altera porro David desperabat se posse evadere a facie Saul itaque Saul et viri eius in modum coronae cingebant David et viros eius ut caperent eos
1SAM|23|27|et nuntius venit ad Saul dicens festina et veni quoniam infuderunt se Philisthim super terram
1SAM|23|28|reversus est ergo Saul desistens persequi David et perrexit in occursum Philisthinorum propter hoc vocaverunt locum illum petram Dividentem
1SAM|24|1|ascendit ergo David inde et habitavit in locis tutissimis Engaddi
1SAM|24|2|cumque reversus esset Saul postquam persecutus est Philistheos nuntiaverunt ei dicentes ecce David in deserto est Engaddi
1SAM|24|3|adsumens ergo Saul tria milia electorum virorum ex omni Israhel perrexit ad investigandum David et viros eius etiam super abruptissimas petras quae solis hibicibus perviae sunt
1SAM|24|4|et venit ad caulas quoque ovium quae se offerebant vianti eratque ibi spelunca quam ingressus est Saul ut purgaret ventrem porro David et viri eius in interiori parte speluncae latebant
1SAM|24|5|et dixerunt servi David ad eum ecce dies de qua locutus est Dominus ad te ego tradam tibi inimicum tuum ut facias ei sicut placuerit in oculis tuis surrexit ergo David et praecidit oram clamydis Saul silenter
1SAM|24|6|post haec percussit cor suum David eo quod abscidisset oram clamydis Saul
1SAM|24|7|dixitque ad viros suos propitius mihi sit Dominus ne faciam hanc rem domino meo christo Domini ut mittam manum meam in eum quoniam christus Domini est
1SAM|24|8|et confregit David viros suos sermonibus et non permisit eos ut consurgerent in Saul porro Saul exsurgens de spelunca pergebat coepto itinere
1SAM|24|9|surrexit autem et David post eum et egressus de spelunca clamavit post tergum Saul dicens domine mi rex et respexit Saul post se et inclinans se David pronus in terram adoravit
1SAM|24|10|dixitque ad Saul quare audis verba hominum loquentium David quaerit malum adversum te
1SAM|24|11|ecce hodie viderunt oculi tui quod tradiderit te Dominus in manu mea in spelunca et cogitavi ut occiderem te sed pepercit tibi oculus meus dixi enim non extendam manum meam in domino meo quia christus Domini est
1SAM|24|12|quin potius pater mi vide et cognosce oram clamydis tuae in manu mea quoniam cum praeciderem summitatem clamydis tuae nolui extendere manum meam in te animadverte et vide quoniam non est in manu mea malum neque iniquitas neque peccavi in te tu autem insidiaris animae meae ut auferas eam
1SAM|24|13|iudicet Dominus inter me et te et ulciscatur me Dominus ex te manus autem mea non sit in te
1SAM|24|14|sicut et in proverbio antiquo dicitur ab impiis egredietur impietas manus ergo mea non sit in te
1SAM|24|15|quem sequeris rex Israhel quem persequeris canem mortuum sequeris et pulicem unum
1SAM|24|16|sit Dominus iudex et iudicet inter me et te et videat et diiudicet causam meam et eruat me de manu tua
1SAM|24|17|cum autem conplesset David loquens sermones huiuscemodi ad Saul dixit Saul numquid vox haec tua est fili mi David et levavit Saul vocem suam et flevit
1SAM|24|18|dixitque ad David iustior tu es quam ego tu enim tribuisti mihi bona ego autem reddidi tibi mala
1SAM|24|19|et tu indicasti hodie quae feceris mihi bona quomodo tradiderit me Dominus in manu tua et non occideris me
1SAM|24|20|quis enim cum invenerit inimicum suum dimittet eum in via bona sed Dominus reddat tibi vicissitudinem hanc pro eo quod hodie operatus es in me
1SAM|24|21|et nunc quia scio quod certissime regnaturus sis et habiturus in manu tua regnum Israhel
1SAM|24|22|iura mihi in Domino ne deleas semen meum post me neque auferas nomen meum de domo patris mei
1SAM|24|23|et iuravit David Sauli abiit ergo Saul in domum suam et David et viri eius ascenderunt ad tutiora loca
1SAM|25|1|mortuus est autem Samuhel et congregatus est universus Israhel et planxerunt eum et sepelierunt in domo sua in Rama consurgensque David descendit in desertum Pharan
1SAM|25|2|erat autem vir quispiam in solitudine Maon et possessio eius in Carmelo et homo ille magnus nimis erantque ei oves tria milia et mille caprae et accidit ut tonderetur grex eius in Carmelo
1SAM|25|3|nomen autem viri illius erat Nabal et nomen uxoris eius Abigail eratque mulier illa prudentissima et speciosa porro vir eius durus et pessimus et malitiosus erat autem de genere Chaleb
1SAM|25|4|cum ergo audisset David in deserto quod tonderet Nabal gregem suum
1SAM|25|5|misit decem iuvenes et dixit eis ascendite in Carmelum et venietis ad Nabal et salutabitis eum ex nomine meo pacifice
1SAM|25|6|et dicetis sic fratribus meis et tibi pax et domui tuae pax et omnibus quaecumque habes sit pax
1SAM|25|7|audivi quod tonderent pastores tui qui erant nobiscum in deserto numquam eis molesti fuimus nec aliquando defuit eis quicquam de grege omni tempore quo fuerunt nobiscum in Carmelo
1SAM|25|8|interroga pueros tuos et indicabunt tibi nunc ergo inveniant pueri gratiam in oculis tuis in die enim bona venimus quodcumque invenerit manus tua da servis tuis et filio tuo David
1SAM|25|9|cumque venissent pueri David locuti sunt ad Nabal omnia verba haec ex nomine David et siluerunt
1SAM|25|10|respondens autem Nabal pueris David ait quis est David et quis est filius Isai hodie increverunt servi qui fugiunt dominos suos
1SAM|25|11|tollam ergo panes meos et aquas meas et carnes pecorum quae occidi tonsoribus meis et dabo viris quos nescio unde sint
1SAM|25|12|regressi sunt itaque pueri David per viam suam et reversi venerunt et nuntiaverunt ei omnia verba quae dixerat
1SAM|25|13|tunc David ait viris suis accingatur unusquisque gladio suo et accincti sunt singuli gladio suo accinctusque est et David ense suo et secuti sunt David quasi quadringenti viri porro ducenti remanserunt ad sarcinas
1SAM|25|14|Abigail autem uxori Nabal nuntiavit unus de pueris dicens ecce misit David nuntios de deserto ut benedicerent domino nostro et aversus est eos
1SAM|25|15|homines isti boni satis fuerunt nobis et non molesti nec quicquam aliquando periit omni tempore quo sumus conversati cum eis in deserto
1SAM|25|16|pro muro erant nobis tam in nocte quam in die omnibus diebus quibus pavimus apud eos greges
1SAM|25|17|quam ob rem considera et recogita quid facias quoniam conpleta est malitia adversum virum tuum et adversus domum tuam et ipse filius est Belial ita ut nemo ei possit loqui
1SAM|25|18|festinavit igitur Abigail et tulit ducentos panes et duos utres vini et quinque arietes coctos et quinque sata pulentae et centum ligaturas uvae passae et ducentas massas caricarum et inposuit super asinos
1SAM|25|19|dixitque pueris suis praecedite me ecce ego post tergum sequar vos viro autem suo Nabal non indicavit
1SAM|25|20|cum ergo ascendisset asinum et descenderet ad radices montis David et viri eius descendebant in occursum eius quibus et illa occurrit
1SAM|25|21|et ait David vere frustra servavi omnia quae huius erant in deserto et non periit quicquam de cunctis quae ad eum pertinebant et reddidit mihi malum pro bono
1SAM|25|22|haec faciat Deus inimicis David et haec addat si reliquero de omnibus quae ad eum pertinent usque mane mingentem ad parietem
1SAM|25|23|cum autem vidisset Abigail David festinavit et descendit de asino et procidit coram David super faciem suam et adoravit super terram
1SAM|25|24|et cecidit ad pedes eius et dixit in me sit domine mi haec iniquitas loquatur obsecro ancilla tua in auribus tuis et audi verba famulae tuae
1SAM|25|25|ne ponat oro dominus meus rex cor suum super virum istum iniquum Nabal quia secundum nomen suum stultus est et est stultitia cum eo ego autem ancilla tua non vidi pueros tuos domine mi quos misisti
1SAM|25|26|nunc ergo domine mi vivit Dominus et vivit anima tua qui prohibuit te ne venires in sanguine et salvavit manum tuam tibi et nunc fiant sicut Nabal inimici tui et qui quaerunt domino meo malum
1SAM|25|27|quapropter suscipe benedictionem hanc quam adtulit ancilla tua tibi domino meo et da pueris qui sequuntur te dominum meum
1SAM|25|28|aufer iniquitatem famulae tuae faciens enim faciet tibi Dominus domino meo domum fidelem quia proelia Domini domine mi tu proeliaris malitia ergo non inveniatur in te omnibus diebus vitae tuae
1SAM|25|29|si enim surrexerit aliquando homo persequens te et quaerens animam tuam erit anima domini mei custodita quasi in fasciculo viventium apud Dominum Deum tuum porro anima inimicorum tuorum rotabitur quasi in impetu et circulo fundae
1SAM|25|30|cum ergo fecerit tibi Dominus domino meo omnia quae locutus est bona de te et constituerit te ducem super Israhel
1SAM|25|31|non erit tibi hoc in singultum et in scrupulum cordis domino meo quod effuderis sanguinem innoxium aut ipse te ultus fueris et cum benefecerit Dominus domino meo recordaberis ancillae tuae
1SAM|25|32|et ait David ad Abigail benedictus Dominus Deus Israhel qui misit te hodie in occursum meum et benedictum eloquium tuum
1SAM|25|33|et benedicta tu quae prohibuisti me hodie ne irem ad sanguinem et ulciscerer me manu mea
1SAM|25|34|alioquin vivit Dominus Deus Israhel qui prohibuit me malum facere tibi nisi cito venisses in occursum mihi non remansisset Nabal usque ad lucem matutinam mingens ad parietem
1SAM|25|35|suscepit ergo David de manu eius omnia quae adtulerat ei dixitque ei vade pacifice in domum tuam ecce audivi vocem tuam et honoravi faciem tuam
1SAM|25|36|venit autem Abigail ad Nabal et ecce erat ei convivium in domo eius quasi convivium regis et cor Nabal iucundum erat enim ebrius nimis et non indicavit ei verbum pusillum aut grande usque in mane
1SAM|25|37|diluculo autem cum digessisset vinum Nabal indicavit ei uxor sua verba haec et emortuum est cor eius intrinsecus et factus est quasi lapis
1SAM|25|38|cumque pertransissent decem dies percussit Dominus Nabal et mortuus est
1SAM|25|39|quod cum audisset David mortuum Nabal ait benedictus Dominus qui iudicavit causam obprobrii mei de manu Nabal et servum suum custodivit a malo et malitiam Nabal reddidit Dominus in caput eius misit ergo David et locutus est ad Abigail ut sumeret eam sibi in uxorem
1SAM|25|40|et venerunt pueri David ad Abigail in Carmelum et locuti sunt ad eam dicentes David misit nos ad te ut accipiat te sibi in uxorem
1SAM|25|41|quae consurgens adoravit prona in terram et ait ecce famula tua sit in ancillam ut lavet pedes servorum domini mei
1SAM|25|42|et festinavit et surrexit Abigail et ascendit super asinum et quinque puellae ierunt cum ea pedisequae eius et secuta est nuntios David et facta est illi uxor
1SAM|25|43|sed et Ahinoem accepit David de Iezrahel et fuit utraque uxor eius
1SAM|25|44|Saul autem dedit Michol filiam suam uxorem David Falti filio Lais qui erat de Gallim
1SAM|26|1|et venerunt Ziphei ad Saul in Gabaa dicentes ecce David absconditus est in colle Achilae quae est ex adverso solitudinis
1SAM|26|2|et surrexit Saul et descendit in desertum Ziph et cum eo tria milia virorum de electis Israhel ut quaereret David in deserto Ziph
1SAM|26|3|et castrametatus est Saul in Gabaa Achilae quae erat ex adverso solitudinis in via David autem habitabat in deserto videns autem quod venisset Saul post se in desertum
1SAM|26|4|misit exploratores et didicit quod venisset certissime
1SAM|26|5|et surrexit David et venit ad locum ubi erat Saul cumque vidisset locum in quo dormiebat Saul et Abner filius Ner princeps militiae eius Saulem dormientem in tentorio et reliquum vulgus per circuitum eius
1SAM|26|6|ait David ad Ahimelech Cettheum et Abisai filium Sarviae fratrem Ioab dicens quis descendet mecum ad Saul in castra dixitque Abisai ego descendam tecum
1SAM|26|7|venerunt ergo David et Abisai ad populum nocte et invenerunt Saul iacentem et dormientem in tentorio et hastam fixam in terra ad caput eius Abner autem et populum dormientes in circuitu eius
1SAM|26|8|dixitque Abisai ad David conclusit Deus hodie inimicum tuum in manus tuas nunc ergo perfodiam eum lancea in terra semel et secundo opus non erit
1SAM|26|9|et dixit David ad Abisai ne interficias eum quis enim extendit manum suam in christum Domini et innocens erit
1SAM|26|10|et dixit David vivit Dominus quia nisi Dominus percusserit eum aut dies eius venerit ut moriatur aut in proelium descendens perierit
1SAM|26|11|propitius mihi sit Dominus ne extendam manum meam in christum Domini nunc igitur tolle hastam quae est ad caput eius et scyphum aquae et abeamus
1SAM|26|12|tulit ergo David hastam et scyphum aquae qui erat ad caput Saul et abierunt et non erat quisquam qui videret et intellegeret et vigilaret sed omnes dormiebant quia sopor Domini inruerat super eos
1SAM|26|13|cumque transisset David ex adverso et stetisset in vertice montis de longe et esset grande intervallum inter eos
1SAM|26|14|clamavit David ad populum et ad Abner filium Ner dicens nonne respondebis Abner et respondens Abner ait quis es tu qui clamas et inquietas regem
1SAM|26|15|et ait David ad Abner numquid non vir tu es et quis alius similis tui in Israhel quare ergo non custodisti dominum tuum regem ingressus est enim unus de turba ut interficeret regem dominum tuum
1SAM|26|16|non est bonum hoc quod fecisti vivit Dominus quoniam filii mortis estis vos qui non custodistis dominum vestrum christum Domini nunc ergo vide ubi sit hasta regis et ubi scyphus aquae qui erat ad caput eius
1SAM|26|17|cognovit autem Saul vocem David et dixit num vox tua est haec fili mi David et David vox mea domine mi rex
1SAM|26|18|et ait quam ob causam dominus meus persequitur servum suum quid feci aut quod est in manu mea malum
1SAM|26|19|nunc ergo audi oro domine mi rex verba servi tui si Dominus incitat te adversum me odoretur sacrificium si autem filii hominum maledicti sunt in conspectu Domini qui eiecerunt me hodie ut non habitem in hereditate Domini dicentes vade servi diis alienis
1SAM|26|20|et nunc non effundatur sanguis meus in terra coram Domino quia egressus est rex Israhel ut quaerat pulicem unum sicut persequitur perdix in montibus
1SAM|26|21|et ait Saul peccavi revertere fili mi David nequaquam enim ultra male tibi faciam eo quod pretiosa fuerit anima mea in oculis tuis hodie apparet quod stulte egerim et ignoraverim multa nimis
1SAM|26|22|et respondens David ait ecce hasta regis transeat unus de pueris et tollat eam
1SAM|26|23|Dominus autem retribuet unicuique secundum iustitiam suam et fidem tradidit enim te Dominus hodie in manu mea et nolui levare manum meam in christum Domini
1SAM|26|24|et sicuti magnificata est anima tua hodie in oculis meis sic magnificetur anima mea in oculis Domini et liberet me de omni angustia
1SAM|26|25|ait ergo Saul ad David benedictus tu fili mi David et quidem faciens facies et potens poteris abiit autem David in viam suam et Saul reversus est in locum suum
1SAM|27|1|et ait David in corde suo aliquando incidam in uno die in manu Saul nonne melius est ut fugiam et salver in terra Philisthinorum ut desperet Saul cessetque me quaerere in cunctis finibus Israhel fugiam ergo manus eius
1SAM|27|2|et surrexit David et abiit ipse et sescenti viri cum eo ad Achis filium Mahoc regem Geth
1SAM|27|3|et habitavit David cum Achis in Geth ipse et viri eius vir et domus eius David et duae uxores eius Ahinoem Iezrahelites et Abigail uxor Nabal Carmeli
1SAM|27|4|et nuntiatum est Saul quod fugisset David in Geth et non addidit ultra ut quaereret eum
1SAM|27|5|dixit autem David ad Achis si inveni gratiam in oculis tuis detur mihi locus in una urbium regionis huius ut habitem ibi cur enim manet servus tuus in civitate regis tecum
1SAM|27|6|dedit itaque ei Achis in die illa Siceleg propter quam causam facta est Siceleg regum Iuda usque in diem hanc
1SAM|27|7|fuit autem numerus dierum quibus habitavit David in regione Philisthinorum quattuor mensuum
1SAM|27|8|et ascendit David et viri eius et agebant praedas de Gesuri et de Gedri et de Amalechitis hii enim pagi habitabantur in terra antiquitus euntibus Sur usque ad terram Aegypti
1SAM|27|9|et percutiebat David omnem terram nec relinquebat viventem virum et mulierem tollensque oves et boves et asinos et camelos et vestes revertebatur et veniebat ad Achis
1SAM|27|10|dicebat autem ei Achis in quem inruisti hodie respondebatque David contra meridiem Iudae et contra meridiem Hiramel et contra meridiem Ceni
1SAM|27|11|virum et mulierem non vivificabat David nec adducebat in Geth dicens ne forte loquantur adversum nos haec fecit David et hoc erat decretum illi omnibus diebus quibus habitavit in regione Philisthinorum
1SAM|27|12|credidit ergo Achis David dicens multa mala operatus est contra populum suum Israhel erit igitur mihi servus sempiternus
1SAM|28|1|factum est autem in diebus illis congregaverunt Philisthim agmina sua ut praepararentur ad bellum contra Israhel dixitque Achis ad David sciens nunc scito quoniam mecum egredieris in castris tu et viri tui
1SAM|28|2|dixitque David ad Achis nunc scies quae facturus est servus tuus et ait Achis ad David et ego custodem capitis mei ponam te cunctis diebus
1SAM|28|3|Samuhel autem mortuus est planxitque eum omnis Israhel et sepelierunt eum in Rama urbe sua et Saul abstulit magos et ariolos de terra
1SAM|28|4|congregatique sunt Philisthim et venerunt et castrametati sunt in Sunam congregavit autem et Saul universum Israhel et venit in Gelboe
1SAM|28|5|et vidit Saul castra Philisthim et timuit et expavit cor eius nimis
1SAM|28|6|consuluitque Dominum et non respondit ei neque per somnia neque per sacerdotes neque per prophetas
1SAM|28|7|dixitque Saul servis suis quaerite mihi mulierem habentem pythonem et vadam ad eam et sciscitabor per illam et dixerunt servi eius ad eum est mulier habens pythonem in Aendor
1SAM|28|8|mutavit ergo habitum suum vestitusque est aliis vestimentis abiit ipse et duo viri cum eo veneruntque ad mulierem nocte et ait divina mihi in pythone et suscita mihi quem dixero tibi
1SAM|28|9|et ait mulier ad eum ecce tu nosti quanta fecerit Saul et quomodo eraserit magos et ariolos de terra quare ergo insidiaris animae meae ut occidar
1SAM|28|10|et iuravit ei Saul in Domino dicens vivit Dominus quia non veniet tibi quicquam mali propter hanc rem
1SAM|28|11|dixitque ei mulier quem suscitabo tibi qui ait Samuhelem suscita mihi
1SAM|28|12|cum autem vidisset mulier Samuhelem exclamavit voce magna et dixit ad Saul quare inposuisti mihi tu es enim Saul
1SAM|28|13|dixitque ei rex noli timere quid vidisti et ait mulier ad Saul deos vidi ascendentes de terra
1SAM|28|14|dixitque ei qualis est forma eius quae ait vir senex ascendit et ipse amictus est pallio intellexit Saul quod Samuhel esset et inclinavit se super faciem suam in terra et adoravit
1SAM|28|15|dixit autem Samuhel ad Saul quare inquietasti me ut suscitarer et ait Saul coartor nimis siquidem Philisthim pugnant adversum me et Deus recessit a me et exaudire me noluit neque in manu prophetarum neque per somnia vocavi ergo te ut ostenderes mihi quid faciam
1SAM|28|16|et ait Samuhel quid interrogas me cum Dominus recesserit a te et transierit ad aemulum tuum
1SAM|28|17|faciet enim Dominus tibi sicut locutus est in manu mea et scindet regnum de manu tua et dabit illud proximo tuo David
1SAM|28|18|quia non oboedisti voci Domini neque fecisti iram furoris eius in Amalech idcirco quod pateris fecit tibi Dominus hodie
1SAM|28|19|et dabit Dominus etiam Israhel tecum in manu Philisthim cras autem tu et filii tui mecum eritis sed et castra Israhel tradet Dominus in manu Philisthim
1SAM|28|20|statimque Saul cecidit porrectus in terram extimuerat enim verba Samuhel et robur non erat in eo quia non comederat panem tota die illa
1SAM|28|21|ingressa est itaque mulier ad Saul et ait conturbatus enim erat valde dixitque ad eum ecce oboedivit ancilla tua voci tuae et posui animam meam in manu mea et audivi sermones tuos quos locutus es ad me
1SAM|28|22|nunc igitur audi et tu vocem ancillae tuae ut ponam coram te buccellam panis et comedens convalescas ut possis iter facere
1SAM|28|23|qui rennuit et ait non comedam coegerunt autem eum servi sui et mulier et tandem audita voce eorum surrexit de terra et sedit super lectum
1SAM|28|24|mulier autem illa habebat vitulum pascualem in domo et festinavit et occidit eum tollensque farinam miscuit eam et coxit azyma
1SAM|28|25|et posuit ante Saul et ante servos eius qui cum comedissent surrexerunt et ambulaverunt per totam noctem illam
1SAM|29|1|congregata sunt ergo Philisthim universa agmina in Afec sed et Israhel castrametatus est super fontem qui erat in Iezrahel
1SAM|29|2|et satrapae quidem Philisthim incedebant in centuriis et milibus David autem et viri eius erant in novissimo agmine cum Achis
1SAM|29|3|dixeruntque principes Philisthim quid sibi volunt Hebraei isti et ait Achis ad principes Philisthim num ignoratis David qui fuit servus Saul regis Israhel et est apud me multis diebus vel annis et non inveni in eo quicquam ex die qua transfugit ad me usque ad diem hanc
1SAM|29|4|irati sunt autem adversus eum principes Philisthim et dixerunt ei revertatur vir et sedeat in loco suo in quo constituisti eum et non descendat nobiscum in proelium ne fiat nobis adversarius cum proeliari coeperimus quomodo enim aliter placare poterit dominum suum nisi in capitibus nostris
1SAM|29|5|nonne iste est David cui cantabant in choro dicentes percussit Saul in milibus suis et David in decem milibus suis
1SAM|29|6|vocavit ergo Achis David et ait ei vivit Dominus quia rectus es tu et bonus in conspectu meo et exitus tuus et introitus tuus mecum est in castris et non inveni in te quicquam mali ex die qua venisti ad me usque ad diem hanc sed satrapis non places
1SAM|29|7|revertere ergo et vade in pace et non offendes oculos satraparum Philisthim
1SAM|29|8|dixitque David ad Achis quid enim feci et quid invenisti in me servo tuo a die qua fui in conspectu tuo usque in diem hanc ut non veniam et pugnem contra inimicos domini mei regis
1SAM|29|9|respondens autem Achis locutus est ad David scio quia bonus es tu in oculis meis sicut angelus Dei sed principes Philisthim dixerunt non ascendet nobiscum in proelium
1SAM|29|10|igitur consurge mane tu et servi domini tui qui venerunt tecum et cum de nocte surrexeritis et coeperit dilucescere pergite
1SAM|29|11|surrexit itaque de nocte David ipse et viri eius ut proficiscerentur mane et reverterentur ad terram Philisthim Philisthim autem ascenderunt in Iezrahel
1SAM|30|1|cumque venissent David et viri eius in Siceleg die tertia Amalechitae impetum fecerant ex parte australi in Siceleg et percusserant Siceleg et succenderant eam igni
1SAM|30|2|et captivas duxerant mulieres ex ea et a minimo usque ad magnum et non interfecerant quemquam sed secum duxerant et pergebant in itinere suo
1SAM|30|3|cum ergo venisset David et viri eius ad civitatem et invenissent eam succensam igni et uxores suas et filios suos et filias ductas esse captivas
1SAM|30|4|levaverunt David et populus qui erat cum eo voces suas et planxerunt donec deficerent in eis lacrimae
1SAM|30|5|siquidem et duae uxores David captivae ductae fuerant Ahinoem Iezrahelites et Abigail uxor Nabal Carmeli
1SAM|30|6|et contristatus est David valde volebat enim eum populus lapidare quia amara erat anima uniuscuiusque viri super filiis suis et filiabus confortatus est autem David in Domino Deo suo
1SAM|30|7|et ait ad Abiathar sacerdotem filium Ahimelech adplica ad me ephod et adplicuit Abiathar ephod ad David
1SAM|30|8|et consuluit David Dominum dicens persequar an non latrunculos hos et conprehendam eos dixitque ei persequere absque dubio enim conprehendes eos et excuties praedam
1SAM|30|9|abiit ergo David ipse et sescenti viri qui erant cum eo et venerunt usque ad torrentem Besor et lassi quidam substiterunt
1SAM|30|10|persecutus est autem David ipse et quadringenti viri substiterant enim ducenti qui lassi transire non poterant torrentem Besor
1SAM|30|11|et invenerunt virum aegyptium in agro et adduxerunt eum ad David dederuntque ei panem ut comederet et ut biberet aquam
1SAM|30|12|sed et fragmen massae caricarum et duas ligaturas uvae passae quae cum comedisset reversus est spiritus eius et refocilatus est non enim comederat panem neque biberat aquam tribus diebus et tribus noctibus
1SAM|30|13|dixit itaque ei David cuius es tu vel unde quo pergis qui ait ei puer aegyptius ego sum servus viri amalechitae dereliquit autem me dominus meus quia aegrotare coepi nudius tertius
1SAM|30|14|siquidem nos erupimus ad australem partem Cerethi et contra Iudam et ad meridiem Chaleb et Siceleg succendimus igni
1SAM|30|15|dixitque ei David potes me ducere ad istum cuneum qui ait iura mihi per Deum quod non occidas me et non tradas me in manu domini mei et ducam te ad cuneum istum
1SAM|30|16|qui cum duxisset eum ecce illi discumbebant super faciem universae terrae comedentes et bibentes et quasi festum celebrantes diem pro cuncta praeda et spoliis quae ceperant de terra Philisthim et de terra Iuda
1SAM|30|17|et percussit eos David a vespere usque ad vesperam alterius diei et non evasit ex eis quisquam nisi quadringenti viri adulescentes qui ascenderant camelos et fugerant
1SAM|30|18|eruit ergo David omnia quae tulerant Amalechitae et duas uxores suas eruit
1SAM|30|19|nec defuit quicquam a parvo usque ad magnum tam de filiis quam de filiabus et de spoliis et quaecumque rapuerant omnia reduxit David
1SAM|30|20|et tulit universos greges et armenta et minavit ante faciem suam dixeruntque haec est praeda David
1SAM|30|21|venit autem David ad ducentos viros qui lassi substiterant nec sequi potuerant David et residere eos iusserat in torrente Besor qui egressi sunt obviam David et populo qui erat cum eo accedens autem David ad populum salutavit eos pacifice
1SAM|30|22|respondensque omnis vir pessimus et iniquus de viris qui ierant cum David dixit quia non venerunt nobiscum non dabimus eis quicquam de praeda quam eruimus sed sufficiat unicuique uxor sua et filii quos cum acceperint recedant
1SAM|30|23|dixit autem David non sic facietis fratres mei de his quae tradidit Dominus nobis et custodivit nos et dedit latrunculos qui eruperant adversum nos in manu nostra
1SAM|30|24|nec audiet vos quisquam super sermone hoc aequa enim pars erit descendentis ad proelium et remanentis ad sarcinas et similiter divident
1SAM|30|25|et factum est hoc ex die illa et deinceps constitutum et praefinitum et quasi lex in Israhel usque ad diem hanc
1SAM|30|26|venit ergo David in Siceleg et misit dona de praeda senioribus Iuda proximis suis dicens accipite benedictionem de praeda hostium Domini
1SAM|30|27|his qui erant in Bethel et qui in Ramoth ad meridiem et qui in Iether
1SAM|30|28|et qui in Aroer et qui in Sefamoth et qui in Esthama
1SAM|30|29|et qui in Rachal et qui in urbibus Ierameli et qui in urbibus Ceni
1SAM|30|30|et qui in Arama et qui in lacu Asan et qui in Athac
1SAM|30|31|et qui in Hebron et reliquis qui erant in his locis in quibus commoratus fuerat David ipse et viri eius
1SAM|31|1|Philisthim autem pugnabant adversum Israhel et fugerunt viri Israhel ante faciem Philisthim et ceciderunt interfecti in monte Gelboe
1SAM|31|2|inrueruntque Philisthim in Saul et filios eius et percusserunt Ionathan et Abinadab et Melchisue filios Saul
1SAM|31|3|totumque pondus proelii versum est in Saul et consecuti sunt eum viri sagittarii et vulneratus est vehementer a sagittariis
1SAM|31|4|dixitque Saul ad armigerum suum evagina gladium tuum et percute me ne forte veniant incircumcisi isti et interficiant me inludentes mihi et noluit armiger eius fuerat enim nimio timore perterritus arripuit itaque Saul gladium et inruit super eum
1SAM|31|5|quod cum vidisset armiger eius videlicet quod mortuus esset Saul inruit etiam ipse super gladium suum et mortuus est cum eo
1SAM|31|6|mortuus est ergo Saul et tres filii eius et armiger illius et universi viri eius in die illa pariter
1SAM|31|7|videntes autem viri Israhel qui erant trans vallem et trans Iordanem quod fugissent viri israhelitae et quod mortuus esset Saul et filii eius reliquerunt civitates suas et fugerunt veneruntque Philisthim et habitaverunt ibi
1SAM|31|8|facta autem die altera venerunt Philisthim ut spoliarent interfectos et invenerunt Saul et tres filios eius iacentes in monte Gelboe
1SAM|31|9|et praeciderunt caput Saul et expoliaverunt eum armis et miserunt in terram Philisthinorum per circuitum ut adnuntiaretur in templo idolorum et in populis
1SAM|31|10|et posuerunt arma eius in templo Astharoth corpus vero eius suspenderunt in muro Bethsan
1SAM|31|11|quod cum audissent habitatores Iabesgalaad quaecumque fecerant Philisthim Saul
1SAM|31|12|surrexerunt omnes viri fortissimi et ambulaverunt tota nocte et tulerunt cadaver Saul et cadavera filiorum eius de muro Bethsan veneruntque Iabes et conbuserunt ea ibi
1SAM|31|13|et tulerunt ossa eorum et sepelierunt in nemore Iabes et ieiunaverunt septem diebus
