HOS|1|1|The word of the LORD that came to Hosea, the son of Beeri, in the days of Uzziah, Jotham, Ahaz, and Hezekiah, kings of Judah, and in the days of Jeroboam the son of Joash, king of Israel.
HOS|1|2|When the LORD first spoke through Hosea, the LORD said to Hosea, "Go, take to yourself a wife of whoredom and have children of whoredom, for the land commits great whoredom by forsaking the LORD."
HOS|1|3|So he went and took Gomer, the daughter of Diblaim, and she conceived and bore him a son.
HOS|1|4|And the LORD said to him, "Call his name Jezreel, for in just a little while I will punish the house of Jehu for the blood of Jezreel, and I will put an end to the kingdom of the house of Israel.
HOS|1|5|And on that day I will break the bow of Israel in the Valley of Jezreel."
HOS|1|6|She conceived again and bore a daughter. And the LORD said to him, "Call her name No Mercy, for I will no more have mercy on the house of Israel, to forgive them at all.
HOS|1|7|But I will have mercy on the house of Judah, and I will save them by the LORD their God. I will not save them by bow or by sword or by war or by horses or by horsemen."
HOS|1|8|When she had weaned No Mercy, she conceived and bore a son.
HOS|1|9|And the LORD said, "Call his name Not My People, for you are not my people, and I am not your God."
HOS|1|10|Yet the number of the children of Israel shall be like the sand of the sea, which cannot be measured or numbered. And in the place where it was said to them, "You are not my people," it shall be said to them, "Children of the living God."
HOS|1|11|And the children of Judah and the children of Israel shall be gathered together, and they shall appoint for themselves one head. And they shall go up from the land, for great shall be the day of Jezreel.
HOS|2|1|Say to your brothers, "You are my people," and to your sisters, "You have received mercy."
HOS|2|2|"Plead with your mother, plead- for she is not my wife, and I am not her husband- that she put away her whoring from her face, and her adultery from between her breasts;
HOS|2|3|lest I strip her naked and make her as in the day she was born, and make her like a wilderness, and make her like a parched land, and kill her with thirst.
HOS|2|4|Upon her children also I will have no mercy, because they are children of whoredom.
HOS|2|5|For their mother has played the whore; she who conceived them has acted shamefully. For she said, 'I will go after my lovers, who give me my bread and my water, my wool and my flax, my oil and my drink.'
HOS|2|6|Therefore I will hedge up her way with thorns, and I will build a wall against her, so that she cannot find her paths.
HOS|2|7|She shall pursue her lovers but not overtake them, and she shall seek them but shall not find them. Then she shall say, 'I will go and return to my first husband, for it was better for me then than now.'
HOS|2|8|And she did not know that it was I who gave her the grain, the wine, and the oil, and who lavished on her silver and gold, which they used for Baal.
HOS|2|9|Therefore I will take back my grain in its time, and my wine in its season, and I will take away my wool and my flax, which were to cover her nakedness.
HOS|2|10|Now I will uncover her lewdness in the sight of her lovers, and no one shall rescue her out of my hand.
HOS|2|11|And I will put an end to all her mirth, her feasts, her new moons, her Sabbaths, and all her appointed feasts.
HOS|2|12|And I will lay waste her vines and her fig trees, of which she said, 'These are my wages, which my lovers have given me.' I will make them a forest, and the beasts of the field shall devour them.
HOS|2|13|And I will punish her for the feast days of the Baals when she burned offerings to them and adorned herself with her ring and jewelry, and went after her lovers and forgot me, declares the LORD.
HOS|2|14|"Therefore, behold, I will allure her, and bring her into the wilderness, and speak tenderly to her.
HOS|2|15|And there I will give her her vineyards and make the Valley of Achor a door of hope. And there she shall answer as in the days of her youth, as at the time when she came out of the land of Egypt.
HOS|2|16|"And in that day, declares the LORD, you will call me 'My Husband,' and no longer will you call me 'My Baal.'
HOS|2|17|For I will remove the names of the Baals from her mouth, and they shall be remembered by name no more.
HOS|2|18|And I will make for them a covenant on that day with the beasts of the field, the birds of the heavens, and the creeping things of the ground. And I will abolish the bow, the sword, and war from the land, and I will make you lie down in safety.
HOS|2|19|And I will betroth you to me forever. I will betroth you to me in righteousness and in justice, in steadfast love and in mercy.
HOS|2|20|I will betroth you to me in faithfulness. And you shall know the LORD.
HOS|2|21|"And in that day I will answer, declares the LORD, I will answer the heavens, and they shall answer the earth,
HOS|2|22|and the earth shall answer the grain, the wine, and the oil, and they shall answer Jezreel,
HOS|2|23|and I will sow her for myself in the land. And I will have mercy on No Mercy, and I will say to Not My People, 'You are my people'; and he shall say, 'You are my God.'"
HOS|3|1|And the LORD said to me, "Go again, love a woman who is loved by another man and is an adulteress, even as the LORD loves the children of Israel, though they turn to other gods and love cakes of raisins."
HOS|3|2|So I bought her for fifteen shekels of silver and a homer and a lethech of barley.
HOS|3|3|And I said to her, "You must dwell as mine for many days. You shall not play the whore, or belong to another man; so will I also be to you."
HOS|3|4|For the children of Israel shall dwell many days without king or prince, without sacrifice or pillar, without ephod or household gods.
HOS|3|5|Afterward the children of Israel shall return and seek the LORD their God, and David their king, and they shall come in fear to the LORD and to his goodness in the latter days.
HOS|4|1|Hear the word of the LORD, O children of Israel, for the LORD has a controversy with the inhabitants of the land. There is no faithfulness or steadfast love, and no knowledge of God in the land;
HOS|4|2|there is swearing, lying, murder, stealing, and committing adultery; they break all bounds, and bloodshed follows bloodshed.
HOS|4|3|Therefore the land mourns, and all who dwell in it languish, and also the beasts of the field and the birds of the heavens, and even the fish of the sea are taken away.
HOS|4|4|Yet let no one contend, and let none accuse, for with you is my contention, O priest.
HOS|4|5|You shall stumble by day; the prophet also shall stumble with you by night; and I will destroy your mother.
HOS|4|6|My people are destroyed for lack of knowledge; because you have rejected knowledge, I reject you from being a priest to me. And since you have forgotten the law of your God, I also will forget your children.
HOS|4|7|The more they increased, the more they sinned against me; I will change their glory into shame.
HOS|4|8|They feed on the sin of my people; they are greedy for their iniquity.
HOS|4|9|And it shall be like people, like priest; I will punish them for their ways and repay them for their deeds.
HOS|4|10|They shall eat, but not be satisfied; they shall play the whore, but not multiply, because they have forsaken the LORD to cherish
HOS|4|11|whoredom, wine, and new wine, which take away the understanding.
HOS|4|12|My people inquire of a piece of wood, and their walking staff gives them oracles. For a spirit of whoredom has led them astray, and they have left their God to play the whore.
HOS|4|13|They sacrifice on the tops of the mountains and burn offerings on the hills, under oak, poplar, and terebinth, because their shade is good. Therefore your daughters play the whore, and your brides commit adultery.
HOS|4|14|I will not punish your daughters when they play the whore, nor your brides when they commit adultery; for the men themselves go aside with prostitutes and sacrifice with cult prostitutes, and a people without understanding shall come to ruin.
HOS|4|15|Though you play the whore, O Israel, let not Judah become guilty. Enter not into Gilgal, nor go up to Beth-aven, and swear not, "As the LORD lives."
HOS|4|16|Like a stubborn heifer, Israel is stubborn; can the LORD now feed them like a lamb in a broad pasture?
HOS|4|17|Ephraim is joined to idols; leave him alone.
HOS|4|18|When their drink is gone, they give themselves to whoring; their rulers dearly love shame.
HOS|4|19|A wind has wrapped them in its wings, and they shall be ashamed because of their sacrifices.
HOS|5|1|Hear this, O priests! Pay attention, O house of Israel! Give ear, O house of the king! For the judgment is for you; for you have been a snare at Mizpah and a net spread upon Tabor.
HOS|5|2|And the revolters have gone deep into slaughter, but I will discipline all of them.
HOS|5|3|I know Ephraim, and Israel is not hidden from me; for now, O Ephraim, you have played the whore; Israel is defiled.
HOS|5|4|Their deeds do not permit them to return to their God. For the spirit of whoredom is within them, and they know not the LORD.
HOS|5|5|The pride of Israel testifies to his face; Israel and Ephraim shall stumble in his guilt; Judah also shall stumble with them.
HOS|5|6|With their flocks and herds they shall go to seek the LORD, but they will not find him; he has withdrawn from them.
HOS|5|7|They have dealt faithlessly with the LORD; for they have borne alien children. Now the new moon shall devour them with their fields.
HOS|5|8|Blow the horn in Gibeah, the trumpet in Ramah. Sound the alarm at Beth-aven; we follow you, O Benjamin!
HOS|5|9|Ephraim shall become a desolation in the day of punishment; among the tribes of Israel I make known what is sure.
HOS|5|10|The princes of Judah have become like those who move the landmark; upon them I will pour out my wrath like water.
HOS|5|11|Ephraim is oppressed, crushed in judgment, because he was determined to go after filth.
HOS|5|12|But I am like a moth to Ephraim, and like dry rot to the house of Judah.
HOS|5|13|When Ephraim saw his sickness, and Judah his wound, then Ephraim went to Assyria, and sent to the great king. But he is not able to cure you or heal your wound.
HOS|5|14|For I will be like a lion to Ephraim, and like a young lion to the house of Judah. I, even I, will tear and go away; I will carry off, and no one shall rescue.
HOS|5|15|I will return again to my place, until they acknowledge their guilt and seek my face, and in their distress earnestly seek me.
HOS|6|1|"Come, let us return to the LORD; for he has torn us, that he may heal us; he has struck us down, and he will bind us up.
HOS|6|2|After two days he will revive us; on the third day he will raise us up, that we may live before him.
HOS|6|3|Let us know; let us press on to know the LORD; his going out is sure as the dawn; he will come to us as the showers, as the spring rains that water the earth."
HOS|6|4|What shall I do with you, O Ephraim? What shall I do with you, O Judah? Your love is like a morning cloud, like the dew that goes early away.
HOS|6|5|Therefore I have hewn them by the prophets; I have slain them by the words of my mouth, and my judgment goes forth as the light.
HOS|6|6|For I desire steadfast love and not sacrifice, the knowledge of God rather than burnt offerings.
HOS|6|7|But like Adam they transgressed the covenant; there they dealt faithlessly with me.
HOS|6|8|Gilead is a city of evildoers, tracked with blood.
HOS|6|9|As robbers lie in wait for a man, so the priests band together; they murder on the way to Shechem; they commit villainy.
HOS|6|10|In the house of Israel I have seen a horrible thing; Ephraim's whoredom is there; Israel is defiled.
HOS|6|11|For you also, O Judah, a harvest is appointed, when I restore the fortunes of my people.
HOS|7|1|When I would heal Israel, the iniquity of Ephraim is revealed, and the evil deeds of Samaria; for they deal falsely; the thief breaks in, and the bandits raid outside.
HOS|7|2|But they do not consider that I remember all their evil. Now their deeds surround them; they are before my face.
HOS|7|3|By their evil they make the king glad, and the princes by their treachery.
HOS|7|4|They are all adulterers; they are like a heated oven whose baker ceases to stir the fire, from the kneading of the dough until it is leavened.
HOS|7|5|On the day of our king, the princes became sick with the heat of wine; he stretched out his hand with mockers.
HOS|7|6|For with hearts like an oven they approach their intrigue; all night their anger smolders; in the morning it blazes like a flaming fire.
HOS|7|7|All of them are hot as an oven, and they devour their rulers. All their kings have fallen, and none of them calls upon me.
HOS|7|8|Ephraim mixes himself with the peoples; Ephraim is a cake not turned.
HOS|7|9|Strangers devour his strength, and he knows it not; gray hairs are sprinkled upon him, and he knows it not.
HOS|7|10|The pride of Israel testifies to his face; yet they do not return to the LORD their God, nor seek him, for all this.
HOS|7|11|Ephraim is like a dove, silly and without sense, calling to Egypt, going to Assyria.
HOS|7|12|As they go, I will spread over them my net; I will bring them down like birds of the heavens; I will discipline them according to the report made to their congregation.
HOS|7|13|Woe to them, for they have strayed from me! Destruction to them, for they have rebelled against me! I would redeem them, but they speak lies against me.
HOS|7|14|They do not cry to me from the heart, but they wail upon their beds; for grain and wine they gash themselves; they rebel against me.
HOS|7|15|Although I trained and strengthened their arms, yet they devise evil against me.
HOS|7|16|They return, but not upwards; they are like a treacherous bow; their princes shall fall by the sword because of the insolence of their tongue. This shall be their derision in the land of Egypt.
HOS|8|1|Set the trumpet to your lips!One like a vulture is over the house of the LORD, because they have transgressed my covenant and rebelled against my law.
HOS|8|2|To me they cry, My God, we- Israel- know you.
HOS|8|3|Israel has spurned the good; the enemy shall pursue him.
HOS|8|4|They made kings, but not through me. They set up princes, but I knew it not. With their silver and gold they made idols for their own destruction.
HOS|8|5|I have spurned your calf, O Samaria. My anger burns against them. How long will they be incapable of innocence?
HOS|8|6|For it is from Israel; a craftsman made it; it is not God. The calf of Samaria shall be broken to pieces.
HOS|8|7|For they sow the wind, and they shall reap the whirlwind. The standing grain has no heads; it shall yield no flour; if it were to yield, strangers would devour it.
HOS|8|8|Israel is swallowed up; already they are among the nations as a useless vessel.
HOS|8|9|For they have gone up to Assyria, a wild donkey wandering alone; Ephraim has hired lovers.
HOS|8|10|Though they hire allies among the nations, I will soon gather them up. And the king and princes shall soon writhe because of the tribute.
HOS|8|11|Because Ephraim has multiplied altars for sinning, they have become to him altars for sinning.
HOS|8|12|Were I to write for him my laws by the ten thousands, they would be regarded as a strange thing.
HOS|8|13|As for my sacrificial offerings, they sacrifice meat and eat it, but the LORD does not accept them. Now he will remember their iniquity and punish their sins; they shall return to Egypt.
HOS|8|14|For Israel has forgotten his Maker and built palaces, and Judah has multiplied fortified cities; so I will send a fire upon his cities, and it shall devour her strongholds.
HOS|9|1|Rejoice not, O Israel!Exult not like the peoples; for you have played the whore, forsaking your God. You have loved a prostitute's wages on all threshing floors.
HOS|9|2|Threshing floor and wine vat shall not feed them, and the new wine shall fail them.
HOS|9|3|They shall not remain in the land of the LORD, but Ephraim shall return to Egypt, and they shall eat unclean food in Assyria.
HOS|9|4|They shall not pour drink offerings of wine to the LORD, and their sacrifices shall not please him. It shall be like mourners' bread to them; all who eat of it shall be defiled; for their bread shall be for their hunger only; it shall not come to the house of the LORD.
HOS|9|5|What will you do on the day of the appointed festival, and on the day of the feast of the LORD?
HOS|9|6|For behold, they are going away from destruction; but Egypt shall gather them; Memphis shall bury them. Nettles shall possess their precious things of silver; thorns shall be in their tents.
HOS|9|7|The days of punishment have come; the days of recompense have come; Israel shall know it. The prophet is a fool; the man of the spirit is mad, because of your great iniquity and great hatred.
HOS|9|8|The prophet is the watchman of Ephraim with my God; yet a fowler's snare is on all his ways, and hatred in the house of his God.
HOS|9|9|They have deeply corrupted themselves as in the days of Gibeah: he will remember their iniquity; he will punish their sins.
HOS|9|10|Like grapes in the wilderness, I found Israel. Like the first fruit on the fig tree in its first season, I saw your fathers. But they came to Baal-peor and consecrated themselves to the thing of shame, and became detestable like the thing they loved.
HOS|9|11|Ephraim's glory shall fly away like a bird- no birth, no pregnancy, no conception!
HOS|9|12|Even if they bring up children, I will bereave them till none is left. Woe to them when I depart from them!
HOS|9|13|Ephraim, as I have seen, was like a young palm planted in a meadow; but Ephraim must lead his children out to slaughter.
HOS|9|14|Give them, O LORD- what will you give? Give them a miscarrying womb and dry breasts.
HOS|9|15|Every evil of theirs is in Gilgal; there I began to hate them. Because of the wickedness of their deeds I will drive them out of my house. I will love them no more; all their princes are rebels.
HOS|9|16|Ephraim is stricken; their root is dried up; they shall bear no fruit. Even though they give birth, I will put their beloved children to death.
HOS|9|17|My God will reject them because they have not listened to him; they shall be wanderers among the nations.
HOS|10|1|Israel is a luxuriant vine that yields its fruit. The more his fruit increased, the more altars he built; as his country improved, he improved his pillars.
HOS|10|2|Their heart is false; now they must bear their guilt. The LORD will break down their altars and destroy their pillars.
HOS|10|3|For now they will say: "We have no king, for we do not fear the LORD; and a king- what could he do for us?"
HOS|10|4|They utter mere words; with empty oaths they make covenants; so judgment springs up like poisonous weeds in the furrows of the field.
HOS|10|5|The inhabitants of Samaria tremble for the calf of Beth-aven. Its people mourn for it, and so do its idolatrous priests- those who rejoiced over it and over its glory- for it has departed from them.
HOS|10|6|The thing itself shall be carried to Assyria as tribute to the great king. Ephraim shall be put to shame, and Israel shall be ashamed of his idol.
HOS|10|7|Samaria's king shall perish like a twig on the face of the waters.
HOS|10|8|The high places of Aven, the sin of Israel, shall be destroyed. Thorn and thistle shall grow up on their altars, and they shall say to the mountains, Cover us, and to the hills, Fall on us.
HOS|10|9|From the days of Gibeah, you have sinned, O Israel; there they have continued. Shall not the war against the unjust overtake them in Gibeah?
HOS|10|10|When I please, I will discipline them, and nations shall be gathered against them when they are bound up for their double iniquity.
HOS|10|11|Ephraim was a trained calf that loved to thresh, and I spared her fair neck; but I will put Ephraim to the yoke; Judah must plow; Jacob must harrow for himself.
HOS|10|12|Sow for yourselves righteousness; reap steadfast love; break up your fallow ground, for it is the time to seek the LORD, that he may come and rain righteousness upon you.
HOS|10|13|You have plowed iniquity; you have reaped injustice; you have eaten the fruit of lies. Because you have trusted in your own way and in the multitude of your warriors,
HOS|10|14|therefore the tumult of war shall arise among your people, and all your fortresses shall be destroyed, as Shalman destroyed Beth-arbel on the day of battle; mothers were dashed in pieces with their children.
HOS|10|15|Thus it shall be done to you, O Bethel, because of your great evil. At dawn the king of Israel shall be utterly cut off.
HOS|11|1|When Israel was a child, I loved him, and out of Egypt I called my son.
HOS|11|2|The more they were called, the more they went away; they kept sacrificing to the Baals and burning offerings to idols.
HOS|11|3|Yet it was I who taught Ephraim to walk; I took them up by their arms, but they did not know that I healed them.
HOS|11|4|I led them with cords of kindness, with the bands of love, and I became to them as one who eases the yoke on their jaws, and I bent down to them and fed them.
HOS|11|5|They shall not return to the land of Egypt, but Assyria shall be their king, because they have refused to return to me.
HOS|11|6|The sword shall rage against their cities, consume the bars of their gates, and devour them because of their own counsels.
HOS|11|7|My people are bent on turning away from me, and though they call out to the Most High, he shall not raise them up at all.
HOS|11|8|How can I give you up, O Ephraim? How can I hand you over, O Israel? How can I make you like Admah? How can I treat you like Zeboiim? My heart recoils within me; my compassion grows warm and tender.
HOS|11|9|I will not execute my burning anger; I will not again destroy Ephraim; for I am God and not a man, the Holy One in your midst, and I will not come in wrath.
HOS|11|10|They shall go after the LORD; he will roar like a lion; when he roars, his children shall come trembling from the west;
HOS|11|11|they shall come trembling like birds from Egypt, and like doves from the land of Assyria, and I will return them to their homes, declares the LORD.
HOS|11|12|Ephraim has surrounded me with lies, and the house of Israel with deceit, but Judah still walks with God and is faithful to the Holy One.
HOS|12|1|Ephraim feeds on the wind and pursues the east wind all day long; they multiply falsehood and violence; they make a covenant with Assyria, and oil is carried to Egypt.
HOS|12|2|The LORD has an indictment against Judah and will punish Jacob according to his ways; he will repay him according to his deeds.
HOS|12|3|In the womb he took his brother by the heel, and in his manhood he strove with God.
HOS|12|4|He strove with the angel and prevailed; he wept and sought his favor. He met God at Bethel, and there God spoke with us-
HOS|12|5|the LORD, the God of hosts, the LORD is his memorial name:
HOS|12|6|"So you, by the help of your God, return, hold fast to love and justice, and wait continually for your God."
HOS|12|7|A merchant, in whose hands are false balances, he loves to oppress.
HOS|12|8|Ephraim has said, "Ah, but I am rich; I have found wealth for myself; in all my labors they cannot find in me iniquity or sin."
HOS|12|9|I am the LORD your God from the land of Egypt; I will again make you dwell in tents, as in the days of the appointed feast.
HOS|12|10|I spoke to the prophets; it was I who multiplied visions, and through the prophets gave parables.
HOS|12|11|If there is iniquity in Gilead, they shall surely come to nothing: in Gilgal they sacrifice bulls; their altars also are like stone heaps on the furrows of the field.
HOS|12|12|Jacob fled to the land of Aram; there Israel served for a wife, and for a wife he guarded sheep.
HOS|12|13|By a prophet the LORD brought Israel up from Egypt, and by a prophet he was guarded.
HOS|12|14|Ephraim has given bitter provocation; so his Lord will leave his bloodguilt on him and will repay him for his disgraceful deeds.
HOS|13|1|When Ephraim spoke, there was trembling; he was exalted in Israel, but he incurred guilt through Baal and died.
HOS|13|2|And now they sin more and more, and make for themselves metal images, idols skillfully made of their silver, all of them the work of craftsmen. It is said of them, "Those who offer human sacrifice kiss calves!"
HOS|13|3|Therefore they shall be like the morning mist or like the dew that goes early away, like the chaff that swirls from the threshing floor or like smoke from a window.
HOS|13|4|But I am the LORD your God from the land of Egypt; you know no God but me, and besides me there is no savior.
HOS|13|5|It was I who knew you in the wilderness, in the land of drought;
HOS|13|6|but when they had grazed, they became full, they were filled, and their heart was lifted up; therefore they forgot me.
HOS|13|7|So I am to them like a lion; like a leopard I will lurk beside the way.
HOS|13|8|I will fall upon them like a bear robbed of her cubs; I will tear open their breast, and there I will devour them like a lion, as a wild beast would rip them open.
HOS|13|9|He destroys you, O Israel, for you are against me, against your helper.
HOS|13|10|Where now is your king, to save you in all your cities? Where are all your rulers- those of whom you said, "Give me a king and princes"?
HOS|13|11|I gave you a king in my anger, and I took him away in my wrath.
HOS|13|12|The iniquity of Ephraim is bound up; his sin is kept in store.
HOS|13|13|The pangs of childbirth come for him, but he is an unwise son, for at the right time he does not present himself at the opening of the womb.
HOS|13|14|Shall I ransom them from the power of Sheol? Shall I redeem them from Death? O Death, where are your plagues? O Sheol, where is your sting? Compassion is hidden from my eyes.
HOS|13|15|Though he may flourish among his brothers, the east wind, the wind of the LORD, shall come, rising from the wilderness, and his fountain shall dry up; his spring shall be parched; it shall strip his treasury of every precious thing.
HOS|13|16|Samaria shall bear her guilt, because she has rebelled against her God; they shall fall by the sword; their little ones shall be dashed in pieces, and their pregnant women ripped open.
HOS|14|1|Return, O Israel, to the LORD your God, for you have stumbled because of your iniquity.
HOS|14|2|Take with you words and return to the LORD; say to him, "Take away all iniquity; accept what is good, and we will pay with bulls the vows of our lips.
HOS|14|3|Assyria shall not save us; we will not ride on horses; and we will say no more, 'Our God,' to the work of our hands. In you the orphan finds mercy."
HOS|14|4|I will heal their apostasy; I will love them freely, for my anger has turned from them.
HOS|14|5|I will be like the dew to Israel; he shall blossom like the lily; he shall take root like the trees of Lebanon;
HOS|14|6|his shoots shall spread out; his beauty shall be like the olive, and his fragrance like Lebanon.
HOS|14|7|They shall return and dwell beneath my shadow; they shall flourish like the grain; they shall blossom like the vine; their fame shall be like the wine of Lebanon.
HOS|14|8|O Ephraim, what have I to do with idols? It is I who answer and look after you. I am like an evergreen cypress; from me comes your fruit.
HOS|14|9|Whoever is wise, let him understand these things; whoever is discerning, let him know them; for the ways of the LORD are right, and the upright walk in them, but transgressors stumble in them.
