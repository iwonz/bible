ROM|1|1|Paul, a servant of Jesus Christ, called to be an apostle, separated unto the gospel of God,
ROM|1|2|(Which he had promised afore by his prophets in the holy scriptures,)
ROM|1|3|Concerning his Son Jesus Christ our Lord, which was made of the seed of David according to the flesh;
ROM|1|4|And declared to be the Son of God with power, according to the spirit of holiness, by the resurrection from the dead:
ROM|1|5|By whom we have received grace and apostleship, for obedience to the faith among all nations, for his name:
ROM|1|6|Among whom are ye also the called of Jesus Christ:
ROM|1|7|To all that be in Rome, beloved of God, called to be saints: Grace to you and peace from God our Father, and the Lord Jesus Christ.
ROM|1|8|First, I thank my God through Jesus Christ for you all, that your faith is spoken of throughout the whole world.
ROM|1|9|For God is my witness, whom I serve with my spirit in the gospel of his Son, that without ceasing I make mention of you always in my prayers;
ROM|1|10|Making request, if by any means now at length I might have a prosperous journey by the will of God to come unto you.
ROM|1|11|For I long to see you, that I may impart unto you some spiritual gift, to the end ye may be established;
ROM|1|12|That is, that I may be comforted together with you by the mutual faith both of you and me.
ROM|1|13|Now I would not have you ignorant, brethren, that oftentimes I purposed to come unto you, (but was let hitherto,) that I might have some fruit among you also, even as among other Gentiles.
ROM|1|14|I am debtor both to the Greeks, and to the Barbarians; both to the wise, and to the unwise.
ROM|1|15|So, as much as in me is, I am ready to preach the gospel to you that are at Rome also.
ROM|1|16|For I am not ashamed of the gospel of Christ: for it is the power of God unto salvation to every one that believeth; to the Jew first, and also to the Greek.
ROM|1|17|For therein is the righteousness of God revealed from faith to faith: as it is written, The just shall live by faith.
ROM|1|18|For the wrath of God is revealed from heaven against all ungodliness and unrighteousness of men, who hold the truth in unrighteousness;
ROM|1|19|Because that which may be known of God is manifest in them; for God hath shewed it unto them.
ROM|1|20|For the invisible things of him from the creation of the world are clearly seen, being understood by the things that are made, even his eternal power and Godhead; so that they are without excuse:
ROM|1|21|Because that, when they knew God, they glorified him not as God, neither were thankful; but became vain in their imaginations, and their foolish heart was darkened.
ROM|1|22|Professing themselves to be wise, they became fools,
ROM|1|23|And changed the glory of the uncorruptible God into an image made like to corruptible man, and to birds, and fourfooted beasts, and creeping things.
ROM|1|24|Wherefore God also gave them up to uncleanness through the lusts of their own hearts, to dishonour their own bodies between themselves:
ROM|1|25|Who changed the truth of God into a lie, and worshipped and served the creature more than the Creator, who is blessed for ever. Amen.
ROM|1|26|For this cause God gave them up unto vile affections: for even their women did change the natural use into that which is against nature:
ROM|1|27|And likewise also the men, leaving the natural use of the woman, burned in their lust one toward another; men with men working that which is unseemly, and receiving in themselves that recompence of their error which was meet.
ROM|1|28|And even as they did not like to retain God in their knowledge, God gave them over to a reprobate mind, to do those things which are not convenient;
ROM|1|29|Being filled with all unrighteousness, fornication, wickedness, covetousness, maliciousness; full of envy, murder, debate, deceit, malignity; whisperers,
ROM|1|30|Backbiters, haters of God, despiteful, proud, boasters, inventors of evil things, disobedient to parents,
ROM|1|31|Without understanding, covenantbreakers, without natural affection, implacable, unmerciful:
ROM|1|32|Who knowing the judgment of God, that they which commit such things are worthy of death, not only do the same, but have pleasure in them that do them.
ROM|2|1|Therefore thou art inexcusable, O man, whosoever thou art that judgest: for wherein thou judgest another, thou condemnest thyself; for thou that judgest doest the same things.
ROM|2|2|But we are sure that the judgment of God is according to truth against them which commit such things.
ROM|2|3|And thinkest thou this, O man, that judgest them which do such things, and doest the same, that thou shalt escape the judgment of God?
ROM|2|4|Or despisest thou the riches of his goodness and forbearance and longsuffering; not knowing that the goodness of God leadeth thee to repentance?
ROM|2|5|But after thy hardness and impenitent heart treasurest up unto thyself wrath against the day of wrath and revelation of the righteous judgment of God;
ROM|2|6|Who will render to every man according to his deeds:
ROM|2|7|To them who by patient continuance in well doing seek for glory and honour and immortality, eternal life:
ROM|2|8|But unto them that are contentious, and do not obey the truth, but obey unrighteousness, indignation and wrath,
ROM|2|9|Tribulation and anguish, upon every soul of man that doeth evil, of the Jew first, and also of the Gentile;
ROM|2|10|But glory, honour, and peace, to every man that worketh good, to the Jew first, and also to the Gentile:
ROM|2|11|For there is no respect of persons with God.
ROM|2|12|For as many as have sinned without law shall also perish without law: and as many as have sinned in the law shall be judged by the law;
ROM|2|13|(For not the hearers of the law are just before God, but the doers of the law shall be justified.
ROM|2|14|For when the Gentiles, which have not the law, do by nature the things contained in the law, these, having not the law, are a law unto themselves:
ROM|2|15|Which shew the work of the law written in their hearts, their conscience also bearing witness, and their thoughts the mean while accusing or else excusing one another;)
ROM|2|16|In the day when God shall judge the secrets of men by Jesus Christ according to my gospel.
ROM|2|17|Behold, thou art called a Jew, and restest in the law, and makest thy boast of God,
ROM|2|18|And knowest his will, and approvest the things that are more excellent, being instructed out of the law;
ROM|2|19|And art confident that thou thyself art a guide of the blind, a light of them which are in darkness,
ROM|2|20|An instructor of the foolish, a teacher of babes, which hast the form of knowledge and of the truth in the law.
ROM|2|21|Thou therefore which teachest another, teachest thou not thyself? thou that preachest a man should not steal, dost thou steal?
ROM|2|22|Thou that sayest a man should not commit adultery, dost thou commit adultery? thou that abhorrest idols, dost thou commit sacrilege?
ROM|2|23|Thou that makest thy boast of the law, through breaking the law dishonourest thou God?
ROM|2|24|For the name of God is blasphemed among the Gentiles through you, as it is written.
ROM|2|25|For circumcision verily profiteth, if thou keep the law: but if thou be a breaker of the law, thy circumcision is made uncircumcision.
ROM|2|26|Therefore if the uncircumcision keep the righteousness of the law, shall not his uncircumcision be counted for circumcision?
ROM|2|27|And shall not uncircumcision which is by nature, if it fulfil the law, judge thee, who by the letter and circumcision dost transgress the law?
ROM|2|28|For he is not a Jew, which is one outwardly; neither is that circumcision, which is outward in the flesh:
ROM|2|29|But he is a Jew, which is one inwardly; and circumcision is that of the heart, in the spirit, and not in the letter; whose praise is not of men, but of God.
ROM|3|1|What advantage then hath the Jew? or what profit is there of circumcision?
ROM|3|2|Much every way: chiefly, because that unto them were committed the oracles of God.
ROM|3|3|For what if some did not believe? shall their unbelief make the faith of God without effect?
ROM|3|4|God forbid: yea, let God be true, but every man a liar; as it is written, That thou mightest be justified in thy sayings, and mightest overcome when thou art judged.
ROM|3|5|But if our unrighteousness commend the righteousness of God, what shall we say? Is God unrighteous who taketh vengeance? (I speak as a man)
ROM|3|6|God forbid: for then how shall God judge the world?
ROM|3|7|For if the truth of God hath more abounded through my lie unto his glory; why yet am I also judged as a sinner?
ROM|3|8|And not rather, (as we be slanderously reported, and as some affirm that we say,) Let us do evil, that good may come? whose damnation is just.
ROM|3|9|What then? are we better than they? No, in no wise: for we have before proved both Jews and Gentiles, that they are all under sin;
ROM|3|10|As it is written, There is none righteous, no, not one:
ROM|3|11|There is none that understandeth, there is none that seeketh after God.
ROM|3|12|They are all gone out of the way, they are together become unprofitable; there is none that doeth good, no, not one.
ROM|3|13|Their throat is an open sepulchre; with their tongues they have used deceit; the poison of asps is under their lips:
ROM|3|14|Whose mouth is full of cursing and bitterness:
ROM|3|15|Their feet are swift to shed blood:
ROM|3|16|Destruction and misery are in their ways:
ROM|3|17|And the way of peace have they not known:
ROM|3|18|There is no fear of God before their eyes.
ROM|3|19|Now we know that what things soever the law saith, it saith to them who are under the law: that every mouth may be stopped, and all the world may become guilty before God.
ROM|3|20|Therefore by the deeds of the law there shall no flesh be justified in his sight: for by the law is the knowledge of sin.
ROM|3|21|But now the righteousness of God without the law is manifested, being witnessed by the law and the prophets;
ROM|3|22|Even the righteousness of God which is by faith of Jesus Christ unto all and upon all them that believe: for there is no difference:
ROM|3|23|For all have sinned, and come short of the glory of God;
ROM|3|24|Being justified freely by his grace through the redemption that is in Christ Jesus:
ROM|3|25|Whom God hath set forth to be a propitiation through faith in his blood, to declare his righteousness for the remission of sins that are past, through the forbearance of God;
ROM|3|26|To declare, I say, at this time his righteousness: that he might be just, and the justifier of him which believeth in Jesus.
ROM|3|27|Where is boasting then? It is excluded. By what law? of works? Nay: but by the law of faith.
ROM|3|28|Therefore we conclude that a man is justified by faith without the deeds of the law.
ROM|3|29|Is he the God of the Jews only? is he not also of the Gentiles? Yes, of the Gentiles also:
ROM|3|30|Seeing it is one God, which shall justify the circumcision by faith, and uncircumcision through faith.
ROM|3|31|Do we then make void the law through faith? God forbid: yea, we establish the law.
ROM|4|1|What shall we say then that Abraham our father, as pertaining to the flesh, hath found?
ROM|4|2|For if Abraham were justified by works, he hath whereof to glory; but not before God.
ROM|4|3|For what saith the scripture? Abraham believed God, and it was counted unto him for righteousness.
ROM|4|4|Now to him that worketh is the reward not reckoned of grace, but of debt.
ROM|4|5|But to him that worketh not, but believeth on him that justifieth the ungodly, his faith is counted for righteousness.
ROM|4|6|Even as David also describeth the blessedness of the man, unto whom God imputeth righteousness without works,
ROM|4|7|Saying, Blessed are they whose iniquities are forgiven, and whose sins are covered.
ROM|4|8|Blessed is the man to whom the Lord will not impute sin.
ROM|4|9|Cometh this blessedness then upon the circumcision only, or upon the uncircumcision also? for we say that faith was reckoned to Abraham for righteousness.
ROM|4|10|How was it then reckoned? when he was in circumcision, or in uncircumcision? Not in circumcision, but in uncircumcision.
ROM|4|11|And he received the sign of circumcision, a seal of the righteousness of the faith which he had yet being uncircumcised: that he might be the father of all them that believe, though they be not circumcised; that righteousness might be imputed unto them also:
ROM|4|12|And the father of circumcision to them who are not of the circumcision only, but who also walk in the steps of that faith of our father Abraham, which he had being yet uncircumcised.
ROM|4|13|For the promise, that he should be the heir of the world, was not to Abraham, or to his seed, through the law, but through the righteousness of faith.
ROM|4|14|For if they which are of the law be heirs, faith is made void, and the promise made of none effect:
ROM|4|15|Because the law worketh wrath: for where no law is, there is no transgression.
ROM|4|16|Therefore it is of faith, that it might be by grace; to the end the promise might be sure to all the seed; not to that only which is of the law, but to that also which is of the faith of Abraham; who is the father of us all,
ROM|4|17|(As it is written, I have made thee a father of many nations,) before him whom he believed, even God, who quickeneth the dead, and calleth those things which be not as though they were.
ROM|4|18|Who against hope believed in hope, that he might become the father of many nations, according to that which was spoken, So shall thy seed be.
ROM|4|19|And being not weak in faith, he considered not his own body now dead, when he was about an hundred years old, neither yet the deadness of Sarah's womb:
ROM|4|20|He staggered not at the promise of God through unbelief; but was strong in faith, giving glory to God;
ROM|4|21|And being fully persuaded that, what he had promised, he was able also to perform.
ROM|4|22|And therefore it was imputed to him for righteousness.
ROM|4|23|Now it was not written for his sake alone, that it was imputed to him;
ROM|4|24|But for us also, to whom it shall be imputed, if we believe on him that raised up Jesus our Lord from the dead;
ROM|4|25|Who was delivered for our offences, and was raised again for our justification.
ROM|5|1|Therefore being justified by faith, we have peace with God through our Lord Jesus Christ:
ROM|5|2|By whom also we have access by faith into this grace wherein we stand, and rejoice in hope of the glory of God.
ROM|5|3|And not only so, but we glory in tribulations also: knowing that tribulation worketh patience;
ROM|5|4|And patience, experience; and experience, hope:
ROM|5|5|And hope maketh not ashamed; because the love of God is shed abroad in our hearts by the Holy Ghost which is given unto us.
ROM|5|6|For when we were yet without strength, in due time Christ died for the ungodly.
ROM|5|7|For scarcely for a righteous man will one die: yet peradventure for a good man some would even dare to die.
ROM|5|8|But God commendeth his love toward us, in that, while we were yet sinners, Christ died for us.
ROM|5|9|Much more then, being now justified by his blood, we shall be saved from wrath through him.
ROM|5|10|For if, when we were enemies, we were reconciled to God by the death of his Son, much more, being reconciled, we shall be saved by his life.
ROM|5|11|And not only so, but we also joy in God through our Lord Jesus Christ, by whom we have now received the atonement.
ROM|5|12|Wherefore, as by one man sin entered into the world, and death by sin; and so death passed upon all men, for that all have sinned:
ROM|5|13|(For until the law sin was in the world: but sin is not imputed when there is no law.
ROM|5|14|Nevertheless death reigned from Adam to Moses, even over them that had not sinned after the similitude of Adam's transgression, who is the figure of him that was to come.
ROM|5|15|But not as the offence, so also is the free gift. For if through the offence of one many be dead, much more the grace of God, and the gift by grace, which is by one man, Jesus Christ, hath abounded unto many.
ROM|5|16|And not as it was by one that sinned, so is the gift: for the judgment was by one to condemnation, but the free gift is of many offences unto justification.
ROM|5|17|For if by one man's offence death reigned by one; much more they which receive abundance of grace and of the gift of righteousness shall reign in life by one, Jesus Christ.)
ROM|5|18|Therefore as by the offence of one judgment came upon all men to condemnation; even so by the righteousness of one the free gift came upon all men unto justification of life.
ROM|5|19|For as by one man's disobedience many were made sinners, so by the obedience of one shall many be made righteous.
ROM|5|20|Moreover the law entered, that the offence might abound. But where sin abounded, grace did much more abound:
ROM|5|21|That as sin hath reigned unto death, even so might grace reign through righteousness unto eternal life by Jesus Christ our Lord.
ROM|6|1|What shall we say then? Shall we continue in sin, that grace may abound?
ROM|6|2|God forbid. How shall we, that are dead to sin, live any longer therein?
ROM|6|3|Know ye not, that so many of us as were baptized into Jesus Christ were baptized into his death?
ROM|6|4|Therefore we are buried with him by baptism into death: that like as Christ was raised up from the dead by the glory of the Father, even so we also should walk in newness of life.
ROM|6|5|For if we have been planted together in the likeness of his death, we shall be also in the likeness of his resurrection:
ROM|6|6|Knowing this, that our old man is crucified with him, that the body of sin might be destroyed, that henceforth we should not serve sin.
ROM|6|7|For he that is dead is freed from sin.
ROM|6|8|Now if we be dead with Christ, we believe that we shall also live with him:
ROM|6|9|Knowing that Christ being raised from the dead dieth no more; death hath no more dominion over him.
ROM|6|10|For in that he died, he died unto sin once: but in that he liveth, he liveth unto God.
ROM|6|11|Likewise reckon ye also yourselves to be dead indeed unto sin, but alive unto God through Jesus Christ our Lord.
ROM|6|12|Let not sin therefore reign in your mortal body, that ye should obey it in the lusts thereof.
ROM|6|13|Neither yield ye your members as instruments of unrighteousness unto sin: but yield yourselves unto God, as those that are alive from the dead, and your members as instruments of righteousness unto God.
ROM|6|14|For sin shall not have dominion over you: for ye are not under the law, but under grace.
ROM|6|15|What then? shall we sin, because we are not under the law, but under grace? God forbid.
ROM|6|16|Know ye not, that to whom ye yield yourselves servants to obey, his servants ye are to whom ye obey; whether of sin unto death, or of obedience unto righteousness?
ROM|6|17|But God be thanked, that ye were the servants of sin, but ye have obeyed from the heart that form of doctrine which was delivered you.
ROM|6|18|Being then made free from sin, ye became the servants of righteousness.
ROM|6|19|I speak after the manner of men because of the infirmity of your flesh: for as ye have yielded your members servants to uncleanness and to iniquity unto iniquity; even so now yield your members servants to righteousness unto holiness.
ROM|6|20|For when ye were the servants of sin, ye were free from righteousness.
ROM|6|21|What fruit had ye then in those things whereof ye are now ashamed? for the end of those things is death.
ROM|6|22|But now being made free from sin, and become servants to God, ye have your fruit unto holiness, and the end everlasting life.
ROM|6|23|For the wages of sin is death; but the gift of God is eternal life through Jesus Christ our Lord.
ROM|7|1|Know ye not, brethren, (for I speak to them that know the law,) how that the law hath dominion over a man as long as he liveth?
ROM|7|2|For the woman which hath an husband is bound by the law to her husband so long as he liveth; but if the husband be dead, she is loosed from the law of her husband.
ROM|7|3|So then if, while her husband liveth, she be married to another man, she shall be called an adulteress: but if her husband be dead, she is free from that law; so that she is no adulteress, though she be married to another man.
ROM|7|4|Wherefore, my brethren, ye also are become dead to the law by the body of Christ; that ye should be married to another, even to him who is raised from the dead, that we should bring forth fruit unto God.
ROM|7|5|For when we were in the flesh, the motions of sins, which were by the law, did work in our members to bring forth fruit unto death.
ROM|7|6|But now we are delivered from the law, that being dead wherein we were held; that we should serve in newness of spirit, and not in the oldness of the letter.
ROM|7|7|What shall we say then? Is the law sin? God forbid. Nay, I had not known sin, but by the law: for I had not known lust, except the law had said, Thou shalt not covet.
ROM|7|8|But sin, taking occasion by the commandment, wrought in me all manner of concupiscence. For without the law sin was dead.
ROM|7|9|For I was alive without the law once: but when the commandment came, sin revived, and I died.
ROM|7|10|And the commandment, which was ordained to life, I found to be unto death.
ROM|7|11|For sin, taking occasion by the commandment, deceived me, and by it slew me.
ROM|7|12|Wherefore the law is holy, and the commandment holy, and just, and good.
ROM|7|13|Was then that which is good made death unto me? God forbid. But sin, that it might appear sin, working death in me by that which is good; that sin by the commandment might become exceeding sinful.
ROM|7|14|For we know that the law is spiritual: but I am carnal, sold under sin.
ROM|7|15|For that which I do I allow not: for what I would, that do I not; but what I hate, that do I.
ROM|7|16|If then I do that which I would not, I consent unto the law that it is good.
ROM|7|17|Now then it is no more I that do it, but sin that dwelleth in me.
ROM|7|18|For I know that in me (that is, in my flesh,) dwelleth no good thing: for to will is present with me; but how to perform that which is good I find not.
ROM|7|19|For the good that I would I do not: but the evil which I would not, that I do.
ROM|7|20|Now if I do that I would not, it is no more I that do it, but sin that dwelleth in me.
ROM|7|21|I find then a law, that, when I would do good, evil is present with me.
ROM|7|22|For I delight in the law of God after the inward man:
ROM|7|23|But I see another law in my members, warring against the law of my mind, and bringing me into captivity to the law of sin which is in my members.
ROM|7|24|O wretched man that I am! who shall deliver me from the body of this death?
ROM|7|25|I thank God through Jesus Christ our Lord. So then with the mind I myself serve the law of God; but with the flesh the law of sin.
ROM|8|1|There is therefore now no condemnation to them which are in Christ Jesus, who walk not after the flesh, but after the Spirit.
ROM|8|2|For the law of the Spirit of life in Christ Jesus hath made me free from the law of sin and death.
ROM|8|3|For what the law could not do, in that it was weak through the flesh, God sending his own Son in the likeness of sinful flesh, and for sin, condemned sin in the flesh:
ROM|8|4|That the righteousness of the law might be fulfilled in us, who walk not after the flesh, but after the Spirit.
ROM|8|5|For they that are after the flesh do mind the things of the flesh; but they that are after the Spirit the things of the Spirit.
ROM|8|6|For to be carnally minded is death; but to be spiritually minded is life and peace.
ROM|8|7|Because the carnal mind is enmity against God: for it is not subject to the law of God, neither indeed can be.
ROM|8|8|So then they that are in the flesh cannot please God.
ROM|8|9|But ye are not in the flesh, but in the Spirit, if so be that the Spirit of God dwell in you. Now if any man have not the Spirit of Christ, he is none of his.
ROM|8|10|And if Christ be in you, the body is dead because of sin; but the Spirit is life because of righteousness.
ROM|8|11|But if the Spirit of him that raised up Jesus from the dead dwell in you, he that raised up Christ from the dead shall also quicken your mortal bodies by his Spirit that dwelleth in you.
ROM|8|12|Therefore, brethren, we are debtors, not to the flesh, to live after the flesh.
ROM|8|13|For if ye live after the flesh, ye shall die: but if ye through the Spirit do mortify the deeds of the body, ye shall live.
ROM|8|14|For as many as are led by the Spirit of God, they are the sons of God.
ROM|8|15|For ye have not received the spirit of bondage again to fear; but ye have received the Spirit of adoption, whereby we cry, Abba, Father.
ROM|8|16|The Spirit itself beareth witness with our spirit, that we are the children of God:
ROM|8|17|And if children, then heirs; heirs of God, and joint-heirs with Christ; if so be that we suffer with him, that we may be also glorified together.
ROM|8|18|For I reckon that the sufferings of this present time are not worthy to be compared with the glory which shall be revealed in us.
ROM|8|19|For the earnest expectation of the creature waiteth for the manifestation of the sons of God.
ROM|8|20|For the creature was made subject to vanity, not willingly, but by reason of him who hath subjected the same in hope,
ROM|8|21|Because the creature itself also shall be delivered from the bondage of corruption into the glorious liberty of the children of God.
ROM|8|22|For we know that the whole creation groaneth and travaileth in pain together until now.
ROM|8|23|And not only they, but ourselves also, which have the firstfruits of the Spirit, even we ourselves groan within ourselves, waiting for the adoption, to wit, the redemption of our body.
ROM|8|24|For we are saved by hope: but hope that is seen is not hope: for what a man seeth, why doth he yet hope for?
ROM|8|25|But if we hope for that we see not, then do we with patience wait for it.
ROM|8|26|Likewise the Spirit also helpeth our infirmities: for we know not what we should pray for as we ought: but the Spirit itself maketh intercession for us with groanings which cannot be uttered.
ROM|8|27|And he that searcheth the hearts knoweth what is the mind of the Spirit, because he maketh intercession for the saints according to the will of God.
ROM|8|28|And we know that all things work together for good to them that love God, to them who are the called according to his purpose.
ROM|8|29|For whom he did foreknow, he also did predestinate to be conformed to the image of his Son, that he might be the firstborn among many brethren.
ROM|8|30|Moreover whom he did predestinate, them he also called: and whom he called, them he also justified: and whom he justified, them he also glorified.
ROM|8|31|What shall we then say to these things? If God be for us, who can be against us?
ROM|8|32|He that spared not his own Son, but delivered him up for us all, how shall he not with him also freely give us all things?
ROM|8|33|Who shall lay any thing to the charge of God's elect? It is God that justifieth.
ROM|8|34|Who is he that condemneth? It is Christ that died, yea rather, that is risen again, who is even at the right hand of God, who also maketh intercession for us.
ROM|8|35|Who shall separate us from the love of Christ? shall tribulation, or distress, or persecution, or famine, or nakedness, or peril, or sword?
ROM|8|36|As it is written, For thy sake we are killed all the day long; we are accounted as sheep for the slaughter.
ROM|8|37|Nay, in all these things we are more than conquerors through him that loved us.
ROM|8|38|For I am persuaded, that neither death, nor life, nor angels, nor principalities, nor powers, nor things present, nor things to come,
ROM|8|39|Nor height, nor depth, nor any other creature, shall be able to separate us from the love of God, which is in Christ Jesus our Lord.
ROM|9|1|I say the truth in Christ, I lie not, my conscience also bearing me witness in the Holy Ghost,
ROM|9|2|That I have great heaviness and continual sorrow in my heart.
ROM|9|3|For I could wish that myself were accursed from Christ for my brethren, my kinsmen according to the flesh:
ROM|9|4|Who are Israelites; to whom pertaineth the adoption, and the glory, and the covenants, and the giving of the law, and the service of God, and the promises;
ROM|9|5|Whose are the fathers, and of whom as concerning the flesh Christ came, who is over all, God blessed for ever. Amen.
ROM|9|6|Not as though the word of God hath taken none effect. For they are not all Israel, which are of Israel:
ROM|9|7|Neither, because they are the seed of Abraham, are they all children: but, In Isaac shall thy seed be called.
ROM|9|8|That is, They which are the children of the flesh, these are not the children of God: but the children of the promise are counted for the seed.
ROM|9|9|For this is the word of promise, At this time will I come, and Sarah shall have a son.
ROM|9|10|And not only this; but when Rebecca also had conceived by one, even by our father Isaac;
ROM|9|11|(For the children being not yet born, neither having done any good or evil, that the purpose of God according to election might stand, not of works, but of him that calleth;)
ROM|9|12|It was said unto her, The elder shall serve the younger.
ROM|9|13|As it is written, Jacob have I loved, but Esau have I hated.
ROM|9|14|What shall we say then? Is there unrighteousness with God? God forbid.
ROM|9|15|For he saith to Moses, I will have mercy on whom I will have mercy, and I will have compassion on whom I will have compassion.
ROM|9|16|So then it is not of him that willeth, nor of him that runneth, but of God that sheweth mercy.
ROM|9|17|For the scripture saith unto Pharaoh, Even for this same purpose have I raised thee up, that I might shew my power in thee, and that my name might be declared throughout all the earth.
ROM|9|18|Therefore hath he mercy on whom he will have mercy, and whom he will he hardeneth.
ROM|9|19|Thou wilt say then unto me, Why doth he yet find fault? For who hath resisted his will?
ROM|9|20|Nay but, O man, who art thou that repliest against God? Shall the thing formed say to him that formed it, Why hast thou made me thus?
ROM|9|21|Hath not the potter power over the clay, of the same lump to make one vessel unto honour, and another unto dishonour?
ROM|9|22|What if God, willing to shew his wrath, and to make his power known, endured with much longsuffering the vessels of wrath fitted to destruction:
ROM|9|23|And that he might make known the riches of his glory on the vessels of mercy, which he had afore prepared unto glory,
ROM|9|24|Even us, whom he hath called, not of the Jews only, but also of the Gentiles?
ROM|9|25|As he saith also in Osee, I will call them my people, which were not my people; and her beloved, which was not beloved.
ROM|9|26|And it shall come to pass, that in the place where it was said unto them, Ye are not my people; there shall they be called the children of the living God.
ROM|9|27|Esaias also crieth concerning Israel, Though the number of the children of Israel be as the sand of the sea, a remnant shall be saved:
ROM|9|28|For he will finish the work, and cut it short in righteousness: because a short work will the Lord make upon the earth.
ROM|9|29|And as Esaias said before, Except the Lord of Sabaoth had left us a seed, we had been as Sodoma, and been made like unto Gomorrha.
ROM|9|30|What shall we say then? That the Gentiles, which followed not after righteousness, have attained to righteousness, even the righteousness which is of faith.
ROM|9|31|But Israel, which followed after the law of righteousness, hath not attained to the law of righteousness.
ROM|9|32|Wherefore? Because they sought it not by faith, but as it were by the works of the law. For they stumbled at that stumblingstone;
ROM|9|33|As it is written, Behold, I lay in Sion a stumblingstone and rock of offence: and whosoever believeth on him shall not be ashamed.
ROM|10|1|Brethren, my heart's desire and prayer to God for Israel is, that they might be saved.
ROM|10|2|For I bear them record that they have a zeal of God, but not according to knowledge.
ROM|10|3|For they being ignorant of God's righteousness, and going about to establish their own righteousness, have not submitted themselves unto the righteousness of God.
ROM|10|4|For Christ is the end of the law for righteousness to every one that believeth.
ROM|10|5|For Moses describeth the righteousness which is of the law, That the man which doeth those things shall live by them.
ROM|10|6|But the righteousness which is of faith speaketh on this wise, Say not in thine heart, Who shall ascend into heaven? (that is, to bring Christ down from above:)
ROM|10|7|Or, Who shall descend into the deep? (that is, to bring up Christ again from the dead.)
ROM|10|8|But what saith it? The word is nigh thee, even in thy mouth, and in thy heart: that is, the word of faith, which we preach;
ROM|10|9|That if thou shalt confess with thy mouth the Lord Jesus, and shalt believe in thine heart that God hath raised him from the dead, thou shalt be saved.
ROM|10|10|For with the heart man believeth unto righteousness; and with the mouth confession is made unto salvation.
ROM|10|11|For the scripture saith, Whosoever believeth on him shall not be ashamed.
ROM|10|12|For there is no difference between the Jew and the Greek: for the same Lord over all is rich unto all that call upon him.
ROM|10|13|For whosoever shall call upon the name of the Lord shall be saved.
ROM|10|14|How then shall they call on him in whom they have not believed? and how shall they believe in him of whom they have not heard? and how shall they hear without a preacher?
ROM|10|15|And how shall they preach, except they be sent? as it is written, How beautiful are the feet of them that preach the gospel of peace, and bring glad tidings of good things!
ROM|10|16|But they have not all obeyed the gospel. For Esaias saith, Lord, who hath believed our report?
ROM|10|17|So then faith cometh by hearing, and hearing by the word of God.
ROM|10|18|But I say, Have they not heard? Yes verily, their sound went into all the earth, and their words unto the ends of the world.
ROM|10|19|But I say, Did not Israel know? First Moses saith, I will provoke you to jealousy by them that are no people, and by a foolish nation I will anger you.
ROM|10|20|But Esaias is very bold, and saith, I was found of them that sought me not; I was made manifest unto them that asked not after me.
ROM|10|21|But to Israel he saith, All day long I have stretched forth my hands unto a disobedient and gainsaying people.
ROM|11|1|I say then, Hath God cast away his people? God forbid. For I also am an Israelite, of the seed of Abraham, of the tribe of Benjamin.
ROM|11|2|God hath not cast away his people which he foreknew. Wot ye not what the scripture saith of Elias? how he maketh intercession to God against Israel saying,
ROM|11|3|Lord, they have killed thy prophets, and digged down thine altars; and I am left alone, and they seek my life.
ROM|11|4|But what saith the answer of God unto him? I have reserved to myself seven thousand men, who have not bowed the knee to the image of Baal.
ROM|11|5|Even so then at this present time also there is a remnant according to the election of grace.
ROM|11|6|And if by grace, then is it no more of works: otherwise grace is no more grace. But if it be of works, then it is no more grace: otherwise work is no more work.
ROM|11|7|What then? Israel hath not obtained that which he seeketh for; but the election hath obtained it, and the rest were blinded.
ROM|11|8|(According as it is written, God hath given them the spirit of slumber, eyes that they should not see, and ears that they should not hear;) unto this day.
ROM|11|9|And David saith, Let their table be made a snare, and a trap, and a stumblingblock, and a recompence unto them:
ROM|11|10|Let their eyes be darkened, that they may not see, and bow down their back alway.
ROM|11|11|I say then, Have they stumbled that they should fall? God forbid: but rather through their fall salvation is come unto the Gentiles, for to provoke them to jealousy.
ROM|11|12|Now if the fall of them be the riches of the world, and the diminishing of them the riches of the Gentiles; how much more their fulness?
ROM|11|13|For I speak to you Gentiles, inasmuch as I am the apostle of the Gentiles, I magnify mine office:
ROM|11|14|If by any means I may provoke to emulation them which are my flesh, and might save some of them.
ROM|11|15|For if the casting away of them be the reconciling of the world, what shall the receiving of them be, but life from the dead?
ROM|11|16|For if the firstfruit be holy, the lump is also holy: and if the root be holy, so are the branches.
ROM|11|17|And if some of the branches be broken off, and thou, being a wild olive tree, wert graffed in among them, and with them partakest of the root and fatness of the olive tree;
ROM|11|18|Boast not against the branches. But if thou boast, thou bearest not the root, but the root thee.
ROM|11|19|Thou wilt say then, The branches were broken off, that I might be graffed in.
ROM|11|20|Well; because of unbelief they were broken off, and thou standest by faith. Be not highminded, but fear:
ROM|11|21|For if God spared not the natural branches, take heed lest he also spare not thee.
ROM|11|22|Behold therefore the goodness and severity of God: on them which fell, severity; but toward thee, goodness, if thou continue in his goodness: otherwise thou also shalt be cut off.
ROM|11|23|And they also, if they abide not still in unbelief, shall be graffed in: for God is able to graff them in again.
ROM|11|24|For if thou wert cut out of the olive tree which is wild by nature, and wert graffed contrary to nature into a good olive tree: how much more shall these, which be the natural branches, be graffed into their own olive tree?
ROM|11|25|For I would not, brethren, that ye should be ignorant of this mystery, lest ye should be wise in your own conceits; that blindness in part is happened to Israel, until the fulness of the Gentiles be come in.
ROM|11|26|And so all Israel shall be saved: as it is written, There shall come out of Sion the Deliverer, and shall turn away ungodliness from Jacob:
ROM|11|27|For this is my covenant unto them, when I shall take away their sins.
ROM|11|28|As concerning the gospel, they are enemies for your sakes: but as touching the election, they are beloved for the father's sakes.
ROM|11|29|For the gifts and calling of God are without repentance.
ROM|11|30|For as ye in times past have not believed God, yet have now obtained mercy through their unbelief:
ROM|11|31|Even so have these also now not believed, that through your mercy they also may obtain mercy.
ROM|11|32|For God hath concluded them all in unbelief, that he might have mercy upon all.
ROM|11|33|O the depth of the riches both of the wisdom and knowledge of God! how unsearchable are his judgments, and his ways past finding out!
ROM|11|34|For who hath known the mind of the Lord? or who hath been his counsellor?
ROM|11|35|Or who hath first given to him, and it shall be recompensed unto him again?
ROM|11|36|For of him, and through him, and to him, are all things: to whom be glory for ever. Amen.
ROM|12|1|I beseech you therefore, brethren, by the mercies of God, that ye present your bodies a living sacrifice, holy, acceptable unto God, which is your reasonable service.
ROM|12|2|And be not conformed to this world: but be ye transformed by the renewing of your mind, that ye may prove what is that good, and acceptable, and perfect, will of God.
ROM|12|3|For I say, through the grace given unto me, to every man that is among you, not to think of himself more highly than he ought to think; but to think soberly, according as God hath dealt to every man the measure of faith.
ROM|12|4|For as we have many members in one body, and all members have not the same office:
ROM|12|5|So we, being many, are one body in Christ, and every one members one of another.
ROM|12|6|Having then gifts differing according to the grace that is given to us, whether prophecy, let us prophesy according to the proportion of faith;
ROM|12|7|Or ministry, let us wait on our ministering: or he that teacheth, on teaching;
ROM|12|8|Or he that exhorteth, on exhortation: he that giveth, let him do it with simplicity; he that ruleth, with diligence; he that sheweth mercy, with cheerfulness.
ROM|12|9|Let love be without dissimulation. Abhor that which is evil; cleave to that which is good.
ROM|12|10|Be kindly affectioned one to another with brotherly love; in honour preferring one another;
ROM|12|11|Not slothful in business; fervent in spirit; serving the Lord;
ROM|12|12|Rejoicing in hope; patient in tribulation; continuing instant in prayer;
ROM|12|13|Distributing to the necessity of saints; given to hospitality.
ROM|12|14|Bless them which persecute you: bless, and curse not.
ROM|12|15|Rejoice with them that do rejoice, and weep with them that weep.
ROM|12|16|Be of the same mind one toward another. Mind not high things, but condescend to men of low estate. Be not wise in your own conceits.
ROM|12|17|Recompense to no man evil for evil. Provide things honest in the sight of all men.
ROM|12|18|If it be possible, as much as lieth in you, live peaceably with all men.
ROM|12|19|Dearly beloved, avenge not yourselves, but rather give place unto wrath: for it is written, Vengeance is mine; I will repay, saith the Lord.
ROM|12|20|Therefore if thine enemy hunger, feed him; if he thirst, give him drink: for in so doing thou shalt heap coals of fire on his head.
ROM|12|21|Be not overcome of evil, but overcome evil with good.
ROM|13|1|Let every soul be subject unto the higher powers. For there is no power but of God: the powers that be are ordained of God.
ROM|13|2|Whosoever therefore resisteth the power, resisteth the ordinance of God: and they that resist shall receive to themselves damnation.
ROM|13|3|For rulers are not a terror to good works, but to the evil. Wilt thou then not be afraid of the power? do that which is good, and thou shalt have praise of the same:
ROM|13|4|For he is the minister of God to thee for good. But if thou do that which is evil, be afraid; for he beareth not the sword in vain: for he is the minister of God, a revenger to execute wrath upon him that doeth evil.
ROM|13|5|Wherefore ye must needs be subject, not only for wrath, but also for conscience sake.
ROM|13|6|For for this cause pay ye tribute also: for they are God's ministers, attending continually upon this very thing.
ROM|13|7|Render therefore to all their dues: tribute to whom tribute is due; custom to whom custom; fear to whom fear; honour to whom honour.
ROM|13|8|Owe no man any thing, but to love one another: for he that loveth another hath fulfilled the law.
ROM|13|9|For this, Thou shalt not commit adultery, Thou shalt not kill, Thou shalt not steal, Thou shalt not bear false witness, Thou shalt not covet; and if there be any other commandment, it is briefly comprehended in this saying, namely, Thou shalt love thy neighbour as thyself.
ROM|13|10|Love worketh no ill to his neighbour: therefore love is the fulfilling of the law.
ROM|13|11|And that, knowing the time, that now it is high time to awake out of sleep: for now is our salvation nearer than when we believed.
ROM|13|12|The night is far spent, the day is at hand: let us therefore cast off the works of darkness, and let us put on the armour of light.
ROM|13|13|Let us walk honestly, as in the day; not in rioting and drunkenness, not in chambering and wantonness, not in strife and envying.
ROM|13|14|But put ye on the Lord Jesus Christ, and make not provision for the flesh, to fulfil the lusts thereof.
ROM|14|1|Him that is weak in the faith receive ye, but not to doubtful disputations.
ROM|14|2|For one believeth that he may eat all things: another, who is weak, eateth herbs.
ROM|14|3|Let not him that eateth despise him that eateth not; and let not him which eateth not judge him that eateth: for God hath received him.
ROM|14|4|Who art thou that judgest another man's servant? to his own master he standeth or falleth. Yea, he shall be holden up: for God is able to make him stand.
ROM|14|5|One man esteemeth one day above another: another esteemeth every day alike. Let every man be fully persuaded in his own mind.
ROM|14|6|He that regardeth the day, regardeth it unto the Lord; and he that regardeth not the day, to the Lord he doth not regard it. He that eateth, eateth to the Lord, for he giveth God thanks; and he that eateth not, to the Lord he eateth not, and giveth God thanks.
ROM|14|7|For none of us liveth to himself, and no man dieth to himself.
ROM|14|8|For whether we live, we live unto the Lord; and whether we die, we die unto the Lord: whether we live therefore, or die, we are the Lord's.
ROM|14|9|For to this end Christ both died, and rose, and revived, that he might be Lord both of the dead and living.
ROM|14|10|But why dost thou judge thy brother? or why dost thou set at nought thy brother? for we shall all stand before the judgment seat of Christ.
ROM|14|11|For it is written, As I live, saith the Lord, every knee shall bow to me, and every tongue shall confess to God.
ROM|14|12|So then every one of us shall give account of himself to God.
ROM|14|13|Let us not therefore judge one another any more: but judge this rather, that no man put a stumblingblock or an occasion to fall in his brother's way.
ROM|14|14|I know, and am persuaded by the Lord Jesus, that there is nothing unclean of itself: but to him that esteemeth any thing to be unclean, to him it is unclean.
ROM|14|15|But if thy brother be grieved with thy meat, now walkest thou not charitably. Destroy not him with thy meat, for whom Christ died.
ROM|14|16|Let not then your good be evil spoken of:
ROM|14|17|For the kingdom of God is not meat and drink; but righteousness, and peace, and joy in the Holy Ghost.
ROM|14|18|For he that in these things serveth Christ is acceptable to God, and approved of men.
ROM|14|19|Let us therefore follow after the things which make for peace, and things wherewith one may edify another.
ROM|14|20|For meat destroy not the work of God. All things indeed are pure; but it is evil for that man who eateth with offence.
ROM|14|21|It is good neither to eat flesh, nor to drink wine, nor any thing whereby thy brother stumbleth, or is offended, or is made weak.
ROM|14|22|Hast thou faith? have it to thyself before God. Happy is he that condemneth not himself in that thing which he alloweth.
ROM|14|23|And he that doubteth is damned if he eat, because he eateth not of faith: for whatsoever is not of faith is sin.
ROM|15|1|We then that are strong ought to bear the infirmities of the weak, and not to please ourselves.
ROM|15|2|Let every one of us please his neighbour for his good to edification.
ROM|15|3|For even Christ pleased not himself; but, as it is written, The reproaches of them that reproached thee fell on me.
ROM|15|4|For whatsoever things were written aforetime were written for our learning, that we through patience and comfort of the scriptures might have hope.
ROM|15|5|Now the God of patience and consolation grant you to be likeminded one toward another according to Christ Jesus:
ROM|15|6|That ye may with one mind and one mouth glorify God, even the Father of our Lord Jesus Christ.
ROM|15|7|Wherefore receive ye one another, as Christ also received us to the glory of God.
ROM|15|8|Now I say that Jesus Christ was a minister of the circumcision for the truth of God, to confirm the promises made unto the fathers:
ROM|15|9|And that the Gentiles might glorify God for his mercy; as it is written, For this cause I will confess to thee among the Gentiles, and sing unto thy name.
ROM|15|10|And again he saith, Rejoice, ye Gentiles, with his people.
ROM|15|11|And again, Praise the Lord, all ye Gentiles; and laud him, all ye people.
ROM|15|12|And again, Esaias saith, There shall be a root of Jesse, and he that shall rise to reign over the Gentiles; in him shall the Gentiles trust.
ROM|15|13|Now the God of hope fill you with all joy and peace in believing, that ye may abound in hope, through the power of the Holy Ghost.
ROM|15|14|And I myself also am persuaded of you, my brethren, that ye also are full of goodness, filled with all knowledge, able also to admonish one another.
ROM|15|15|Nevertheless, brethren, I have written the more boldly unto you in some sort, as putting you in mind, because of the grace that is given to me of God,
ROM|15|16|That I should be the minister of Jesus Christ to the Gentiles, ministering the gospel of God, that the offering up of the Gentiles might be acceptable, being sanctified by the Holy Ghost.
ROM|15|17|I have therefore whereof I may glory through Jesus Christ in those things which pertain to God.
ROM|15|18|For I will not dare to speak of any of those things which Christ hath not wrought by me, to make the Gentiles obedient, by word and deed,
ROM|15|19|Through mighty signs and wonders, by the power of the Spirit of God; so that from Jerusalem, and round about unto Illyricum, I have fully preached the gospel of Christ.
ROM|15|20|Yea, so have I strived to preach the gospel, not where Christ was named, lest I should build upon another man's foundation:
ROM|15|21|But as it is written, To whom he was not spoken of, they shall see: and they that have not heard shall understand.
ROM|15|22|For which cause also I have been much hindered from coming to you.
ROM|15|23|But now having no more place in these parts, and having a great desire these many years to come unto you;
ROM|15|24|Whensoever I take my journey into Spain, I will come to you: for I trust to see you in my journey, and to be brought on my way thitherward by you, if first I be somewhat filled with your company.
ROM|15|25|But now I go unto Jerusalem to minister unto the saints.
ROM|15|26|For it hath pleased them of Macedonia and Achaia to make a certain contribution for the poor saints which are at Jerusalem.
ROM|15|27|It hath pleased them verily; and their debtors they are. For if the Gentiles have been made partakers of their spiritual things, their duty is also to minister unto them in carnal things.
ROM|15|28|When therefore I have performed this, and have sealed to them this fruit, I will come by you into Spain.
ROM|15|29|And I am sure that, when I come unto you, I shall come in the fulness of the blessing of the gospel of Christ.
ROM|15|30|Now I beseech you, brethren, for the Lord Jesus Christ's sake, and for the love of the Spirit, that ye strive together with me in your prayers to God for me;
ROM|15|31|That I may be delivered from them that do not believe in Judaea; and that my service which I have for Jerusalem may be accepted of the saints;
ROM|15|32|That I may come unto you with joy by the will of God, and may with you be refreshed.
ROM|15|33|Now the God of peace be with you all. Amen.
ROM|16|1|I commend unto you Phebe our sister, which is a servant of the church which is at Cenchrea:
ROM|16|2|That ye receive her in the Lord, as becometh saints, and that ye assist her in whatsoever business she hath need of you: for she hath been a succourer of many, and of myself also.
ROM|16|3|Greet Priscilla and Aquila my helpers in Christ Jesus:
ROM|16|4|Who have for my life laid down their own necks: unto whom not only I give thanks, but also all the churches of the Gentiles.
ROM|16|5|Likewise greet the church that is in their house. Salute my well-beloved Epaenetus, who is the firstfruits of Achaia unto Christ.
ROM|16|6|Greet Mary, who bestowed much labour on us.
ROM|16|7|Salute Andronicus and Junia, my kinsmen, and my fellow-prisoners, who are of note among the apostles, who also were in Christ before me.
ROM|16|8|Greet Amplias my beloved in the Lord.
ROM|16|9|Salute Urbane, our helper in Christ, and Stachys my beloved.
ROM|16|10|Salute Apelles approved in Christ. Salute them which are of Aristobulus' household.
ROM|16|11|Salute Herodion my kinsman. Greet them that be of the household of Narcissus, which are in the Lord.
ROM|16|12|Salute Tryphena and Tryphosa, who labour in the Lord. Salute the beloved Persis, which laboured much in the Lord.
ROM|16|13|Salute Rufus chosen in the Lord, and his mother and mine.
ROM|16|14|Salute Asyncritus, Phlegon, Hermas, Patrobas, Hermes, and the brethren which are with them.
ROM|16|15|Salute Philologus, and Julia, Nereus, and his sister, and Olympas, and all the saints which are with them.
ROM|16|16|Salute one another with an holy kiss. The churches of Christ salute you.
ROM|16|17|Now I beseech you, brethren, mark them which cause divisions and offences contrary to the doctrine which ye have learned; and avoid them.
ROM|16|18|For they that are such serve not our Lord Jesus Christ, but their own belly; and by good words and fair speeches deceive the hearts of the simple.
ROM|16|19|For your obedience is come abroad unto all men. I am glad therefore on your behalf: but yet I would have you wise unto that which is good, and simple concerning evil.
ROM|16|20|And the God of peace shall bruise Satan under your feet shortly. The grace of our Lord Jesus Christ be with you. Amen.
ROM|16|21|Timotheus my workfellow, and Lucius, and Jason, and Sosipater, my kinsmen, salute you.
ROM|16|22|I Tertius, who wrote this epistle, salute you in the Lord.
ROM|16|23|Gaius mine host, and of the whole church, saluteth you. Erastus the chamberlain of the city saluteth you, and Quartus a brother.
ROM|16|24|The grace of our Lord Jesus Christ be with you all. Amen.
ROM|16|25|Now to him that is of power to stablish you according to my gospel, and the preaching of Jesus Christ, according to the revelation of the mystery, which was kept secret since the world began,
ROM|16|26|But now is made manifest, and by the scriptures of the prophets, according to the commandment of the everlasting God, made known to all nations for the obedience of faith:
ROM|16|27|To God only wise, be glory through Jesus Christ for ever. Amen.
