1PET|1|1|Петр, Апостол Иисуса Христа, пришельцам, рассеянным в Понте, Галатии, Каппадокии, Асии и Вифинии, избранным,
1PET|1|2|по предведению Бога Отца, при освящении от Духа, к послушанию и окроплению Кровию Иисуса Христа: благодать вам и мир да умножится.
1PET|1|3|Благословен Бог и Отец Господа нашего Иисуса Христа, по великой Своей милости возродивший нас воскресением Иисуса Христа из мертвых к упованию живому,
1PET|1|4|к наследству нетленному, чистому, неувядаемому, хранящемуся на небесах для вас,
1PET|1|5|силою Божиею через веру соблюдаемых ко спасению, готовому открыться в последнее время.
1PET|1|6|О сем радуйтесь, поскорбев теперь немного, если нужно, от различных искушений,
1PET|1|7|дабы испытанная вера ваша оказалась драгоценнее гибнущего, хотя и огнем испытываемого золота, к похвале и чести и славе в явление Иисуса Христа,
1PET|1|8|Которого, не видев, любите, и Которого доселе не видя, но веруя в Него, радуетесь радостью неизреченною и преславною,
1PET|1|9|достигая наконец верою вашею спасения душ.
1PET|1|10|К сему–то спасению относились изыскания и исследования пророков, которые предсказывали о назначенной вам благодати,
1PET|1|11|исследывая, на которое и на какое время указывал сущий в них Дух Христов, когда Он предвозвещал Христовы страдания и последующую за ними славу.
1PET|1|12|Им открыто было, что не им самим, а нам служило то, что ныне проповедано вам благовествовавшими Духом Святым, посланным с небес, во что желают проникнуть Ангелы.
1PET|1|13|Посему, (возлюбленные), препоясав чресла ума вашего, бодрствуя, совершенно уповайте на подаваемую вам благодать в явлении Иисуса Христа.
1PET|1|14|Как послушные дети, не сообразуйтесь с прежними похотями, бывшими в неведении вашем,
1PET|1|15|но, по примеру призвавшего вас Святаго, и сами будьте святы во всех поступках.
1PET|1|16|Ибо написано: будьте святы, потому что Я свят.
1PET|1|17|И если вы называете Отцем Того, Который нелицеприятно судит каждого по делам, то со страхом проводите время странствования вашего,
1PET|1|18|зная, что не тленным серебром или золотом искуплены вы от суетной жизни, преданной вам от отцов,
1PET|1|19|но драгоценною Кровию Христа, как непорочного и чистого Агнца,
1PET|1|20|предназначенного еще прежде создания мира, но явившегося в последние времена для вас,
1PET|1|21|уверовавших чрез Него в Бога, Который воскресил Его из мертвых и дал Ему славу, чтобы вы имели веру и упование на Бога.
1PET|1|22|Послушанием истине чрез Духа, очистив души ваши к нелицемерному братолюбию, постоянно любите друг друга от чистого сердца,
1PET|1|23|[как] возрожденные не от тленного семени, но от нетленного, от слова Божия, живаго и пребывающего вовек.
1PET|1|24|Ибо всякая плоть – как трава, и всякая слава человеческая – как цвет на траве: засохла трава, и цвет ее опал;
1PET|1|25|но слово Господне пребывает вовек; а это есть то слово, которое вам проповедано.
1PET|2|1|Итак, отложив всякую злобу и всякое коварство, и лицемерие, и зависть, и всякое злословие,
1PET|2|2|как новорожденные младенцы, возлюбите чистое словесное молоко, дабы от него возрасти вам во спасение;
1PET|2|3|ибо вы вкусили, что благ Господь.
1PET|2|4|Приступая к Нему, камню живому, человеками отверженному, но Богом избранному, драгоценному,
1PET|2|5|и сами, как живые камни, устрояйте из себя дом духовный, священство святое, чтобы приносить духовные жертвы, благоприятные Богу Иисусом Христом.
1PET|2|6|Ибо сказано в Писании: вот, Я полагаю в Сионе камень краеугольный, избранный, драгоценный; и верующий в Него не постыдится.
1PET|2|7|Итак Он для вас, верующих, драгоценность, а для неверующих камень, который отвергли строители, но который сделался главою угла, камень претыкания и камень соблазна,
1PET|2|8|о который они претыкаются, не покоряясь слову, на что они и оставлены.
1PET|2|9|Но вы – род избранный, царственное священство, народ святой, люди, взятые в удел, дабы возвещать совершенства Призвавшего вас из тьмы в чудный Свой свет;
1PET|2|10|некогда не народ, а ныне народ Божий; [некогда] непомилованные, а ныне помилованы.
1PET|2|11|Возлюбленные! прошу вас, как пришельцев и странников, удаляться от плотских похотей, восстающих на душу,
1PET|2|12|и провождать добродетельную жизнь между язычниками, дабы они за то, за что злословят вас, как злодеев, увидя добрые дела ваши, прославили Бога в день посещения.
1PET|2|13|Итак будьте покорны всякому человеческому начальству, для Господа: царю ли, как верховной власти,
1PET|2|14|правителям ли, как от него посылаемым для наказания преступников и для поощрения делающих добро, –
1PET|2|15|ибо такова есть воля Божия, чтобы мы, делая добро, заграждали уста невежеству безумных людей, –
1PET|2|16|как свободные, не как употребляющие свободу для прикрытия зла, но как рабы Божии.
1PET|2|17|Всех почитайте, братство любите, Бога бойтесь, царя чтите.
1PET|2|18|Слуги, со всяким страхом повинуйтесь господам, не только добрым и кротким, но и суровым.
1PET|2|19|Ибо то угодно Богу, если кто, помышляя о Боге, переносит скорби, страдая несправедливо.
1PET|2|20|Ибо что за похвала, если вы терпите, когда вас бьют за проступки? Но если, делая добро и страдая, терпите, это угодно Богу.
1PET|2|21|Ибо вы к тому призваны, потому что и Христос пострадал за нас, оставив нам пример, дабы мы шли по следам Его.
1PET|2|22|Он не сделал никакого греха, и не было лести в устах Его.
1PET|2|23|Будучи злословим, Он не злословил взаимно; страдая, не угрожал, но предавал то Судии Праведному.
1PET|2|24|Он грехи наши Сам вознес телом Своим на древо, дабы мы, избавившись от грехов, жили для правды: ранами Его вы исцелились.
1PET|2|25|Ибо вы были, как овцы блуждающие (не имея пастыря), но возвратились ныне к Пастырю и Блюстителю душ ваших.
1PET|3|1|Также и вы, жены, повинуйтесь своим мужьям, чтобы те из них, которые не покоряются слову, житием жен своих без слова приобретаемы были,
1PET|3|2|когда увидят ваше чистое, богобоязненное житие.
1PET|3|3|Да будет украшением вашим не внешнее плетение волос, не золотые уборы или нарядность в одежде,
1PET|3|4|но сокровенный сердца человек в нетленной [красоте] кроткого и молчаливого духа, что драгоценно пред Богом.
1PET|3|5|Так некогда и святые жены, уповавшие на Бога, украшали себя, повинуясь своим мужьям.
1PET|3|6|Так Сарра повиновалась Аврааму, называя его господином. Вы – дети ее, если делаете добро и не смущаетесь ни от какого страха.
1PET|3|7|Также и вы, мужья, обращайтесь благоразумно с женами, как с немощнейшим сосудом, оказывая им честь, как сонаследницам благодатной жизни, дабы не было вам препятствия в молитвах.
1PET|3|8|Наконец будьте все единомысленны, сострадательны, братолюбивы, милосерды, дружелюбны, смиренномудры;
1PET|3|9|не воздавайте злом за зло или ругательством за ругательство; напротив, благословляйте, зная, что вы к тому призваны, чтобы наследовать благословение.
1PET|3|10|Ибо, кто любит жизнь и хочет видеть добрые дни, тот удерживай язык свой от зла и уста свои от лукавых речей;
1PET|3|11|уклоняйся от зла и делай добро; ищи мира и стремись к нему,
1PET|3|12|потому что очи Господа [обращены] к праведным и уши Его к молитве их, но лице Господне против делающих зло, (чтобы истребить их с земли).
1PET|3|13|И кто сделает вам зло, если вы будете ревнителями доброго?
1PET|3|14|Но если и страдаете за правду, то вы блаженны; а страха их не бойтесь и не смущайтесь.
1PET|3|15|Господа Бога святите в сердцах ваших; [будьте] всегда готовы всякому, требующему у вас отчета в вашем уповании, дать ответ с кротостью и благоговением.
1PET|3|16|Имейте добрую совесть, дабы тем, за что злословят вас, как злодеев, были постыжены порицающие ваше доброе житие во Христе.
1PET|3|17|Ибо, если угодно воле Божией, лучше пострадать за добрые дела, нежели за злые;
1PET|3|18|потому что и Христос, чтобы привести нас к Богу, однажды пострадал за грехи наши, праведник за неправедных, быв умерщвлен по плоти, но ожив духом,
1PET|3|19|которым Он и находящимся в темнице духам, сойдя, проповедал,
1PET|3|20|некогда непокорным ожидавшему их Божию долготерпению, во дни Ноя, во время строения ковчега, в котором немногие, то есть восемь душ, спаслись от воды.
1PET|3|21|Так и нас ныне подобное сему образу крещение, не плотской нечистоты омытие, но обещание Богу доброй совести, спасает воскресением Иисуса Христа,
1PET|3|22|Который, восшед на небо, пребывает одесную Бога и Которому покорились Ангелы и Власти и Силы.
1PET|4|1|Итак, как Христос пострадал за нас плотию, то и вы вооружитесь тою же мыслью; ибо страдающий плотию перестает грешить,
1PET|4|2|чтобы остальное во плоти время жить уже не по человеческим похотям, но по воле Божией.
1PET|4|3|Ибо довольно, что вы в прошедшее время жизни поступали по воле языческой, предаваясь нечистотам, похотям (мужеложству, скотоложству, помыслам), пьянству, излишеству в пище и питии и нелепому идолослужению;
1PET|4|4|почему они и дивятся, что вы не участвуете с ними в том же распутстве, и злословят вас.
1PET|4|5|Они дадут ответ Имеющему вскоре судить живых и мертвых.
1PET|4|6|Ибо для того и мертвым было благовествуемо, чтобы они, подвергшись суду по человеку плотию, жили по Богу духом.
1PET|4|7|Впрочем близок всему конец. Итак будьте благоразумны и бодрствуйте в молитвах.
1PET|4|8|Более же всего имейте усердную любовь друг ко другу, потому что любовь покрывает множество грехов.
1PET|4|9|Будьте страннолюбивы друг ко другу без ропота.
1PET|4|10|Служите друг другу, каждый тем даром, какой получил, как добрые домостроители многоразличной благодати Божией.
1PET|4|11|Говорит ли кто, [говори] как слова Божии; служит ли кто, [служи] по силе, какую дает Бог, дабы во всем прославлялся Бог через Иисуса Христа, Которому слава и держава во веки веков. Аминь.
1PET|4|12|Возлюбленные! огненного искушения, для испытания вам посылаемого, не чуждайтесь, как приключения для вас странного,
1PET|4|13|но как вы участвуете в Христовых страданиях, радуйтесь, да и в явление славы Его возрадуетесь и восторжествуете.
1PET|4|14|Если злословят вас за имя Христово, то вы блаженны, ибо Дух Славы, Дух Божий почивает на вас. Теми Он хулится, а вами прославляется.
1PET|4|15|Только бы не пострадал кто из вас, как убийца, или вор, или злодей, или как посягающий на чужое;
1PET|4|16|а если как Христианин, то не стыдись, но прославляй Бога за такую участь.
1PET|4|17|Ибо время начаться суду с дома Божия; если же прежде с нас [начнется], то какой конец непокоряющимся Евангелию Божию?
1PET|4|18|И если праведник едва спасается, то нечестивый и грешный где явится?
1PET|4|19|Итак страждущие по воле Божией да предадут Ему, как верному Создателю, души свои, делая добро.
1PET|5|1|Пастырей ваших умоляю я, сопастырь и свидетель страданий Христовых и соучастник в славе, которая должна открыться:
1PET|5|2|пасите Божие стадо, какое у вас, надзирая за ним не принужденно, но охотно и богоугодно, не для гнусной корысти, но из усердия,
1PET|5|3|и не господствуя над наследием [Божиим], но подавая пример стаду;
1PET|5|4|и когда явится Пастыреначальник, вы получите неувядающий венец славы.
1PET|5|5|Также и младшие, повинуйтесь пастырям; все же, подчиняясь друг другу, облекитесь смиренномудрием, потому что Бог гордым противится, а смиренным дает благодать.
1PET|5|6|Итак смиритесь под крепкую руку Божию, да вознесет вас в свое время.
1PET|5|7|Все заботы ваши возложите на Него, ибо Он печется о вас.
1PET|5|8|Трезвитесь, бодрствуйте, потому что противник ваш диавол ходит, как рыкающий лев, ища, кого поглотить.
1PET|5|9|Противостойте ему твердою верою, зная, что такие же страдания случаются и с братьями вашими в мире.
1PET|5|10|Бог же всякой благодати, призвавший нас в вечную славу Свою во Христе Иисусе, Сам, по кратковременном страдании вашем, да совершит вас, да утвердит, да укрепит, да соделает непоколебимыми.
1PET|5|11|Ему слава и держава во веки веков. Аминь.
1PET|5|12|Сие кратко написал я вам чрез Силуана, верного, как думаю, вашего брата, чтобы уверить вас, утешая и свидетельствуя, что это истинная благодать Божия, в которой вы стоите.
1PET|5|13|Приветствует вас избранная, подобно [вам, церковь] в Вавилоне и Марк, сын мой.
1PET|5|14|Приветствуйте друг друга лобзанием любви. Мир вам всем во Христе Иисусе. Аминь.
