MAL|1|1|An oracle: The word of the LORD to Israel through Malachi.
MAL|1|2|"I have loved you," says the LORD. "But you ask, 'How have you loved us?'"Was not Esau Jacob's brother?" the LORD says. "Yet I have loved Jacob,
MAL|1|3|but Esau I have hated, and I have turned his mountains into a wasteland and left his inheritance to the desert jackals."
MAL|1|4|Edom may say, "Though we have been crushed, we will rebuild the ruins." But this is what the LORD Almighty says: "They may build, but I will demolish. They will be called the Wicked Land, a people always under the wrath of the LORD.
MAL|1|5|You will see it with your own eyes and say, 'Great is the LORD -even beyond the borders of Israel!'
MAL|1|6|"A son honors his father, and a servant his master. If I am a father, where is the honor due me? If I am a master, where is the respect due me?" says the LORD Almighty. "It is you, O priests, who show contempt for my name. "But you ask, 'How have we shown contempt for your name?'
MAL|1|7|"You place defiled food on my altar. "But you ask, 'How have we defiled you?'"By saying that the LORD's table is contemptible.
MAL|1|8|When you bring blind animals for sacrifice, is that not wrong? When you sacrifice crippled or diseased animals, is that not wrong? Try offering them to your governor! Would he be pleased with you? Would he accept you?" says the LORD Almighty.
MAL|1|9|"Now implore God to be gracious to us. With such offerings from your hands, will he accept you?"-says the LORD Almighty.
MAL|1|10|"Oh, that one of you would shut the temple doors, so that you would not light useless fires on my altar! I am not pleased with you," says the LORD Almighty, "and I will accept no offering from your hands.
MAL|1|11|My name will be great among the nations, from the rising to the setting of the sun. In every place incense and pure offerings will be brought to my name, because my name will be great among the nations," says the LORD Almighty.
MAL|1|12|"But you profane it by saying of the Lord's table, 'It is defiled,' and of its food, 'It is contemptible.'
MAL|1|13|And you say, 'What a burden!' and you sniff at it contemptuously," says the LORD Almighty. "When you bring injured, crippled or diseased animals and offer them as sacrifices, should I accept them from your hands?" says the LORD.
MAL|1|14|"Cursed is the cheat who has an acceptable male in his flock and vows to give it, but then sacrifices a blemished animal to the Lord. For I am a great king," says the LORD Almighty, "and my name is to be feared among the nations.
MAL|2|1|"And now this admonition is for you, O priests.
MAL|2|2|If you do not listen, and if you do not set your heart to honor my name," says the LORD Almighty, "I will send a curse upon you, and I will curse your blessings. Yes, I have already cursed them, because you have not set your heart to honor me.
MAL|2|3|"Because of you I will rebuke your descendants; I will spread on your faces the offal from your festival sacrifices, and you will be carried off with it.
MAL|2|4|And you will know that I have sent you this admonition so that my covenant with Levi may continue," says the LORD Almighty.
MAL|2|5|"My covenant was with him, a covenant of life and peace, and I gave them to him; this called for reverence and he revered me and stood in awe of my name.
MAL|2|6|True instruction was in his mouth and nothing false was found on his lips. He walked with me in peace and uprightness, and turned many from sin.
MAL|2|7|"For the lips of a priest ought to preserve knowledge, and from his mouth men should seek instruction-because he is the messenger of the LORD Almighty.
MAL|2|8|But you have turned from the way and by your teaching have caused many to stumble; you have violated the covenant with Levi," says the LORD Almighty.
MAL|2|9|"So I have caused you to be despised and humiliated before all the people, because you have not followed my ways but have shown partiality in matters of the law."
MAL|2|10|Have we not all one Father? Did not one God create us? Why do we profane the covenant of our fathers by breaking faith with one another?
MAL|2|11|Judah has broken faith. A detestable thing has been committed in Israel and in Jerusalem: Judah has desecrated the sanctuary the LORD loves, by marrying the daughter of a foreign god.
MAL|2|12|As for the man who does this, whoever he may be, may the LORD cut him off from the tents of Jacob -even though he brings offerings to the LORD Almighty.
MAL|2|13|Another thing you do: You flood the LORD's altar with tears. You weep and wail because he no longer pays attention to your offerings or accepts them with pleasure from your hands.
MAL|2|14|You ask, "Why?" It is because the LORD is acting as the witness between you and the wife of your youth, because you have broken faith with her, though she is your partner, the wife of your marriage covenant.
MAL|2|15|Has not the LORD made them one? In flesh and spirit they are his. And why one? Because he was seeking godly offspring. So guard yourself in your spirit, and do not break faith with the wife of your youth.
MAL|2|16|"I hate divorce," says the LORD God of Israel, "and I hate a man's covering himself with violence as well as with his garment," says the LORD Almighty. So guard yourself in your spirit, and do not break faith.
MAL|2|17|You have wearied the LORD with your words. "How have we wearied him?" you ask. By saying, "All who do evil are good in the eyes of the LORD, and he is pleased with them" or "Where is the God of justice?"
MAL|3|1|"See, I will send my messenger, who will prepare the way before me. Then suddenly the Lord you are seeking will come to his temple; the messenger of the covenant, whom you desire, will come," says the LORD Almighty.
MAL|3|2|But who can endure the day of his coming? Who can stand when he appears? For he will be like a refiner's fire or a launderer's soap.
MAL|3|3|He will sit as a refiner and purifier of silver; he will purify the Levites and refine them like gold and silver. Then the LORD will have men who will bring offerings in righteousness,
MAL|3|4|and the offerings of Judah and Jerusalem will be acceptable to the LORD, as in days gone by, as in former years.
MAL|3|5|"So I will come near to you for judgment. I will be quick to testify against sorcerers, adulterers and perjurers, against those who defraud laborers of their wages, who oppress the widows and the fatherless, and deprive aliens of justice, but do not fear me," says the LORD Almighty.
MAL|3|6|"I the LORD do not change. So you, O descendants of Jacob, are not destroyed.
MAL|3|7|Ever since the time of your forefathers you have turned away from my decrees and have not kept them. Return to me, and I will return to you," says the LORD Almighty. "But you ask, 'How are we to return?'
MAL|3|8|"Will a man rob God? Yet you rob me. "But you ask, 'How do we rob you?'"In tithes and offerings.
MAL|3|9|You are under a curse-the whole nation of you-because you are robbing me.
MAL|3|10|Bring the whole tithe into the storehouse, that there may be food in my house. Test me in this," says the LORD Almighty, "and see if I will not throw open the floodgates of heaven and pour out so much blessing that you will not have room enough for it.
MAL|3|11|I will prevent pests from devouring your crops, and the vines in your fields will not cast their fruit," says the LORD Almighty.
MAL|3|12|"Then all the nations will call you blessed, for yours will be a delightful land," says the LORD Almighty.
MAL|3|13|"You have said harsh things against me," says the LORD. "Yet you ask, 'What have we said against you?'
MAL|3|14|"You have said, 'It is futile to serve God. What did we gain by carrying out his requirements and going about like mourners before the LORD Almighty?
MAL|3|15|But now we call the arrogant blessed. Certainly the evildoers prosper, and even those who challenge God escape.'"
MAL|3|16|Then those who feared the LORD talked with each other, and the LORD listened and heard. A scroll of remembrance was written in his presence concerning those who feared the LORD and honored his name.
MAL|3|17|"They will be mine," says the LORD Almighty, "in the day when I make up my treasured possession. I will spare them, just as in compassion a man spares his son who serves him.
MAL|3|18|And you will again see the distinction between the righteous and the wicked, between those who serve God and those who do not.
MAL|4|1|"Surely the day is coming; it will burn like a furnace. All the arrogant and every evildoer will be stubble, and that day that is coming will set them on fire," says the LORD Almighty. "Not a root or a branch will be left to them.
MAL|4|2|But for you who revere my name, the sun of righteousness will rise with healing in its wings. And you will go out and leap like calves released from the stall.
MAL|4|3|Then you will trample down the wicked; they will be ashes under the soles of your feet on the day when I do these things," says the LORD Almighty.
MAL|4|4|"Remember the law of my servant Moses, the decrees and laws I gave him at Horeb for all Israel.
MAL|4|5|"See, I will send you the prophet Elijah before that great and dreadful day of the LORD comes.
MAL|4|6|He will turn the hearts of the fathers to their children, and the hearts of the children to their fathers; or else I will come and strike the land with a curse."
