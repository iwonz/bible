GAL|1|1|Павел Апостол, [избранный] не человеками и не через человека, но Иисусом Христом и Богом Отцем, воскресившим Его из мертвых,
GAL|1|2|и все находящиеся со мною братия – церквам Галатийским:
GAL|1|3|благодать вам и мир от Бога Отца и Господа нашего Иисуса Христа,
GAL|1|4|Который отдал Себя Самого за грехи наши, чтобы избавить нас от настоящего лукавого века, по воле Бога и Отца нашего;
GAL|1|5|Ему слава во веки веков. Аминь.
GAL|1|6|Удивляюсь, что вы от призвавшего вас благодатью Христовою так скоро переходите к иному благовествованию,
GAL|1|7|которое [впрочем] не иное, а только есть люди, смущающие вас и желающие превратить благовествование Христово.
GAL|1|8|Но если бы даже мы или Ангел с неба стал благовествовать вам не то, что мы благовествовали вам, да будет анафема.
GAL|1|9|Как прежде мы сказали, [так] и теперь еще говорю: кто благовествует вам не то, что вы приняли, да будет анафема.
GAL|1|10|У людей ли я ныне ищу благоволения, или у Бога? людям ли угождать стараюсь? Если бы я и поныне угождал людям, то не был бы рабом Христовым.
GAL|1|11|Возвещаю вам, братия, что Евангелие, которое я благовествовал, не есть человеческое,
GAL|1|12|ибо и я принял его и научился не от человека, но через откровение Иисуса Христа.
GAL|1|13|Вы слышали о моем прежнем образе жизни в Иудействе, что я жестоко гнал Церковь Божию, и опустошал ее,
GAL|1|14|и преуспевал в Иудействе более многих сверстников в роде моем, будучи неумеренным ревнителем отеческих моих преданий.
GAL|1|15|Когда же Бог, избравший меня от утробы матери моей и призвавший благодатью Своею, благоволил
GAL|1|16|открыть во мне Сына Своего, чтобы я благовествовал Его язычникам, – я не стал тогда же советоваться с плотью и кровью,
GAL|1|17|и не пошел в Иерусалим к предшествовавшим мне Апостолам, а пошел в Аравию, и опять возвратился в Дамаск.
GAL|1|18|Потом, спустя три года, ходил я в Иерусалим видеться с Петром и пробыл у него дней пятнадцать.
GAL|1|19|Другого же из Апостолов я не видел [никого], кроме Иакова, брата Господня.
GAL|1|20|А в том, что пишу вам, пред Богом, не лгу.
GAL|1|21|После сего отошел я в страны Сирии и Киликии.
GAL|1|22|Церквам Христовым в Иудее лично я не был известен,
GAL|1|23|а только слышали они, что гнавший их некогда ныне благовествует веру, которую прежде истреблял, –
GAL|1|24|и прославляли за меня Бога.
GAL|2|1|Потом, через четырнадцать лет, опять ходил я в Иерусалим с Варнавою, взяв с собою и Тита.
GAL|2|2|Ходил же по откровению, и предложил там, и особо знаменитейшим, благовествование, проповедуемое мною язычникам, не напрасно ли я подвизаюсь или подвизался.
GAL|2|3|Но они и Тита, бывшего со мною, хотя и Еллина, не принуждали обрезаться,
GAL|2|4|а вкравшимся лжебратиям, скрытно приходившим подсмотреть за нашею свободою, которую мы имеем во Христе Иисусе, чтобы поработить нас,
GAL|2|5|мы ни на час не уступили и не покорились, дабы истина благовествования сохранилась у вас.
GAL|2|6|И в знаменитых чем–либо, какими бы ни были они когда–либо, для меня нет ничего особенного: Бог не взирает на лице человека. И знаменитые не возложили на меня ничего более.
GAL|2|7|Напротив того, увидев, что мне вверено благовестие для необрезанных, как Петру для обрезанных –
GAL|2|8|ибо Содействовавший Петру в апостольстве у обрезанных содействовал и мне у язычников, –
GAL|2|9|и, узнав о благодати, данной мне, Иаков и Кифа и Иоанн, почитаемые столпами, подали мне и Варнаве руку общения, чтобы нам [идти] к язычникам, а им к обрезанным,
GAL|2|10|только чтобы мы помнили нищих, что и старался я исполнять в точности.
GAL|2|11|Когда же Петр пришел в Антиохию, то я лично противостал ему, потому что он подвергался нареканию.
GAL|2|12|Ибо, до прибытия некоторых от Иакова, ел вместе с язычниками; а когда те пришли, стал таиться и устраняться, опасаясь обрезанных.
GAL|2|13|Вместе с ним лицемерили и прочие Иудеи, так что даже Варнава был увлечен их лицемерием.
GAL|2|14|Но когда я увидел, что они не прямо поступают по истине Евангельской, то сказал Петру при всех: если ты, будучи Иудеем, живешь по–язычески, а не по–иудейски, то для чего язычников принуждаешь жить по–иудейски?
GAL|2|15|Мы по природе Иудеи, а не из язычников грешники;
GAL|2|16|однако же, узнав, что человек оправдывается не делами закона, а только верою в Иисуса Христа, и мы уверовали во Христа Иисуса, чтобы оправдаться верою во Христа, а не делами закона; ибо делами закона не оправдается никакая плоть.
GAL|2|17|Если же, ища оправдания во Христе, мы и сами оказались грешниками, то неужели Христос есть служитель греха? Никак.
GAL|2|18|Ибо если я снова созидаю, что разрушил, то сам себя делаю преступником.
GAL|2|19|Законом я умер для закона, чтобы жить для Бога. Я сораспялся Христу,
GAL|2|20|и уже не я живу, но живет во мне Христос. А что ныне живу во плоти, то живу верою в Сына Божия, возлюбившего меня и предавшего Себя за меня.
GAL|2|21|Не отвергаю благодати Божией; а если законом оправдание, то Христос напрасно умер.
GAL|3|1|О, несмысленные Галаты! кто прельстил вас не покоряться истине, [вас], у которых перед глазами предначертан был Иисус Христос, [как] [бы] у вас распятый?
GAL|3|2|Сие только хочу знать от вас: через дела ли закона вы получили Духа, или через наставление в вере?
GAL|3|3|Так ли вы несмысленны, что, начав духом, теперь оканчиваете плотью?
GAL|3|4|Столь многое потерпели вы неужели без пользы? О, если бы только без пользы!
GAL|3|5|Подающий вам Духа и совершающий между вами чудеса через дела ли закона [сие производит], или через наставление в вере?
GAL|3|6|Так Авраам поверил Богу, и это вменилось ему в праведность.
GAL|3|7|Познайте же, что верующие суть сыны Авраама.
GAL|3|8|И Писание, провидя, что Бог верою оправдает язычников, предвозвестило Аврааму: в тебе благословятся все народы.
GAL|3|9|Итак верующие благословляются с верным Авраамом,
GAL|3|10|а все, утверждающиеся на делах закона, находятся под клятвою. Ибо написано: проклят всяк, кто не исполняет постоянно всего, что написано в книге закона.
GAL|3|11|А что законом никто не оправдывается пред Богом, это ясно, потому что праведный верою жив будет.
GAL|3|12|А закон не по вере; но кто исполняет его, тот жив будет им.
GAL|3|13|Христос искупил нас от клятвы закона, сделавшись за нас клятвою – ибо написано: проклят всяк, висящий на древе, –
GAL|3|14|дабы благословение Авраамово через Христа Иисуса распространилось на язычников, чтобы нам получить обещанного Духа верою.
GAL|3|15|Братия! говорю по [рассуждению] человеческому: даже человеком утвержденного завещания никто не отменяет и не прибавляет [к нему].
GAL|3|16|Но Аврааму даны были обетования и семени его. Не сказано: и потомкам, как бы о многих, но как об одном: и семени твоему, которое есть Христос.
GAL|3|17|Я говорю то, что завета о Христе, прежде Богом утвержденного, закон, явившийся спустя четыреста тридцать лет, не отменяет так, чтобы обетование потеряло силу.
GAL|3|18|Ибо если по закону наследство, то уже не по обетованию; но Аврааму Бог даровал [оное] по обетованию.
GAL|3|19|Для чего же закон? Он дан после по причине преступлений, до времени пришествия семени, к которому [относится] обетование, и преподан через Ангелов, рукою посредника.
GAL|3|20|Но посредник при одном не бывает, а Бог один.
GAL|3|21|Итак закон противен обетованиям Божиим? Никак! Ибо если бы дан был закон, могущий животворить, то подлинно праведность была бы от закона;
GAL|3|22|но Писание всех заключило под грехом, дабы обетование верующим дано было по вере в Иисуса Христа.
GAL|3|23|А до пришествия веры мы заключены были под стражею закона, до того [времени], как надлежало открыться вере.
GAL|3|24|Итак закон был для нас детоводителем ко Христу, дабы нам оправдаться верою;
GAL|3|25|по пришествии же веры, мы уже не под [руководством] детоводителя.
GAL|3|26|Ибо все вы сыны Божии по вере во Христа Иисуса;
GAL|3|27|все вы, во Христа крестившиеся, во Христа облеклись.
GAL|3|28|Нет уже Иудея, ни язычника; нет раба, ни свободного; нет мужеского пола, ни женского: ибо все вы одно во Христе Иисусе.
GAL|3|29|Если же вы Христовы, то вы семя Авраамово и по обетованию наследники.
GAL|4|1|Еще скажу: наследник, доколе в детстве, ничем не отличается от раба, хотя и господин всего:
GAL|4|2|он подчинен попечителям и домоправителям до срока, отцом [назначенного].
GAL|4|3|Так и мы, доколе были в детстве, были порабощены вещественным началам мира;
GAL|4|4|но когда пришла полнота времени, Бог послал Сына Своего (Единородного), Который родился от жены, подчинился закону,
GAL|4|5|чтобы искупить подзаконных, дабы нам получить усыновление.
GAL|4|6|А как вы – сыны, то Бог послал в сердца ваши Духа Сына Своего, вопиющего: "Авва, Отче!"
GAL|4|7|Посему ты уже не раб, но сын; а если сын, то и наследник Божий через Иисуса Христа.
GAL|4|8|Но тогда, не знав Бога, вы служили [богам], которые в существе не боги.
GAL|4|9|Ныне же, познав Бога, или, лучше, получив познание от Бога, для чего возвращаетесь опять к немощным и бедным вещественным началам и хотите еще снова поработить себя им?
GAL|4|10|Наблюдаете дни, месяцы, времена и годы.
GAL|4|11|Боюсь за вас, не напрасно ли я трудился у вас.
GAL|4|12|Прошу вас, братия, будьте, как я, потому что и я, как вы. Вы ничем не обидели меня:
GAL|4|13|знаете, что, [хотя] я в немощи плоти благовествовал вам в первый раз,
GAL|4|14|но вы не презрели искушения моего во плоти моей и не возгнушались [им], а приняли меня, как Ангела Божия, как Христа Иисуса.
GAL|4|15|Как вы были блаженны! Свидетельствую о вас, что, если бы возможно было, вы исторгли бы очи свои и отдали мне.
GAL|4|16|Итак, неужели я сделался врагом вашим, говоря вам истину?
GAL|4|17|Ревнуют по вас нечисто, а хотят вас отлучить, чтобы вы ревновали по них.
GAL|4|18|Хорошо ревновать в добром всегда, а не в моем только присутствии у вас.
GAL|4|19|Дети мои, для которых я снова в муках рождения, доколе не изобразится в вас Христос!
GAL|4|20|Хотел бы я теперь быть у вас и изменить голос мой, потому что я в недоумении о вас.
GAL|4|21|Скажите мне вы, желающие быть под законом: разве вы не слушаете закона?
GAL|4|22|Ибо написано: Авраам имел двух сынов, одного от рабы, а другого от свободной.
GAL|4|23|Но который от рабы, тот рожден по плоти; а который от свободной, тот по обетованию.
GAL|4|24|В этом есть иносказание. Это два завета: один от горы Синайской, рождающий в рабство, который есть Агарь,
GAL|4|25|ибо Агарь означает гору Синай в Аравии и соответствует нынешнему Иерусалиму, потому что он с детьми своими в рабстве;
GAL|4|26|а вышний Иерусалим свободен: он – матерь всем нам.
GAL|4|27|Ибо написано: возвеселись, неплодная, нерождающая; воскликни и возгласи, не мучившаяся родами; потому что у оставленной гораздо более детей, нежели у имеющей мужа.
GAL|4|28|Мы, братия, дети обетования по Исааку.
GAL|4|29|Но, как тогда рожденный по плоти гнал [рожденного] по духу, так и ныне.
GAL|4|30|Что же говорит Писание? Изгони рабу и сына ее, ибо сын рабы не будет наследником вместе с сыном свободной.
GAL|4|31|Итак, братия, мы дети не рабы, но свободной.
GAL|5|1|Итак стойте в свободе, которую даровал нам Христос, и не подвергайтесь опять игу рабства.
GAL|5|2|Вот, я, Павел, говорю вам: если вы обрезываетесь, не будет вам никакой пользы от Христа.
GAL|5|3|Еще свидетельствую всякому человеку обрезывающемуся, что он должен исполнить весь закон.
GAL|5|4|Вы, оправдывающие себя законом, остались без Христа, отпали от благодати,
GAL|5|5|а мы духом ожидаем и надеемся праведности от веры.
GAL|5|6|Ибо во Христе Иисусе не имеет силы ни обрезание, ни необрезание, но вера, действующая любовью.
GAL|5|7|Вы шли хорошо: кто остановил вас, чтобы вы не покорялись истине?
GAL|5|8|Такое убеждение не от Призывающего вас.
GAL|5|9|Малая закваска заквашивает все тесто.
GAL|5|10|Я уверен о вас в Господе, что вы не будете мыслить иначе; а смущающий вас, кто бы он ни был, понесет на себе осуждение.
GAL|5|11|За что же гонят меня, братия, если я и теперь проповедую обрезание? Тогда соблазн креста прекратился бы.
GAL|5|12|О, если бы удалены были возмущающие вас!
GAL|5|13|К свободе призваны вы, братия, только бы свобода ваша не была поводом к [угождению] плоти, но любовью служите друг другу.
GAL|5|14|Ибо весь закон в одном слове заключается: люби ближнего твоего, как самого себя.
GAL|5|15|Если же друг друга угрызаете и съедаете, берегитесь, чтобы вы не были истреблены друг другом.
GAL|5|16|Я говорю: поступайте по духу, и вы не будете исполнять вожделений плоти,
GAL|5|17|ибо плоть желает противного духу, а дух – противного плоти: они друг другу противятся, так что вы не то делаете, что хотели бы.
GAL|5|18|Если же вы духом водитесь, то вы не под законом.
GAL|5|19|Дела плоти известны; они суть: прелюбодеяние, блуд, нечистота, непотребство,
GAL|5|20|идолослужение, волшебство, вражда, ссоры, зависть, гнев, распри, разногласия, (соблазны), ереси,
GAL|5|21|ненависть, убийства, пьянство, бесчинство и тому подобное. Предваряю вас, как и прежде предварял, что поступающие так Царствия Божия не наследуют.
GAL|5|22|Плод же духа: любовь, радость, мир, долготерпение, благость, милосердие, вера,
GAL|5|23|кротость, воздержание. На таковых нет закона.
GAL|5|24|Но те, которые Христовы, распяли плоть со страстями и похотями.
GAL|5|25|Если мы живем духом, то по духу и поступать должны.
GAL|5|26|Не будем тщеславиться, друг друга раздражать, друг другу завидовать.
GAL|6|1|Братия! если и впадет человек в какое согрешение, вы, духовные, исправляйте такового в духе кротости, наблюдая каждый за собою, чтобы не быть искушенным.
GAL|6|2|Носите бремена друг друга, и таким образом исполните закон Христов.
GAL|6|3|Ибо кто почитает себя чем–нибудь, будучи ничто, тот обольщает сам себя.
GAL|6|4|Каждый да испытывает свое дело, и тогда будет иметь похвалу только в себе, а не в другом,
GAL|6|5|ибо каждый понесет свое бремя.
GAL|6|6|Наставляемый словом, делись всяким добром с наставляющим.
GAL|6|7|Не обманывайтесь: Бог поругаем не бывает. Что посеет человек, то и пожнет:
GAL|6|8|сеющий в плоть свою от плоти пожнет тление, а сеющий в дух от духа пожнет жизнь вечную.
GAL|6|9|Делая добро, да не унываем, ибо в свое время пожнем, если не ослабеем.
GAL|6|10|Итак, доколе есть время, будем делать добро всем, а наипаче своим по вере.
GAL|6|11|Видите, как много написал я вам своею рукою.
GAL|6|12|Желающие хвалиться по плоти принуждают вас обрезываться только для того, чтобы не быть гонимыми за крест Христов,
GAL|6|13|ибо и сами обрезывающиеся не соблюдают закона, но хотят, чтобы вы обрезывались, дабы похвалиться в вашей плоти.
GAL|6|14|А я не желаю хвалиться, разве только крестом Господа нашего Иисуса Христа, которым для меня мир распят, и я для мира.
GAL|6|15|Ибо во Христе Иисусе ничего не значит ни обрезание, ни необрезание, а новая тварь.
GAL|6|16|Тем, которые поступают по сему правилу, мир им и милость, и Израилю Божию.
GAL|6|17|Впрочем никто не отягощай меня, ибо я ношу язвы Господа Иисуса на теле моем.
GAL|6|18|Благодать Господа нашего Иисуса Христа со духом вашим, братия. Аминь.
