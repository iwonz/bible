2KGS|1|1|Then Moab rebelled against Israel after the death of Ahab.
2KGS|1|2|And Ahaziah fell down through a lattice in his upper chamber that was in Samaria, and was sick: and he sent messengers, and said unto them, Go, enquire of Baalzebub the god of Ekron whether I shall recover of this disease.
2KGS|1|3|But the angel of the LORD said to Elijah the Tishbite, Arise, go up to meet the messengers of the king of Samaria, and say unto them, Is it not because there is not a God in Israel, that ye go to enquire of Baalzebub the god of Ekron?
2KGS|1|4|Now therefore thus saith the LORD, Thou shalt not come down from that bed on which thou art gone up, but shalt surely die. And Elijah departed.
2KGS|1|5|And when the messengers turned back unto him, he said unto them, Why are ye now turned back?
2KGS|1|6|And they said unto him, There came a man up to meet us, and said unto us, Go, turn again unto the king that sent you, and say unto him, Thus saith the LORD, Is it not because there is not a God in Israel, that thou sendest to enquire of Baalzebub the god of Ekron? therefore thou shalt not come down from that bed on which thou art gone up, but shalt surely die.
2KGS|1|7|And he said unto them, What manner of man was he which came up to meet you, and told you these words?
2KGS|1|8|And they answered him, He was an hairy man, and girt with a girdle of leather about his loins. And he said, It is Elijah the Tishbite.
2KGS|1|9|Then the king sent unto him a captain of fifty with his fifty. And he went up to him: and, behold, he sat on the top of an hill. And he spake unto him, Thou man of God, the king hath said, Come down.
2KGS|1|10|And Elijah answered and said to the captain of fifty, If I be a man of God, then let fire come down from heaven, and consume thee and thy fifty. And there came down fire from heaven, and consumed him and his fifty.
2KGS|1|11|Again also he sent unto him another captain of fifty with his fifty. And he answered and said unto him, O man of God, thus hath the king said, Come down quickly.
2KGS|1|12|And Elijah answered and said unto them, If I be a man of God, let fire come down from heaven, and consume thee and thy fifty. And the fire of God came down from heaven, and consumed him and his fifty.
2KGS|1|13|And he sent again a captain of the third fifty with his fifty. And the third captain of fifty went up, and came and fell on his knees before Elijah, and besought him, and said unto him, O man of God, I pray thee, let my life, and the life of these fifty thy servants, be precious in thy sight.
2KGS|1|14|Behold, there came fire down from heaven, and burnt up the two captains of the former fifties with their fifties: therefore let my life now be precious in thy sight.
2KGS|1|15|And the angel of the LORD said unto Elijah, Go down with him: be not afraid of him. And he arose, and went down with him unto the king.
2KGS|1|16|And he said unto him, Thus saith the LORD, Forasmuch as thou hast sent messengers to enquire of Baalzebub the god of Ekron, is it not because there is no God in Israel to enquire of his word? therefore thou shalt not come down off that bed on which thou art gone up, but shalt surely die.
2KGS|1|17|So he died according to the word of the LORD which Elijah had spoken. And Jehoram reigned in his stead in the second year of Jehoram the son of Jehoshaphat king of Judah; because he had no son.
2KGS|1|18|Now the rest of the acts of Ahaziah which he did, are they not written in the book of the chronicles of the kings of Israel?
2KGS|2|1|And it came to pass, when the LORD would take up Elijah into heaven by a whirlwind, that Elijah went with Elisha from Gilgal.
2KGS|2|2|And Elijah said unto Elisha, Tarry here, I pray thee; for the LORD hath sent me to Bethel. And Elisha said unto him, As the LORD liveth, and as thy soul liveth, I will not leave thee. So they went down to Bethel.
2KGS|2|3|And the sons of the prophets that were at Bethel came forth to Elisha, and said unto him, Knowest thou that the LORD will take away thy master from thy head to day? And he said, Yea, I know it; hold ye your peace.
2KGS|2|4|And Elijah said unto him, Elisha, tarry here, I pray thee; for the LORD hath sent me to Jericho. And he said, As the LORD liveth, and as thy soul liveth, I will not leave thee. So they came to Jericho.
2KGS|2|5|And the sons of the prophets that were at Jericho came to Elisha, and said unto him, Knowest thou that the LORD will take away thy master from thy head to day? And he answered, Yea, I know it; hold ye your peace.
2KGS|2|6|And Elijah said unto him, Tarry, I pray thee, here; for the LORD hath sent me to Jordan. And he said, As the LORD liveth, and as thy soul liveth, I will not leave thee. And they two went on.
2KGS|2|7|And fifty men of the sons of the prophets went, and stood to view afar off: and they two stood by Jordan.
2KGS|2|8|And Elijah took his mantle, and wrapped it together, and smote the waters, and they were divided hither and thither, so that they two went over on dry ground.
2KGS|2|9|And it came to pass, when they were gone over, that Elijah said unto Elisha, Ask what I shall do for thee, before I be taken away from thee. And Elisha said, I pray thee, let a double portion of thy spirit be upon me.
2KGS|2|10|And he said, Thou hast asked a hard thing: nevertheless, if thou see me when I am taken from thee, it shall be so unto thee; but if not, it shall not be so.
2KGS|2|11|And it came to pass, as they still went on, and talked, that, behold, there appeared a chariot of fire, and horses of fire, and parted them both asunder; and Elijah went up by a whirlwind into heaven.
2KGS|2|12|And Elisha saw it, and he cried, My father, my father, the chariot of Israel, and the horsemen thereof. And he saw him no more: and he took hold of his own clothes, and rent them in two pieces.
2KGS|2|13|He took up also the mantle of Elijah that fell from him, and went back, and stood by the bank of Jordan;
2KGS|2|14|And he took the mantle of Elijah that fell from him, and smote the waters, and said, Where is the LORD God of Elijah? and when he also had smitten the waters, they parted hither and thither: and Elisha went over.
2KGS|2|15|And when the sons of the prophets which were to view at Jericho saw him, they said, The spirit of Elijah doth rest on Elisha. And they came to meet him, and bowed themselves to the ground before him.
2KGS|2|16|And they said unto him, Behold now, there be with thy servants fifty strong men; let them go, we pray thee, and seek thy master: lest peradventure the Spirit of the LORD hath taken him up, and cast him upon some mountain, or into some valley. And he said, Ye shall not send.
2KGS|2|17|And when they urged him till he was ashamed, he said, Send. They sent therefore fifty men; and they sought three days, but found him not.
2KGS|2|18|And when they came again to him, (for he tarried at Jericho,) he said unto them, Did I not say unto you, Go not?
2KGS|2|19|And the men of the city said unto Elisha, Behold, I pray thee, the situation of this city is pleasant, as my lord seeth: but the water is naught, and the ground barren.
2KGS|2|20|And he said, Bring me a new cruse, and put salt therein. And they brought it to him.
2KGS|2|21|And he went forth unto the spring of the waters, and cast the salt in there, and said, Thus saith the LORD, I have healed these waters; there shall not be from thence any more death or barren land.
2KGS|2|22|So the waters were healed unto this day, according to the saying of Elisha which he spake.
2KGS|2|23|And he went up from thence unto Bethel: and as he was going up by the way, there came forth little children out of the city, and mocked him, and said unto him, Go up, thou bald head; go up, thou bald head.
2KGS|2|24|And he turned back, and looked on them, and cursed them in the name of the LORD. And there came forth two she bears out of the wood, and tare forty and two children of them.
2KGS|2|25|And he went from thence to mount Carmel, and from thence he returned to Samaria.
2KGS|3|1|Now Jehoram the son of Ahab began to reign over Israel in Samaria the eighteenth year of Jehoshaphat king of Judah, and reigned twelve years.
2KGS|3|2|And he wrought evil in the sight of the LORD; but not like his father, and like his mother: for he put away the image of Baal that his father had made.
2KGS|3|3|Nevertheless he cleaved unto the sins of Jeroboam the son of Nebat, which made Israel to sin; he departed not therefrom.
2KGS|3|4|And Mesha king of Moab was a sheepmaster, and rendered unto the king of Israel an hundred thousand lambs, and an hundred thousand rams, with the wool.
2KGS|3|5|But it came to pass, when Ahab was dead, that the king of Moab rebelled against the king of Israel.
2KGS|3|6|And king Jehoram went out of Samaria the same time, and numbered all Israel.
2KGS|3|7|And he went and sent to Jehoshaphat the king of Judah, saying, The king of Moab hath rebelled against me: wilt thou go with me against Moab to battle? And he said, I will go up: I am as thou art, my people as thy people, and my horses as thy horses.
2KGS|3|8|And he said, Which way shall we go up? And he answered, The way through the wilderness of Edom.
2KGS|3|9|So the king of Israel went, and the king of Judah, and the king of Edom: and they fetched a compass of seven days' journey: and there was no water for the host, and for the cattle that followed them.
2KGS|3|10|And the king of Israel said, Alas! that the LORD hath called these three kings together, to deliver them into the hand of Moab!
2KGS|3|11|But Jehoshaphat said, Is there not here a prophet of the LORD, that we may enquire of the LORD by him? And one of the king of Israel's servants answered and said, Here is Elisha the son of Shaphat, which poured water on the hands of Elijah.
2KGS|3|12|And Jehoshaphat said, The word of the LORD is with him. So the king of Israel and Jehoshaphat and the king of Edom went down to him.
2KGS|3|13|And Elisha said unto the king of Israel, What have I to do with thee? get thee to the prophets of thy father, and to the prophets of thy mother. And the king of Israel said unto him, Nay: for the LORD hath called these three kings together, to deliver them into the hand of Moab.
2KGS|3|14|And Elisha said, As the LORD of hosts liveth, before whom I stand, surely, were it not that I regard the presence of Jehoshaphat the king of Judah, I would not look toward thee, nor see thee.
2KGS|3|15|But now bring me a minstrel. And it came to pass, when the minstrel played, that the hand of the LORD came upon him.
2KGS|3|16|And he said, Thus saith the LORD, Make this valley full of ditches.
2KGS|3|17|For thus saith the LORD, Ye shall not see wind, neither shall ye see rain; yet that valley shall be filled with water, that ye may drink, both ye, and your cattle, and your beasts.
2KGS|3|18|And this is but a light thing in the sight of the LORD: he will deliver the Moabites also into your hand.
2KGS|3|19|And ye shall smite every fenced city, and every choice city, and shall fell every good tree, and stop all wells of water, and mar every good piece of land with stones.
2KGS|3|20|And it came to pass in the morning, when the meat offering was offered, that, behold, there came water by the way of Edom, and the country was filled with water.
2KGS|3|21|And when all the Moabites heard that the kings were come up to fight against them, they gathered all that were able to put on armor, and upward, and stood in the border.
2KGS|3|22|And they rose up early in the morning, and the sun shone upon the water, and the Moabites saw the water on the other side as red as blood:
2KGS|3|23|And they said, This is blood: the kings are surely slain, and they have smitten one another: now therefore, Moab, to the spoil.
2KGS|3|24|And when they came to the camp of Israel, the Israelites rose up and smote the Moabites, so that they fled before them: but they went forward smiting the Moabites, even in their country.
2KGS|3|25|And they beat down the cities, and on every good piece of land cast every man his stone, and filled it; and they stopped all the wells of water, and felled all the good trees: only in Kirharaseth left they the stones thereof; howbeit the slingers went about it, and smote it.
2KGS|3|26|And when the king of Moab saw that the battle was too sore for him, he took with him seven hundred men that drew swords, to break through even unto the king of Edom: but they could not.
2KGS|3|27|Then he took his eldest son that should have reigned in his stead, and offered him for a burnt offering upon the wall. And there was great indignation against Israel: and they departed from him, and returned to their own land.
2KGS|4|1|Now there cried a certain woman of the wives of the sons of the prophets unto Elisha, saying, Thy servant my husband is dead; and thou knowest that thy servant did fear the LORD: and the creditor is come to take unto him my two sons to be bondmen.
2KGS|4|2|And Elisha said unto her, What shall I do for thee? tell me, what hast thou in the house? And she said, Thine handmaid hath not any thing in the house, save a pot of oil.
2KGS|4|3|Then he said, Go, borrow thee vessels abroad of all thy neighbors, even empty vessels; borrow not a few.
2KGS|4|4|And when thou art come in, thou shalt shut the door upon thee and upon thy sons, and shalt pour out into all those vessels, and thou shalt set aside that which is full.
2KGS|4|5|So she went from him, and shut the door upon her and upon her sons, who brought the vessels to her; and she poured out.
2KGS|4|6|And it came to pass, when the vessels were full, that she said unto her son, Bring me yet a vessel. And he said unto her, There is not a vessel more. And the oil stayed.
2KGS|4|7|Then she came and told the man of God. And he said, Go, sell the oil, and pay thy debt, and live thou and thy children of the rest.
2KGS|4|8|And it fell on a day, that Elisha passed to Shunem, where was a great woman; and she constrained him to eat bread. And so it was, that as oft as he passed by, he turned in thither to eat bread.
2KGS|4|9|And she said unto her husband, Behold now, I perceive that this is an holy man of God, which passeth by us continually.
2KGS|4|10|Let us make a little chamber, I pray thee, on the wall; and let us set for him there a bed, and a table, and a stool, and a candlestick: and it shall be, when he cometh to us, that he shall turn in thither.
2KGS|4|11|And it fell on a day, that he came thither, and he turned into the chamber, and lay there.
2KGS|4|12|And he said to Gehazi his servant, Call this Shunammite. And when he had called her, she stood before him.
2KGS|4|13|And he said unto him, Say now unto her, Behold, thou hast been careful for us with all this care; what is to be done for thee? wouldest thou be spoken for to the king, or to the captain of the host? And she answered, I dwell among mine own people.
2KGS|4|14|And he said, What then is to be done for her? And Gehazi answered, Verily she hath no child, and her husband is old.
2KGS|4|15|And he said, Call her. And when he had called her, she stood in the door.
2KGS|4|16|And he said, About this season, according to the time of life, thou shalt embrace a son. And she said, Nay, my lord, thou man of God, do not lie unto thine handmaid.
2KGS|4|17|And the woman conceived, and bare a son at that season that Elisha had said unto her, according to the time of life.
2KGS|4|18|And when the child was grown, it fell on a day, that he went out to his father to the reapers.
2KGS|4|19|And he said unto his father, My head, my head. And he said to a lad, Carry him to his mother.
2KGS|4|20|And when he had taken him, and brought him to his mother, he sat on her knees till noon, and then died.
2KGS|4|21|And she went up, and laid him on the bed of the man of God, and shut the door upon him, and went out.
2KGS|4|22|And she called unto her husband, and said, Send me, I pray thee, one of the young men, and one of the asses, that I may run to the man of God, and come again.
2KGS|4|23|And he said, Wherefore wilt thou go to him to day? it is neither new moon, nor sabbath. And she said, It shall be well.
2KGS|4|24|Then she saddled an ass, and said to her servant, Drive, and go forward; slack not thy riding for me, except I bid thee.
2KGS|4|25|So she went and came unto the man of God to mount Carmel. And it came to pass, when the man of God saw her afar off, that he said to Gehazi his servant, Behold, yonder is that Shunammite:
2KGS|4|26|Run now, I pray thee, to meet her, and say unto her, Is it well with thee? is it well with thy husband? is it well with the child? And she answered, It is well:
2KGS|4|27|And when she came to the man of God to the hill, she caught him by the feet: but Gehazi came near to thrust her away. And the man of God said, Let her alone; for her soul is vexed within her: and the LORD hath hid it from me, and hath not told me.
2KGS|4|28|Then she said, Did I desire a son of my lord? did I not say, Do not deceive me?
2KGS|4|29|Then he said to Gehazi, Gird up thy loins, and take my staff in thine hand, and go thy way: if thou meet any man, salute him not; and if any salute thee, answer him not again: and lay my staff upon the face of the child.
2KGS|4|30|And the mother of the child said, As the LORD liveth, and as thy soul liveth, I will not leave thee. And he arose, and followed her.
2KGS|4|31|And Gehazi passed on before them, and laid the staff upon the face of the child; but there was neither voice, nor hearing. Wherefore he went again to meet him, and told him, saying, The child is not awaked.
2KGS|4|32|And when Elisha was come into the house, behold, the child was dead, and laid upon his bed.
2KGS|4|33|He went in therefore, and shut the door upon them twain, and prayed unto the LORD.
2KGS|4|34|And he went up, and lay upon the child, and put his mouth upon his mouth, and his eyes upon his eyes, and his hands upon his hands: and stretched himself upon the child; and the flesh of the child waxed warm.
2KGS|4|35|Then he returned, and walked in the house to and fro; and went up, and stretched himself upon him: and the child sneezed seven times, and the child opened his eyes.
2KGS|4|36|And he called Gehazi, and said, Call this Shunammite. So he called her. And when she was come in unto him, he said, Take up thy son.
2KGS|4|37|Then she went in, and fell at his feet, and bowed herself to the ground, and took up her son, and went out.
2KGS|4|38|And Elisha came again to Gilgal: and there was a dearth in the land; and the sons of the prophets were sitting before him: and he said unto his servant, Set on the great pot, and seethe pottage for the sons of the prophets.
2KGS|4|39|And one went out into the field to gather herbs, and found a wild vine, and gathered thereof wild gourds his lap full, and came and shred them into the pot of pottage: for they knew them not.
2KGS|4|40|So they poured out for the men to eat. And it came to pass, as they were eating of the pottage, that they cried out, and said, O thou man of God, there is death in the pot. And they could not eat thereof.
2KGS|4|41|But he said, Then bring meal. And he cast it into the pot; and he said, Pour out for the people, that they may eat. And there was no harm in the pot.
2KGS|4|42|And there came a man from Baalshalisha, and brought the man of God bread of the firstfruits, twenty loaves of barley, and full ears of corn in the husk thereof. And he said, Give unto the people, that they may eat.
2KGS|4|43|And his servitor said, What, should I set this before an hundred men? He said again, Give the people, that they may eat: for thus saith the LORD, They shall eat, and shall leave thereof.
2KGS|4|44|So he set it before them, and they did eat, and left thereof, according to the word of the LORD.
2KGS|5|1|Now Naaman, captain of the host of the king of Syria, was a great man with his master, and honorable, because by him the LORD had given deliverance unto Syria: he was also a mighty man in valor, but he was a leper.
2KGS|5|2|And the Syrians had gone out by companies, and had brought away captive out of the land of Israel a little maid; and she waited on Naaman's wife.
2KGS|5|3|And she said unto her mistress, Would God my lord were with the prophet that is in Samaria! for he would recover him of his leprosy.
2KGS|5|4|And one went in, and told his lord, saying, Thus and thus said the maid that is of the land of Israel.
2KGS|5|5|And the king of Syria said, Go to, go, and I will send a letter unto the king of Israel. And he departed, and took with him ten talents of silver, and six thousand pieces of gold, and ten changes of raiment.
2KGS|5|6|And he brought the letter to the king of Israel, saying, Now when this letter is come unto thee, behold, I have therewith sent Naaman my servant to thee, that thou mayest recover him of his leprosy.
2KGS|5|7|And it came to pass, when the king of Israel had read the letter, that he rent his clothes, and said, Am I God, to kill and to make alive, that this man doth send unto me to recover a man of his leprosy? wherefore consider, I pray you, and see how he seeketh a quarrel against me.
2KGS|5|8|And it was so, when Elisha the man of God had heard that the king of Israel had rent his clothes, that he sent to the king, saying, Wherefore hast thou rent thy clothes? let him come now to me, and he shall know that there is a prophet in Israel.
2KGS|5|9|So Naaman came with his horses and with his chariot, and stood at the door of the house of Elisha.
2KGS|5|10|And Elisha sent a messenger unto him, saying, Go and wash in Jordan seven times, and thy flesh shall come again to thee, and thou shalt be clean.
2KGS|5|11|But Naaman was wroth, and went away, and said, Behold, I thought, He will surely come out to me, and stand, and call on the name of the LORD his God, and strike his hand over the place, and recover the leper.
2KGS|5|12|Are not Abana and Pharpar, rivers of Damascus, better than all the waters of Israel? may I not wash in them, and be clean? So he turned and went away in a rage.
2KGS|5|13|And his servants came near, and spake unto him, and said, My father, if the prophet had bid thee do some great thing, wouldest thou not have done it? how much rather then, when he saith to thee, Wash, and be clean?
2KGS|5|14|Then went he down, and dipped himself seven times in Jordan, according to the saying of the man of God: and his flesh came again like unto the flesh of a little child, and he was clean.
2KGS|5|15|And he returned to the man of God, he and all his company, and came, and stood before him: and he said, Behold, now I know that there is no God in all the earth, but in Israel: now therefore, I pray thee, take a blessing of thy servant.
2KGS|5|16|But he said, As the LORD liveth, before whom I stand, I will receive none. And he urged him to take it; but he refused.
2KGS|5|17|And Naaman said, Shall there not then, I pray thee, be given to thy servant two mules' burden of earth? for thy servant will henceforth offer neither burnt offering nor sacrifice unto other gods, but unto the LORD.
2KGS|5|18|In this thing the LORD pardon thy servant, that when my master goeth into the house of Rimmon to worship there, and he leaneth on my hand, and I bow myself in the house of Rimmon: when I bow down myself in the house of Rimmon, the LORD pardon thy servant in this thing.
2KGS|5|19|And he said unto him, Go in peace. So he departed from him a little way.
2KGS|5|20|But Gehazi, the servant of Elisha the man of God, said, Behold, my master hath spared Naaman this Syrian, in not receiving at his hands that which he brought: but, as the LORD liveth, I will run after him, and take somewhat of him.
2KGS|5|21|So Gehazi followed after Naaman. And when Naaman saw him running after him, he lighted down from the chariot to meet him, and said, Is all well?
2KGS|5|22|And he said, All is well. My master hath sent me, saying, Behold, even now there be come to me from mount Ephraim two young men of the sons of the prophets: give them, I pray thee, a talent of silver, and two changes of garments.
2KGS|5|23|And Naaman said, Be content, take two talents. And he urged him, and bound two talents of silver in two bags, with two changes of garments, and laid them upon two of his servants; and they bare them before him.
2KGS|5|24|And when he came to the tower, he took them from their hand, and bestowed them in the house: and he let the men go, and they departed.
2KGS|5|25|But he went in, and stood before his master. And Elisha said unto him, Whence comest thou, Gehazi? And he said, Thy servant went no whither.
2KGS|5|26|And he said unto him, Went not mine heart with thee, when the man turned again from his chariot to meet thee? Is it a time to receive money, and to receive garments, and oliveyards, and vineyards, and sheep, and oxen, and menservants, and maidservants?
2KGS|5|27|The leprosy therefore of Naaman shall cleave unto thee, and unto thy seed for ever. And he went out from his presence a leper as white as snow.
2KGS|6|1|And the sons of the prophets said unto Elisha, Behold now, the place where we dwell with thee is too strait for us.
2KGS|6|2|Let us go, we pray thee, unto Jordan, and take thence every man a beam, and let us make us a place there, where we may dwell. And he answered, Go ye.
2KGS|6|3|And one said, Be content, I pray thee, and go with thy servants. And he answered, I will go.
2KGS|6|4|So he went with them. And when they came to Jordan, they cut down wood.
2KGS|6|5|But as one was felling a beam, the axe head fell into the water: and he cried, and said, Alas, master! for it was borrowed.
2KGS|6|6|And the man of God said, Where fell it? And he showed him the place. And he cut down a stick, and cast it in thither; and the iron did swim.
2KGS|6|7|Therefore said he, Take it up to thee. And he put out his hand, and took it.
2KGS|6|8|Then the king of Syria warred against Israel, and took counsel with his servants, saying, In such and such a place shall be my camp.
2KGS|6|9|And the man of God sent unto the king of Israel, saying, Beware that thou pass not such a place; for thither the Syrians are come down.
2KGS|6|10|And the king of Israel sent to the place which the man of God told him and warned him of, and saved himself there, not once nor twice.
2KGS|6|11|Therefore the heart of the king of Syria was sore troubled for this thing; and he called his servants, and said unto them, Will ye not show me which of us is for the king of Israel?
2KGS|6|12|And one of his servants said, None, my lord, O king: but Elisha, the prophet that is in Israel, telleth the king of Israel the words that thou speakest in thy bedchamber.
2KGS|6|13|And he said, Go and spy where he is, that I may send and fetch him. And it was told him, saying, Behold, he is in Dothan.
2KGS|6|14|Therefore sent he thither horses, and chariots, and a great host: and they came by night, and compassed the city about.
2KGS|6|15|And when the servant of the man of God was risen early, and gone forth, behold, an host compassed the city both with horses and chariots. And his servant said unto him, Alas, my master! how shall we do?
2KGS|6|16|And he answered, Fear not: for they that be with us are more than they that be with them.
2KGS|6|17|And Elisha prayed, and said, LORD, I pray thee, open his eyes, that he may see. And the LORD opened the eyes of the young man; and he saw: and, behold, the mountain was full of horses and chariots of fire round about Elisha.
2KGS|6|18|And when they came down to him, Elisha prayed unto the LORD, and said, Smite this people, I pray thee, with blindness. And he smote them with blindness according to the word of Elisha.
2KGS|6|19|And Elisha said unto them, This is not the way, neither is this the city: follow me, and I will bring you to the man whom ye seek. But he led them to Samaria.
2KGS|6|20|And it came to pass, when they were come into Samaria, that Elisha said, LORD, open the eyes of these men, that they may see. And the LORD opened their eyes, and they saw; and, behold, they were in the midst of Samaria.
2KGS|6|21|And the king of Israel said unto Elisha, when he saw them, My father, shall I smite them? shall I smite them?
2KGS|6|22|And he answered, Thou shalt not smite them: wouldest thou smite those whom thou hast taken captive with thy sword and with thy bow? set bread and water before them, that they may eat and drink, and go to their master.
2KGS|6|23|And he prepared great provision for them: and when they had eaten and drunk, he sent them away, and they went to their master. So the bands of Syria came no more into the land of Israel.
2KGS|6|24|And it came to pass after this, that Benhadad king of Syria gathered all his host, and went up, and besieged Samaria.
2KGS|6|25|And there was a great famine in Samaria: and, behold, they besieged it, until an ass's head was sold for fourscore pieces of silver, and the fourth part of a cab of dove's dung for five pieces of silver.
2KGS|6|26|And as the king of Israel was passing by upon the wall, there cried a woman unto him, saying, Help, my lord, O king.
2KGS|6|27|And he said, If the LORD do not help thee, whence shall I help thee? out of the barnfloor, or out of the winepress?
2KGS|6|28|And the king said unto her, What aileth thee? And she answered, This woman said unto me, Give thy son, that we may eat him to day, and we will eat my son to morrow.
2KGS|6|29|So we boiled my son, and did eat him: and I said unto her on the next day, Give thy son, that we may eat him: and she hath hid her son.
2KGS|6|30|And it came to pass, when the king heard the words of the woman, that he rent his clothes; and he passed by upon the wall, and the people looked, and, behold, he had sackcloth within upon his flesh.
2KGS|6|31|Then he said, God do so and more also to me, if the head of Elisha the son of Shaphat shall stand on him this day.
2KGS|6|32|But Elisha sat in his house, and the elders sat with him; and the king sent a man from before him: but ere the messenger came to him, he said to the elders, See ye how this son of a murderer hath sent to take away mine head? look, when the messenger cometh, shut the door, and hold him fast at the door: is not the sound of his master's feet behind him?
2KGS|6|33|And while he yet talked with them, behold, the messenger came down unto him: and he said, Behold, this evil is of the LORD; what should I wait for the LORD any longer?
2KGS|7|1|Then Elisha said, Hear ye the word of the LORD; Thus saith the LORD, To morrow about this time shall a measure of fine flour be sold for a shekel, and two measures of barley for a shekel, in the gate of Samaria.
2KGS|7|2|Then a lord on whose hand the king leaned answered the man of God, and said, Behold, if the LORD would make windows in heaven, might this thing be? And he said, Behold, thou shalt see it with thine eyes, but shalt not eat thereof.
2KGS|7|3|And there were four leprous men at the entering in of the gate: and they said one to another, Why sit we here until we die?
2KGS|7|4|If we say, We will enter into the city, then the famine is in the city, and we shall die there: and if we sit still here, we die also. Now therefore come, and let us fall unto the host of the Syrians: if they save us alive, we shall live; and if they kill us, we shall but die.
2KGS|7|5|And they rose up in the twilight, to go unto the camp of the Syrians: and when they were come to the uttermost part of the camp of Syria, behold, there was no man there.
2KGS|7|6|For the LORD had made the host of the Syrians to hear a noise of chariots, and a noise of horses, even the noise of a great host: and they said one to another, Lo, the king of Israel hath hired against us the kings of the Hittites, and the kings of the Egyptians, to come upon us.
2KGS|7|7|Wherefore they arose and fled in the twilight, and left their tents, and their horses, and their asses, even the camp as it was, and fled for their life.
2KGS|7|8|And when these lepers came to the uttermost part of the camp, they went into one tent, and did eat and drink, and carried thence silver, and gold, and raiment, and went and hid it; and came again, and entered into another tent, and carried thence also, and went and hid it.
2KGS|7|9|Then they said one to another, We do not well: this day is a day of good tidings, and we hold our peace: if we tarry till the morning light, some mischief will come upon us: now therefore come, that we may go and tell the king's household.
2KGS|7|10|So they came and called unto the porter of the city: and they told them, saying, We came to the camp of the Syrians, and, behold, there was no man there, neither voice of man, but horses tied, and asses tied, and the tents as they were.
2KGS|7|11|And he called the porters; and they told it to the king's house within.
2KGS|7|12|And the king arose in the night, and said unto his servants, I will now show you what the Syrians have done to us. They know that we be hungry; therefore are they gone out of the camp to hide themselves in the field, saying, When they come out of the city, we shall catch them alive, and get into the city.
2KGS|7|13|And one of his servants answered and said, Let some take, I pray thee, five of the horses that remain, which are left in the city, (behold, they are as all the multitude of Israel that are left in it: behold, I say, they are even as all the multitude of the Israelites that are consumed:) and let us send and see.
2KGS|7|14|They took therefore two chariot horses; and the king sent after the host of the Syrians, saying, Go and see.
2KGS|7|15|And they went after them unto Jordan: and, lo, all the way was full of garments and vessels, which the Syrians had cast away in their haste. And the messengers returned, and told the king.
2KGS|7|16|And the people went out, and spoiled the tents of the Syrians. So a measure of fine flour was sold for a shekel, and two measures of barley for a shekel, according to the word of the LORD.
2KGS|7|17|And the king appointed the lord on whose hand he leaned to have the charge of the gate: and the people trode upon him in the gate, and he died, as the man of God had said, who spake when the king came down to him.
2KGS|7|18|And it came to pass as the man of God had spoken to the king, saying, Two measures of barley for a shekel, and a measure of fine flour for a shekel, shall be to morrow about this time in the gate of Samaria:
2KGS|7|19|And that lord answered the man of God, and said, Now, behold, if the LORD should make windows in heaven, might such a thing be? And he said, Behold, thou shalt see it with thine eyes, but shalt not eat thereof.
2KGS|7|20|And so it fell out unto him: for the people trode upon him in the gate, and he died.
2KGS|8|1|Then spake Elisha unto the woman, whose son he had restored to life, saying, Arise, and go thou and thine household, and sojourn wheresoever thou canst sojourn: for the LORD hath called for a famine; and it shall also come upon the land seven years.
2KGS|8|2|And the woman arose, and did after the saying of the man of God: and she went with her household, and sojourned in the land of the Philistines seven years.
2KGS|8|3|And it came to pass at the seven years' end, that the woman returned out of the land of the Philistines: and she went forth to cry unto the king for her house and for her land.
2KGS|8|4|And the king talked with Gehazi the servant of the man of God, saying, Tell me, I pray thee, all the great things that Elisha hath done.
2KGS|8|5|And it came to pass, as he was telling the king how he had restored a dead body to life, that, behold, the woman, whose son he had restored to life, cried to the king for her house and for her land. And Gehazi said, My lord, O king, this is the woman, and this is her son, whom Elisha restored to life.
2KGS|8|6|And when the king asked the woman, she told him. So the king appointed unto her a certain officer, saying, Restore all that was hers, and all the fruits of the field since the day that she left the land, even until now.
2KGS|8|7|And Elisha came to Damascus; and Benhadad the king of Syria was sick; and it was told him, saying, The man of God is come hither.
2KGS|8|8|And the king said unto Hazael, Take a present in thine hand, and go, meet the man of God, and enquire of the LORD by him, saying, Shall I recover of this disease?
2KGS|8|9|So Hazael went to meet him, and took a present with him, even of every good thing of Damascus, forty camels' burden, and came and stood before him, and said, Thy son Benhadad king of Syria hath sent me to thee, saying, Shall I recover of this disease?
2KGS|8|10|And Elisha said unto him, Go, say unto him, Thou mayest certainly recover: howbeit the LORD hath showed me that he shall surely die.
2KGS|8|11|And he settled his countenance stedfastly, until he was ashamed: and the man of God wept.
2KGS|8|12|And Hazael said, Why weepeth my lord? And he answered, Because I know the evil that thou wilt do unto the children of Israel: their strong holds wilt thou set on fire, and their young men wilt thou slay with the sword, and wilt dash their children, and rip up their women with child.
2KGS|8|13|And Hazael said, But what, is thy servant a dog, that he should do this great thing? And Elisha answered, The LORD hath showed me that thou shalt be king over Syria.
2KGS|8|14|So he departed from Elisha, and came to his master; who said to him, What said Elisha to thee? And he answered, He told me that thou shouldest surely recover.
2KGS|8|15|And it came to pass on the morrow, that he took a thick cloth, and dipped it in water, and spread it on his face, so that he died: and Hazael reigned in his stead.
2KGS|8|16|And in the fifth year of Joram the son of Ahab king of Israel, Jehoshaphat being then king of Judah, Jehoram the son of Jehoshaphat king of Judah began to reign.
2KGS|8|17|Thirty and two years old was he when he began to reign; and he reigned eight years in Jerusalem.
2KGS|8|18|And he walked in the way of the kings of Israel, as did the house of Ahab: for the daughter of Ahab was his wife: and he did evil in the sight of the LORD.
2KGS|8|19|Yet the LORD would not destroy Judah for David his servant's sake, as he promised him to give him alway a light, and to his children.
2KGS|8|20|In his days Edom revolted from under the hand of Judah, and made a king over themselves.
2KGS|8|21|So Joram went over to Zair, and all the chariots with him: and he rose by night, and smote the Edomites which compassed him about, and the captains of the chariots: and the people fled into their tents.
2KGS|8|22|Yet Edom revolted from under the hand of Judah unto this day. Then Libnah revolted at the same time.
2KGS|8|23|And the rest of the acts of Joram, and all that he did, are they not written in the book of the chronicles of the kings of Judah?
2KGS|8|24|And Joram slept with his fathers, and was buried with his fathers in the city of David: and Ahaziah his son reigned in his stead.
2KGS|8|25|In the twelfth year of Joram the son of Ahab king of Israel did Ahaziah the son of Jehoram king of Judah begin to reign.
2KGS|8|26|Two and twenty years old was Ahaziah when he began to reign; and he reigned one year in Jerusalem. And his mother's name was Athaliah, the daughter of Omri king of Israel.
2KGS|8|27|And he walked in the way of the house of Ahab, and did evil in the sight of the LORD, as did the house of Ahab: for he was the son in law of the house of Ahab.
2KGS|8|28|And he went with Joram the son of Ahab to the war against Hazael king of Syria in Ramothgilead; and the Syrians wounded Joram.
2KGS|8|29|And king Joram went back to be healed in Jezreel of the wounds which the Syrians had given him at Ramah, when he fought against Hazael king of Syria. And Ahaziah the son of Jehoram king of Judah went down to see Joram the son of Ahab in Jezreel, because he was sick.
2KGS|9|1|And Elisha the prophet called one of the children of the prophets, and said unto him, Gird up thy loins, and take this box of oil in thine hand, and go to Ramothgilead:
2KGS|9|2|And when thou comest thither, look out there Jehu the son of Jehoshaphat the son of Nimshi, and go in, and make him arise up from among his brethren, and carry him to an inner chamber;
2KGS|9|3|Then take the box of oil, and pour it on his head, and say, Thus saith the LORD, I have anointed thee king over Israel. Then open the door, and flee, and tarry not.
2KGS|9|4|So the young man, even the young man the prophet, went to Ramothgilead.
2KGS|9|5|And when he came, behold, the captains of the host were sitting; and he said, I have an errand to thee, O captain. And Jehu said, Unto which of all us? And he said, To thee, O captain.
2KGS|9|6|And he arose, and went into the house; and he poured the oil on his head, and said unto him, Thus saith the LORD God of Israel, I have anointed thee king over the people of the LORD, even over Israel.
2KGS|9|7|And thou shalt smite the house of Ahab thy master, that I may avenge the blood of my servants the prophets, and the blood of all the servants of the LORD, at the hand of Jezebel.
2KGS|9|8|For the whole house of Ahab shall perish: and I will cut off from Ahab him that pisseth against the wall, and him that is shut up and left in Israel:
2KGS|9|9|And I will make the house of Ahab like the house of Jeroboam the son of Nebat, and like the house of Baasha the son of Ahijah:
2KGS|9|10|And the dogs shall eat Jezebel in the portion of Jezreel, and there shall be none to bury her. And he opened the door, and fled.
2KGS|9|11|Then Jehu came forth to the servants of his lord: and one said unto him, Is all well? wherefore came this mad fellow to thee? And he said unto them, Ye know the man, and his communication.
2KGS|9|12|And they said, It is false; tell us now. And he said, Thus and thus spake he to me, saying, Thus saith the LORD, I have anointed thee king over Israel.
2KGS|9|13|Then they hasted, and took every man his garment, and put it under him on the top of the stairs, and blew with trumpets, saying, Jehu is king.
2KGS|9|14|So Jehu the son of Jehoshaphat the son of Nimshi conspired against Joram. (Now Joram had kept Ramothgilead, he and all Israel, because of Hazael king of Syria.
2KGS|9|15|But king Joram was returned to be healed in Jezreel of the wounds which the Syrians had given him, when he fought with Hazael king of Syria.) And Jehu said, If it be your minds, then let none go forth nor escape out of the city to go to tell it in Jezreel.
2KGS|9|16|So Jehu rode in a chariot, and went to Jezreel; for Joram lay there. And Ahaziah king of Judah was come down to see Joram.
2KGS|9|17|And there stood a watchman on the tower in Jezreel, and he spied the company of Jehu as he came, and said, I see a company. And Joram said, Take an horseman, and send to meet them, and let him say, Is it peace?
2KGS|9|18|So there went one on horseback to meet him, and said, Thus saith the king, Is it peace? And Jehu said, What hast thou to do with peace? turn thee behind me. And the watchman told, saying, The messenger came to them, but he cometh not again.
2KGS|9|19|Then he sent out a second on horseback, which came to them, and said, Thus saith the king, Is it peace? And Jehu answered, What hast thou to do with peace? turn thee behind me.
2KGS|9|20|And the watchman told, saying, He came even unto them, and cometh not again: and the driving is like the driving of Jehu the son of Nimshi; for he driveth furiously.
2KGS|9|21|And Joram said, Make ready. And his chariot was made ready. And Joram king of Israel and Ahaziah king of Judah went out, each in his chariot, and they went out against Jehu, and met him in the portion of Naboth the Jezreelite.
2KGS|9|22|And it came to pass, when Joram saw Jehu, that he said, Is it peace, Jehu? And he answered, What peace, so long as the whoredoms of thy mother Jezebel and her witchcrafts are so many?
2KGS|9|23|And Joram turned his hands, and fled, and said to Ahaziah, There is treachery, O Ahaziah.
2KGS|9|24|And Jehu drew a bow with his full strength, and smote Jehoram between his arms, and the arrow went out at his heart, and he sunk down in his chariot.
2KGS|9|25|Then said Jehu to Bidkar his captain, Take up, and cast him in the portion of the field of Naboth the Jezreelite: for remember how that, when I and thou rode together after Ahab his father, the LORD laid this burden upon him;
2KGS|9|26|Surely I have seen yesterday the blood of Naboth, and the blood of his sons, saith the LORD; and I will requite thee in this plat, saith the LORD. Now therefore take and cast him into the plat of ground, according to the word of the LORD.
2KGS|9|27|But when Ahaziah the king of Judah saw this, he fled by the way of the garden house. And Jehu followed after him, and said, Smite him also in the chariot. And they did so at the going up to Gur, which is by Ibleam. And he fled to Megiddo, and died there.
2KGS|9|28|And his servants carried him in a chariot to Jerusalem, and buried him in his sepulchre with his fathers in the city of David.
2KGS|9|29|And in the eleventh year of Joram the son of Ahab began Ahaziah to reign over Judah.
2KGS|9|30|And when Jehu was come to Jezreel, Jezebel heard of it; and she painted her face, and tired her head, and looked out at a window.
2KGS|9|31|And as Jehu entered in at the gate, she said, Had Zimri peace, who slew his master?
2KGS|9|32|And he lifted up his face to the window, and said, Who is on my side? who? And there looked out to him two or three eunuchs.
2KGS|9|33|And he said, Throw her down. So they threw her down: and some of her blood was sprinkled on the wall, and on the horses: and he trode her under foot.
2KGS|9|34|And when he was come in, he did eat and drink, and said, Go, see now this cursed woman, and bury her: for she is a king's daughter.
2KGS|9|35|And they went to bury her: but they found no more of her than the skull, and the feet, and the palms of her hands.
2KGS|9|36|Wherefore they came again, and told him. And he said, This is the word of the LORD, which he spake by his servant Elijah the Tishbite, saying, In the portion of Jezreel shall dogs eat the flesh of Jezebel:
2KGS|9|37|And the carcass of Jezebel shall be as dung upon the face of the field in the portion of Jezreel; so that they shall not say, This is Jezebel.
2KGS|10|1|And Ahab had seventy sons in Samaria. And Jehu wrote letters, and sent to Samaria, unto the rulers of Jezreel, to the elders, and to them that brought up Ahab's children, saying,
2KGS|10|2|Now as soon as this letter cometh to you, seeing your master's sons are with you, and there are with you chariots and horses, a fenced city also, and armor;
2KGS|10|3|Look even out the best and meetest of your master's sons, and set him on his father's throne, and fight for your master's house.
2KGS|10|4|But they were exceedingly afraid, and said, Behold, two kings stood not before him: how then shall we stand?
2KGS|10|5|And he that was over the house, and he that was over the city, the elders also, and the bringers up of the children, sent to Jehu, saying, We are thy servants, and will do all that thou shalt bid us; we will not make any king: do thou that which is good in thine eyes.
2KGS|10|6|Then he wrote a letter the second time to them, saying, If ye be mine, and if ye will hearken unto my voice, take ye the heads of the men your master's sons, and come to me to Jezreel by to morrow this time. Now the king's sons, being seventy persons, were with the great men of the city, which brought them up.
2KGS|10|7|And it came to pass, when the letter came to them, that they took the king's sons, and slew seventy persons, and put their heads in baskets, and sent him them to Jezreel.
2KGS|10|8|And there came a messenger, and told him, saying, They have brought the heads of the king's sons. And he said, Lay ye them in two heaps at the entering in of the gate until the morning.
2KGS|10|9|And it came to pass in the morning, that he went out, and stood, and said to all the people, Ye be righteous: behold, I conspired against my master, and slew him: but who slew all these?
2KGS|10|10|Know now that there shall fall unto the earth nothing of the word of the LORD, which the LORD spake concerning the house of Ahab: for the LORD hath done that which he spake by his servant Elijah.
2KGS|10|11|So Jehu slew all that remained of the house of Ahab in Jezreel, and all his great men, and his kinsfolk, and his priests, until he left him none remaining.
2KGS|10|12|And he arose and departed, and came to Samaria. And as he was at the shearing house in the way,
2KGS|10|13|Jehu met with the brethren of Ahaziah king of Judah, and said, Who are ye? And they answered, We are the brethren of Ahaziah; and we go down to salute the children of the king and the children of the queen.
2KGS|10|14|And he said, Take them alive. And they took them alive, and slew them at the pit of the shearing house, even two and forty men; neither left he any of them.
2KGS|10|15|And when he was departed thence, he lighted on Jehonadab the son of Rechab coming to meet him: and he saluted him, and said to him, Is thine heart right, as my heart is with thy heart? And Jehonadab answered, It is. If it be, give me thine hand. And he gave him his hand; and he took him up to him into the chariot.
2KGS|10|16|And he said, Come with me, and see my zeal for the LORD. So they made him ride in his chariot.
2KGS|10|17|And when he came to Samaria, he slew all that remained unto Ahab in Samaria, till he had destroyed him, according to the saying of the LORD, which he spake to Elijah.
2KGS|10|18|And Jehu gathered all the people together, and said unto them, Ahab served Baal a little; but Jehu shall serve him much.
2KGS|10|19|Now therefore call unto me all the prophets of Baal, all his servants, and all his priests; let none be wanting: for I have a great sacrifice to do to Baal; whosoever shall be wanting, he shall not live. But Jehu did it in subtilty, to the intent that he might destroy the worshippers of Baal.
2KGS|10|20|And Jehu said, Proclaim a solemn assembly for Baal. And they proclaimed it.
2KGS|10|21|And Jehu sent through all Israel: and all the worshippers of Baal came, so that there was not a man left that came not. And they came into the house of Baal; and the house of Baal was full from one end to another.
2KGS|10|22|And he said unto him that was over the vestry, Bring forth vestments for all the worshippers of Baal. And he brought them forth vestments.
2KGS|10|23|And Jehu went, and Jehonadab the son of Rechab, into the house of Baal, and said unto the worshippers of Baal, Search, and look that there be here with you none of the servants of the LORD, but the worshippers of Baal only.
2KGS|10|24|And when they went in to offer sacrifices and burnt offerings, Jehu appointed fourscore men without, and said, If any of the men whom I have brought into your hands escape, he that letteth him go, his life shall be for the life of him.
2KGS|10|25|And it came to pass, as soon as he had made an end of offering the burnt offering, that Jehu said to the guard and to the captains, Go in, and slay them; let none come forth. And they smote them with the edge of the sword; and the guard and the captains cast them out, and went to the city of the house of Baal.
2KGS|10|26|And they brought forth the images out of the house of Baal, and burned them.
2KGS|10|27|And they brake down the image of Baal, and brake down the house of Baal, and made it a draught house unto this day.
2KGS|10|28|Thus Jehu destroyed Baal out of Israel.
2KGS|10|29|Howbeit from the sins of Jeroboam the son of Nebat, who made Israel to sin, Jehu departed not from after them, to wit, the golden calves that were in Bethel, and that were in Dan.
2KGS|10|30|And the LORD said unto Jehu, Because thou hast done well in executing that which is right in mine eyes, and hast done unto the house of Ahab according to all that was in mine heart, thy children of the fourth generation shall sit on the throne of Israel.
2KGS|10|31|But Jehu took no heed to walk in the law of the LORD God of Israel with all his heart: for he departed not from the sins of Jeroboam, which made Israel to sin.
2KGS|10|32|In those days the LORD began to cut Israel short: and Hazael smote them in all the coasts of Israel;
2KGS|10|33|From Jordan eastward, all the land of Gilead, the Gadites, and the Reubenites, and the Manassites, from Aroer, which is by the river Arnon, even Gilead and Bashan.
2KGS|10|34|Now the rest of the acts of Jehu, and all that he did, and all his might, are they not written in the book of the chronicles of the kings of Israel?
2KGS|10|35|And Jehu slept with his fathers: and they buried him in Samaria. And Jehoahaz his son reigned in his stead.
2KGS|10|36|And the time that Jehu reigned over Israel in Samaria was twenty and eight years.
2KGS|11|1|And when Athaliah the mother of Ahaziah saw that her son was dead, she arose and destroyed all the seed royal.
2KGS|11|2|But Jehosheba, the daughter of king Joram, sister of Ahaziah, took Joash the son of Ahaziah, and stole him from among the king's sons which were slain; and they hid him, even him and his nurse, in the bedchamber from Athaliah, so that he was not slain.
2KGS|11|3|And he was with her hid in the house of the LORD six years. And Athaliah did reign over the land.
2KGS|11|4|And the seventh year Jehoiada sent and fetched the rulers over hundreds, with the captains and the guard, and brought them to him into the house of the LORD, and made a covenant with them, and took an oath of them in the house of the LORD, and showed them the king's son.
2KGS|11|5|And he commanded them, saying, This is the thing that ye shall do; A third part of you that enter in on the sabbath shall even be keepers of the watch of the king's house;
2KGS|11|6|And a third part shall be at the gate of Sur; and a third part at the gate behind the guard: so shall ye keep the watch of the house, that it be not broken down.
2KGS|11|7|And two parts of all you that go forth on the sabbath, even they shall keep the watch of the house of the LORD about the king.
2KGS|11|8|And ye shall compass the king round about, every man with his weapons in his hand: and he that cometh within the ranges, let him be slain: and be ye with the king as he goeth out and as he cometh in.
2KGS|11|9|And the captains over the hundreds did according to all things that Jehoiada the priest commanded: and they took every man his men that were to come in on the sabbath, with them that should go out on the sabbath, and came to Jehoiada the priest.
2KGS|11|10|And to the captains over hundreds did the priest give king David's spears and shields, that were in the temple of the LORD.
2KGS|11|11|And the guard stood, every man with his weapons in his hand, round about the king, from the right corner of the temple to the left corner of the temple, along by the altar and the temple.
2KGS|11|12|And he brought forth the king's son, and put the crown upon him, and gave him the testimony; and they made him king, and anointed him; and they clapped their hands, and said, God save the king.
2KGS|11|13|And when Athaliah heard the noise of the guard and of the people, she came to the people into the temple of the LORD.
2KGS|11|14|And when she looked, behold, the king stood by a pillar, as the manner was, and the princes and the trumpeters by the king, and all the people of the land rejoiced, and blew with trumpets: and Athaliah rent her clothes, and cried, Treason, Treason.
2KGS|11|15|But Jehoiada the priest commanded the captains of the hundreds, the officers of the host, and said unto them, Have her forth without the ranges: and him that followeth her kill with the sword. For the priest had said, Let her not be slain in the house of the LORD.
2KGS|11|16|And they laid hands on her; and she went by the way by the which the horses came into the king's house: and there was she slain.
2KGS|11|17|And Jehoiada made a covenant between the LORD and the king and the people, that they should be the LORD's people; between the king also and the people.
2KGS|11|18|And all the people of the land went into the house of Baal, and brake it down; his altars and his images brake they in pieces thoroughly, and slew Mattan the priest of Baal before the altars. And the priest appointed officers over the house of the LORD.
2KGS|11|19|And he took the rulers over hundreds, and the captains, and the guard, and all the people of the land; and they brought down the king from the house of the LORD, and came by the way of the gate of the guard to the king's house. And he sat on the throne of the kings.
2KGS|11|20|And all the people of the land rejoiced, and the city was in quiet: and they slew Athaliah with the sword beside the king's house.
2KGS|11|21|Seven years old was Jehoash when he began to reign.
2KGS|12|1|In the seventh year of Jehu Jehoash began to reign; and forty years reigned he in Jerusalem. And his mother's name was Zibiah of Beersheba.
2KGS|12|2|And Jehoash did that which was right in the sight of the LORD all his days wherein Jehoiada the priest instructed him.
2KGS|12|3|But the high places were not taken away: the people still sacrificed and burnt incense in the high places.
2KGS|12|4|And Jehoash said to the priests, All the money of the dedicated things that is brought into the house of the LORD, even the money of every one that passeth the account, the money that every man is set at, and all the money that cometh into any man's heart to bring into the house of the LORD,
2KGS|12|5|Let the priests take it to them, every man of his acquaintance: and let them repair the breaches of the house, wheresoever any breach shall be found.
2KGS|12|6|But it was so, that in the three and twentieth year of king Jehoash the priests had not repaired the breaches of the house.
2KGS|12|7|Then king Jehoash called for Jehoiada the priest, and the other priests, and said unto them, Why repair ye not the breaches of the house? now therefore receive no more money of your acquaintance, but deliver it for the breaches of the house.
2KGS|12|8|And the priests consented to receive no more money of the people, neither to repair the breaches of the house.
2KGS|12|9|But Jehoiada the priest took a chest, and bored a hole in the lid of it, and set it beside the altar, on the right side as one cometh into the house of the LORD: and the priests that kept the door put therein all the money that was brought into the house of the LORD.
2KGS|12|10|And it was so, when they saw that there was much money in the chest, that the king's scribe and the high priest came up, and they put up in bags, and told the money that was found in the house of the LORD.
2KGS|12|11|And they gave the money, being told, into the hands of them that did the work, that had the oversight of the house of the LORD: and they laid it out to the carpenters and builders, that wrought upon the house of the LORD,
2KGS|12|12|And to masons, and hewers of stone, and to buy timber and hewed stone to repair the breaches of the house of the LORD, and for all that was laid out for the house to repair it.
2KGS|12|13|Howbeit there were not made for the house of the LORD bowls of silver, snuffers, basins, trumpets, any vessels of gold, or vessels of silver, of the money that was brought into the house of the LORD:
2KGS|12|14|But they gave that to the workmen, and repaired therewith the house of the LORD.
2KGS|12|15|Moreover they reckoned not with the men, into whose hand they delivered the money to be bestowed on workmen: for they dealt faithfully.
2KGS|12|16|The trespass money and sin money was not brought into the house of the LORD: it was the priests'.
2KGS|12|17|Then Hazael king of Syria went up, and fought against Gath, and took it: and Hazael set his face to go up to Jerusalem.
2KGS|12|18|And Jehoash king of Judah took all the hallowed things that Jehoshaphat, and Jehoram, and Ahaziah, his fathers, kings of Judah, had dedicated, and his own hallowed things, and all the gold that was found in the treasures of the house of the LORD, and in the king's house, and sent it to Hazael king of Syria: and he went away from Jerusalem.
2KGS|12|19|And the rest of the acts of Joash, and all that he did, are they not written in the book of the chronicles of the kings of Judah?
2KGS|12|20|And his servants arose, and made a conspiracy, and slew Joash in the house of Millo, which goeth down to Silla.
2KGS|12|21|For Jozachar the son of Shimeath, and Jehozabad the son of Shomer, his servants, smote him, and he died; and they buried him with his fathers in the city of David: and Amaziah his son reigned in his stead.
2KGS|13|1|In the three and twentieth year of Joash the son of Ahaziah king of Judah Jehoahaz the son of Jehu began to reign over Israel in Samaria, and reigned seventeen years.
2KGS|13|2|And he did that which was evil in the sight of the LORD, and followed the sins of Jeroboam the son of Nebat, which made Israel to sin; he departed not therefrom.
2KGS|13|3|And the anger of the LORD was kindled against Israel, and he delivered them into the hand of Hazael king of Syria, and into the hand of Benhadad the son of Hazael, all their days.
2KGS|13|4|And Jehoahaz besought the LORD, and the LORD hearkened unto him: for he saw the oppression of Israel, because the king of Syria oppressed them.
2KGS|13|5|(And the LORD gave Israel a saviour, so that they went out from under the hand of the Syrians: and the children of Israel dwelt in their tents, as beforetime.
2KGS|13|6|Nevertheless they departed not from the sins of the house of Jeroboam, who made Israel sin, but walked therein: and there remained the grove also in Samaria.)
2KGS|13|7|Neither did he leave of the people to Jehoahaz but fifty horsemen, and ten chariots, and ten thousand footmen; for the king of Syria had destroyed them, and had made them like the dust by threshing.
2KGS|13|8|Now the rest of the acts of Jehoahaz, and all that he did, and his might, are they not written in the book of the chronicles of the kings of Israel?
2KGS|13|9|And Jehoahaz slept with his fathers; and they buried him in Samaria: and Joash his son reigned in his stead.
2KGS|13|10|In the thirty and seventh year of Joash king of Judah began Jehoash the son of Jehoahaz to reign over Israel in Samaria, and reigned sixteen years.
2KGS|13|11|And he did that which was evil in the sight of the LORD; he departed not from all the sins of Jeroboam the son of Nebat, who made Israel sin: but he walked therein.
2KGS|13|12|And the rest of the acts of Joash, and all that he did, and his might wherewith he fought against Amaziah king of Judah, are they not written in the book of the chronicles of the kings of Israel?
2KGS|13|13|And Joash slept with his fathers; and Jeroboam sat upon his throne: and Joash was buried in Samaria with the kings of Israel.
2KGS|13|14|Now Elisha was fallen sick of his sickness whereof he died. And Joash the king of Israel came down unto him, and wept over his face, and said, O my father, my father, the chariot of Israel, and the horsemen thereof.
2KGS|13|15|And Elisha said unto him, Take bow and arrows. And he took unto him bow and arrows.
2KGS|13|16|And he said to the king of Israel, Put thine hand upon the bow. And he put his hand upon it: and Elisha put his hands upon the king's hands.
2KGS|13|17|And he said, Open the window eastward. And he opened it. Then Elisha said, Shoot. And he shot. And he said, The arrow of the LORD's deliverance, and the arrow of deliverance from Syria: for thou shalt smite the Syrians in Aphek, till thou have consumed them.
2KGS|13|18|And he said, Take the arrows. And he took them. And he said unto the king of Israel, Smite upon the ground. And he smote thrice, and stayed.
2KGS|13|19|And the man of God was wroth with him, and said, Thou shouldest have smitten five or six times; then hadst thou smitten Syria till thou hadst consumed it: whereas now thou shalt smite Syria but thrice.
2KGS|13|20|And Elisha died, and they buried him. And the bands of the Moabites invaded the land at the coming in of the year.
2KGS|13|21|And it came to pass, as they were burying a man, that, behold, they spied a band of men; and they cast the man into the sepulchre of Elisha: and when the man was let down, and touched the bones of Elisha, he revived, and stood up on his feet.
2KGS|13|22|But Hazael king of Syria oppressed Israel all the days of Jehoahaz.
2KGS|13|23|And the LORD was gracious unto them, and had compassion on them, and had respect unto them, because of his covenant with Abraham, Isaac, and Jacob, and would not destroy them, neither cast he them from his presence as yet.
2KGS|13|24|So Hazael king of Syria died; and Benhadad his son reigned in his stead.
2KGS|13|25|And Jehoash the son of Jehoahaz took again out of the hand of Benhadad the son of Hazael the cities, which he had taken out of the hand of Jehoahaz his father by war. Three times did Joash beat him, and recovered the cities of Israel.
2KGS|14|1|In the second year of Joash son of Jehoahaz king of Israel reigned Amaziah the son of Joash king of Judah.
2KGS|14|2|He was twenty and five years old when he began to reign, and reigned twenty and nine years in Jerusalem. And his mother's name was Jehoaddan of Jerusalem.
2KGS|14|3|And he did that which was right in the sight of the LORD, yet not like David his father: he did according to all things as Joash his father did.
2KGS|14|4|Howbeit the high places were not taken away: as yet the people did sacrifice and burnt incense on the high places.
2KGS|14|5|And it came to pass, as soon as the kingdom was confirmed in his hand, that he slew his servants which had slain the king his father.
2KGS|14|6|But the children of the murderers he slew not: according unto that which is written in the book of the law of Moses, wherein the LORD commanded, saying, The fathers shall not be put to death for the children, nor the children be put to death for the fathers; but every man shall be put to death for his own sin.
2KGS|14|7|He slew of Edom in the valley of salt ten thousand, and took Selah by war, and called the name of it Joktheel unto this day.
2KGS|14|8|Then Amaziah sent messengers to Jehoash, the son of Jehoahaz son of Jehu, king of Israel, saying, Come, let us look one another in the face.
2KGS|14|9|And Jehoash the king of Israel sent to Amaziah king of Judah, saying, The thistle that was in Lebanon sent to the cedar that was in Lebanon, saying, Give thy daughter to my son to wife: and there passed by a wild beast that was in Lebanon, and trode down the thistle.
2KGS|14|10|Thou hast indeed smitten Edom, and thine heart hath lifted thee up: glory of this, and tarry at home: for why shouldest thou meddle to thy hurt, that thou shouldest fall, even thou, and Judah with thee?
2KGS|14|11|But Amaziah would not hear. Therefore Jehoash king of Israel went up; and he and Amaziah king of Judah looked one another in the face at Bethshemesh, which belongeth to Judah.
2KGS|14|12|And Judah was put to the worse before Israel; and they fled every man to their tents.
2KGS|14|13|And Jehoash king of Israel took Amaziah king of Judah, the son of Jehoash the son of Ahaziah, at Bethshemesh, and came to Jerusalem, and brake down the wall of Jerusalem from the gate of Ephraim unto the corner gate, four hundred cubits.
2KGS|14|14|And he took all the gold and silver, and all the vessels that were found in the house of the LORD, and in the treasures of the king's house, and hostages, and returned to Samaria.
2KGS|14|15|Now the rest of the acts of Jehoash which he did, and his might, and how he fought with Amaziah king of Judah, are they not written in the book of the chronicles of the kings of Israel?
2KGS|14|16|And Jehoash slept with his fathers, and was buried in Samaria with the kings of Israel; and Jeroboam his son reigned in his stead.
2KGS|14|17|And Amaziah the son of Joash king of Judah lived after the death of Jehoash son of Jehoahaz king of Israel fifteen years.
2KGS|14|18|And the rest of the acts of Amaziah, are they not written in the book of the chronicles of the kings of Judah?
2KGS|14|19|Now they made a conspiracy against him in Jerusalem: and he fled to Lachish; but they sent after him to Lachish, and slew him there.
2KGS|14|20|And they brought him on horses: and he was buried at Jerusalem with his fathers in the city of David.
2KGS|14|21|And all the people of Judah took Azariah, which was sixteen years old, and made him king instead of his father Amaziah.
2KGS|14|22|He built Elath, and restored it to Judah, after that the king slept with his fathers.
2KGS|14|23|In the fifteenth year of Amaziah the son of Joash king of Judah Jeroboam the son of Joash king of Israel began to reign in Samaria, and reigned forty and one years.
2KGS|14|24|And he did that which was evil in the sight of the LORD: he departed not from all the sins of Jeroboam the son of Nebat, who made Israel to sin.
2KGS|14|25|He restored the coast of Israel from the entering of Hamath unto the sea of the plain, according to the word of the LORD God of Israel, which he spake by the hand of his servant Jonah, the son of Amittai, the prophet, which was of Gathhepher.
2KGS|14|26|For the LORD saw the affliction of Israel, that it was very bitter: for there was not any shut up, nor any left, nor any helper for Israel.
2KGS|14|27|And the LORD said not that he would blot out the name of Israel from under heaven: but he saved them by the hand of Jeroboam the son of Joash.
2KGS|14|28|Now the rest of the acts of Jeroboam, and all that he did, and his might, how he warred, and how he recovered Damascus, and Hamath, which belonged to Judah, for Israel, are they not written in the book of the chronicles of the kings of Israel?
2KGS|14|29|And Jeroboam slept with his fathers, even with the kings of Israel; and Zachariah his son reigned in his stead.
2KGS|15|1|In the twenty and seventh year of Jeroboam king of Israel began Azariah son of Amaziah king of Judah to reign.
2KGS|15|2|Sixteen years old was he when he began to reign, and he reigned two and fifty years in Jerusalem. And his mother's name was Jecholiah of Jerusalem.
2KGS|15|3|And he did that which was right in the sight of the LORD, according to all that his father Amaziah had done;
2KGS|15|4|Save that the high places were not removed: the people sacrificed and burnt incense still on the high places.
2KGS|15|5|And the LORD smote the king, so that he was a leper unto the day of his death, and dwelt in a several house. And Jotham the king's son was over the house, judging the people of the land.
2KGS|15|6|And the rest of the acts of Azariah, and all that he did, are they not written in the book of the chronicles of the kings of Judah?
2KGS|15|7|So Azariah slept with his fathers; and they buried him with his fathers in the city of David: and Jotham his son reigned in his stead.
2KGS|15|8|In the thirty and eighth year of Azariah king of Judah did Zachariah the son of Jeroboam reign over Israel in Samaria six months.
2KGS|15|9|And he did that which was evil in the sight of the LORD, as his fathers had done: he departed not from the sins of Jeroboam the son of Nebat, who made Israel to sin.
2KGS|15|10|And Shallum the son of Jabesh conspired against him, and smote him before the people, and slew him, and reigned in his stead.
2KGS|15|11|And the rest of the acts of Zachariah, behold, they are written in the book of the chronicles of the kings of Israel.
2KGS|15|12|This was the word of the LORD which he spake unto Jehu, saying, Thy sons shall sit on the throne of Israel unto the fourth generation. And so it came to pass.
2KGS|15|13|Shallum the son of Jabesh began to reign in the nine and thirtieth year of Uzziah king of Judah; and he reigned a full month in Samaria.
2KGS|15|14|For Menahem the son of Gadi went up from Tirzah, and came to Samaria, and smote Shallum the son of Jabesh in Samaria, and slew him, and reigned in his stead.
2KGS|15|15|And the rest of the acts of Shallum, and his conspiracy which he made, behold, they are written in the book of the chronicles of the kings of Israel.
2KGS|15|16|Then Menahem smote Tiphsah, and all that were therein, and the coasts thereof from Tirzah: because they opened not to him, therefore he smote it; and all the women therein that were with child he ripped up.
2KGS|15|17|In the nine and thirtieth year of Azariah king of Judah began Menahem the son of Gadi to reign over Israel, and reigned ten years in Samaria.
2KGS|15|18|And he did that which was evil in the sight of the LORD: he departed not all his days from the sins of Jeroboam the son of Nebat, who made Israel to sin.
2KGS|15|19|And Pul the king of Assyria came against the land: and Menahem gave Pul a thousand talents of silver, that his hand might be with him to confirm the kingdom in his hand.
2KGS|15|20|And Menahem exacted the money of Israel, even of all the mighty men of wealth, of each man fifty shekels of silver, to give to the king of Assyria. So the king of Assyria turned back, and stayed not there in the land.
2KGS|15|21|And the rest of the acts of Menahem, and all that he did, are they not written in the book of the chronicles of the kings of Israel?
2KGS|15|22|And Menahem slept with his fathers; and Pekahiah his son reigned in his stead.
2KGS|15|23|In the fiftieth year of Azariah king of Judah Pekahiah the son of Menahem began to reign over Israel in Samaria, and reigned two years.
2KGS|15|24|And he did that which was evil in the sight of the LORD: he departed not from the sins of Jeroboam the son of Nebat, who made Israel to sin.
2KGS|15|25|But Pekah the son of Remaliah, a captain of his, conspired against him, and smote him in Samaria, in the palace of the king's house, with Argob and Arieh, and with him fifty men of the Gileadites: and he killed him, and reigned in his room.
2KGS|15|26|And the rest of the acts of Pekahiah, and all that he did, behold, they are written in the book of the chronicles of the kings of Israel.
2KGS|15|27|In the two and fiftieth year of Azariah king of Judah Pekah the son of Remaliah began to reign over Israel in Samaria, and reigned twenty years.
2KGS|15|28|And he did that which was evil in the sight of the LORD: he departed not from the sins of Jeroboam the son of Nebat, who made Israel to sin.
2KGS|15|29|In the days of Pekah king of Israel came Tiglathpileser king of Assyria, and took Ijon, and Abelbethmaachah, and Janoah, and Kedesh, and Hazor, and Gilead, and Galilee, all the land of Naphtali, and carried them captive to Assyria.
2KGS|15|30|And Hoshea the son of Elah made a conspiracy against Pekah the son of Remaliah, and smote him, and slew him, and reigned in his stead, in the twentieth year of Jotham the son of Uzziah.
2KGS|15|31|And the rest of the acts of Pekah, and all that he did, behold, they are written in the book of the chronicles of the kings of Israel.
2KGS|15|32|In the second year of Pekah the son of Remaliah king of Israel began Jotham the son of Uzziah king of Judah to reign.
2KGS|15|33|Five and twenty years old was he when he began to reign, and he reigned sixteen years in Jerusalem. And his mother's name was Jerusha, the daughter of Zadok.
2KGS|15|34|And he did that which was right in the sight of the LORD: he did according to all that his father Uzziah had done.
2KGS|15|35|Howbeit the high places were not removed: the people sacrificed and burned incense still in the high places. He built the higher gate of the house of the LORD.
2KGS|15|36|Now the rest of the acts of Jotham, and all that he did, are they not written in the book of the chronicles of the kings of Judah?
2KGS|15|37|In those days the LORD began to send against Judah Rezin the king of Syria, and Pekah the son of Remaliah.
2KGS|15|38|And Jotham slept with his fathers, and was buried with his fathers in the city of David his father: and Ahaz his son reigned in his stead.
2KGS|16|1|In the seventeenth year of Pekah the son of Remaliah Ahaz the son of Jotham king of Judah began to reign.
2KGS|16|2|Twenty years old was Ahaz when he began to reign, and reigned sixteen years in Jerusalem, and did not that which was right in the sight of the LORD his God, like David his father.
2KGS|16|3|But he walked in the way of the kings of Israel, yea, and made his son to pass through the fire, according to the abominations of the heathen, whom the LORD cast out from before the children of Israel.
2KGS|16|4|And he sacrificed and burnt incense in the high places, and on the hills, and under every green tree.
2KGS|16|5|Then Rezin king of Syria and Pekah son of Remaliah king of Israel came up to Jerusalem to war: and they besieged Ahaz, but could not overcome him.
2KGS|16|6|At that time Rezin king of Syria recovered Elath to Syria, and drave the Jews from Elath: and the Syrians came to Elath, and dwelt there unto this day.
2KGS|16|7|So Ahaz sent messengers to Tiglathpileser king of Assyria, saying, I am thy servant and thy son: come up, and save me out of the hand of the king of Syria, and out of the hand of the king of Israel, which rise up against me.
2KGS|16|8|And Ahaz took the silver and gold that was found in the house of the LORD, and in the treasures of the king's house, and sent it for a present to the king of Assyria.
2KGS|16|9|And the king of Assyria hearkened unto him: for the king of Assyria went up against Damascus, and took it, and carried the people of it captive to Kir, and slew Rezin.
2KGS|16|10|And king Ahaz went to Damascus to meet Tiglathpileser king of Assyria, and saw an altar that was at Damascus: and king Ahaz sent to Urijah the priest the fashion of the altar, and the pattern of it, according to all the workmanship thereof.
2KGS|16|11|And Urijah the priest built an altar according to all that king Ahaz had sent from Damascus: so Urijah the priest made it against king Ahaz came from Damascus.
2KGS|16|12|And when the king was come from Damascus, the king saw the altar: and the king approached to the altar, and offered thereon.
2KGS|16|13|And he burnt his burnt offering and his meat offering, and poured his drink offering, and sprinkled the blood of his peace offerings, upon the altar.
2KGS|16|14|And he brought also the brazen altar, which was before the LORD, from the forefront of the house, from between the altar and the house of the LORD, and put it on the north side of the altar.
2KGS|16|15|And king Ahaz commanded Urijah the priest, saying, Upon the great altar burn the morning burnt offering, and the evening meat offering, and the king's burnt sacrifice, and his meat offering, with the burnt offering of all the people of the land, and their meat offering, and their drink offerings; and sprinkle upon it all the blood of the burnt offering, and all the blood of the sacrifice: and the brazen altar shall be for me to enquire by.
2KGS|16|16|Thus did Urijah the priest, according to all that king Ahaz commanded.
2KGS|16|17|And king Ahaz cut off the borders of the bases, and removed the laver from off them; and took down the sea from off the brazen oxen that were under it, and put it upon the pavement of stones.
2KGS|16|18|And the covert for the sabbath that they had built in the house, and the king's entry without, turned he from the house of the LORD for the king of Assyria.
2KGS|16|19|Now the rest of the acts of Ahaz which he did, are they not written in the book of the chronicles of the kings of Judah?
2KGS|16|20|And Ahaz slept with his fathers, and was buried with his fathers in the city of David: and Hezekiah his son reigned in his stead.
2KGS|17|1|In the twelfth year of Ahaz king of Judah began Hoshea the son of Elah to reign in Samaria over Israel nine years.
2KGS|17|2|And he did that which was evil in the sight of the LORD, but not as the kings of Israel that were before him.
2KGS|17|3|Against him came up Shalmaneser king of Assyria; and Hoshea became his servant, and gave him presents.
2KGS|17|4|And the king of Assyria found conspiracy in Hoshea: for he had sent messengers to So king of Egypt, and brought no present to the king of Assyria, as he had done year by year: therefore the king of Assyria shut him up, and bound him in prison.
2KGS|17|5|Then the king of Assyria came up throughout all the land, and went up to Samaria, and besieged it three years.
2KGS|17|6|In the ninth year of Hoshea the king of Assyria took Samaria, and carried Israel away into Assyria, and placed them in Halah and in Habor by the river of Gozan, and in the cities of the Medes.
2KGS|17|7|For so it was, that the children of Israel had sinned against the LORD their God, which had brought them up out of the land of Egypt, from under the hand of Pharaoh king of Egypt, and had feared other gods,
2KGS|17|8|And walked in the statutes of the heathen, whom the LORD cast out from before the children of Israel, and of the kings of Israel, which they had made.
2KGS|17|9|And the children of Israel did secretly those things that were not right against the LORD their God, and they built them high places in all their cities, from the tower of the watchmen to the fenced city.
2KGS|17|10|And they set them up images and groves in every high hill, and under every green tree:
2KGS|17|11|And there they burnt incense in all the high places, as did the heathen whom the LORD carried away before them; and wrought wicked things to provoke the LORD to anger:
2KGS|17|12|For they served idols, whereof the LORD had said unto them, Ye shall not do this thing.
2KGS|17|13|Yet the LORD testified against Israel, and against Judah, by all the prophets, and by all the seers, saying, Turn ye from your evil ways, and keep my commandments and my statutes, according to all the law which I commanded your fathers, and which I sent to you by my servants the prophets.
2KGS|17|14|Notwithstanding they would not hear, but hardened their necks, like to the neck of their fathers, that did not believe in the LORD their God.
2KGS|17|15|And they rejected his statutes, and his covenant that he made with their fathers, and his testimonies which he testified against them; and they followed vanity, and became vain, and went after the heathen that were round about them, concerning whom the LORD had charged them, that they should not do like them.
2KGS|17|16|And they left all the commandments of the LORD their God, and made them molten images, even two calves, and made a grove, and worshipped all the host of heaven, and served Baal.
2KGS|17|17|And they caused their sons and their daughters to pass through the fire, and used divination and enchantments, and sold themselves to do evil in the sight of the LORD, to provoke him to anger.
2KGS|17|18|Therefore the LORD was very angry with Israel, and removed them out of his sight: there was none left but the tribe of Judah only.
2KGS|17|19|Also Judah kept not the commandments of the LORD their God, but walked in the statutes of Israel which they made.
2KGS|17|20|And the LORD rejected all the seed of Israel, and afflicted them, and delivered them into the hand of spoilers, until he had cast them out of his sight.
2KGS|17|21|For he rent Israel from the house of David; and they made Jeroboam the son of Nebat king: and Jeroboam drave Israel from following the LORD, and made them sin a great sin.
2KGS|17|22|For the children of Israel walked in all the sins of Jeroboam which he did; they departed not from them;
2KGS|17|23|Until the LORD removed Israel out of his sight, as he had said by all his servants the prophets. So was Israel carried away out of their own land to Assyria unto this day.
2KGS|17|24|And the king of Assyria brought men from Babylon, and from Cuthah, and from Ava, and from Hamath, and from Sepharvaim, and placed them in the cities of Samaria instead of the children of Israel: and they possessed Samaria, and dwelt in the cities thereof.
2KGS|17|25|And so it was at the beginning of their dwelling there, that they feared not the LORD: therefore the LORD sent lions among them, which slew some of them.
2KGS|17|26|Wherefore they spake to the king of Assyria, saying, The nations which thou hast removed, and placed in the cities of Samaria, know not the manner of the God of the land: therefore he hath sent lions among them, and, behold, they slay them, because they know not the manner of the God of the land.
2KGS|17|27|Then the king of Assyria commanded, saying, Carry thither one of the priests whom ye brought from thence; and let them go and dwell there, and let him teach them the manner of the God of the land.
2KGS|17|28|Then one of the priests whom they had carried away from Samaria came and dwelt in Bethel, and taught them how they should fear the LORD.
2KGS|17|29|Howbeit every nation made gods of their own, and put them in the houses of the high places which the Samaritans had made, every nation in their cities wherein they dwelt.
2KGS|17|30|And the men of Babylon made Succothbenoth, and the men of Cuth made Nergal, and the men of Hamath made Ashima,
2KGS|17|31|And the Avites made Nibhaz and Tartak, and the Sepharvites burnt their children in fire to Adrammelech and Anammelech, the gods of Sepharvaim.
2KGS|17|32|So they feared the LORD, and made unto themselves of the lowest of them priests of the high places, which sacrificed for them in the houses of the high places.
2KGS|17|33|They feared the LORD, and served their own gods, after the manner of the nations whom they carried away from thence.
2KGS|17|34|Unto this day they do after the former manners: they fear not the LORD, neither do they after their statutes, or after their ordinances, or after the law and commandment which the LORD commanded the children of Jacob, whom he named Israel;
2KGS|17|35|With whom the LORD had made a covenant, and charged them, saying, Ye shall not fear other gods, nor bow yourselves to them, nor serve them, nor sacrifice to them:
2KGS|17|36|But the LORD, who brought you up out of the land of Egypt with great power and a stretched out arm, him shall ye fear, and him shall ye worship, and to him shall ye do sacrifice.
2KGS|17|37|And the statutes, and the ordinances, and the law, and the commandment, which he wrote for you, ye shall observe to do for evermore; and ye shall not fear other gods.
2KGS|17|38|And the covenant that I have made with you ye shall not forget; neither shall ye fear other gods.
2KGS|17|39|But the LORD your God ye shall fear; and he shall deliver you out of the hand of all your enemies.
2KGS|17|40|Howbeit they did not hearken, but they did after their former manner.
2KGS|17|41|So these nations feared the LORD, and served their graven images, both their children, and their children's children: as did their fathers, so do they unto this day.
2KGS|18|1|Now it came to pass in the third year of Hoshea son of Elah king of Israel, that Hezekiah the son of Ahaz king of Judah began to reign.
2KGS|18|2|Twenty and five years old was he when he began to reign; and he reigned twenty and nine years in Jerusalem. His mother's name also was Abi, the daughter of Zachariah.
2KGS|18|3|And he did that which was right in the sight of the LORD, according to all that David his father did.
2KGS|18|4|He removed the high places, and brake the images, and cut down the groves, and brake in pieces the brazen serpent that Moses had made: for unto those days the children of Israel did burn incense to it: and he called it Nehushtan.
2KGS|18|5|He trusted in the LORD God of Israel; so that after him was none like him among all the kings of Judah, nor any that were before him.
2KGS|18|6|For he clave to the LORD, and departed not from following him, but kept his commandments, which the LORD commanded Moses.
2KGS|18|7|And the LORD was with him; and he prospered whithersoever he went forth: and he rebelled against the king of Assyria, and served him not.
2KGS|18|8|He smote the Philistines, even unto Gaza, and the borders thereof, from the tower of the watchmen to the fenced city.
2KGS|18|9|And it came to pass in the fourth year of king Hezekiah, which was the seventh year of Hoshea son of Elah king of Israel, that Shalmaneser king of Assyria came up against Samaria, and besieged it.
2KGS|18|10|And at the end of three years they took it: even in the sixth year of Hezekiah, that is in the ninth year of Hoshea king of Israel, Samaria was taken.
2KGS|18|11|And the king of Assyria did carry away Israel unto Assyria, and put them in Halah and in Habor by the river of Gozan, and in the cities of the Medes:
2KGS|18|12|Because they obeyed not the voice of the LORD their God, but transgressed his covenant, and all that Moses the servant of the LORD commanded, and would not hear them, nor do them.
2KGS|18|13|Now in the fourteenth year of king Hezekiah did Sennacherib king of Assyria come up against all the fenced cities of Judah, and took them.
2KGS|18|14|And Hezekiah king of Judah sent to the king of Assyria to Lachish, saying, I have offended; return from me: that which thou puttest on me will I bear. And the king of Assyria appointed unto Hezekiah king of Judah three hundred talents of silver and thirty talents of gold.
2KGS|18|15|And Hezekiah gave him all the silver that was found in the house of the LORD, and in the treasures of the king's house.
2KGS|18|16|At that time did Hezekiah cut off the gold from the doors of the temple of the LORD, and from the pillars which Hezekiah king of Judah had overlaid, and gave it to the king of Assyria.
2KGS|18|17|And the king of Assyria sent Tartan and Rabsaris and Rabshakeh from Lachish to king Hezekiah with a great host against Jerusalem. And they went up and came to Jerusalem. And when they were come up, they came and stood by the conduit of the upper pool, which is in the highway of the fuller's field.
2KGS|18|18|And when they had called to the king, there came out to them Eliakim the son of Hilkiah, which was over the household, and Shebna the scribe, and Joah the son of Asaph the recorder.
2KGS|18|19|And Rabshakeh said unto them, Speak ye now to Hezekiah, Thus saith the great king, the king of Assyria, What confidence is this wherein thou trustest?
2KGS|18|20|Thou sayest, (but they are but vain words,) I have counsel and strength for the war. Now on whom dost thou trust, that thou rebellest against me?
2KGS|18|21|Now, behold, thou trustest upon the staff of this bruised reed, even upon Egypt, on which if a man lean, it will go into his hand, and pierce it: so is Pharaoh king of Egypt unto all that trust on him.
2KGS|18|22|But if ye say unto me, We trust in the LORD our God: is not that he, whose high places and whose altars Hezekiah hath taken away, and hath said to Judah and Jerusalem, Ye shall worship before this altar in Jerusalem?
2KGS|18|23|Now therefore, I pray thee, give pledges to my lord the king of Assyria, and I will deliver thee two thousand horses, if thou be able on thy part to set riders upon them.
2KGS|18|24|How then wilt thou turn away the face of one captain of the least of my master's servants, and put thy trust on Egypt for chariots and for horsemen?
2KGS|18|25|Am I now come up without the LORD against this place to destroy it? The LORD said to me, Go up against this land, and destroy it.
2KGS|18|26|Then said Eliakim the son of Hilkiah, and Shebna, and Joah, unto Rabshakeh, Speak, I pray thee, to thy servants in the Syrian language; for we understand it: and talk not with us in the Jews' language in the ears of the people that are on the wall.
2KGS|18|27|But Rabshakeh said unto them, Hath my master sent me to thy master, and to thee, to speak these words? hath he not sent me to the men which sit on the wall, that they may eat their own dung, and drink their own piss with you?
2KGS|18|28|Then Rabshakeh stood and cried with a loud voice in the Jews' language, and spake, saying, Hear the word of the great king, the king of Assyria:
2KGS|18|29|Thus saith the king, Let not Hezekiah deceive you: for he shall not be able to deliver you out of his hand:
2KGS|18|30|Neither let Hezekiah make you trust in the LORD, saying, The LORD will surely deliver us, and this city shall not be delivered into the hand of the king of Assyria.
2KGS|18|31|Hearken not to Hezekiah: for thus saith the king of Assyria, Make an agreement with me by a present, and come out to me, and then eat ye every man of his own vine, and every one of his fig tree, and drink ye every one the waters of his cistern:
2KGS|18|32|Until I come and take you away to a land like your own land, a land of corn and wine, a land of bread and vineyards, a land of oil olive and of honey, that ye may live, and not die: and hearken not unto Hezekiah, when he persuadeth you, saying, The LORD will deliver us.
2KGS|18|33|Hath any of the gods of the nations delivered at all his land out of the hand of the king of Assyria?
2KGS|18|34|Where are the gods of Hamath, and of Arpad? where are the gods of Sepharvaim, Hena, and Ivah? have they delivered Samaria out of mine hand?
2KGS|18|35|Who are they among all the gods of the countries, that have delivered their country out of mine hand, that the LORD should deliver Jerusalem out of mine hand?
2KGS|18|36|But the people held their peace, and answered him not a word: for the king's commandment was, saying, Answer him not.
2KGS|18|37|Then came Eliakim the son of Hilkiah, which was over the household, and Shebna the scribe, and Joah the son of Asaph the recorder, to Hezekiah with their clothes rent, and told him the words of Rabshakeh.
2KGS|19|1|And it came to pass, when king Hezekiah heard it, that he rent his clothes, and covered himself with sackcloth, and went into the house of the LORD.
2KGS|19|2|And he sent Eliakim, which was over the household, and Shebna the scribe, and the elders of the priests, covered with sackcloth, to Isaiah the prophet the son of Amoz.
2KGS|19|3|And they said unto him, Thus saith Hezekiah, This day is a day of trouble, and of rebuke, and blasphemy; for the children are come to the birth, and there is not strength to bring forth.
2KGS|19|4|It may be the LORD thy God will hear all the words of Rabshakeh, whom the king of Assyria his master hath sent to reproach the living God; and will reprove the words which the LORD thy God hath heard: wherefore lift up thy prayer for the remnant that are left.
2KGS|19|5|So the servants of king Hezekiah came to Isaiah.
2KGS|19|6|And Isaiah said unto them, Thus shall ye say to your master, Thus saith the LORD, Be not afraid of the words which thou hast heard, with which the servants of the king of Assyria have blasphemed me.
2KGS|19|7|Behold, I will send a blast upon him, and he shall hear a rumor, and shall return to his own land; and I will cause him to fall by the sword in his own land.
2KGS|19|8|So Rabshakeh returned, and found the king of Assyria warring against Libnah: for he had heard that he was departed from Lachish.
2KGS|19|9|And when he heard say of Tirhakah king of Ethiopia, Behold, he is come out to fight against thee: he sent messengers again unto Hezekiah, saying,
2KGS|19|10|Thus shall ye speak to Hezekiah king of Judah, saying, Let not thy God in whom thou trustest deceive thee, saying, Jerusalem shall not be delivered into the hand of the king of Assyria.
2KGS|19|11|Behold, thou hast heard what the kings of Assyria have done to all lands, by destroying them utterly: and shalt thou be delivered?
2KGS|19|12|Have the gods of the nations delivered them which my fathers have destroyed; as Gozan, and Haran, and Rezeph, and the children of Eden which were in Thelasar?
2KGS|19|13|Where is the king of Hamath, and the king of Arpad, and the king of the city of Sepharvaim, of Hena, and Ivah?
2KGS|19|14|And Hezekiah received the letter of the hand of the messengers, and read it: and Hezekiah went up into the house of the LORD, and spread it before the LORD.
2KGS|19|15|And Hezekiah prayed before the LORD, and said, O LORD God of Israel, which dwellest between the cherubim, thou art the God, even thou alone, of all the kingdoms of the earth; thou hast made heaven and earth.
2KGS|19|16|LORD, bow down thine ear, and hear: open, LORD, thine eyes, and see: and hear the words of Sennacherib, which hath sent him to reproach the living God.
2KGS|19|17|Of a truth, LORD, the kings of Assyria have destroyed the nations and their lands,
2KGS|19|18|And have cast their gods into the fire: for they were no gods, but the work of men's hands, wood and stone: therefore they have destroyed them.
2KGS|19|19|Now therefore, O LORD our God, I beseech thee, save thou us out of his hand, that all the kingdoms of the earth may know that thou art the LORD God, even thou only.
2KGS|19|20|Then Isaiah the son of Amoz sent to Hezekiah, saying, Thus saith the LORD God of Israel, That which thou hast prayed to me against Sennacherib king of Assyria I have heard.
2KGS|19|21|This is the word that the LORD hath spoken concerning him; The virgin the daughter of Zion hath despised thee, and laughed thee to scorn; the daughter of Jerusalem hath shaken her head at thee.
2KGS|19|22|Whom hast thou reproached and blasphemed? and against whom hast thou exalted thy voice, and lifted up thine eyes on high? even against the Holy One of Israel.
2KGS|19|23|By thy messengers thou hast reproached the LORD, and hast said, With the multitude of my chariots I am come up to the height of the mountains, to the sides of Lebanon, and will cut down the tall cedar trees thereof, and the choice fir trees thereof: and I will enter into the lodgings of his borders, and into the forest of his Carmel.
2KGS|19|24|I have digged and drunk strange waters, and with the sole of my feet have I dried up all the rivers of besieged places.
2KGS|19|25|Hast thou not heard long ago how I have done it, and of ancient times that I have formed it? now have I brought it to pass, that thou shouldest be to lay waste fenced cities into ruinous heaps.
2KGS|19|26|Therefore their inhabitants were of small power, they were dismayed and confounded; they were as the grass of the field, and as the green herb, as the grass on the house tops, and as corn blasted before it be grown up.
2KGS|19|27|But I know thy abode, and thy going out, and thy coming in, and thy rage against me.
2KGS|19|28|Because thy rage against me and thy tumult is come up into mine ears, therefore I will put my hook in thy nose, and my bridle in thy lips, and I will turn thee back by the way by which thou camest.
2KGS|19|29|And this shall be a sign unto thee, Ye shall eat this year such things as grow of themselves, and in the second year that which springeth of the same; and in the third year sow ye, and reap, and plant vineyards, and eat the fruits thereof.
2KGS|19|30|And the remnant that is escaped of the house of Judah shall yet again take root downward, and bear fruit upward.
2KGS|19|31|For out of Jerusalem shall go forth a remnant, and they that escape out of mount Zion: the zeal of the LORD of hosts shall do this.
2KGS|19|32|Therefore thus saith the LORD concerning the king of Assyria, He shall not come into this city, nor shoot an arrow there, nor come before it with shield, nor cast a bank against it.
2KGS|19|33|By the way that he came, by the same shall he return, and shall not come into this city, saith the LORD.
2KGS|19|34|For I will defend this city, to save it, for mine own sake, and for my servant David's sake.
2KGS|19|35|And it came to pass that night, that the angel of the LORD went out, and smote in the camp of the Assyrians an hundred fourscore and five thousand: and when they arose early in the morning, behold, they were all dead corpses.
2KGS|19|36|So Sennacherib king of Assyria departed, and went and returned, and dwelt at Nineveh.
2KGS|19|37|And it came to pass, as he was worshipping in the house of Nisroch his god, that Adrammelech and Sharezer his sons smote him with the sword: and they escaped into the land of Armenia. And Esarhaddon his son reigned in his stead.
2KGS|20|1|In those days was Hezekiah sick unto death. And the prophet Isaiah the son of Amoz came to him, and said unto him, Thus saith the LORD, Set thine house in order; for thou shalt die, and not live.
2KGS|20|2|Then he turned his face to the wall, and prayed unto the LORD, saying,
2KGS|20|3|I beseech thee, O LORD, remember now how I have walked before thee in truth and with a perfect heart, and have done that which is good in thy sight. And Hezekiah wept sore.
2KGS|20|4|And it came to pass, afore Isaiah was gone out into the middle court, that the word of the LORD came to him, saying,
2KGS|20|5|Turn again, and tell Hezekiah the captain of my people, Thus saith the LORD, the God of David thy father, I have heard thy prayer, I have seen thy tears: behold, I will heal thee: on the third day thou shalt go up unto the house of the LORD.
2KGS|20|6|And I will add unto thy days fifteen years; and I will deliver thee and this city out of the hand of the king of Assyria; and I will defend this city for mine own sake, and for my servant David's sake.
2KGS|20|7|And Isaiah said, Take a lump of figs. And they took and laid it on the boil, and he recovered.
2KGS|20|8|And Hezekiah said unto Isaiah, What shall be the sign that the LORD will heal me, and that I shall go up into the house of the LORD the third day?
2KGS|20|9|And Isaiah said, This sign shalt thou have of the LORD, that the LORD will do the thing that he hath spoken: shall the shadow go forward ten degrees, or go back ten degrees?
2KGS|20|10|And Hezekiah answered, It is a light thing for the shadow to go down ten degrees: nay, but let the shadow return backward ten degrees.
2KGS|20|11|And Isaiah the prophet cried unto the LORD: and he brought the shadow ten degrees backward, by which it had gone down in the dial of Ahaz.
2KGS|20|12|At that time Berodachbaladan, the son of Baladan, king of Babylon, sent letters and a present unto Hezekiah: for he had heard that Hezekiah had been sick.
2KGS|20|13|And Hezekiah hearkened unto them, and showed them all the house of his precious things, the silver, and the gold, and the spices, and the precious ointment, and all the house of his armor, and all that was found in his treasures: there was nothing in his house, nor in all his dominion, that Hezekiah showed them not.
2KGS|20|14|Then came Isaiah the prophet unto king Hezekiah, and said unto him, What said these men? and from whence came they unto thee? And Hezekiah said, They are come from a far country, even from Babylon.
2KGS|20|15|And he said, What have they seen in thine house? And Hezekiah answered, All the things that are in mine house have they seen: there is nothing among my treasures that I have not showed them.
2KGS|20|16|And Isaiah said unto Hezekiah, Hear the word of the LORD.
2KGS|20|17|Behold, the days come, that all that is in thine house, and that which thy fathers have laid up in store unto this day, shall be carried into Babylon: nothing shall be left, saith the LORD.
2KGS|20|18|And of thy sons that shall issue from thee, which thou shalt beget, shall they take away; and they shall be eunuchs in the palace of the king of Babylon.
2KGS|20|19|Then said Hezekiah unto Isaiah, Good is the word of the LORD which thou hast spoken. And he said, Is it not good, if peace and truth be in my days?
2KGS|20|20|And the rest of the acts of Hezekiah, and all his might, and how he made a pool, and a conduit, and brought water into the city, are they not written in the book of the chronicles of the kings of Judah?
2KGS|20|21|And Hezekiah slept with his fathers: and Manasseh his son reigned in his stead.
2KGS|21|1|Manasseh was twelve years old when he began to reign, and reigned fifty and five years in Jerusalem. And his mother's name was Hephzibah.
2KGS|21|2|And he did that which was evil in the sight of the LORD, after the abominations of the heathen, whom the LORD cast out before the children of Israel.
2KGS|21|3|For he built up again the high places which Hezekiah his father had destroyed; and he reared up altars for Baal, and made a grove, as did Ahab king of Israel; and worshipped all the host of heaven, and served them.
2KGS|21|4|And he built altars in the house of the LORD, of which the LORD said, In Jerusalem will I put my name.
2KGS|21|5|And he built altars for all the host of heaven in the two courts of the house of the LORD.
2KGS|21|6|And he made his son pass through the fire, and observed times, and used enchantments, and dealt with familiar spirits and wizards: he wrought much wickedness in the sight of the LORD, to provoke him to anger.
2KGS|21|7|And he set a graven image of the grove that he had made in the house, of which the LORD said to David, and to Solomon his son, In this house, and in Jerusalem, which I have chosen out of all tribes of Israel, will I put my name for ever:
2KGS|21|8|Neither will I make the feet of Israel move any more out of the land which I gave their fathers; only if they will observe to do according to all that I have commanded them, and according to all the law that my servant Moses commanded them.
2KGS|21|9|But they hearkened not: and Manasseh seduced them to do more evil than did the nations whom the LORD destroyed before the children of Israel.
2KGS|21|10|And the LORD spake by his servants the prophets, saying,
2KGS|21|11|Because Manasseh king of Judah hath done these abominations, and hath done wickedly above all that the Amorites did, which were before him, and hath made Judah also to sin with his idols:
2KGS|21|12|Therefore thus saith the LORD God of Israel, Behold, I am bringing such evil upon Jerusalem and Judah, that whosoever heareth of it, both his ears shall tingle.
2KGS|21|13|And I will stretch over Jerusalem the line of Samaria, and the plummet of the house of Ahab: and I will wipe Jerusalem as a man wipeth a dish, wiping it, and turning it upside down.
2KGS|21|14|And I will forsake the remnant of mine inheritance, and deliver them into the hand of their enemies; and they shall become a prey and a spoil to all their enemies;
2KGS|21|15|Because they have done that which was evil in my sight, and have provoked me to anger, since the day their fathers came forth out of Egypt, even unto this day.
2KGS|21|16|Moreover Manasseh shed innocent blood very much, till he had filled Jerusalem from one end to another; beside his sin wherewith he made Judah to sin, in doing that which was evil in the sight of the LORD.
2KGS|21|17|Now the rest of the acts of Manasseh, and all that he did, and his sin that he sinned, are they not written in the book of the chronicles of the kings of Judah?
2KGS|21|18|And Manasseh slept with his fathers, and was buried in the garden of his own house, in the garden of Uzza: and Amon his son reigned in his stead.
2KGS|21|19|Amon was twenty and two years old when he began to reign, and he reigned two years in Jerusalem. And his mother's name was Meshullemeth, the daughter of Haruz of Jotbah.
2KGS|21|20|And he did that which was evil in the sight of the LORD, as his father Manasseh did.
2KGS|21|21|And he walked in all the way that his father walked in, and served the idols that his father served, and worshipped them:
2KGS|21|22|And he forsook the LORD God of his fathers, and walked not in the way of the LORD.
2KGS|21|23|And the servants of Amon conspired against him, and slew the king in his own house.
2KGS|21|24|And the people of the land slew all them that had conspired against king Amon; and the people of the land made Josiah his son king in his stead.
2KGS|21|25|Now the rest of the acts of Amon which he did, are they not written in the book of the chronicles of the kings of Judah?
2KGS|21|26|And he was buried in his sepulchre in the garden of Uzza: and Josiah his son reigned in his stead.
2KGS|22|1|Josiah was eight years old when he began to reign, and he reigned thirty and one years in Jerusalem. And his mother's name was Jedidah, the daughter of Adaiah of Boscath.
2KGS|22|2|And he did that which was right in the sight of the LORD, and walked in all the way of David his father, and turned not aside to the right hand or to the left.
2KGS|22|3|And it came to pass in the eighteenth year of king Josiah, that the king sent Shaphan the son of Azaliah, the son of Meshullam, the scribe, to the house of the LORD, saying,
2KGS|22|4|Go up to Hilkiah the high priest, that he may sum the silver which is brought into the house of the LORD, which the keepers of the door have gathered of the people:
2KGS|22|5|And let them deliver it into the hand of the doers of the work, that have the oversight of the house of the LORD: and let them give it to the doers of the work which is in the house of the LORD, to repair the breaches of the house,
2KGS|22|6|Unto carpenters, and builders, and masons, and to buy timber and hewn stone to repair the house.
2KGS|22|7|Howbeit there was no reckoning made with them of the money that was delivered into their hand, because they dealt faithfully.
2KGS|22|8|And Hilkiah the high priest said unto Shaphan the scribe, I have found the book of the law in the house of the LORD. And Hilkiah gave the book to Shaphan, and he read it.
2KGS|22|9|And Shaphan the scribe came to the king, and brought the king word again, and said, Thy servants have gathered the money that was found in the house, and have delivered it into the hand of them that do the work, that have the oversight of the house of the LORD.
2KGS|22|10|And Shaphan the scribe showed the king, saying, Hilkiah the priest hath delivered me a book. And Shaphan read it before the king.
2KGS|22|11|And it came to pass, when the king had heard the words of the book of the law, that he rent his clothes.
2KGS|22|12|And the king commanded Hilkiah the priest, and Ahikam the son of Shaphan, and Achbor the son of Michaiah, and Shaphan the scribe, and Asahiah a servant of the king's, saying,
2KGS|22|13|Go ye, enquire of the LORD for me, and for the people, and for all Judah, concerning the words of this book that is found: for great is the wrath of the LORD that is kindled against us, because our fathers have not hearkened unto the words of this book, to do according unto all that which is written concerning us.
2KGS|22|14|So Hilkiah the priest, and Ahikam, and Achbor, and Shaphan, and Asahiah, went unto Huldah the prophetess, the wife of Shallum the son of Tikvah, the son of Harhas, keeper of the wardrobe; (now she dwelt in Jerusalem in the college;) and they communed with her.
2KGS|22|15|And she said unto them, Thus saith the LORD God of Israel, Tell the man that sent you to me,
2KGS|22|16|Thus saith the LORD, Behold, I will bring evil upon this place, and upon the inhabitants thereof, even all the words of the book which the king of Judah hath read:
2KGS|22|17|Because they have forsaken me, and have burned incense unto other gods, that they might provoke me to anger with all the works of their hands; therefore my wrath shall be kindled against this place, and shall not be quenched.
2KGS|22|18|But to the king of Judah which sent you to enquire of the LORD, thus shall ye say to him, Thus saith the LORD God of Israel, As touching the words which thou hast heard;
2KGS|22|19|Because thine heart was tender, and thou hast humbled thyself before the LORD, when thou heardest what I spake against this place, and against the inhabitants thereof, that they should become a desolation and a curse, and hast rent thy clothes, and wept before me; I also have heard thee, saith the LORD.
2KGS|22|20|Behold therefore, I will gather thee unto thy fathers, and thou shalt be gathered into thy grave in peace; and thine eyes shall not see all the evil which I will bring upon this place. And they brought the king word again.
2KGS|23|1|And the king sent, and they gathered unto him all the elders of Judah and of Jerusalem.
2KGS|23|2|And the king went up into the house of the LORD, and all the men of Judah and all the inhabitants of Jerusalem with him, and the priests, and the prophets, and all the people, both small and great: and he read in their ears all the words of the book of the covenant which was found in the house of the LORD.
2KGS|23|3|And the king stood by a pillar, and made a covenant before the LORD, to walk after the LORD, and to keep his commandments and his testimonies and his statutes with all their heart and all their soul, to perform the words of this covenant that were written in this book. And all the people stood to the covenant.
2KGS|23|4|And the king commanded Hilkiah the high priest, and the priests of the second order, and the keepers of the door, to bring forth out of the temple of the LORD all the vessels that were made for Baal, and for the grove, and for all the host of heaven: and he burned them without Jerusalem in the fields of Kidron, and carried the ashes of them unto Bethel.
2KGS|23|5|And he put down the idolatrous priests, whom the kings of Judah had ordained to burn incense in the high places in the cities of Judah, and in the places round about Jerusalem; them also that burned incense unto Baal, to the sun, and to the moon, and to the planets, and to all the host of heaven.
2KGS|23|6|And he brought out the grove from the house of the LORD, without Jerusalem, unto the brook Kidron, and burned it at the brook Kidron, and stamped it small to powder, and cast the powder thereof upon the graves of the children of the people.
2KGS|23|7|And he brake down the houses of the sodomites, that were by the house of the LORD, where the women wove hangings for the grove.
2KGS|23|8|And he brought all the priests out of the cities of Judah, and defiled the high places where the priests had burned incense, from Geba to Beersheba, and brake down the high places of the gates that were in the entering in of the gate of Joshua the governor of the city, which were on a man's left hand at the gate of the city.
2KGS|23|9|Nevertheless the priests of the high places came not up to the altar of the LORD in Jerusalem, but they did eat of the unleavened bread among their brethren.
2KGS|23|10|And he defiled Topheth, which is in the valley of the children of Hinnom, that no man might make his son or his daughter to pass through the fire to Molech.
2KGS|23|11|And he took away the horses that the kings of Judah had given to the sun, at the entering in of the house of the LORD, by the chamber of Nathanmelech the chamberlain, which was in the suburbs, and burned the chariots of the sun with fire.
2KGS|23|12|And the altars that were on the top of the upper chamber of Ahaz, which the kings of Judah had made, and the altars which Manasseh had made in the two courts of the house of the LORD, did the king beat down, and brake them down from thence, and cast the dust of them into the brook Kidron.
2KGS|23|13|And the high places that were before Jerusalem, which were on the right hand of the mount of corruption, which Solomon the king of Israel had builded for Ashtoreth the abomination of the Zidonians, and for Chemosh the abomination of the Moabites, and for Milcom the abomination of the children of Ammon, did the king defile.
2KGS|23|14|And he brake in pieces the images, and cut down the groves, and filled their places with the bones of men.
2KGS|23|15|Moreover the altar that was at Bethel, and the high place which Jeroboam the son of Nebat, who made Israel to sin, had made, both that altar and the high place he brake down, and burned the high place, and stamped it small to powder, and burned the grove.
2KGS|23|16|And as Josiah turned himself, he spied the sepulchres that were there in the mount, and sent, and took the bones out of the sepulchres, and burned them upon the altar, and polluted it, according to the word of the LORD which the man of God proclaimed, who proclaimed these words.
2KGS|23|17|Then he said, What title is that that I see? And the men of the city told him, It is the sepulchre of the man of God, which came from Judah, and proclaimed these things that thou hast done against the altar of Bethel.
2KGS|23|18|And he said, Let him alone; let no man move his bones. So they let his bones alone, with the bones of the prophet that came out of Samaria.
2KGS|23|19|And all the houses also of the high places that were in the cities of Samaria, which the kings of Israel had made to provoke the Lord to anger, Josiah took away, and did to them according to all the acts that he had done in Bethel.
2KGS|23|20|And he slew all the priests of the high places that were there upon the altars, and burned men's bones upon them, and returned to Jerusalem.
2KGS|23|21|And the king commanded all the people, saying, Keep the passover unto the LORD your God, as it is written in the book of this covenant.
2KGS|23|22|Surely there was not holden such a passover from the days of the judges that judged Israel, nor in all the days of the kings of Israel, nor of the kings of Judah;
2KGS|23|23|But in the eighteenth year of king Josiah, wherein this passover was holden to the LORD in Jerusalem.
2KGS|23|24|Moreover the workers with familiar spirits, and the wizards, and the images, and the idols, and all the abominations that were spied in the land of Judah and in Jerusalem, did Josiah put away, that he might perform the words of the law which were written in the book that Hilkiah the priest found in the house of the LORD.
2KGS|23|25|And like unto him was there no king before him, that turned to the LORD with all his heart, and with all his soul, and with all his might, according to all the law of Moses; neither after him arose there any like him.
2KGS|23|26|Notwithstanding the LORD turned not from the fierceness of his great wrath, wherewith his anger was kindled against Judah, because of all the provocations that Manasseh had provoked him withal.
2KGS|23|27|And the LORD said, I will remove Judah also out of my sight, as I have removed Israel, and will cast off this city Jerusalem which I have chosen, and the house of which I said, My name shall be there.
2KGS|23|28|Now the rest of the acts of Josiah, and all that he did, are they not written in the book of the chronicles of the kings of Judah?
2KGS|23|29|In his days Pharaohnechoh king of Egypt went up against the king of Assyria to the river Euphrates: and king Josiah went against him; and he slew him at Megiddo, when he had seen him.
2KGS|23|30|And his servants carried him in a chariot dead from Megiddo, and brought him to Jerusalem, and buried him in his own sepulchre. And the people of the land took Jehoahaz the son of Josiah, and anointed him, and made him king in his father's stead.
2KGS|23|31|Jehoahaz was twenty and three years old when he began to reign; and he reigned three months in Jerusalem. And his mother's name was Hamutal, the daughter of Jeremiah of Libnah.
2KGS|23|32|And he did that which was evil in the sight of the LORD, according to all that his fathers had done.
2KGS|23|33|And Pharaohnechoh put him in bands at Riblah in the land of Hamath, that he might not reign in Jerusalem; and put the land to a tribute of an hundred talents of silver, and a talent of gold.
2KGS|23|34|And Pharaohnechoh made Eliakim the son of Josiah king in the room of Josiah his father, and turned his name to Jehoiakim, and took Jehoahaz away: and he came to Egypt, and died there.
2KGS|23|35|And Jehoiakim gave the silver and the gold to Pharaoh; but he taxed the land to give the money according to the commandment of Pharaoh: he exacted the silver and the gold of the people of the land, of every one according to his taxation, to give it unto Pharaohnechoh.
2KGS|23|36|Jehoiakim was twenty and five years old when he began to reign; and he reigned eleven years in Jerusalem. And his mother's name was Zebudah, the daughter of Pedaiah of Rumah.
2KGS|23|37|And he did that which was evil in the sight of the LORD, according to all that his fathers had done.
2KGS|24|1|In his days Nebuchadnezzar king of Babylon came up, and Jehoiakim became his servant three years: then he turned and rebelled against him.
2KGS|24|2|And the LORD sent against him bands of the Chaldees, and bands of the Syrians, and bands of the Moabites, and bands of the children of Ammon, and sent them against Judah to destroy it, according to the word of the LORD, which he spake by his servants the prophets.
2KGS|24|3|Surely at the commandment of the LORD came this upon Judah, to remove them out of his sight, for the sins of Manasseh, according to all that he did;
2KGS|24|4|And also for the innocent blood that he shed: for he filled Jerusalem with innocent blood; which the LORD would not pardon.
2KGS|24|5|Now the rest of the acts of Jehoiakim, and all that he did, are they not written in the book of the chronicles of the kings of Judah?
2KGS|24|6|So Jehoiakim slept with his fathers: and Jehoiachin his son reigned in his stead.
2KGS|24|7|And the king of Egypt came not again any more out of his land: for the king of Babylon had taken from the river of Egypt unto the river Euphrates all that pertained to the king of Egypt.
2KGS|24|8|Jehoiachin was eighteen years old when he began to reign, and he reigned in Jerusalem three months. And his mother's name was Nehushta, the daughter of Elnathan of Jerusalem.
2KGS|24|9|And he did that which was evil in the sight of the LORD, according to all that his father had done.
2KGS|24|10|At that time the servants of Nebuchadnezzar king of Babylon came up against Jerusalem, and the city was besieged.
2KGS|24|11|And Nebuchadnezzar king of Babylon came against the city, and his servants did besiege it.
2KGS|24|12|And Jehoiachin the king of Judah went out to the king of Babylon, he, and his mother, and his servants, and his princes, and his officers: and the king of Babylon took him in the eighth year of his reign.
2KGS|24|13|And he carried out thence all the treasures of the house of the LORD, and the treasures of the king's house, and cut in pieces all the vessels of gold which Solomon king of Israel had made in the temple of the LORD, as the LORD had said.
2KGS|24|14|And he carried away all Jerusalem, and all the princes, and all the mighty men of valor, even ten thousand captives, and all the craftsmen and smiths: none remained, save the poorest sort of the people of the land.
2KGS|24|15|And he carried away Jehoiachin to Babylon, and the king's mother, and the king's wives, and his officers, and the mighty of the land, those carried he into captivity from Jerusalem to Babylon.
2KGS|24|16|And all the men of might, even seven thousand, and craftsmen and smiths a thousand, all that were strong and apt for war, even them the king of Babylon brought captive to Babylon.
2KGS|24|17|And the king of Babylon made Mattaniah his father's brother king in his stead, and changed his name to Zedekiah.
2KGS|24|18|Zedekiah was twenty and one years old when he began to reign, and he reigned eleven years in Jerusalem. And his mother's name was Hamutal, the daughter of Jeremiah of Libnah.
2KGS|24|19|And he did that which was evil in the sight of the LORD, according to all that Jehoiakim had done.
2KGS|24|20|For through the anger of the LORD it came to pass in Jerusalem and Judah, until he had cast them out from his presence, that Zedekiah rebelled against the king of Babylon.
2KGS|25|1|And it came to pass in the ninth year of his reign, in the tenth month, in the tenth day of the month, that Nebuchadnezzar king of Babylon came, he, and all his host, against Jerusalem, and pitched against it; and they built forts against it round about.
2KGS|25|2|And the city was besieged unto the eleventh year of king Zedekiah.
2KGS|25|3|And on the ninth day of the fourth month the famine prevailed in the city, and there was no bread for the people of the land.
2KGS|25|4|And the city was broken up, and all the men of war fled by night by the way of the gate between two walls, which is by the king's garden: (now the Chaldees were against the city round about:) and the king went the way toward the plain.
2KGS|25|5|And the army of the Chaldees pursued after the king, and overtook him in the plains of Jericho: and all his army were scattered from him.
2KGS|25|6|So they took the king, and brought him up to the king of Babylon to Riblah; and they gave judgment upon him.
2KGS|25|7|And they slew the sons of Zedekiah before his eyes, and put out the eyes of Zedekiah, and bound him with fetters of brass, and carried him to Babylon.
2KGS|25|8|And in the fifth month, on the seventh day of the month, which is the nineteenth year of king Nebuchadnezzar king of Babylon, came Nebuzaradan, captain of the guard, a servant of the king of Babylon, unto Jerusalem:
2KGS|25|9|And he burnt the house of the LORD, and the king's house, and all the houses of Jerusalem, and every great man's house burnt he with fire.
2KGS|25|10|And all the army of the Chaldees, that were with the captain of the guard, brake down the walls of Jerusalem round about.
2KGS|25|11|Now the rest of the people that were left in the city, and the fugitives that fell away to the king of Babylon, with the remnant of the multitude, did Nebuzaradan the captain of the guard carry away.
2KGS|25|12|But the captain of the guard left of the door of the poor of the land to be vinedressers and husbandmen.
2KGS|25|13|And the pillars of brass that were in the house of the LORD, and the bases, and the brazen sea that was in the house of the LORD, did the Chaldees break in pieces, and carried the brass of them to Babylon.
2KGS|25|14|And the pots, and the shovels, and the snuffers, and the spoons, and all the vessels of brass wherewith they ministered, took they away.
2KGS|25|15|And the firepans, and the bowls, and such things as were of gold, in gold, and of silver, in silver, the captain of the guard took away.
2KGS|25|16|The two pillars, one sea, and the bases which Solomon had made for the house of the LORD; the brass of all these vessels was without weight.
2KGS|25|17|The height of the one pillar was eighteen cubits, and the chapiter upon it was brass: and the height of the chapiter three cubits; and the wreathed work, and pomegranates upon the chapiter round about, all of brass: and like unto these had the second pillar with wreathed work.
2KGS|25|18|And the captain of the guard took Seraiah the chief priest, and Zephaniah the second priest, and the three keepers of the door:
2KGS|25|19|And out of the city he took an officer that was set over the men of war, and five men of them that were in the king's presence, which were found in the city, and the principal scribe of the host, which mustered the people of the land, and threescore men of the people of the land that were found in the city:
2KGS|25|20|And Nebuzaradan captain of the guard took these, and brought them to the king of Babylon to Riblah:
2KGS|25|21|And the king of Babylon smote them, and slew them at Riblah in the land of Hamath. So Judah was carried away out of their land.
2KGS|25|22|And as for the people that remained in the land of Judah, whom Nebuchadnezzar king of Babylon had left, even over them he made Gedaliah the son of Ahikam, the son of Shaphan, ruler.
2KGS|25|23|And when all the captains of the armies, they and their men, heard that the king of Babylon had made Gedaliah governor, there came to Gedaliah to Mizpah, even Ishmael the son of Nethaniah, and Johanan the son of Careah, and Seraiah the son of Tanhumeth the Netophathite, and Jaazaniah the son of a Maachathite, they and their men.
2KGS|25|24|And Gedaliah sware to them, and to their men, and said unto them, Fear not to be the servants of the Chaldees: dwell in the land, and serve the king of Babylon; and it shall be well with you.
2KGS|25|25|But it came to pass in the seventh month, that Ishmael the son of Nethaniah, the son of Elishama, of the seed royal, came, and ten men with him, and smote Gedaliah, that he died, and the Jews and the Chaldees that were with him at Mizpah.
2KGS|25|26|And all the people, both small and great, and the captains of the armies, arose, and came to Egypt: for they were afraid of the Chaldees.
2KGS|25|27|And it came to pass in the seven and thirtieth year of the captivity of Jehoiachin king of Judah, in the twelfth month, on the seven and twentieth day of the month, that Evilmerodach king of Babylon in the year that he began to reign did lift up the head of Jehoiachin king of Judah out of prison;
2KGS|25|28|And he spake kindly to him, and set his throne above the throne of the kings that were with him in Babylon;
2KGS|25|29|And changed his prison garments: and he did eat bread continually before him all the days of his life.
2KGS|25|30|And his allowance was a continual allowance given him of the king, a daily rate for every day, all the days of his life.
