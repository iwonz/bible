2SAM|1|1|掃羅 死後， 大衛 擊殺 亞瑪力 人回來，在 洗革拉 住了兩天。
2SAM|1|2|第三天，看哪，有一人從 掃羅 的營裏出來，衣服撕裂，頭蒙灰塵，到 大衛 面前伏地叩拜。
2SAM|1|3|大衛 對他說：「你從哪裏來？」他說：「我從 以色列 的營裏逃來。」
2SAM|1|4|大衛 又對他說：「事情怎麼樣？請你告訴我。」他說：「士兵從陣上逃跑，也有許多士兵仆倒死亡， 掃羅 和他兒子 約拿單 也死了。」
2SAM|1|5|大衛 問報信的青年說：「你怎麼知道 掃羅 和他兒子 約拿單 死了呢？」
2SAM|1|6|報信的青年說：「我恰巧到 基利波山 ，看哪， 掃羅 靠在自己的槍上，看哪，有戰車、騎兵緊緊地追他。
2SAM|1|7|他回頭看見我，就呼叫我。我說：『我在這裏。』
2SAM|1|8|他問我說：『你是甚麼人？』我說：『我是 亞瑪力 人。』
2SAM|1|9|他對我說：『請你站到我這裏來，把我殺死，因為我非常痛苦，只剩下一口氣。』
2SAM|1|10|我就站到他那裏，殺了他，因為我知道他一倒下就活不了。然後，我把他頭上的冠冕和臂上的鐲子拿到我主這裏來。」
2SAM|1|11|大衛 就抓著自己的衣服，把衣服撕裂，所有跟隨他的人也都如此。
2SAM|1|12|他們為 掃羅 和他兒子 約拿單 ，以及耶和華的百姓和 以色列 家的人悲哀哭泣，禁食到晚上，因為他們都倒在刀下。
2SAM|1|13|大衛 問報信的青年說：「你是哪裏人？」他說：「我是一個寄居者的兒子，是 亞瑪力 人。」
2SAM|1|14|大衛 對他說：「你動手殺害耶和華的受膏者，怎麼不畏懼呢？」
2SAM|1|15|大衛 叫了一個僕人來，說：「來，殺了他！」僕人擊殺他，他就死了。
2SAM|1|16|大衛 對他說：「你的血歸到你自己頭上，因為你親口作證控訴自己，說：『我殺了耶和華的受膏者。』」
2SAM|1|17|大衛 作了這首哀歌，哀悼 掃羅 和他兒子 約拿單 ，
2SAM|1|18|並吩咐人把這首「弓歌」教導 猶大 人，看哪，它寫在《雅煞珥書》上：
2SAM|1|19|以色列 啊，尊榮者在你的高處被殺！ 大英雄竟然仆倒！
2SAM|1|20|不要在 迦特 報告， 不要在 亞實基倫 街上傳揚， 免得 非利士 的女子歡喜， 免得未受割禮之人的女子歡樂。
2SAM|1|21|基利波山 哪，願你那裏沒有雨，沒有露！ 願你的田地無土產可作供物！ 因為英雄的盾牌在那裏受辱， 掃羅 的盾牌沒有抹油。
2SAM|1|22|在被殺者的血前， 在勇士的脂肪前， 約拿單 的弓絕不退縮， 掃羅 的刀斷不虛回。
2SAM|1|23|掃羅 和 約拿單 生時相悅相愛， 死時也不分離。 他們比鷹更快， 比獅子還強。
2SAM|1|24|以色列 的女子啊，當為 掃羅 哭泣！ 他曾使你們穿朱紅色的美衣， 使你們衣服有黃金的妝飾。
2SAM|1|25|英雄竟然在陣上仆倒！ 約拿單 竟然在你的高處被殺！
2SAM|1|26|我兄 約拿單 哪，我為你悲傷！ 我甚喜愛你！ 你對我的愛何等奇妙， 過於婦女的愛情。
2SAM|1|27|英雄竟然仆倒！ 兵器竟然廢棄！
2SAM|2|1|此後， 大衛 求問耶和華說：「我可以上 猶大 的一個城去嗎？」耶和華對他說：「可以上去。」 大衛 說：「我上哪一個城去呢？」耶和華說：「 希伯崙 。」
2SAM|2|2|於是 大衛 和他的兩個妻子，一個是 耶斯列 人 亞希暖 ，一個是作過 迦密 人 拿八 妻子的 亞比該 ，都上那裏去了。
2SAM|2|3|大衛 也把跟隨他的人和他們各人的眷屬一同帶上去，住在 希伯崙 的城鎮中。
2SAM|2|4|猶大 人來，在那裏膏 大衛 作 猶大 家的王。 有人告訴 大衛 說：「埋葬 掃羅 的是 基列 的 雅比 人。」
2SAM|2|5|大衛 就派使者到 基列 的 雅比 人那裏，對他們說：「願耶和華賜福給你們！因為你們忠心對待你們的主 掃羅 ，埋葬了他。
2SAM|2|6|你們既做了這事，願耶和華以慈愛和信實待你們，我也要為此厚待你們。
2SAM|2|7|現在，你們的主 掃羅 死了， 猶大 家也已經膏我作他們的王，你們的手要堅強，要作英勇的人。」
2SAM|2|8|掃羅 軍隊的元帥， 尼珥 的兒子 押尼珥 ，曾將 掃羅 的兒子 伊施．波設 帶過河，到 瑪哈念 ，
2SAM|2|9|立他作王，治理 基列 、 亞書利 、 耶斯列 、 以法蓮 、 便雅憫 和 以色列 眾人。
2SAM|2|10|掃羅 的兒子 伊施．波設 登基的時候年四十歲，作 以色列 王二年，但是 猶大 家卻隨從 大衛 。
2SAM|2|11|大衛 在 希伯崙 作 猶大 家的王，共七年六個月。
2SAM|2|12|尼珥 的兒子 押尼珥 和 掃羅 的兒子 伊施．波設 的僕人從 瑪哈念 出來，往 基遍 去。
2SAM|2|13|洗魯雅 的兒子 約押 和 大衛 的僕人也出來，在 基遍 池旁與他們相遇；一隊坐在池的這邊，一隊坐在池的那邊。
2SAM|2|14|押尼珥 對 約押 說：「讓年輕人起來，在我們面前較量一下吧！」 約押 說：「讓他們起來吧。」
2SAM|2|15|他們就起來，點了人數過來：屬 掃羅 兒子 伊施．波設 的有 便雅憫 人十二名， 大衛 的僕人也有十二名。
2SAM|2|16|每人抓住對方的頭，用刀刺對方的肋旁，一同仆倒。所以，那地叫做 希利甲‧哈素林 ，就在 基遍 。
2SAM|2|17|那日戰況激烈， 押尼珥 和 以色列 人敗在 大衛 的僕人面前。
2SAM|2|18|在那裏有 洗魯雅 的三個兒子： 約押 、 亞比篩 、 亞撒黑 。 亞撒黑 的腳快如野地裏的羚羊；
2SAM|2|19|亞撒黑 追趕 押尼珥 ，直追趕他不偏左右。
2SAM|2|20|押尼珥 回頭說：「 亞撒黑 ，是你嗎？」他說：「是我。」
2SAM|2|21|押尼珥 對他說：「你轉左或轉右，去抓一個年輕人，剝去他的戰衣吧。」 亞撒黑 卻不肯轉開而不追趕他。
2SAM|2|22|押尼珥 又對 亞撒黑 說：「轉開，不要再追我了！我何必把你擊殺在地上呢？我若殺了你，怎麼有臉見你哥哥 約押 呢？」
2SAM|2|23|亞撒黑 仍不肯轉開， 押尼珥 就用回馬槍 刺入他的肚腹，甚至槍從背後穿出， 亞撒黑 就仆倒在那裏，當場死了。眾人趕到 亞撒黑 仆倒而死的地方，就都站住。
2SAM|2|24|約押 和 亞比篩 追趕 押尼珥 。日落的時候，他們到了通往 基遍 曠野的路旁， 基亞 對面的 亞瑪山 。
2SAM|2|25|便雅憫 人聚集在 押尼珥 後面，成為一隊，站在一座山頂上。
2SAM|2|26|押尼珥 呼叫 約押 說：「刀劍豈可永遠吞噬呢？你豈不知，結局必是痛苦的嗎？你要等到何時才叫百姓回去，不追趕他們的弟兄呢？」
2SAM|2|27|約押 說：「我指著永生的上帝起誓：你若沒有這麼說，百姓就必繼續追趕弟兄，直到早晨 。」
2SAM|2|28|於是 約押 吹角，眾百姓就站住，不再追趕 以色列 人，也不再打仗了。
2SAM|2|29|押尼珥 和他的人整夜行過 亞拉巴 。他們過了 約旦河 ，走過 畢倫 ，到了 瑪哈念 。
2SAM|2|30|約押 追趕 押尼珥 回來，聚集眾百姓， 大衛 的僕人中缺少了十九個人和 亞撒黑 。
2SAM|2|31|但 大衛 的僕人殺了 押尼珥 的人， 便雅憫 人三百六十名。
2SAM|2|32|他們把 亞撒黑 送到 伯利恆 ，葬在他父親的墳墓裏。 約押 和他的人走了一整夜，天亮的時候他們才到 希伯崙 。
2SAM|3|1|掃羅 家和 大衛 家爭戰許久。 大衛 家日見強盛， 掃羅 家卻日見衰弱。
2SAM|3|2|大衛 在 希伯崙 生了幾個兒子：長子 暗嫩 是 耶斯列 人 亞希暖 所生的；
2SAM|3|3|次子 基利押 是作過 迦密 人 拿八 的妻子 亞比該 所生的；三子 押沙龍 是 基述 王 達買 的女兒 瑪迦 所生的；
2SAM|3|4|四子 亞多尼雅 是 哈及 所生的；五子 示法提雅 是 亞比她 所生的；
2SAM|3|5|六子 以特念 是 大衛 的妻子 以格拉 所生的。 大衛 這六個兒子都是在 希伯崙 生的。
2SAM|3|6|掃羅 家和 大衛 家爭戰的時候， 押尼珥 在 掃羅 家大有權勢。
2SAM|3|7|掃羅 有一妃子，名叫 利斯巴 ，是 愛亞 的女兒。一日， 伊施．波設 對 押尼珥 說：「你為甚麼與我父的妃子同寢呢？」
2SAM|3|8|押尼珥 因 伊施．波設 的話非常生氣，說：「我豈是狗的頭，向著 猶大 呢？我今日忠心對待你父 掃羅 的家和他的弟兄、朋友，不將你交在 大衛 手裏，今日你竟為這婦人責備我嗎？
2SAM|3|9|願上帝重重懲罰 押尼珥 ！我要照著耶和華起誓應許 大衛 的話為他成就，
2SAM|3|10|廢去 掃羅 家的國度，建立 大衛 的王位，使他治理 以色列 和 猶大 ，從 但 直到 別是巴 。」
2SAM|3|11|伊施．波設 懼怕 押尼珥 ，一句話也不能回答。
2SAM|3|12|押尼珥 派使者到 大衛 所在的地方 ，說：「這地歸誰呢？」又說：「你與我立約，看哪，我必幫助你，使全 以色列 都擁護你。」
2SAM|3|13|大衛 說：「好！我與你立約。但有一件事我要求你，你來見我面的時候，除非把 掃羅 的女兒 米甲 帶來，就不必來見我的面了。」
2SAM|3|14|大衛 派使者到 掃羅 的兒子 伊施．波設 那裏，說：「你要把我的妻子 米甲 歸還我；她是我從前用一百 非利士 人的包皮所聘定的。」
2SAM|3|15|伊施．波設 就派人去，把 米甲 從 拉億 的兒子，她丈夫 帕鐵 那裏帶來。
2SAM|3|16|米甲 的丈夫跟著她，一面走一面哭，直跟到 巴戶琳 。 押尼珥 對他說：「你回去吧！」 帕鐵 就回去了。
2SAM|3|17|押尼珥 與 以色列 長老商議，說：「從前你們企盼 大衛 作王治理你們，
2SAM|3|18|現在你們可以這樣做了。因為耶和華曾論到 大衛 說：『我必藉我僕人 大衛 的手，救我民 以色列 脫離 非利士 人和眾仇敵的手。』」
2SAM|3|19|押尼珥 也說給 便雅憫 人聽。 押尼珥 又到 希伯崙 ，把 以色列 人和 便雅憫 全家所看為好的，說給 大衛 聽。
2SAM|3|20|押尼珥 帶著二十個人來到 希伯崙大衛 那裏， 大衛 就為 押尼珥 和他帶來的人擺設宴席。
2SAM|3|21|押尼珥 對 大衛 說：「我要起身去召集全 以色列 ，來到我主我王這裏，與你立約，你就可以照你的心願作王，統治一切。」於是 大衛 送走 押尼珥 ，他就平安地去了。
2SAM|3|22|看哪， 大衛 的僕人和 約押 突擊回來，帶回許多掠物。那時 押尼珥 不在 希伯崙大衛 那裏，因 大衛 已經送他走，他也平安地去了。
2SAM|3|23|約押 和跟隨他的全軍到了，有人告訴 約押 說：「 尼珥 的兒子 押尼珥 來到王這裏，王送走他，他也平安地去了。」
2SAM|3|24|約押 到王那裏，說：「你這是做甚麼呢？看哪， 押尼珥 來到你這裏，你為何送他走，讓他去了呢？
2SAM|3|25|你知道， 尼珥 的兒子 押尼珥 來，是要騙你，要打聽你的出入，知道你一切所行的事。」
2SAM|3|26|約押 從 大衛 那裏出來，派些使者去追 押尼珥 ，從 西拉井 那裏帶他回來， 大衛 卻不知道。
2SAM|3|27|押尼珥 回到 希伯崙 ， 約押 領他到城門中間，要與他私下交談，就在那裏刺穿了他的肚腹。他就死了，因為他流了 約押 兄弟 亞撒黑 的血。
2SAM|3|28|這事以後， 大衛 聽見了，說：「流 尼珥 兒子 押尼珥 的血，我和我的國在耶和華面前永遠是無辜的。
2SAM|3|29|願這血歸到 約押 頭上和他父的全家；又願 約押 家不斷有患漏症的，長痲瘋 的，架柺杖而行的 ，仆倒在刀下的，缺乏食物的。」
2SAM|3|30|約押 和他弟弟 亞比篩 殺了 押尼珥 ，是因為在 基遍 戰爭的時候， 押尼珥 殺了他們的弟弟 亞撒黑 。
2SAM|3|31|大衛 對 約押 和跟隨他的眾百姓說：「你們當撕裂衣服，腰束麻布，在 押尼珥 前面哀哭。」 大衛 王也跟在棺木後面。
2SAM|3|32|他們把 押尼珥 葬在 希伯崙 。王在 押尼珥 的墓旁放聲大哭，眾百姓也都哭了。
2SAM|3|33|王為 押尼珥 舉哀，說： 押尼珥 怎麼會像愚頑人一樣地死呢？
2SAM|3|34|你手未曾被捆綁，腳未曾被腳鐐鎖住。 你仆倒，如仆倒在兇惡之子手下一樣。 於是眾百姓又為 押尼珥 哀哭。
2SAM|3|35|白天的時候，眾百姓來勸 大衛 吃飯，但 大衛 起誓說：「我若在太陽未下山以前吃飯，或吃任何東西，願上帝重重懲罰我！」
2SAM|3|36|眾百姓知道了就看為好。凡王所做的，眾百姓都看為好。
2SAM|3|37|那日， 以色列 眾百姓才知道殺 尼珥 的兒子 押尼珥 並非出於王意。
2SAM|3|38|王對臣僕說：「你們豈不知今日在 以色列 中倒了一個作元帥的大人物嗎？
2SAM|3|39|我雖然受膏為王，今日還是軟弱。 洗魯雅 的兩個兒子，這些人比我強硬。願耶和華照著惡人所行的惡報應他。」
2SAM|4|1|掃羅 的兒子 伊施．波設 聽見 押尼珥 死在 希伯崙 ，手就發軟，全 以色列 也都驚惶。
2SAM|4|2|掃羅 的兒子 伊施．波設 有兩個軍官，一個叫 巴拿 ，第二個叫 利甲 ，都是 便雅憫 支派 比錄 人 臨門 的兒子；因為 比錄 也算是屬於 便雅憫 的。
2SAM|4|3|比錄 人先前逃到 基他音 ，在那裏寄居，直到今日。
2SAM|4|4|掃羅 的兒子 約拿單 有一個兒子，名叫 米非波設 ，是瘸腿的。 掃羅 和 約拿單 的消息從 耶斯列 傳來的時候，他才五歲。他的奶媽抱著他逃跑；因為跑得太急，孩子掉在地上，腿就瘸了。
2SAM|4|5|比錄 人 臨門 的兩個兒子 利甲 和 巴拿 出去，天正熱的時候到了 伊施．波設 的家。那時， 伊施．波設 在睡午覺。
2SAM|4|6|婦人進到房子中間，要取麥子。 利甲 和他的哥哥 巴拿 刺穿了 伊施．波設 的肚腹，然後逃跑了。
2SAM|4|7|他們進到房子的時候， 伊施．波設 正躺在臥房的床上，他們就把他殺死，割了他的首級，拿著首級在 亞拉巴 的路上走了一整夜。
2SAM|4|8|他們把 伊施．波設 的首級拿到 希伯崙 大衛 那裏，對王說：「王的仇敵 掃羅 曾尋索你的性命。看哪，這是他兒子 伊施．波設 的首級；耶和華今日為我主我王在 掃羅 和他後裔身上報了仇。」
2SAM|4|9|大衛 回答 比錄 人 臨門 的兒子 利甲 和他哥哥 巴拿 說：「我指著救我性命脫離一切苦難、永生的耶和華起誓：
2SAM|4|10|從前有人告訴我說：『看哪， 掃羅 死了。』他自以為報好消息，我就拿住他，把他殺在 洗革拉 ，作為他報消息的賞賜。
2SAM|4|11|更何況惡人把義人殺在他家的床上，我豈不從你們手中追討他的血，從地上除滅你們嗎？」
2SAM|4|12|於是 大衛 吩咐僕人把他們殺了，砍斷他們的手腳，掛在 希伯崙 的池旁。然後，他們把 伊施．波設 的首級葬在 希伯崙押尼珥 的墳墓裏。
2SAM|5|1|以色列 眾支派來到 希伯崙 見 大衛 ，說：「看哪，我們是你的骨肉。
2SAM|5|2|從前 掃羅 作我們王的時候，率領 以色列 人出入的是你。耶和華也曾對你說：『你必牧養我的百姓 以色列 ，你必作 以色列 的君王。』」
2SAM|5|3|於是 以色列 的眾長老都來到 希伯崙 見王 。 大衛 在 希伯崙 ，在耶和華面前與他們立約，他們就膏 大衛 作 以色列 的王。
2SAM|5|4|大衛 登基的時候年三十歲，作王四十年。
2SAM|5|5|他在 希伯崙 作 猶大 王七年六個月，在 耶路撒冷 作 以色列 和 猶大 王三十三年。
2SAM|5|6|王和他的人到了 耶路撒冷 ，要攻打住那地方的 耶布斯 人。 耶布斯 人對 大衛 說：「你必不能進到這裏，就是盲人、瘸子都可以把你擊退。」就是說：「 大衛 絕不能進到這裏。」
2SAM|5|7|然而 大衛 攻取了 錫安 的堡壘，就是 大衛 的城。
2SAM|5|8|當日， 大衛 說：「誰攻打 耶布斯 人，就要從水道上去，攻打我心裏所恨惡的 瘸子、盲人。」因此有人說：「盲人和瘸子不得進殿裏去。」
2SAM|5|9|大衛 住在堡壘裏，給它起名叫 大衛城 。 大衛 又從 米羅 往內，周圍建築。
2SAM|5|10|大衛 日見強大，耶和華－萬軍之上帝與他同在。
2SAM|5|11|推羅 王 希蘭 派使者把香柏木運到 大衛 那裏，又派木匠和石匠給 大衛 建造宮殿。
2SAM|5|12|大衛 知道耶和華堅立他作 以色列 王，又為自己百姓 以色列 的緣故，使他的國興盛。
2SAM|5|13|大衛 離開 希伯崙 之後，在 耶路撒冷 又立后妃，又生兒女。
2SAM|5|14|在 耶路撒冷 所生的孩子的名字是 沙母亞 、 朔罷 、 拿單 、 所羅門 、
2SAM|5|15|益轄 、 以利書亞 、 尼斐 、 雅非亞 、
2SAM|5|16|以利沙瑪 、 以利雅大 、 以利法列 。
2SAM|5|17|非利士 人聽見 大衛 受膏作 以色列 王， 非利士 眾人就上來尋索 大衛 。 大衛 聽見了，就下到堡壘去。
2SAM|5|18|非利士 人來了，散佈在 利乏音谷 。
2SAM|5|19|大衛 求問耶和華說：「我可以上去攻打 非利士 人嗎？你將他們交在我手裏嗎？」耶和華對 大衛 說：「你可以上去，我必將 非利士 人交在你手裏。」
2SAM|5|20|大衛 來到 巴力‧毗拉心 ，在那裏擊敗了 非利士 人。他說：「耶和華在我面前沖破敵人，如水沖破一樣。」因此他稱那地方為 巴力‧毗拉心 。
2SAM|5|21|非利士 人把偶像拋棄在那裏， 大衛 和他的人拿去了。
2SAM|5|22|非利士 人又上來，散佈在 利乏音谷 。
2SAM|5|23|大衛 求問耶和華；耶和華說：「不要直上，要繞到他們後頭，從桑樹林對面攻打他們。
2SAM|5|24|你聽見桑樹梢上有腳步的聲音，就要急速前去，因為那時耶和華已經出去，在你前頭攻打 非利士 人的軍隊了。」
2SAM|5|25|大衛 就遵照耶和華所吩咐的去做，攻打 非利士 人，從 迦巴 直到 基色 。
2SAM|6|1|大衛 又聚集 以色列 中所有挑選的人，共三萬名。
2SAM|6|2|大衛 起身，和跟隨他的眾百姓前往，要從 巴拉‧猶大 那裏將上帝的約櫃接上來；這約櫃是以坐在二基路伯上萬軍之耶和華的名所命名的。
2SAM|6|3|他們將上帝的約櫃從山岡上 亞比拿達 的家裏抬出來，放在新車上； 亞比拿達 的兒子 烏撒 和 亞希約 趕這新車。
2SAM|6|4|他們將上帝的約櫃從山岡上 亞比拿達 家裏抬出來 ， 亞希約 在約櫃前行走。
2SAM|6|5|大衛 和 以色列 全家在耶和華面前，隨著松木製造的各樣樂器 和琴、瑟、鼓、鈸、鑼跳舞。
2SAM|6|6|到了 拿艮 的禾場，因為牛失前蹄 ， 烏撒 就伸手扶住上帝的約櫃。
2SAM|6|7|耶和華的怒氣向 烏撒 發作；上帝因這冒犯在那裏擊打他，他就死在那裏，在上帝的約櫃旁。
2SAM|6|8|大衛 因耶和華突然衝出撞死 烏撒 就生氣，稱那地方為 毗列斯‧烏撒 ，直到今日。
2SAM|6|9|那日， 大衛 懼怕耶和華，說：「耶和華的約櫃怎可到我這裏來呢？」
2SAM|6|10|於是 大衛 不願將耶和華的約櫃接進 大衛城 他自己的地方，卻轉送到 迦特 人 俄別‧以東 的家中。
2SAM|6|11|耶和華的約櫃停在 迦特 人 俄別‧以東 家中三個月，耶和華賜福給 俄別‧以東 和他的全家。
2SAM|6|12|有人告訴 大衛 王說：「耶和華因約櫃的緣故賜福給 俄別‧以東 的家和一切屬他的。」 大衛 就去，歡歡喜喜地將上帝的約櫃從 俄別‧以東 家中接上來，到 大衛城 裏。
2SAM|6|13|抬耶和華約櫃的人走了六步， 大衛 就獻牛與肥畜為祭。
2SAM|6|14|大衛 穿著細麻布以弗得，在耶和華面前極力跳舞。
2SAM|6|15|這樣， 大衛 和 以色列 全家歡呼吹角，將耶和華的約櫃接了上來。
2SAM|6|16|耶和華的約櫃進 大衛城 的時候， 掃羅 的女兒 米甲 從窗戶裏往外觀看，見 大衛 王在耶和華面前踴躍跳舞，心裏就輕視他。
2SAM|6|17|眾人將耶和華的約櫃請進去，安放在所預備的地方，就是 大衛 為它搭的帳幕中。 大衛 在耶和華面前獻燔祭和平安祭。
2SAM|6|18|大衛 獻完了燔祭和平安祭，就奉萬軍之耶和華的名祝福百姓，
2SAM|6|19|並且分給 以色列 眾人，所有的百姓，無論男女，每人一個餅，一個棗子餅 ，一個葡萄餅。眾人就各自回家去了。
2SAM|6|20|大衛 回去要為家裏的人祝福， 掃羅 的女兒 米甲 出來迎接他，說：「 以色列 王今日有好大的榮耀啊！他今日在臣僕的使女眼前露體，如同一個無賴赤身露體一樣，」
2SAM|6|21|大衛 對 米甲 說：「這是在耶和華面前的。耶和華已揀選我，在你父和你父的全家之上，立我作耶和華百姓 以色列 的君王，所以我在耶和華面前跳舞，
2SAM|6|22|我也必更加卑微，自己看為低賤 。至於你所說的那些使女，她們反而尊重我。」
2SAM|6|23|掃羅 的女兒 米甲 ，直到死的那日沒有孩子。
2SAM|7|1|王住在自己宮中，耶和華使他平靜，不被四圍的仇敵擾亂。
2SAM|7|2|王對 拿單 先知說：「你看，我住在香柏木的宮中，上帝的約櫃卻停在幔子裏。」
2SAM|7|3|拿單 對王說：「你可以完全照你的心意去做，因為耶和華與你同在。」
2SAM|7|4|當夜耶和華的話臨到 拿單 ，說：
2SAM|7|5|「你去對我僕人 大衛 說：『耶和華如此說：你要建造殿宇給我居住嗎？
2SAM|7|6|自從我領 以色列 人從 埃及 上來，直到今日，我未曾住過殿宇，卻在會幕和帳幕中行走。
2SAM|7|7|凡我同 以色列 人所走的地方，我何曾向 以色列 任何一個領袖 ，就是我吩咐牧養我百姓 以色列 的，說過這話：你們為何不給我建造香柏木的殿宇呢？』
2SAM|7|8|現在，你要對我僕人 大衛這樣 說：『萬軍之耶和華如此說：我從羊圈中將你召來，叫你不再牧放羊群，立你作我百姓 以色列 的君王。
2SAM|7|9|你無論往哪裏去，我都與你同在，剪除你所有的仇敵。我必使你得大名，好像世上偉人的名一樣。
2SAM|7|10|我必為我百姓 以色列 選定一個地方，栽植他們，使他們住自己的地方，不再受攪擾；兇惡之子也不像從前那樣苦待他們，
2SAM|7|11|並不像我命令士師治理我百姓 以色列 的日子。我必使你平靜，不受任何仇敵攪擾，並且耶和華應許你，耶和華必為你建立家室。
2SAM|7|12|當你壽數滿足、與你祖先同睡的時候，我必使你身所生的後裔接續你；我也必堅定他的國。
2SAM|7|13|他必為我的名建造殿宇，我必堅定他國度的王位，直到永遠。
2SAM|7|14|我要作他的父，他要作我的子；他若犯了罪，我必用人的杖，用世人的鞭責罰他。
2SAM|7|15|但我的慈愛仍不離開他，像離開在你面前所廢的 掃羅 一樣。
2SAM|7|16|你的家和你的國必在你 面前永遠堅立，你的王位也必堅定，直到永遠。』」
2SAM|7|17|拿單 就按這一切話，照這一切異象告訴 大衛 。
2SAM|7|18|於是 大衛 王進去，坐在耶和華面前，說：「主耶和華啊，我是誰，我的家算甚麼，你竟帶領我到這地步呢？
2SAM|7|19|主耶和華啊，這在你眼中還看為小，你又說到你僕人的家將來的情況。主耶和華啊，這豈是人的常理嗎？
2SAM|7|20|大衛 還有甚麼可以對你說呢？主耶和華啊，你是知道你僕人的。
2SAM|7|21|你行這一切大事，使你的僕人明白，是因你應許的緣故，也照著你的心意。
2SAM|7|22|因此，主耶和華啊，你本為大；照我們耳中一切所聽見的，沒有可比你的，除你以外再沒有上帝。
2SAM|7|23|誰像你的百姓 以色列 呢？上帝親自去救贖世上的一國 ，作自己的子民，顯出他的大名；為了你的地，從列國和他們的神明中，在你親自從埃及贖出來的子民面前，為自己行了大而可畏的事 。
2SAM|7|24|你曾堅立你的百姓 以色列 作你的子民，直到永遠；你－耶和華也作他們的上帝。
2SAM|7|25|現在，耶和華上帝啊，你所應許僕人和僕人家的話，求你堅定，直到永遠；求你照你所說的而行。
2SAM|7|26|願人永遠尊你的名為大，說：『萬軍之耶和華是治理 以色列 的上帝。』這樣，你僕人 大衛 的家必在你面前堅立。
2SAM|7|27|萬軍之耶和華－ 以色列 的上帝啊，因你啟示你的僕人說：『我必為你建立家室』，所以僕人大膽向你如此祈禱。
2SAM|7|28|現在，主耶和華啊，惟有你是上帝！你的話是真實的，你也應許將這福氣賜給僕人。
2SAM|7|29|現在，求你賜福給你僕人的家，可以永存在你面前。主耶和華啊，因為這是你所應許的。願你的福分永遠賜給你僕人的家，使之蒙福！」
2SAM|8|1|此後， 大衛 攻打 非利士 人，制伏了他們。 大衛 從 非利士 人手中奪取了京城的治理權 。
2SAM|8|2|他又攻打 摩押 人，使他們躺臥在地上，用繩來量，量二繩的殺了，量一繩的活著。 摩押 人就臣服 大衛 ，向他進貢。
2SAM|8|3|利合 的兒子 瑣巴 王 哈大底謝 往 幼發拉底河 去，要奪回他的國權， 大衛 就攻打他，
2SAM|8|4|俘擄了他的騎兵一千七百人，步兵二萬人。 大衛 把所有戰馬的蹄筋砍斷，只留下一百輛戰車。
2SAM|8|5|大馬士革 的 亞蘭 人來幫助 瑣巴 王 哈大底謝 ， 大衛 殺了 亞蘭 人二萬二千。
2SAM|8|6|於是 大衛 在 大馬士革 的 亞蘭 設立軍營， 亞蘭 人就臣服 大衛 ，向他進貢。 大衛 無論往哪裏去，耶和華都使他得勝。
2SAM|8|7|大衛奪了 哈大底謝 臣僕擁有的金盾牌，帶到 耶路撒冷 。
2SAM|8|8|大衛 王又從 哈大底謝 的 比他 和 比羅他 二城奪取了許多的銅。
2SAM|8|9|哈馬 王 陀以 聽見 大衛 擊敗 哈大底謝 的全軍，
2SAM|8|10|就派他兒子 約蘭 到 大衛 王那裏，向他請安，為他祝福，因他與 哈大底謝 爭戰，並且擊敗了他；原來 哈大底謝 與 陀以 常常爭戰。 約蘭 手裏帶了金銀銅的器皿來。
2SAM|8|11|大衛 王把這些器皿分別為聖，連同他制伏各國所分別為聖的金銀，獻給耶和華，
2SAM|8|12|就是從 亞蘭 、 摩押 、 亞捫 人、 非利士 人、 亞瑪力 人，以及從 利合 的兒子 瑣巴 王 哈大底謝 所掠之物。
2SAM|8|13|大衛 得了名聲。當他回來的時候，在 鹽谷 擊殺了一萬八千 以東 人。
2SAM|8|14|大衛 在 以東 設立軍營；他在全 以東 設立軍營， 以東 人就都臣服他。 大衛 無論往哪裏去，耶和華都使他得勝。
2SAM|8|15|大衛 作全 以色列 的王，又向眾百姓秉公行義。
2SAM|8|16|洗魯雅 的兒子 約押 作元帥； 亞希律 的兒子 約沙法 作史官；
2SAM|8|17|亞希突 的兒子 撒督 和 亞比亞他 的兒子 亞希米勒 作祭司； 西萊雅 作書記；
2SAM|8|18|耶何耶大 的兒子 比拿雅 管轄 基利提 人和 比利提 人。 大衛 的眾子都作祭司。
2SAM|9|1|大衛 說：「 掃羅 家還有剩下的人沒有？我要因 約拿單 的緣故向他施恩。」
2SAM|9|2|掃羅 家有一個僕人名叫 洗巴 ，有人叫他來到 大衛 那裏。王對他說：「你是 洗巴 嗎？」他說：「僕人是。」
2SAM|9|3|王說：「 掃羅 家還有沒有剩下的人？我要照上帝的慈愛恩待他。」 洗巴 對王說：「還有 約拿單 的一個兒子，雙腿是瘸的。」
2SAM|9|4|王對他說：「他在哪裏？」 洗巴 對王說：「看哪，他在 羅‧底巴 ， 亞米利 的兒子 瑪吉 家裏。」
2SAM|9|5|於是 大衛 王派人去，從 羅‧底巴 ， 亞米利 的兒子 瑪吉 家裏召了他來。
2SAM|9|6|掃羅 的孫子， 約拿單 的兒子 米非波設 來到 大衛 那裏，臉伏於地叩拜。 大衛 說：「 米非波設 ！」 米非波設 說：「看哪，僕人在此。」
2SAM|9|7|大衛 對他說：「你不要懼怕，我必因你父親 約拿單 的緣故向你施恩，把你祖父 掃羅 的一切田地都歸還你，你也可以常與我同席吃飯。」
2SAM|9|8|米非波設 叩拜，說：「你的僕人算甚麼，不過如死狗一般，竟蒙你這樣眷顧！」
2SAM|9|9|王召了 掃羅 的僕人 洗巴 來，對他說：「我已把屬 掃羅 和他的一切家產都賜給你主人的兒子了。
2SAM|9|10|你，你的眾子和僕人要為你主人的兒子耕種田地，把所收穫的拿來供他食用；你主人的兒子 米非波設 卻要常與我同席吃飯。」 洗巴 有十五個兒子和二十個僕人。
2SAM|9|11|洗巴 對王說：「凡我主我王吩咐僕人的，僕人都必遵行。」於是 米非波設 與王 同席吃飯，如王的兒子一樣。
2SAM|9|12|米非波設 有一個小兒子，名叫 米迦 。凡住在 洗巴 家裏的人都作了 米非波設 的僕人。
2SAM|9|13|米非波設 住在 耶路撒冷 ，常與王同席吃飯。他兩腿都是瘸的。
2SAM|10|1|此後， 亞捫 人的王死了，他兒子 哈嫩 接續他作王。
2SAM|10|2|大衛 說：「 哈嫩 的父親 拿轄 怎樣向我施恩，我也要怎樣向 哈嫩 施恩。」於是 大衛 派臣僕為他的父親安慰他。當 大衛 的臣僕到了 亞捫 人的境內，
2SAM|10|3|亞捫 人的領袖對他們的主 哈嫩 說：「 大衛 派人來安慰你，你看他是要尊敬你父親嗎？ 大衛 派臣僕到你這裏，不是為了要窺探偵察，而傾覆這城嗎？」
2SAM|10|4|哈嫩 就抓住 大衛 的臣僕，把他們的鬍鬚剃去一半，又割斷他們下半截的袍子，露出下體，然後放了他們。
2SAM|10|5|有人告訴 大衛 ，他就派人去迎接他們，因為這些人覺得很羞恥。王說：「可以住在 耶利哥 ，等到鬍鬚長出來再回來。」
2SAM|10|6|亞捫 人看到 大衛 憎惡他們，就派人去雇用 伯‧利合 的 亞蘭 人和 瑣巴 的 亞蘭 人，步兵二萬，以及 瑪迦 王的人一千、 陀伯 人一萬二千。
2SAM|10|7|大衛 聽見了，就派 約押 和所有勇猛的軍隊出去。
2SAM|10|8|亞捫 人出來，在城門前擺陣； 瑣巴 與 利合 的 亞蘭 人、 陀伯 人，以及 瑪迦 人另外在郊野擺陣。
2SAM|10|9|約押 看見戰陣對著他前後擺列，就把從 以色列 所有精兵中挑選出來的，擺陣迎戰 亞蘭 人。
2SAM|10|10|他把其餘的兵交在他兄弟 亞比篩 手裏， 亞比篩 就擺陣迎戰 亞捫 人。
2SAM|10|11|約押 對 亞比篩說：「 亞蘭 人若強過我，你就來幫助我； 亞捫 人若強過你，我就去幫助你。
2SAM|10|12|你要剛強，我們要為自己的百姓，為我們上帝的城鎮奮勇。願耶和華照他所看為好的去做！」
2SAM|10|13|於是， 約押 和跟隨他的士兵前進攻打 亞蘭 人； 亞蘭 人在他面前逃跑。
2SAM|10|14|亞捫 人見 亞蘭 人逃跑，他們也在 亞比篩 面前逃跑進城。 約押 就離開 亞捫 人，回 耶路撒冷 去了。
2SAM|10|15|亞蘭 人見自己被 以色列 打敗，就集合起來。
2SAM|10|16|哈大底謝 派人去，把 大河 那邊的 亞蘭 人調來；他們到了 希蘭 ，由 哈大底謝 的將軍 朔法 在他們前面率領。
2SAM|10|17|有人告訴 大衛 ，他就聚集 以色列 眾人過 約旦河 ，來到 希蘭 。 亞蘭 人迎著 大衛 擺陣，與他打仗。
2SAM|10|18|亞蘭 人在 以色列 人面前逃跑。 大衛 殺了 亞蘭 七百輛戰車的士兵，四萬騎兵 ，又擊殺 亞蘭 的將軍 朔法 ，他就死在那裏。
2SAM|10|19|哈大底謝 屬下的諸王見自己被 以色列 打敗，就與 以色列 講和，臣服他們。於是 亞蘭 人害怕，不再幫助 亞捫 人了。
2SAM|11|1|過了一年，正是諸王出戰的時候， 大衛 派 約押 率領臣僕和 以色列 眾人出去。他們打敗 亞捫 人，圍攻 拉巴 。 大衛 仍然留在 耶路撒冷 。
2SAM|11|2|黃昏的時候， 大衛 從床上起來，在王宮的平頂上散步。他從平頂上看見一個婦人沐浴，這婦人容貌非常美麗。
2SAM|11|3|大衛 派人打聽那婦人是誰。有人說：「她不是 以連 的女兒， 赫 人 烏利亞 的妻子 拔示巴 嗎？」
2SAM|11|4|大衛 派使者去把婦人接來；她來到大衛那裏，那時她的月經剛潔淨， 大衛 與她同寢。她就回家去了。
2SAM|11|5|那婦人懷了孕，派人去告訴 大衛 說：「我懷孕了。」
2SAM|11|6|大衛 派人告訴 約押 ：「你派 赫 人 烏利亞 到我這裏來。」 約押 就派 烏利亞 到 大衛 那裏。
2SAM|11|7|烏利亞 來到 大衛那裏， 大衛 問 約押 好，也問士兵好，又問戰爭的情況。
2SAM|11|8|大衛 對 烏利亞 說：「下到你家去，洗洗腳吧！」 烏利亞 出了王宮，隨後王送他一份禮物。
2SAM|11|9|烏利亞 卻和他主人所有的僕人一同睡在王宮門口，沒有下到他家去。
2SAM|11|10|有人告訴 大衛 說：「 烏利亞 沒有下到他的家。」 大衛 就對 烏利亞 說：「你不是從遠路上來嗎？為甚麼不下到你家去呢？」
2SAM|11|11|烏利亞 對 大衛 說：「約櫃， 以色列 和 猶大 都留在棚裏，我主 約押 和我主的僕人都在田野安營，我豈可回家吃喝，與妻子同房呢？我指著王和王的性命起誓：『我絕不做這事！』」
2SAM|11|12|大衛 對 烏利亞 說：「你今日仍留在這裏，明日我打發你去。」於是 烏利亞 那日留在 耶路撒冷 。次日，
2SAM|11|13|大衛 召了 烏利亞 來，叫他在自己面前吃喝，使他喝醉。黃昏的時候， 烏利亞 出去，躺臥在自己的床上；與他主的僕人在一起，並沒有下到他的家去。
2SAM|11|14|早晨， 大衛 寫信給 約押 ，交 烏利亞 親手帶去。
2SAM|11|15|他在信內寫著說：「要派 烏利亞 到戰爭激烈的前線去，然後你們撤退離開他，使他被擊殺而死。」
2SAM|11|16|約押 偵察城的時候，知道敵人哪裏有勇士，就派 烏利亞 到那地方。
2SAM|11|17|城裏的人出來和 約押 打仗， 大衛 的僕人中有幾個士兵被殺， 赫 人 烏利亞 也死了。
2SAM|11|18|於是， 約押 派人去將戰爭的一切事奏告 大衛 ，
2SAM|11|19|又吩咐使者說：「你把戰爭的一切事對王說完了，
2SAM|11|20|王若發怒，對你說：『你們打仗為甚麼挨近城呢？豈不知敵人會從城牆上射箭嗎？
2SAM|11|21|從前擊殺 耶路比設 的兒子 亞比米勒 的是誰呢？豈不是一個婦人從城牆上拋下一塊上磨石來，打在他身上，他就死在 提備斯 嗎？你們為甚麼挨近城牆呢？』你就說：『你的僕人 赫 人 烏利亞 也死了。』」
2SAM|11|22|使者就去，照著 約押 所吩咐的一切話來奏告 大衛 。
2SAM|11|23|使者對 大衛 說：「敵人強過我們，出到郊外攻打我們，我們把他們趕回到城門口。
2SAM|11|24|弓箭手從城牆上射你的僕人，射死幾個王的僕人，你的僕人 赫 人 烏利亞 也死了。」
2SAM|11|25|大衛 向使者說：「你對 約押 這樣說：『不要為這事難過，因為刀劍可能吞滅這人或那人。你只管竭力攻城，將城傾覆。』你要勉勵 約押 。」
2SAM|11|26|烏利亞 的妻聽見丈夫 烏利亞 死了，就為丈夫哀哭。
2SAM|11|27|居喪的日子過了， 大衛 派人把她接到宮裏，她就作了 大衛 的妻子，給 大衛 生了一個兒子。但 大衛 做的這事，耶和華的眼中看為惡。
2SAM|12|1|耶和華差遣 拿單 到 大衛 那裏。 拿單 到了他那裏，對他說：「在一座城裏有兩個人，一個是富翁，一個是窮人。
2SAM|12|2|富翁有極多的牛群羊群；
2SAM|12|3|窮人除了所買來養活的一隻小母羊之外，一無所有。小羊在他家裏和他兒女一同長大，吃他所吃的，喝他所喝的，睡在他懷中，在他看來如同女兒一樣。
2SAM|12|4|有一客人來到這富翁那裏，富翁捨不得從自己的牛群羊群中取一隻招待來到他那裏的旅客，卻取了窮人的小母羊，招待來到他那裏的人。」
2SAM|12|5|大衛 就非常惱怒那人，對 拿單 說：「我指著永生的耶和華起誓，做這事的人該死！
2SAM|12|6|他必須償還小母羊四倍，因為他做這事，沒有憐憫的心。」
2SAM|12|7|拿單 對 大衛 說：「你就是那人！耶和華－ 以色列 的上帝如此說：『我膏你作 以色列 的王，我救你脫離 掃羅 的手；
2SAM|12|8|我將你主人的家業賜給你，將你主人的妃嬪交在你懷裏，又將 以色列 和 猶大 家賜給你；若還嫌少，我也會如此這般加倍賜給你。
2SAM|12|9|你為甚麼藐視耶和華的命令，做他眼中看為惡的事呢？你用刀擊殺 赫 人 烏利亞 ，又娶了他的妻子為妻，借 亞捫 人的刀殺死他。
2SAM|12|10|現在刀劍必永不離開你的家，因你藐視我，娶了 赫 人 烏利亞 的妻子為妻。』
2SAM|12|11|耶和華如此說：『看哪，我必從你家中興起災禍攻擊你；我必在你眼前把你的妃嬪賜給你身邊的人，他要在光天化日下與你的妃嬪同寢。
2SAM|12|12|你在暗中做那事，我卻要在 以色列 眾人面前，在日光之下做這事。』」
2SAM|12|13|大衛 對 拿單 說：「我得罪耶和華了！」 拿單 說：「耶和華已經除去你的罪，你必不至於死。
2SAM|12|14|只是在這事上，你大大藐視耶和華 ，因此，你生的孩子必定要死。」
2SAM|12|15|拿單 就回家去了。 耶和華擊打 烏利亞 的妻子為 大衛 生的孩子，他就得了重病。
2SAM|12|16|大衛 為這孩子懇求上帝。 大衛 刻苦禁食，到裏面去，躺在地上過夜。
2SAM|12|17|他家中的老臣來到他旁邊，要把他從地上扶起來，他卻不肯，也不同他們吃飯。
2SAM|12|18|到第七日，孩子死了。 大衛 的臣僕不敢告訴他孩子死了，因他們說：「看哪，孩子還活著的時候，我們勸他，他尚且不聽我們的話，我們怎麼能告訴他孩子死了，讓他做出不好的事呢？」
2SAM|12|19|大衛 見臣僕彼此低聲說話，就知道孩子死了。他問臣僕說：「孩子死了嗎？」他們說：「死了。」
2SAM|12|20|大衛 就從地上起來，沐浴，抹膏，換了衣服，進耶和華的殿敬拜。然後他回宮，吩咐人為他擺飯，他就吃了。
2SAM|12|21|臣僕對他說：「你所做的是甚麼事呢？孩子活著的時候，你為他禁食哭泣；孩子死了，你卻起來吃飯。」
2SAM|12|22|大衛 說：「孩子還活著，我禁食哭泣，因為我想，或許耶和華憐憫我，會讓孩子活下來。
2SAM|12|23|現在孩子死了，我何必禁食呢？我能使他回來嗎？我必往他那裏去，他卻不能回到我這裏來。」
2SAM|12|24|大衛 安慰他的妻子 拔示巴 ，與她同房，她就生了兒子，給他起名叫 所羅門 。耶和華喜愛他，
2SAM|12|25|就藉 拿單 先知賜他一個名字，叫 耶底底亞 ；這是為了耶和華的緣故。
2SAM|12|26|約押 攻打 亞捫 人的 拉巴 ，攻佔了京城。
2SAM|12|27|約押 派使者到 大衛 那裏，說：「我攻打 拉巴 ， 也攻佔了水城。
2SAM|12|28|現在你要召集其餘的軍兵，安營圍攻這城，攻佔它，免得我攻佔這城，人就以我的名叫這城。」
2SAM|12|29|於是 大衛 召集全軍，往 拉巴 去攻城，就攻佔了它。
2SAM|12|30|他也奪了 米勒公 頭上所戴的冠冕，其上的金子重一他連得，又嵌著寶石。這冠冕就戴在 大衛 頭上。 大衛 又從城裏奪了許多財物，
2SAM|12|31|把城裏的百姓拉出來，叫他們用鋸，用鐵耙，用鐵斧做工，派他們在磚窯中服役； 大衛 待 亞捫 各城的居民都是如此。於是， 大衛 和全軍都回 耶路撒冷 去了。
2SAM|13|1|後來發生了一件事。 大衛 的兒子 押沙龍 有一個美貌的妹妹，名叫 她瑪 。 大衛 的兒子 暗嫩 愛上了她。
2SAM|13|2|暗嫩 為他妹妹 她瑪 苦戀成疾，因為 她瑪 還是處女， 暗嫩 眼看難以向她行事。
2SAM|13|3|暗嫩 有一個密友，名叫 約拿達 ，是 大衛 長兄 示米亞 的兒子。這 約拿達 為人極其狡猾。
2SAM|13|4|他對 暗嫩 說：「王的兒子啊，你何不告訴我，為何你一天比一天憔悴呢？」 暗嫩 對他說：「我愛上了我兄弟 押沙龍 的妹妹 她瑪 。」
2SAM|13|5|約拿達 對他說：「你躺在床上裝病，等你父親來看你，就對他說：『請讓我妹妹 她瑪 來，給我東西吃，在我眼前預備食物，使我可以看見，好從她手裏接過來吃。』」
2SAM|13|6|於是 暗嫩 躺著裝病，王來看他。 暗嫩 對王說：「請讓我妹妹 她瑪 來，在我眼前為我做兩個餅，我好從她手裏接過來吃。」
2SAM|13|7|大衛 就派人去宮裏，到 她瑪 那裏，說：「你到你哥哥 暗嫩 的屋裏去，為他預備食物。」
2SAM|13|8|她瑪 就到她哥哥 暗嫩 的屋裏，那時 暗嫩 正躺著。 她瑪 拿了麵團揉麵，在他眼前做餅，把餅烤熟了。
2SAM|13|9|她瑪 拿了鍋子，在他面前把餅倒出來，他卻不肯吃。 暗嫩 說：「每一個人都離開我，出去吧！」眾人就都離開他，出去了。
2SAM|13|10|暗嫩 對 她瑪 說：「你把食物拿進臥房，我好從你手裏接過來吃。」 她瑪 就把所做的餅拿進臥房，到她哥哥 暗嫩 那裏。
2SAM|13|11|她瑪 上前去給他吃，他就拉住 她瑪 ，對她說：「我妹妹，你來與我同寢。」
2SAM|13|12|她瑪 對他說：「哥哥，不可以！不要玷辱我！ 以色列 中不可以這樣做，你不要做這醜事！
2SAM|13|13|我蒙受恥辱，該往那裏去呢？至於你，你在 以色列 中也成了一個愚頑人。現在你可以求王，他必不禁止我歸你。」
2SAM|13|14|但 暗嫩 不肯聽她的話，因他比她更有力，就玷辱她，與她同寢。
2SAM|13|15|隨後， 暗嫩 極其恨她，恨她的心比先前愛她的心更甚，就對她說：「你起來，去吧！」
2SAM|13|16|她瑪 對 暗嫩 說：「不要這樣！你趕我出去的這惡比你剛才向我所做的更嚴重！」但 暗嫩 不肯聽她，
2SAM|13|17|就叫伺候自己的僕人來，說：「把這女子從我這裏趕出去！她一出去，你就閂上門。」
2SAM|13|18|那時 她瑪 穿著彩衣，因為沒有出嫁的公主都穿這樣的外袍。 暗嫩 的僕人把她趕出去，她一出去，僕人就閂上門。
2SAM|13|19|她瑪 把灰塵撒在頭上，撕裂所穿的彩衣，以手抱頭，一面走一面哭喊。
2SAM|13|20|她胞兄 押沙龍 對她說：「你哥哥 暗嫩 與你親近了嗎？妹妹，現在暫且不要作聲，他是你的哥哥，不要把這事放在心上。」 她瑪 就孤孤單單地住在她胞兄 押沙龍 的家裏。
2SAM|13|21|大衛 王聽見這一切的事，就非常憤怒。
2SAM|13|22|押沙龍 卻不和 暗嫩 說好說歹；因為 暗嫩 玷辱他妹妹 她瑪 ，所以 押沙龍 恨惡他。
2SAM|13|23|過了二年，有人在靠近 以法蓮 的 巴力‧夏瑣 為 押沙龍 剪羊毛。 押沙龍 請了王所有的兒子來。
2SAM|13|24|押沙龍 來到王那裏，說：「看哪，有人正為你的僕人剪羊毛，請王和王的臣僕與你的僕人同去。」
2SAM|13|25|王對 押沙龍 說：「不，我兒，我們不必都去，免得成了你的負擔。」 押沙龍 再三請王，王仍是不肯去，只為他祝福。
2SAM|13|26|押沙龍 說：「王若不去，請讓我哥哥 暗嫩 與我們同去。」王對他說：「為何要他與你同去呢？」
2SAM|13|27|押沙龍 再三求王，王就派 暗嫩 和王所有的兒子與他同去。
2SAM|13|28|押沙龍 吩咐僕人說：「你們注意， 暗嫩 開懷暢飲的時候，我對你們說擊殺 暗嫩 ，你們就殺他。不要懼怕，這不是我吩咐你們的嗎？你們要剛強，作勇士！」
2SAM|13|29|押沙龍 的僕人就照 押沙龍 所吩咐的，向 暗嫩 行了。王所有的兒子都起來，各人騎上騾子逃跑了。
2SAM|13|30|他們還在路上，就有風聲傳到 大衛 那裏，說：「 押沙龍 擊殺了王所有的兒子，沒有留下一個。」
2SAM|13|31|王就起來，撕裂衣服，躺在地上。王的臣僕全都撕裂衣服，站在旁邊。
2SAM|13|32|大衛 的長兄 示米亞 的兒子 約拿達 說：「我主，不要以為他們把所有的年輕人，就是王的兒子都殺了，只有 暗嫩 一個人死了。自從 暗嫩 玷辱了 押沙龍 的妹妹 她瑪 那日， 押沙龍 已經決定這事了。
2SAM|13|33|現在，我主我王，不要把這事放在心上，以為王所有的兒子都死了。其實，只有 暗嫩 一人死了。」
2SAM|13|34|押沙龍 逃跑了。守望的年輕人舉目觀看，看哪，有許多人從 何羅念 山坡的路上來。
2SAM|13|35|約拿達 對王說：「看哪，王的兒子都來了，正如你僕人所說的，事情就這樣發生了。」
2SAM|13|36|話剛說完，看哪，王的兒子都到了，放聲大哭。王和他的眾臣僕也都號咷痛哭。
2SAM|13|37|押沙龍 逃到 亞米忽 的兒子 基述 王 達買 那裏去了。 大衛 天天為他兒子悲哀。
2SAM|13|38|押沙龍 逃到 基述 去了，在那裏住了三年。
2SAM|13|39|王想要出去對付 押沙龍 的心化解了 ，因為王對 暗嫩 之死這事已經得了安慰。
2SAM|14|1|洗魯雅 的兒子 約押 知道王心裏想念 押沙龍 。
2SAM|14|2|他派人往 提哥亞 去，從那裏叫了一個有智慧的婦人來，對她說：「請你裝作居喪的人，穿上喪服，不用膏抹身，裝作為死者悲哀多日的婦人。
2SAM|14|3|你到王那裏，對王如此如此說。」於是 約押 把當說的話放在她口中。
2SAM|14|4|提哥亞 婦人到王面前 ，臉伏於地叩拜，說：「王啊，求你拯救！」
2SAM|14|5|王對她說：「你有甚麼事呢？」她說：「我實在是個寡婦，我丈夫死了。
2SAM|14|6|婢女有兩個兒子，二人在田間打架，沒有人從中勸解，一個擊殺另一個，把他打死了。
2SAM|14|7|看哪，全家族都起來攻擊婢女，說：『把那打死兄弟的交出來，我們好處死他，為他所打死的兄弟償命，滅絕那承受家業的。』這樣，他們要把我剩下的炭火滅盡，不給我丈夫留名或留後在地面上。」
2SAM|14|8|王對婦人說：「你回家去吧！我必為你下個命令。」
2SAM|14|9|提哥亞 婦人又對王說：「我主我王，願這罪孽歸我和我的父家，與王和王的位無關。」
2SAM|14|10|王說：「有人說話難為你，你就帶他到我這裏來，他必不再攪擾你。」
2SAM|14|11|婦人說：「願王對耶和華－你的上帝發誓，不許報血仇的人施行毀滅，免得他們滅絕我的兒子。」王說：「我指著永生的耶和華起誓：你的兒子連一根頭髮也不致落在地上。」
2SAM|14|12|婦人說：「求我主我王容許婢女再說一句話。」王說：「你說吧！」
2SAM|14|13|婦人說：「王為何起意做這事，要害上帝的百姓呢？王不使那逃亡的人回來，王說這話就證實自己錯了！
2SAM|14|14|我們都必死，如同水潑在地上，不能收回。上帝不會讓人不死，但仍設法 使逃亡的人不致成為趕出、回不來的人。
2SAM|14|15|現在我來將這話告訴我主我王，是因百姓使我懼怕。婢女想：『不如告訴王，或者王會成就使女所求的。
2SAM|14|16|人要把我和我兒子從上帝的地業上一同除滅，王必應允救使女脫離他的手。』
2SAM|14|17|婢女想：『我主我王的話必安慰我』；因為我主我王能辨別是非，如同上帝的使者一樣。惟願耶和華－你的上帝與你同在！」
2SAM|14|18|王回答婦人說：「我問你一句話，你一點也不可瞞我。」婦人說：「我主我王，請說。」
2SAM|14|19|王說：「這一切莫非是 約押 的手指使你的嗎？」婦人回答說：「我敢在我主我王面前起誓：我主我王所說的一切不偏左右，這是王的僕人 約押 吩咐我的，這一切話是他放在婢女口中的。
2SAM|14|20|王的僕人 約押 做這事，為要扭轉局面。我主的智慧卻如上帝使者的智慧，能知地上一切的事。」
2SAM|14|21|王對 約押 說：「看哪，我應允這事。你去，把那年輕人 押沙龍 帶回來。」
2SAM|14|22|約押 臉伏於地叩拜，為王祝福，說：「王既應允僕人這件事，僕人今日知道在我主我王眼前蒙恩寵了。」
2SAM|14|23|於是 約押 起身往 基述 去，把 押沙龍 帶回 耶路撒冷 。
2SAM|14|24|王說：「讓他回自己的家去，不要來見我的面。」 押沙龍 就回自己的家去，沒有見王的面。
2SAM|14|25|全 以色列 中，無人像 押沙龍 那樣俊美，得人稱讚，從腳底到頭頂毫無瑕疵。
2SAM|14|26|他的頭髮很重，每到年底剪髮一次，所剪下來的，按王的秤稱一稱，重二百舍客勒。
2SAM|14|27|押沙龍 生了三個兒子，一個女兒。女兒名叫 她瑪 ，是個容貌美麗的女子。
2SAM|14|28|押沙龍 住在 耶路撒冷 ，足足有二年沒有見王的面。
2SAM|14|29|押沙龍 派人去叫 約押 來，要託他到王那裏去， 約押 卻不肯來。 押沙龍 第二次派人去叫他，他仍不肯來。
2SAM|14|30|於是 押沙龍 對僕人說：「你們看， 約押 有一塊田靠近我的田，其中有大麥，你們去放火把它燒了。」 押沙龍 的僕人就去放火燒了那田。
2SAM|14|31|於是 約押 起來，到了 押沙龍 家裏，對他說：「你的僕人為何放火燒我的田呢？」
2SAM|14|32|押沙龍 對 約押 說：「看哪，我派人去請你來，好託你到王那裏去，說：『我為何從 基述 回來呢？我仍在那裏比較好。』現在讓我去見王的面；我若有罪孽，就任憑王殺了我吧。」
2SAM|14|33|於是 約押 到王那裏，奏告王，王就叫 押沙龍 來。 押沙龍 到王那裏，在王面前臉伏於地，王就親吻 押沙龍 。
2SAM|15|1|此後， 押沙龍 為自己預備車馬，又派五十人在他前頭奔跑。
2SAM|15|2|押沙龍 常常早晨起來，站在城門的路旁，任何人有爭訟要去求王判決， 押沙龍 就叫他過來，說：「你是哪一城的人？」他說：「僕人是 以色列 某支派的人。」
2SAM|15|3|押沙龍 就對他說：「看，你的案件合情合理，無奈王沒有委派人聽你申訴。」
2SAM|15|4|押沙龍 又說：「恨不得我作這地的審判官！ 凡有爭訟的人可以到我這裏來，我必秉公判斷。」
2SAM|15|5|若有人近前來要拜 押沙龍 ， 押沙龍 就伸手拉住他，親吻他。
2SAM|15|6|以色列 中，凡到王那裏求判決的， 押沙龍 都這麼做。這樣， 押沙龍 暗中贏得了 以色列 人的心。
2SAM|15|7|過了四年 ， 押沙龍 對王說：「求你准我往 希伯崙 去，還我向耶和華所許的願。
2SAM|15|8|因為僕人住在 亞蘭 的 基述 時，曾許願說：『耶和華若使我再回 耶路撒冷 ，我必事奉他 。』」
2SAM|15|9|王對他說：「你平安地去吧！」 押沙龍 就動身，往 希伯崙 去了。
2SAM|15|10|押沙龍 派密使走遍 以色列 各支派，說：「你們一聽見角聲就說：『 押沙龍 在 希伯崙 作王了！』」
2SAM|15|11|押沙龍 在 耶路撒冷 請了二百人與他同去，都是誠心誠意去的，一點也不知道實情。
2SAM|15|12|押沙龍 獻祭的時候，派人去把 大衛 的謀士， 基羅 人 亞希多弗 從他本城 基羅 請來 。於是叛亂越發強大，因為隨從 押沙龍 的百姓日漸增多。
2SAM|15|13|報信的人來到 大衛 那裏，說：「 以色列 人的心都歸向 押沙龍 了！」
2SAM|15|14|大衛 就對 耶路撒冷 所有跟隨他的臣僕說：「起來，我們逃吧！否則，我們來不及逃避 押沙龍 。要快點離開，免得他很快追上我們，加害於我們，用刀擊殺城裏的人。」
2SAM|15|15|王的臣僕對王說：「我主我王所決定的一切，看哪，僕人都願遵行。」
2SAM|15|16|於是王出去了，他的全家都跟隨他，但留下十個妃嬪看守宮殿。
2SAM|15|17|王出去，眾百姓都跟隨他；到了最後一座屋子 ，他們就停下來。
2SAM|15|18|王的眾臣僕都在他旁邊過去。 基利提 人、 比利提 人，和從 迦特 跟隨王來的六百個 迦特 人，也都在王面前過去。
2SAM|15|19|王對 迦特 人 以太 說：「你是外邦人，從你本地逃來的，為甚麼與我們同去呢？你回去留在新王那裏吧！
2SAM|15|20|你昨天才到，我今日怎好叫你與我們一同流亡，而我卻要到處飄流呢？回去吧，你帶你的弟兄回去吧！願主用慈愛信實待你 。」
2SAM|15|21|以太 回答王說：「我指著永生的耶和華起誓，又敢在王面前起誓：無論生死，王在哪裏，你的僕人也必在哪裏。」
2SAM|15|22|大衛 對 以太 說：「去，過去吧！」於是 迦特 人 以太 帶著所有跟隨他的人和孩子過去了。
2SAM|15|23|眾百姓過去時，當地的人全都放聲大哭。王過了 汲淪溪 ，眾百姓就往曠野的路上去了。
2SAM|15|24|看哪， 撒督 和所有抬上帝約櫃的 利未 人也一同來了。他們將上帝的約櫃放下， 亞比亞他 上來 ，直到眾百姓從城裏出來走過去為止。
2SAM|15|25|王對 撒督 說：「你將上帝的約櫃請回城去。我若在耶和華眼前蒙恩，他必使我回來，再見到約櫃和他的居所。
2SAM|15|26|倘若他說：『我不喜愛你』；我在這裏，就照他眼中看為好的待我！」
2SAM|15|27|王對 撒督 祭司說：「你不是先見嗎？你可以平安地回城，你兒子 亞希瑪斯 和 亞比亞他 的兒子 約拿單 ，你們二人的兒子可以與你們同去。
2SAM|15|28|看，我在曠野的渡口那裏等，直到你們來報信給我。」
2SAM|15|29|於是 撒督 和 亞比亞他 將上帝的約櫃請回 耶路撒冷 ，他們就留在那裏。
2SAM|15|30|大衛 蒙頭赤腳走上 橄欖山 的斜坡，一面上一面哭。所有跟隨他的百姓也都各自蒙頭哭著上去；
2SAM|15|31|有人告訴 大衛 說 ：「 亞希多弗 也在叛黨之中，隨從 押沙龍 。」 大衛 說：「耶和華啊，求你使 亞希多弗 的計謀變為愚拙！」
2SAM|15|32|大衛 到了山頂，敬拜上帝的地方，看哪， 亞基 人 戶篩 衣服撕裂，頭蒙灰塵來迎見他。
2SAM|15|33|大衛 對他說：「你若與我一同過去，必拖累我；
2SAM|15|34|你若回城去，對 押沙龍 說：『王啊，我願作你的僕人。我向來作你父親的僕人，現在我也願意作你的僕人。』你就可以為我破壞 亞希多弗 的計謀。
2SAM|15|35|撒督 和 亞比亞他 二位祭司豈不都在你那裏嗎？你在王宮裏聽見甚麼，就要告訴 撒督 和 亞比亞他 二位祭司。
2SAM|15|36|看哪， 撒督 的兒子 亞希瑪斯 ， 亞比亞他 的兒子 約拿單 ，也跟二位祭司在那裏。凡你們所聽見的事，可以託這二人來向我報告。」
2SAM|15|37|於是， 大衛 的朋友 戶篩 進了城， 押沙龍 也進了 耶路撒冷 。
2SAM|16|1|大衛 剛過山頂，看哪， 米非波設 的僕人 洗巴 拉著裝好鞍子的兩匹驢，驢上馱著二百個麵餅，一百個葡萄餅，一百個夏天的果餅，一皮袋酒來迎接他。
2SAM|16|2|王對 洗巴 說：「你的這些東西是甚麼意思呢？」 洗巴 說：「驢是給王的家眷騎的，麵餅和夏天的果餅是給年輕人吃的，酒是給在曠野疲乏的人喝的。」
2SAM|16|3|王說：「你主人的兒子在哪裏呢？」 洗巴 對王說：「看哪，他留在 耶路撒冷 ，因他說：『 以色列 家今日必將我父的國歸還我。』」
2SAM|16|4|王對 洗巴 說：「看哪，凡屬 米非波設 的都是你的了。」 洗巴 說：「我叩拜我主我王，願我在你眼前蒙恩寵。」
2SAM|16|5|大衛 王到了 巴戶琳 ，看哪，有一個人從那裏出來，是 掃羅 家族中 基拉 的兒子，名叫 示每 。他一面走一面咒罵，
2SAM|16|6|又向 大衛 王和王的眾臣僕扔石頭；眾百姓和勇士都在王的左右。
2SAM|16|7|示每 這樣咒罵說：「你這好流人血的，你這無賴，滾吧！滾吧！
2SAM|16|8|你流了 掃羅 全家的血，接續他作王，耶和華把這罪歸在你身上。耶和華將這國交在你兒子 押沙龍 的手中。看哪，你咎由自取，因為你是好流人血的人。」
2SAM|16|9|洗魯雅 的兒子 亞比篩 對王說：「這死狗為何咒罵我主我王呢？讓我過去，割下他的頭來。」
2SAM|16|10|王說：「 洗魯雅 的兒子，我與你們有何相干呢？他這樣咒罵是因耶和華吩咐他：『你要咒罵 大衛 。』如此，誰敢說：『你為甚麼這樣做呢？』」
2SAM|16|11|大衛 又對 亞比篩 和眾臣僕說：「看哪，我親生的兒子尚且尋索我的性命，何況現在這 便雅憫 人呢？由他咒罵吧！因為這是耶和華吩咐他的。
2SAM|16|12|或者耶和華見我遭難 ，因我今日被這人咒罵而向我施恩。」
2SAM|16|13|於是 大衛 和他的人在路上走。 示每 走在 大衛 對面的山坡，一面走一面咒罵，又向他扔石頭，揚起塵土。
2SAM|16|14|王和跟隨他的眾百姓來了，非常疲乏，就在那裏歇息。
2SAM|16|15|押沙龍 和 以色列 眾百姓來到 耶路撒冷 ， 亞希多弗 也與他同來。
2SAM|16|16|大衛 的朋友 亞基 人 戶篩 來到 押沙龍 那裏，對他說：「願王萬歲！願王萬歲！」
2SAM|16|17|押沙龍 對 戶篩 說：「你這樣做是忠誠對待你的朋友嗎？為甚麼不與你的朋友同去呢？」
2SAM|16|18|戶篩 對 押沙龍 說：「不，誰是耶和華和這百姓，以及 以色列 眾人所揀選的，我必歸順他，留在他那裏。
2SAM|16|19|再者，我當服事誰呢？豈不是前王的兒子嗎？我怎樣服事你父親，也必照樣服事你。」
2SAM|16|20|押沙龍 對 亞希多弗 說：「你們出個主意，我們該怎麼做？」
2SAM|16|21|亞希多弗 對 押沙龍 說：「你父親所留下看守宮殿的妃嬪，你可以與她們親近。 以色列 眾人聽見你敢惹你父親憎惡你，凡歸順你人的手就更堅強了。」
2SAM|16|22|於是他們為 押沙龍 在屋頂上支搭帳棚， 押沙龍 就在 以色列 眾人眼前，與他父親的妃嬪親近。
2SAM|16|23|那時 亞希多弗 所出的主意好像人從上帝求問得來的話一樣；他給 大衛 ，給 押沙龍 所出的一切主意，都是這樣。
2SAM|17|1|亞希多弗 對 押沙龍 說：「請讓我挑選一萬二千人，今夜起身追趕 大衛 。
2SAM|17|2|我必趁他疲乏手軟的時候追上他，使他驚惶。跟隨他的眾百姓必都逃跑，我就只殺王一個人。
2SAM|17|3|我必使眾百姓都歸順你，正如眾人歸順你所追殺的人一樣 ，眾百姓就都平安無事了。」
2SAM|17|4|這話在 押沙龍 和 以色列 眾長老的眼中都看為好。
2SAM|17|5|押沙龍 說：「把 亞基 人 戶篩 也召來，我們也要聽他怎麼說。」
2SAM|17|6|戶篩 到了 押沙龍 那裏， 押沙龍 向他說：「 亞希多弗 說了這樣的話，我們要照他的話做嗎？若不可，你就說吧！」
2SAM|17|7|戶篩 對 押沙龍 說：「 亞希多弗 這次所出的主意不好。」
2SAM|17|8|戶篩 又說：「你知道，你父親和他的人都是勇士，他們心裏惱怒，如同田野中失去小熊的母熊一樣；而且你父親是個戰士，必不和百姓一同住宿。
2SAM|17|9|看哪，他現今或藏在一個坑中或在別處，若我們 有人首先被殺，聽見的必說：『跟隨 押沙龍 的百姓被殺了。』
2SAM|17|10|雖有勇士膽大如獅子，他的心也必定融化，因為全 以色列 都知道你父親是英雄，跟隨他的人都是勇士。
2SAM|17|11|依我之計，要把如同海邊的沙那樣多的 以色列 眾人，從 但 直到 別是巴 ，聚集到你這裏來，由你親自率領他們出戰。
2SAM|17|12|我們到他那裏，在任何地方遇見他，就突然臨到他，如同露水滴在泥土上。這樣，他和所有跟隨他的人，一個也不留。
2SAM|17|13|他若撤退到一座城， 以色列 眾人必帶繩子去那城，把城拉到河裏，甚至連一塊小石子也找不到。」
2SAM|17|14|押沙龍 和 以色列 眾人都說：「 亞基 人 戶篩 的計謀比 亞希多弗 的更好！」這是因為耶和華定意破壞 亞希多弗 的良謀，為的是耶和華要降禍給 押沙龍 。
2SAM|17|15|戶篩 對 撒督 和 亞比亞他 二位祭司說：「 亞希多弗 為 押沙龍 和 以色列 的長老出的主意是如此如此，我出的主意是如此如此。
2SAM|17|16|現在你們要急速派人去告訴 大衛 說：『今夜不可在曠野的渡口住宿，務要過河，免得王和所有跟隨他的百姓都被吞滅。』」
2SAM|17|17|約拿單 和 亞希瑪斯 在 隱‧羅結 等候，不敢進城，恐怕被人看見。有一個婢女出來，把這話告訴他們，他們就去報信給 大衛 王。
2SAM|17|18|然而有一個僮僕看見他們，就去告訴 押沙龍 。他們二人急忙離開，跑到 巴戶琳 一個人的家裏。那人院中有一口井，他們就下到那裏。
2SAM|17|19|那家的婦人用蓋蓋上井口，又在上頭鋪上碎麥，事情就沒有洩漏。
2SAM|17|20|押沙龍 的僕人來到婦人的家，說：「 亞希瑪斯 和 約拿單 在哪裏？」婦人對他們說：「他們過了河了。」僕人搜尋，卻找不著，就回 耶路撒冷 去了。
2SAM|17|21|他們走後，二人從井裏上來，去告訴 大衛 王。他們對 大衛 說：「 亞希多弗 出這樣的主意要害你，你們起來，快快過河。」
2SAM|17|22|於是 大衛 和所有跟隨他的百姓都起來，過 約旦河 。到了天亮，無一人不過 約旦河 的。
2SAM|17|23|亞希多弗 見他的計謀不被接納，就備上驢，動身歸回本城，到了自己的家。他留下遺囑給他的家，就上吊死了，葬在他父親的墳墓裏。
2SAM|17|24|大衛 到了 瑪哈念 ， 押沙龍 和跟隨他的 以色列 眾人也都過了 約旦河 。
2SAM|17|25|押沙龍 立 亞瑪撒 作元帥，取代 約押 。 亞瑪撒 是 以實瑪利 人 以特拉 的兒子。 以特拉 曾與 拿轄 的女兒 亞比該 親近；這 亞比該 與 約押 的母親 洗魯雅 是姊妹。
2SAM|17|26|押沙龍 和 以色列 人安營在 基列 地。
2SAM|17|27|大衛 到了 瑪哈念 ， 亞捫 族的 拉巴 人 拿轄 的兒子 朔比 ， 羅‧底巴 人 亞米利 的兒子 瑪吉 ，來自 羅基琳 的 基列 人 巴西萊 ，
2SAM|17|28|帶著被褥、盆、瓦器，還有小麥、大麥、麥麵、烤熟的穀穗、豆子、紅豆、炒豆、
2SAM|17|29|蜂蜜、奶油、綿羊、奶餅，供給 大衛 和跟隨他的人吃，因為他們想：「百姓在曠野中，必定又飢渴又疲乏。」
2SAM|18|1|大衛 數點跟隨他的百姓，立千夫長、百夫長率領他們。
2SAM|18|2|大衛 把軍兵分為三隊 ：三分之一在 約押 手下，三分之一在 洗魯雅 的兒子 約押 弟弟 亞比篩 手下，三分之一在 迦特 人 以太 手下。王對軍兵說：「我必與你們一同出戰。」
2SAM|18|3|軍兵卻說：「你不可出戰。若是我們逃跑，敵人不會把心放在我們身上；我們陣亡一半，敵人也不會把心放在我們身上。但現在你一人抵過我們萬人，所以你最好留在城裏支援我們。」
2SAM|18|4|王對他們說：「你們看怎樣好，我就怎樣做。」於是王站在城門旁，所有的軍兵成百成千地挨次出戰去了。
2SAM|18|5|王囑咐 約押 、 亞比篩 、 以太 說：「你們要為我的緣故寬待那年輕人 押沙龍 。」王為 押沙龍 的事囑咐眾將領的話，所有的軍兵都聽見了。
2SAM|18|6|軍兵出到田野迎戰 以色列 ，在 以法蓮 的樹林裏交戰。
2SAM|18|7|在那裏， 以色列 百姓敗在 大衛 的臣僕面前。那日在那裏陣亡的很多，共有二萬人。
2SAM|18|8|戰爭蔓延到整個地面，那日被樹林吞噬的軍兵比被刀劍吞噬的更多。
2SAM|18|9|押沙龍 剛好遇見了 大衛 的臣僕。 押沙龍 騎著騾子，從大橡樹密枝底下經過，他的頭被橡樹夾住，懸掛在空中 ，所騎的騾子就離他去了。
2SAM|18|10|有個人看見，就告訴 約押 說：「看哪，我看見 押沙龍 掛在橡樹上了。」
2SAM|18|11|約押 對報信的人說：「看哪，你既看見了，為甚麼不當場把他擊殺在地呢？我必賞你十個銀子和一條帶子。」
2SAM|18|12|那人對 約押 說：「即使我手裏得了一千銀子，也不敢伸手害王的兒子，因為我們聽見王囑咐你、 亞比篩 、 以太 說：『你們要謹慎，不可害那年輕人 押沙龍 。』
2SAM|18|13|我若冒著生命危險做這傻事 ，無論何事都瞞不過王，你自己也必遠遠站在一旁。」
2SAM|18|14|約押 說：「我不能在你面前這樣耗下去！」 約押 手拿三枝短槍，趁 押沙龍 在橡樹上 還活著，就刺透他的心。
2SAM|18|15|給 約押 拿兵器的十個青年圍著 押沙龍 ，擊殺他，將他殺死。
2SAM|18|16|約押 吹角，軍兵就回來，不去追趕 以色列 人，因為 約押 制止了軍兵。
2SAM|18|17|他們拿下 押沙龍 ，把他丟在樹林中一個大坑裏，上頭堆起一大堆石頭。 以色列 眾人都逃跑，各回自己的帳棚去了。
2SAM|18|18|押沙龍 活著的時候，曾在 王谷 立了一根柱子，因他說：「我沒有兒子為我留名。」他就以自己的名字稱那柱子為 押沙龍碑 ，直到今日。
2SAM|18|19|撒督 的兒子 亞希瑪斯 說：「讓我跑去報信給王，耶和華已經為王伸冤，使他脫離仇敵的手了。」
2SAM|18|20|約押 對他說：「你今日不可作報信的人，改日再去報信；因為今日王的兒子死了，所以你不可去報信。」
2SAM|18|21|約押 對 古實 人說：「你去把你所看見的告訴王。」 古實 人向 約押 叩拜後，就跑去了。
2SAM|18|22|撒督 的兒子 亞希瑪斯 又對 約押 說：「無論怎樣，讓我隨著 古實 人跑去吧！」 約押 說：「我兒，你報這信息，既不得賞賜，何必要跑去呢？」
2SAM|18|23|他說：「無論怎樣，我要跑去。」 約押 對他說：「你跑去吧！」 亞希瑪斯 就從平原的路往前跑，越過了 古實 人。
2SAM|18|24|大衛 正坐在內外城門之間。守望的人上到城牆，在城門的頂上舉目觀看，看哪，有一個人獨自跑來。
2SAM|18|25|守望的人就大聲告訴王。王說：「他若獨自來，必是報口信的。」那人跑得越來越近了。
2SAM|18|26|守望的人又見一人跑來，就對守城門的人喊說：「看哪，又有一人獨自跑來。」王說：「這也是報信的。」
2SAM|18|27|守望的人說：「我看前面那人的跑法，好像 撒督 的兒子 亞希瑪斯 的跑法。」王說：「他是個好人，是來報好消息的。」
2SAM|18|28|亞希瑪斯 向王呼叫說：「平安了！」他就臉伏於地向王叩拜，說：「耶和華－你的上帝是應當稱頌的，他已把些那舉手攻擊我主我王的人交出來了。」
2SAM|18|29|王說：「年輕人 押沙龍 平安嗎？」 亞希瑪斯 說：「 約押 派王的僕人，就是你的僕人時，我看見一陣大騷動，卻不知道是甚麼事。」
2SAM|18|30|王說：「你退去，站在這裏。」他就退去，站著。
2SAM|18|31|看哪， 古實 人也來到，說：「有信息報給我主我王！耶和華今日為你伸冤，使你脫離一切起來攻擊你之人的手。」
2SAM|18|32|王對 古實 人說：「年輕人 押沙龍 平安嗎？」 古實 人說：「願我主我王的仇敵，和一切起來惡意要害你的人，都像那年輕人一樣。」
2SAM|18|33|王戰抖，就上城門的樓房去痛哭，一面走一面說：「我兒 押沙龍 啊！我兒，我兒 押沙龍 啊！我恨不得替你死， 押沙龍 啊，我兒！我兒！」
2SAM|19|1|有人告訴 約押 ：「看哪，王為 押沙龍 悲哀哭泣。」
2SAM|19|2|那日眾軍兵聽說王為他兒子悲傷，他們得勝的日子變成悲哀了。
2SAM|19|3|那日軍兵暗暗地進城，如同戰場上逃跑、羞愧的士兵一般。
2SAM|19|4|王蒙著臉，大聲哭號說：「我兒 押沙龍 啊！ 押沙龍 ，我兒，我兒啊！」
2SAM|19|5|約押 進了宮到王那裏，說：「你今日使你眾臣僕的臉面羞愧了！他們今日救了你的性命和你兒女妻妾的性命，
2SAM|19|6|你卻愛那些恨你的人，恨那些愛你的人。今日你擺明了不以將帥、臣僕為念。我今日看得出，若 押沙龍 活著，我們今日全都死了，你就高興了。
2SAM|19|7|現在你要起來，出去安慰你臣僕的心。我指著耶和華起誓：你若不出去，今夜必沒有一人跟你在一起了。這禍患比你從幼年到如今所遭受的更嚴重！」
2SAM|19|8|於是王起來，坐在城門口。有人告訴眾軍兵說：「看哪，王坐在城門口。」眾軍兵就都到王的面前。 那時， 以色列 人已經逃跑，各回自己的帳棚去了。
2SAM|19|9|以色列 眾支派的百姓都議論紛紛，說：「王曾救我們脫離仇敵的手，又救我們脫離 非利士 人的手，現在他為了 押沙龍 逃離這地了。
2SAM|19|10|我們所膏治理我們的 押沙龍 已經陣亡。現在你們為甚麼沉默，不請王回來呢？」
2SAM|19|11|大衛 王派人到 撒督 和 亞比亞他 二位祭司那裏，說：「你們當向 猶大 長老說：『 以色列 眾人已經有話到了王那裏 ，你們為甚麼最後才請王回宮呢？
2SAM|19|12|你們是我的弟兄，是我的骨肉，為甚麼最後才請王回來呢？』
2SAM|19|13|你們要對 亞瑪撒 說：『你不是我的骨肉嗎？我若不立你在我面前取代 約押 永久作元帥，願上帝重重懲罰我！』」
2SAM|19|14|這樣，他挽回了 猶大 眾人的心，如同一人。他們就派人到王那裏，說：「請王和王的眾臣僕回來。」
2SAM|19|15|王回來了，到 約旦河 。 猶大 人來到 吉甲 ，去迎接王，請王過 約旦河 。
2SAM|19|16|來自 巴戶琳 的 便雅憫 人 基拉 的兒子 示每 急忙與 猶大 人一同下去迎接 大衛 王。
2SAM|19|17|跟從 示每 的有一千個 便雅憫 人，還有 掃羅 家的僕人 洗巴 和他十五個兒子、二十個隨從僕人，他們都趕緊過 約旦河 到王的面前。
2SAM|19|18|渡船就渡王的家眷過河 ，照王看為好的去做。 王過 約旦河 的時候， 基拉 的兒子 示每 俯伏在王面前，
2SAM|19|19|對王說：「我主我王離開 耶路撒冷 的那日，僕人行了悖逆的事，現在求我主不要因此加罪於僕人，不要記得，也不要放在心上。
2SAM|19|20|僕人明知自己有罪，看哪， 約瑟 全家之中，今日我首先下來迎接我主我王。」
2SAM|19|21|洗魯雅 的兒子 亞比篩 回答說：「 示每 既然咒罵耶和華的受膏者，不應當為這緣故處死他嗎？」
2SAM|19|22|大衛 說：「 洗魯雅 的兒子，我與你們有何相干，你們今日要跟我作對嗎？今日在 以色列 中豈可把任何人處死呢？我豈不知今日我是 以色列 的王嗎？」
2SAM|19|23|於是王對 示每 說：「你必不死。」王就向他起誓。
2SAM|19|24|掃羅 的孫子 米非波設 也下去迎接王。他自從王離開的那一日，直到王平安回 耶路撒冷 的日子，沒有修腳，沒有剃鬍鬚，也沒有洗衣服。
2SAM|19|25|他來迎接王的時候 ，王對他說：「 米非波設 ，你為甚麼沒有與我同去呢？」
2SAM|19|26|他說：「我主我王啊，我的僕人欺騙了我。那日僕人想要備驢騎上，與王同去，因為僕人是瘸腿的。
2SAM|19|27|他卻在我主我王面前毀謗僕人。然而我主我王如同上帝的使者一樣，你看怎樣好，就怎樣做吧！
2SAM|19|28|因為我祖全家的人，在我主我王面前不過是該死的人，王卻使僕人列在王的席上吃飯的人當中，我現在還有甚麼權利能向王請求呢？」
2SAM|19|29|王對他說：「你何必再提你的事呢？我說，你與 洗巴 要平分土地。」
2SAM|19|30|米非波設 對王說：「我主我王既然平安地回宮，甚至讓 洗巴 全都拿去也沒關係。」
2SAM|19|31|基列 人 巴西萊 從 羅基琳 下來，要護送王過 約旦河 ，就跟王一同過 約旦河 。
2SAM|19|32|巴西萊 年紀老邁，已經八十歲了。王住在 瑪哈念 的時候，他拿食物來供給王，因他是個大富翁。
2SAM|19|33|王對 巴西萊 說：「你與我一同渡過去，我要在 耶路撒冷 我的身邊奉養你。」
2SAM|19|34|巴西萊 對王說：「我還能活多少年日，可以與王一同上 耶路撒冷 呢？
2SAM|19|35|今日我已八十歲了，還能辨別美醜嗎？僕人還能嘗出飲食的滋味嗎？還能聽男女歌唱的聲音嗎？僕人何必拖累我主我王呢？
2SAM|19|36|僕人護送王過 約旦河 只是一件小事，王何必用這樣的賞賜來報答我呢？
2SAM|19|37|請讓我回去，死在我本城，葬在我父母的墓旁。看哪，這裏有 金罕 作王的僕人，讓他同我主我王過去，你看怎樣好，就怎樣對待他吧。」
2SAM|19|38|王說：「 金罕 可以與我一同過去，我必照你看為好的待他。你要我做的，我都會為你做。」
2SAM|19|39|於是眾百姓過了 約旦河 ，王也過去了。王親吻 巴西萊 ，為他祝福， 巴西萊 就回自己的地方去了。
2SAM|19|40|王渡過去 ，到了 吉甲 ， 金罕 也跟他過去。 猶大 眾百姓和 以色列 百姓的一半也都送王過去。
2SAM|19|41|看哪， 以色列 眾人來到王那裏，對王說：「我們的弟兄 猶大 人為甚麼暗暗地送王和王的家眷，以及所有跟隨王的人，過 約旦河 呢？」
2SAM|19|42|猶大 眾人回答 以色列 人說：「因為王與我們是親屬，你們為何因這事發怒呢？我們靠王吃了甚麼呢？王真正給了我們甚麼賞賜呢？」
2SAM|19|43|以色列 人回答 猶大 人說：「我們與王有十倍的關係，就是在 大衛 身上，我們也比你們更有權利 。你們為何藐視我們呢？我們不是最先提議請王回來的嗎？」但 猶大 人的話比 以色列 人的話更強硬。
2SAM|20|1|在那裏恰巧有一個無賴，名叫 示巴 ，是 便雅憫 人 比基利 的兒子。他吹角，說： 「我們與 大衛 無份， 與 耶西 的兒子無關。 以色列 啊，各回自己的帳棚去吧！」
2SAM|20|2|於是 以色列 眾人都離棄 大衛 去跟隨 比基利 的兒子 示巴 ，但 猶大 人從 約旦河 直到 耶路撒冷 ，都緊緊跟隨他們的王。
2SAM|20|3|大衛 王來到 耶路撒冷 ，進了宮，就把從前留下看守宮殿的十個妃嬪軟禁在冷宮，養活她們，卻不與她們親近。她們被關起來，活著如同寡婦，直到死的日子。
2SAM|20|4|王對 亞瑪撒 說：「你要在三日之內召集 猶大 人到我這裏來，你自己也要留在這裏。」
2SAM|20|5|亞瑪撒 就去召集 猶大 人，不過他卻耽延，過了王所定的期限。
2SAM|20|6|大衛 對 亞比篩 說：「現在 比基利 的兒子 示巴 對我們的危害恐怕比 押沙龍 更大。你要帶領你主的一些僕人追趕他，免得他得了堅固的城鎮，在我們眼前逃脫 。」
2SAM|20|7|約押 的人和 基利提 人、 比利提 人，以及所有的勇士都跟著 亞比篩 ，從 耶路撒冷 出去追趕 比基利 的兒子 示巴 。
2SAM|20|8|他們到了 基遍 的大石頭那裏， 亞瑪撒 來迎接他們。那時 約押 穿著戰衣，腰束佩刀的帶子，刀在鞘內。 約押 前行時，刀從鞘內掉出來。
2SAM|20|9|約押 對 亞瑪撒 說：「我的弟兄，你平安嗎？」他就用右手抓住 亞瑪撒 的鬍子，要親吻他。
2SAM|20|10|亞瑪撒 沒有防備 約押 手裏拿著的刀； 約押 用刀刺入他的肚腹，他的腸子流在地上， 約押 沒有再刺，他就死了。 約押 和他弟弟 亞比篩 往前追趕 比基利 的兒子 示巴 。
2SAM|20|11|有 約押 的一個僕人站在 亞瑪撒 屍體的旁邊，說：「誰喜愛 約押 ，誰歸順 大衛 ，就當跟隨 約押 。」
2SAM|20|12|亞瑪撒 渾身是血，躺在路中間。那人見眾百姓都站住，就把 亞瑪撒 的屍體從路上移到田間，把衣服蓋在他身上，因為他看見眾人經過時都站住。
2SAM|20|13|屍體從路上移走之後，眾人就都跟隨 約押 去追趕 比基利 的兒子 示巴 。
2SAM|20|14|示巴 走遍 以色列 各支派，直到 伯‧瑪迦 的 亞比拉 ；所有精選的人 都聚集跟隨他。
2SAM|20|15|跟隨 約押 的眾百姓到了 伯‧瑪迦 的 亞比拉 ，圍困 示巴 ，對著城建土堆，與城郭相對。他們猛撞城牆，要使城倒塌。
2SAM|20|16|一個有智慧的婦人從城上呼叫：「聽啊，聽啊，請你們告訴 約押 ：『近前來到這裏，我好與你說話。』」
2SAM|20|17|約押 就近前到她那裏，婦人對他說：「你是 約押 嗎？」他說：「我是。」婦人對他說：「請你聽使女的話。」 約押 說：「我正在聽。」
2SAM|20|18|婦人說：「古時有話說，當在 亞比拉 求問，事情就可以解決。
2SAM|20|19|我在 以色列 中是和平、忠誠的。你現在想要毀壞這城， 以色列 的根源 ，為何你要吞滅耶和華的產業呢？」
2SAM|20|20|約押 回答說：「不，我絕不吞滅和毀壞！
2SAM|20|21|話不是這麼說的，只是因為有一個 以法蓮 山區的人，就是 比基利 的兒子名叫 示巴 ，他舉手攻擊 大衛 王；你們只要把他一人交出來，我就離城而去。」婦人對 約押 說：「看哪，他的首級必從城牆上丟給你。」
2SAM|20|22|婦人憑她的智慧去勸眾百姓，他們就割下 比基利 的兒子 示巴 的首級，丟給 約押 。 約押 吹角，眾人就離城散開，各回自己的帳棚去了。 約押 回 耶路撒冷 ，到王那裏。
2SAM|20|23|約押 統管 以色列 全軍； 耶何耶大 的兒子 比拿雅 統管 基利提 人和 比利提 人；
2SAM|20|24|亞多蘭 管理勞役的人； 亞希律 的兒子 約沙法 作史官；
2SAM|20|25|示法 作書記； 撒督 和 亞比亞他 作祭司；
2SAM|20|26|睚珥 人 以拉 也作 大衛 的祭司。
2SAM|21|1|大衛 在位年間有饑荒，一連三年， 大衛 求問耶和華，耶和華說：「 掃羅 和他家犯了流人血之罪，因為他殺死了 基遍 人。」
2SAM|21|2|大衛 王召了 基遍 人來，跟他們說話。 基遍 人不是 以色列 人，而是 亞摩利 人中所剩下的人。 以色列 人曾向他們起誓， 掃羅 卻為 以色列 人和 猶大 人大發熱心，追殺他們，為了要消滅他們。
2SAM|21|3|大衛 對 基遍 人說：「我當為你們做甚麼呢？要用甚麼贖這罪，使你們為耶和華的產業祝福呢？」
2SAM|21|4|基遍 人對他說：「我們和 掃羅 以及他家的事與金銀無關，也不要因我們的緣故殺任何 以色列 人。」 大衛 說：「你們怎樣說，我就為你們怎樣做。」
2SAM|21|5|他們對王說：「那謀害我們、要消滅我們、使我們不得住 以色列 境內的人，
2SAM|21|6|請把他的子孫七人交給我們，我們好在耶和華面前，把他們懸掛在 基比亞 ，就是耶和華揀選 掃羅 的地方。」王說：「我必交給你們。」
2SAM|21|7|王顧惜 掃羅 的孫子， 約拿單 的兒子 米非波設 ，因為在 大衛 和 掃羅 的兒子 約拿單 之間，有指著耶和華的誓言。
2SAM|21|8|王卻把 愛亞 的女兒 利斯巴 為 掃羅 所生的兩個兒子 亞摩尼 和 米非波設 ，以及 掃羅 的女兒 米拉 為 米何拉 人 巴西萊 兒子 亞得列 所生的五個兒子
2SAM|21|9|交在 基遍 人的手裏。 基遍 人在耶和華面前把他們懸掛在山上，這七人就一起死了。他們被殺的時候正是收割的頭幾天，就是開始收割大麥的時候。
2SAM|21|10|愛亞 的女兒 利斯巴 用麻布舖在磐石上搭棚，從收割的開始直到天降雨在屍體上，她白日不許空中的飛鳥落在屍體上，夜間不讓田野的走獸前來。
2SAM|21|11|有人把 掃羅 的妃子 愛亞 女兒 利斯巴 所做的事告訴 大衛 。
2SAM|21|12|大衛 就去，從 基列 的 雅比 人那裏把 掃羅 和他兒子 約拿單 的骸骨搬來。先前 非利士 人在 基利波 殺了 掃羅 ，把屍體懸掛在 伯‧珊 的廣場上，後來 基列 的 雅比 人把屍體偷走。
2SAM|21|13|大衛 把 掃羅 和他兒子 約拿單 的骸骨從那裏搬上來，又收殮了被懸掛的那些人的骸骨。
2SAM|21|14|他們將 掃羅 和他兒子 約拿單 的骸骨葬在 便雅憫 的 洗拉 ，在 掃羅 父親 基士 的墳墓裏。他們遵照王所吩咐的一切做了。此後上帝垂聽了為那地的祈求。
2SAM|21|15|非利士 人與 以色列 人打仗。 大衛 帶領僕人下去，與 非利士 人交戰， 大衛 就疲乏了。
2SAM|21|16|巨人族的後裔 以實‧比諾 說要殺 大衛 ；他的銅槍重三百舍客勒，腰間又佩著新刀 。
2SAM|21|17|但 洗魯雅 的兒子 亞比篩 幫助 大衛 攻擊 非利士 人，殺死了他。當日， 大衛 的人向 大衛 起誓說：「你不可再與我們一同出戰，免得 以色列 的燈熄滅了。」
2SAM|21|18|後來，在 歌伯 又與 非利士 人打仗，那時 戶沙 人 西比該 殺了巨人族的後裔 撒弗 。
2SAM|21|19|他們又在 歌伯 與 非利士 人打仗， 伯利恆 人 雅雷 的兒子 伊勒哈難 殺了 迦特 人 歌利亞 ；這人的槍桿粗如織布機的軸。
2SAM|21|20|又有一次，他們在 迦特 打仗。那裏有一個身材高大的人，雙手各有六根手指，雙腳各有六根腳趾，共有二十四根；他也是巨人族的後裔。
2SAM|21|21|他向 以色列 罵陣， 大衛 的哥哥 示米亞 的兒子 約拿單 就殺了他。
2SAM|21|22|這四個人是 迦特 巨人族的後裔，都仆倒在 大衛 和他僕人的手下。
2SAM|22|1|當耶和華救 大衛 脫離所有仇敵和 掃羅 之手的日子，他用這詩的歌詞向耶和華說話。
2SAM|22|2|他說： 耶和華是我的巖石、我的山寨、我的救主、
2SAM|22|3|我的上帝、我的磐石、我所投靠的。 他是我的盾牌，是拯救我的角， 是我的碉堡，是我的避難所， 是我的救主，救我脫離兇暴的。
2SAM|22|4|我要求告當讚美的耶和華， 我必從仇敵手中被救出來。
2SAM|22|5|死亡的波浪環繞我， 毀滅的急流驚嚇我，
2SAM|22|6|陰間的繩索纏繞我， 死亡的圈套臨到我。
2SAM|22|7|我在急難中求告耶和華， 向我的上帝呼求。 他從殿中聽了我的聲音； 我的呼求進入他的耳中。
2SAM|22|8|那時，因他發怒地就搖撼震動； 天的根基也戰抖搖撼。
2SAM|22|9|他的鼻孔冒煙上騰； 他的口發火焚燒，連煤炭也燒著了。
2SAM|22|10|他使天下垂，親自降臨； 黑雲在他腳下。
2SAM|22|11|他乘坐基路伯飛行， 在風的翅膀上顯現。
2SAM|22|12|他以黑暗和聚集的水、 天空的密雲為四圍的行宮。
2SAM|22|13|因他發出光輝， 火炭都燒著了。
2SAM|22|14|耶和華在天上打雷； 至高者發出聲音。
2SAM|22|15|他射出箭來，使仇敵四散； 發出閃電，擊潰他們。
2SAM|22|16|耶和華的斥責一發，鼻孔的氣一出， 海底就顯現，大地的根基也暴露。
2SAM|22|17|他從高天伸手抓住我， 把我從大水中拉上來。
2SAM|22|18|他救我脫離我的強敵， 脫離那些恨我的人， 因為他們比我強盛。
2SAM|22|19|我遭遇災難的日子，他們來攻擊我； 但耶和華是我的倚靠。
2SAM|22|20|他領我到寬闊之處， 他救拔我，因他喜愛我。
2SAM|22|21|耶和華必按我的公義報答我， 按我手中的清潔賞賜我。
2SAM|22|22|因為我遵守耶和華的道， 未曾作惡離開我的上帝。
2SAM|22|23|他的一切典章在我面前， 他的律例我也未曾丟棄。
2SAM|22|24|我在他面前作了完全人， 我也持守自己遠離罪孽。
2SAM|22|25|所以耶和華按我的公義， 在他眼前按我的清潔賞賜我。
2SAM|22|26|慈愛的人，你以慈愛待他； 完全的人，你以完善待他；
2SAM|22|27|清潔的人，你以清潔待他； 歪曲的人，你以彎曲待他。
2SAM|22|28|困苦的百姓，你必拯救； 但你的眼目察看高傲的人，使他們降卑。
2SAM|22|29|耶和華啊，你是我的燈； 耶和華必照明我的黑暗。
2SAM|22|30|我藉著你衝入敵軍， 藉著我的上帝跳過城牆。
2SAM|22|31|至於上帝，他的道是完全的； 耶和華的話是純淨的。 凡投靠他的，他就作他們的盾牌。
2SAM|22|32|除了耶和華，誰是上帝呢？ 除了我們的上帝，誰是磐石呢？
2SAM|22|33|上帝是我堅固的保障， 他為我開完全的路。
2SAM|22|34|他使我的腳快如母鹿， 使我站穩在高處。
2SAM|22|35|他教導我的手能爭戰， 我的膀臂能開銅造的弓。
2SAM|22|36|你賜救恩給我作盾牌， 你的庇護 使我為大。
2SAM|22|37|你使我腳步寬闊， 我的腳踝未曾滑跌。
2SAM|22|38|我追趕我的仇敵，消滅他們； 若不將他們滅絕，我總不歸回。
2SAM|22|39|我滅絕了他們， 打傷了他們，使他們站不起來； 他們都倒在我的腳下。
2SAM|22|40|你曾以力量束我的腰，使我能爭戰； 也曾使那起來攻擊我的，都服在我以下。
2SAM|22|41|你又使我的仇敵在我面前轉身逃跑， 使我能殲滅那恨我的人。
2SAM|22|42|他們仰望，卻無人拯救； 就是呼求耶和華，他也不應允。
2SAM|22|43|我搗碎他們，如同地上的灰塵； 踐踏壓碎他們，如同街上的泥土。
2SAM|22|44|你救我脫離我百姓 的紛爭， 保護我作列國的元首； 我素不認識的百姓必事奉我。
2SAM|22|45|外邦人要向我投降， 一聽見我的名聲就必順從我。
2SAM|22|46|外邦人要喪膽， 戰戰兢兢地出營寨。
2SAM|22|47|耶和華永遠活著。 願我的磐石被稱頌， 願上帝－救我的磐石受尊崇。
2SAM|22|48|這位上帝為我伸冤， 使萬民服在我以下。
2SAM|22|49|他救我脫離仇敵， 又把我舉起，高過那些起來攻擊我的人， 救我脫離殘暴的人。
2SAM|22|50|耶和華啊，因此我要在列國中稱謝你， 歌頌你的名。
2SAM|22|51|耶和華賜極大的救恩給他所立的王， 施慈愛給他的受膏者， 就是給 大衛 和他的後裔，直到永遠！
2SAM|23|1|以下是 大衛 末了的話： 「 耶西 的兒子 大衛 的話， 得居高位的， 雅各 的上帝所膏的， 以色列 所喜愛的詩人的話。
2SAM|23|2|耶和華的靈藉著我說話， 他的言語在我的舌頭上。
2SAM|23|3|以色列 的上帝說， 以色列 的磐石向我說： 『那以公義治理人， 以敬畏上帝來治理的，
2SAM|23|4|他必像晨光， 如無雲清晨的日出， 如雨後的光輝， 在嫩草地上。』
2SAM|23|5|我的家在上帝面前不是如此嗎？ 上帝與我立永遠的約， 這約既全備又穩妥。 我的一切救恩和我一切所想望的， 他豈不成全嗎？
2SAM|23|6|但無賴全都像被丟棄的荊棘； 它們不能用手去拿；
2SAM|23|7|碰它們的人必須用鐵器和槍桿， 它們必在那裏被火燒盡。」
2SAM|23|8|大衛 勇士的名字如下： 哈革摩尼 人 約設‧巴設 ，他是三勇士之首；他又名叫 伊斯尼 人 亞底挪 ，曾一次就殺了八百人 。
2SAM|23|9|跟隨 大衛 的三勇士中，其次是 亞何亞 人 朵多 的兒子 以利亞撒 。從前 非利士 人聚集要打仗，他們向 非利士 人罵陣。 以色列 人上去的時候，
2SAM|23|10|他起來擊殺 非利士 人，直到手臂疲乏，手黏住刀把。那日耶和華大獲全勝，百姓跟在 以利亞撒 後面只顧奪取掠物。
2SAM|23|11|再其次是 哈拉 人 亞基 的兒子 沙瑪 。一次， 非利士 人聚集在 利希 ，在一塊長滿紅豆的田裏，百姓在 非利士 人面前逃跑。
2SAM|23|12|沙瑪 卻站在那田的中間，防守那田，擊敗了 非利士 人。耶和華大獲全勝。
2SAM|23|13|開始收割的時候，三個 侍衛 下到 亞杜蘭洞 ，到 大衛 那裏。 非利士 的軍兵在 利乏音谷 安營。
2SAM|23|14|那時 大衛 在山寨， 非利士 人的駐軍在 伯利恆 。
2SAM|23|15|大衛 渴想著說：「但願有人從 伯利恆 城門旁的井裏打水來給我喝！」
2SAM|23|16|這三個勇士就闖過 非利士 人的軍營，從 伯利恆 城門旁的井裏打水，拿來給 大衛 喝。他卻不肯喝，將水澆在耶和華面前，
2SAM|23|17|說：「耶和華啊，我絕不做這事！這三個人冒生命的危險，這不是他們的血嗎？」 大衛 不肯喝這水。這是三個勇士所做的事。
2SAM|23|18|洗魯雅 的兒子， 約押 的兄弟 亞比篩 是這三個勇士的領袖；他曾舉槍殺了三百人，就在三個勇士中得了名。
2SAM|23|19|他在這三個 勇士中是最有名望的，所以作他們的領袖，只是不及前三個勇士。
2SAM|23|20|耶何耶大 的兒子 比拿雅 是來自 甲薛 的勇士，曾行了大事。他殺了 摩押 人 亞利伊勒 的兩個兒子，又在下雪的時候下到坑裏去，殺了一隻獅子。
2SAM|23|21|他又殺了一個魁梧的 埃及 人； 埃及 人手裏拿著槍。 比拿雅 只拿著棍子下到他那裏去，從 埃及 人手裏奪過槍來，用那槍殺死了他。
2SAM|23|22|這些是 耶何耶大 的兒子 比拿雅 所做的事，就在三個勇士裏得了名。
2SAM|23|23|他比那三十個勇士 更有名望，只是不及前三個勇士。 大衛 立他作護衛長。
2SAM|23|24|三十個勇士中有 約押 的兄弟 亞撒黑 ， 伯利恆 人 朵多 的兒子 伊勒哈難 ，
2SAM|23|25|哈律 人 沙瑪 ， 哈律 人 以利加 ，
2SAM|23|26|帕勒提 人 希利斯 ， 提哥亞 人 益吉 的兒子 以拉 ，
2SAM|23|27|亞拿突 人 亞比以謝 ， 戶沙 人 米本乃 ，
2SAM|23|28|亞何亞 人 撒們 ， 尼陀法 人 瑪哈萊 ，
2SAM|23|29|尼陀法 人 巴拿 的兒子 希立 ， 便雅憫 族 基比亞 人 利拜 的兒子 以太 ，
2SAM|23|30|比拉頓 人 比拿雅 ， 迦實溪 人 希太 ，
2SAM|23|31|亞拉巴 人 亞比‧亞本 ， 巴魯米 人 押斯瑪弗 ，
2SAM|23|32|沙本 人 以利雅哈巴 ， 雅善 兒子中的 約拿單 ，
2SAM|23|33|哈拉 人 沙瑪 ， 哈拉 人 沙拉 的兒子 亞希暗 ，
2SAM|23|34|瑪迦 人 亞哈拜 的兒子 以利法列 ， 基羅 人 亞希多弗 的兒子 以連 ，
2SAM|23|35|迦密 人 希斯萊 ， 亞巴 人 帕萊 ，
2SAM|23|36|瑣巴 人 拿單 的兒子 以甲 ， 迦得 人 巴尼 ，
2SAM|23|37|亞捫 人 洗勒 ， 比錄 人 拿哈萊 ，是給 洗魯雅 的兒子 約押 拿兵器的，
2SAM|23|38|以帖 人 以拉 ， 以帖 人 迦立 ，
2SAM|23|39|赫 人 烏利亞 ，共三十七人。
2SAM|24|1|耶和華的怒氣又向 以色列 發作，激起 大衛 來對付他們，說：「去，數點 以色列 人和 猶大 人。」
2SAM|24|2|大衛 對跟隨他的 約押 元帥說：「你來回走遍 以色列 眾支派，從 但 直到 別是巴 ，數點百姓，我好知道百姓的數目。」
2SAM|24|3|約押 對王說：「願耶和華－你的上帝使百姓的數目增加百倍，使我主我王親眼得見。我主我王何必要做這事呢？」
2SAM|24|4|但王堅持他對 約押 和眾軍官的命令。 約押 和眾軍官就從王面前出去，數點 以色列 的百姓。
2SAM|24|5|他們過 約旦河 ，在 迦得谷 中、城的右邊 亞羅珥 安營，與 雅謝 相對。
2SAM|24|6|他們來到 基列 ，到了 他停‧合示 地 ，又來到 但‧雅安 ，繞到 西頓 。
2SAM|24|7|他們來到 推羅 的堡壘，以及 希未 人和 迦南 人的各城，又出來，到 猶大尼革夫 的 別是巴 。
2SAM|24|8|他們來回走遍全地，過了九個月又二十天，就回到 耶路撒冷 。
2SAM|24|9|約押 向王報告百姓的總數： 以色列 拿刀的勇士有八十萬； 猶大 有五十萬人。
2SAM|24|10|大衛 數點百姓以後，心中自責。大衛向耶和華說：「我做這事大大有罪了。耶和華啊，現在求你除掉僕人的罪孽，因我所做的非常愚昧。」
2SAM|24|11|大衛 早晨起來，耶和華的話臨到 迦得 先知，就是 大衛 的先見，說：
2SAM|24|12|「你去告訴 大衛 ：『耶和華如此說：我向你提出三樣，隨你選擇一樣，我好降給你。』」
2SAM|24|13|於是 迦得 來到 大衛 那裏告訴他，問他：「你要國中有七 年的饑荒呢？或是你在敵人面前逃跑，被追趕三個月呢？或是在你國中有三日的瘟疫呢？現在你要考慮思量，我怎樣去回覆那差我來的。」
2SAM|24|14|大衛 對 迦得 說：「我很為難。我們寧願落在耶和華的手裏，因為他有豐盛的憐憫；我不願落在人的手裏。」
2SAM|24|15|於是，耶和華降瘟疫給 以色列 。自早晨到所定的時候，從 但 直到 別是巴 ，百姓中死了七萬人。
2SAM|24|16|天使向 耶路撒冷 伸手要毀滅這城的時候，耶和華改變心意，不降那災難，就對那在百姓中施行毀滅的天使說：「夠了！住手吧！」耶和華的使者正在 耶布斯 人 亞勞拿 的禾場那裏。
2SAM|24|17|大衛 看見那在百姓中施行毀滅的天使，就向耶和華說：「看哪，我犯了罪，行了惡，但這群羊做了甚麼呢？願你的手攻擊我和我的父家。」
2SAM|24|18|當日， 迦得 來到 大衛 那裏，對他說：「你上去，在 耶布斯 人 亞勞拿 的禾場上為耶和華立一座壇。」
2SAM|24|19|大衛 就照著 迦得 的話，照著耶和華所吩咐的上去了。
2SAM|24|20|亞勞拿 觀看，看見王和臣僕向他走過來。 亞勞拿 就出去，臉伏於地，向王下拜。
2SAM|24|21|亞勞拿 說：「我主我王為何來到僕人這裏呢？」 大衛 說：「我要買你這禾場，為耶和華築一座壇，使瘟疫在百姓中停止。」
2SAM|24|22|亞勞拿 對 大衛 說：「我主我王，你眼中看為好，就拿去獻祭。看，這裏有牛可以作燔祭，有打糧的器具和套牛的軛可以當作柴。
2SAM|24|23|王啊，這一切， 亞勞拿 都獻給王。」 亞勞拿 又對王說：「願耶和華－你的上帝悅納你。」
2SAM|24|24|王對 亞勞拿 說：「不，我一定要按價錢向你買；我不能用白白得來的東西作燔祭獻給耶和華－我的上帝。」 大衛 就用五十舍客勒銀子買了那禾場與牛。
2SAM|24|25|大衛 在那裏為耶和華築了一座壇，獻燔祭和平安祭。耶和華垂聽了為那地的祈求，瘟疫就在 以色列 中停止了。
