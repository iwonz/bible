EZRA|1|1|А першого року Кіра, царя перського, щоб сповнилось слово Господнє, проречене устами Єреміїними, збудив Господь духа Кіра, царя перського, і він оголосив по всьому царству своєму, а також на письмі, говорячи:
EZRA|1|2|Так говорить Кір, цар перський: Усі земні царства дав мені Господь, Бог Небесний, і Він наказав мені збудувати Йому храма в Єрусалимі, що в Юдеї.
EZRA|1|3|Хто між вами з усього Його народу, нехай буде Бог його з ним, і нехай він іде до Єрусалиму, що в Юдеї, і нехай будує дім Господа, Бога Ізраїлевого. Це той Бог, що в Єрусалимі.
EZRA|1|4|А кожному позосталому по всіх тих містах, хто мешкає там, нехай допоможуть йому люди його місця сріблом, і золотом, і маєтком, і худобою, з добровільною жертвою для дому Божого, що в Єрусалимі.
EZRA|1|5|І повставали голови батьківських родів Юди та Веніямина, і священики, і Левити, аж до всякого, що Бог збудив духа його, щоб піти будувати дім Господа, що в Єрусалимі.
EZRA|1|6|А все їхнє довкілля зміцнило їм руки речами срібними та золотими, маєтком, і худобою, і коштовностями, окрім того, що хто пожертвував був добровільно.
EZRA|1|7|А цар Кір повиносив речі Господнього дому, які забрав був Навуходоносор з Єрусалиму, і дав їх до дому бога свого,
EZRA|1|8|і повиносив їх Кір, цар перський, рукою скарбника Мітредата, а той відрахував їх Шешбаццарові, Юдиному начальникові.
EZRA|1|9|І оце їхнє число: мисок золотих тридцять, мисок срібних тисяча, ножів двадцять і дев'ять,
EZRA|1|10|келіхів золотих тридцять, келіхів срібних подвійних чотири сотні й десять, посуду іншого тисяча.
EZRA|1|11|Усього золотого й срібного посуду п'ять тисяч і чотири сотні. Усе це завіз Шешбаццар, коли вигнанці верталися з Вавилону до Єрусалиму.
EZRA|2|1|А оце виходьки з округи, що прийшли з полону вигнання, яких вигнав був Навуходоносор, цар вавилонський, до Вавилону, і вони повернулися до Єрусалиму та Юдеї, кожен до міста свого,
EZRA|2|2|ті, що прийшли були з Зоровавелем, Ісусом, Неємією, Сераєю, Реелаєю, Мордехаєм, Білшаном, Міспаром, Біґваєм, Рехумом, Бааною. Число людей Ізраїлевого народу:
EZRA|2|3|синів Пар'ошових дві тисячі сто сімдесят і два,
EZRA|2|4|синів Шефатіїних три сотні сімдесят і два,
EZRA|2|5|синів Арахових сім сотень сімдесят і п'ять,
EZRA|2|6|синів Пахат-Моавових, із синів Ісусових та Йоавових дві тисячі вісім сотень і дванадцять,
EZRA|2|7|синів Еламових тисяча двісті п'ятдесят і чотири,
EZRA|2|8|синів Заттуєвих дев'ять сотень і сорок і п'ять,
EZRA|2|9|синів Заккеєвих сім сотень і шістдесят,
EZRA|2|10|синів Банієвих шість сотень сорок і два,
EZRA|2|11|синів Беваєвих шість сотень двадцять і три,
EZRA|2|12|синів Азґадових тисяча двісті двадцять і два,
EZRA|2|13|синів Адонікамових шість сотень шістдесят і шість,
EZRA|2|14|синів Біґваєвих дві тисячі п'ятдесят і шість,
EZRA|2|15|синів Адінових чотири сотні п'ятдесят і чотири,
EZRA|2|16|синів Атерових, від Єзекії дев'ятдесят і вісім,
EZRA|2|17|синів Бецаєвих три сотні двадцять і три,
EZRA|2|18|синів Йориних сто й дванадцять,
EZRA|2|19|синів Хашумових двісті двадцять і три,
EZRA|2|20|синів Ґіббарових дев'ятдесят і п'ять,
EZRA|2|21|виходьків з Віфлеєму сто двадцять і три,
EZRA|2|22|людей з Нетофи п'ятдесят і шість,
EZRA|2|23|людей з Анатоту сто двадцять і вісім,
EZRA|2|24|виходьків з Азмавету сорок і два,
EZRA|2|25|виходьків з Кір'ят-Аріму, Кефіри та Беероту сім сотень і сорок і три,
EZRA|2|26|виходьків з Рами та Ґеви: шість сотень двадцять і один,
EZRA|2|27|людей з Міхмасу сто двадцять і два,
EZRA|2|28|людей з Бет-Елу та Аю двісті двадцять і три,
EZRA|2|29|виходьків з Нево п'ятдесят і два,
EZRA|2|30|виходьків з Маґбішу сто п'ятдесят і шість,
EZRA|2|31|виходьків з Еламу Другого тисяча двісті п'ятдесят і чотири,
EZRA|2|32|виходьків з Харіму три сотні й двадцять,
EZRA|2|33|виходьків з Лоду, Хадіду та Оно сім сотень двадцять і п'ять,
EZRA|2|34|виходьків з Єрихону три сотні сорок і п'ять,
EZRA|2|35|виходьків з Сенаї три тисячі і шість сотень і тридцять.
EZRA|2|36|Священиків: синів Єдаєвих з Ісусового дому дев'ять сотень сімдесят і три,
EZRA|2|37|синів Іммерових тисяча п'ятдесят і два,
EZRA|2|38|синів Пашхурових тисяча двісті сорок і сім,
EZRA|2|39|синів Харімових тисяча й сімнадцять.
EZRA|2|40|Левитів: синів Ісусових і Кадміїлових, з синів Гадавії сімдесят і чотири.
EZRA|2|41|Співаків: синів Асафових сто двадцять і вісім.
EZRA|2|42|Синів придверних: синів Шаллумових, синів Атерових, синів Талмонових, синів Аккувових, синів Хатітиних, синів Шоваєвих, усіх сто тридцять і дев'ять.
EZRA|2|43|Храмових підданців: синів Ціхіних, синів Хасуфіних, синів Таббаотових,
EZRA|2|44|синів Керосових, синів Сіагіних, синів Падонових,
EZRA|2|45|синів Леваниних, синів Хаґавиних, синів Аккувових,
EZRA|2|46|синів Хаґавових, синів Самлаєвих, синів Хананових,
EZRA|2|47|синів Ґідделових, синів Ґахарових, синів Реаїних,
EZRA|2|48|синів Рецінових, синів Некодиних, синів Ґаззамових,
EZRA|2|49|синів Уззиних, синів Пасеахових, синів Бесаєвих,
EZRA|2|50|синів Асниних, синів Меунімових, синів Нефусімових,
EZRA|2|51|синів Бакбукових, синів Хакуфиних, синів Хархурових,
EZRA|2|52|синів Бацлутових, синів Мехідиних, синів Харшиних,
EZRA|2|53|синів Баркосових, синів Сісриних, синів Темахових,
EZRA|2|54|синів Незіхових, синів Хатіфиних,
EZRA|2|55|синів Соломонових рабів: синів Сотаєвих, синів Соферетових, синів Терудиних,
EZRA|2|56|Синів Яалиних, синів Дарконових, синів Ґідделових,
EZRA|2|57|синів Шефатіїних, синів Хаттілових, синів Похерет-Гаццеваїмових, синів Амієвих,
EZRA|2|58|усього цих храмових підданців та синів Соломонових рабів три сотні дев'ятдесят і два.
EZRA|2|59|А оце ті, що прийшли з Тел-Мелаху, з Тел-Харші, Керув-Аддану та Іммеру, та не могли довести роду батьків своїх та свого насіння, чи вони з Ізраїля:
EZRA|2|60|синів Делаїних, синів Товійїних, синів Некодиних шість сотень п'ятдесят і два.
EZRA|2|61|І з синів священичих: сини Ховайїні, сини Коцові, сини Барзіллая, що взяв жінку з дочок ґілеадянина Барзіллая, і звався їхнім ім'ям.
EZRA|2|62|Вони шукали свого запису родоводу, та не знайшли, і були вони вилучені зо священства,
EZRA|2|63|а намісник сказав їм, щоб вони не їли зо Святого Святих, аж поки не стане священик до уріму та тумміму.
EZRA|2|64|Усього збору разом сорок дві тисячі три сотні шістдесят,
EZRA|2|65|окрім їхніх рабів та невільниць, цих було сім тисяч три сотні тридцять і сім; а їхніх співаків та співачок двісті.
EZRA|2|66|Їхніх коней було сім сотень тридцять і шість, їхніх мулів двісті сорок і п'ять,
EZRA|2|67|їхніх верблюдів чотири сотні тридцять і п'ять, ослів шість тисяч сім сотень і двадцять.
EZRA|2|68|А з голів батьківських родів, коли вони прийшли до Господнього дому, що в Єрусалимі, то вони жертвували до Божого дому, щоб поставити його на його становищі.
EZRA|2|69|За своєю спроможністю вони дали до скарбу на працю: золота шістдесят одну тисячу дарейків, а срібла п'ять тисяч мін, а священичих убрань сто.
EZRA|2|70|І осілися священики й Левити, та з народу, і співаки, і придверні, і храмові підданці по своїх містах, і ввесь Ізраїль по своїх містах.
EZRA|3|1|А коли настав сьомий місяць, і Ізраїлеві сини були по містах, то зібрався народ, як один чоловік, до Єрусалиму.
EZRA|3|2|І встав Ісус, син Йоцадаків, та брати його священики, і Зоровавель, син Шеалтіїлів, та брати його, і збудували жертівника Бога Ізраїля, щоб приносити на ньому цілопалення, як написано в Законі Мойсея, Божого чоловіка.
EZRA|3|3|І поставили міцно жертівника на його основі, бо були вони в страху від народів країв, і приносили на ньому цілопалення для Господа, цілопалення на ранок та на вечір.
EZRA|3|4|І справили свято Кучок, як написано, і щоденні цілопалення в кількості за постановою щодо жертов на кожен день,
EZRA|3|5|а по тому цілопалення стале, і на молодики, і на всі присвячені Господеві свята, і для кожного, хто жертвує добровільну жертву для Господа.
EZRA|3|6|Від першого дня сьомого місяця зачали приносити цілопалення для Господа. А під Господній храм не були ще покладені основи.
EZRA|3|7|І дали срібла каменярам та теслям, і їжі, і питва та оливи, сидонянам та тирянам, щоб достачали кедрові дерева з Ливану до Яфського моря за дозволом їм Кіра, царя перського.
EZRA|3|8|А другого року по своєму приході до Божого дому до Єрусалиму, другого місяця, почали робити Зоровавель, син Шеалтіїлів, і Ісус, син Йоцадаків, і решта їхніх братів, священики та Левити, і всі, хто поприходив з неволі в Єрусалим, а Левитів від віку двадцяти років і вище поставили керувати над працею Господнього дому.
EZRA|3|9|І став Ісус, сини його та брати його, Кадміїл та сини його, сини Юдині, як один чоловік, на догляд над робітниками праці в Божому домі, сини Хенададові, сини їх та їхні брати, Левити.
EZRA|3|10|А коли клали основу Господнього храму, то поставили облаченних священиків із сурмами, а Левитів, Асафових синів, із цимбалами, щоб славити Господа за уставом Давида, Ізраїлевого царя.
EZRA|3|11|І відповіли вони хвалою та подякою Господеві, Добрий бо Він, бо навіки Його милосердя на Ізраїля. А ввесь народ викликував гучним покликом, славлячи Господа за основу Господнього дому!
EZRA|3|12|А багато-хто зо священиків і Левитів та з голів батьківських родів, старші, що бачили перший храм, при заснуванні його, того храму, своїми очима, плакали ревним голосом, а багато-хто покликували піднесеним голосом у радості...
EZRA|3|13|І не міг народ розпізнати голосу поклику радости від голосу плачу народу, бо народ сильно викликував, а голос був чутий аж далеко...
EZRA|4|1|І почули Юдині та Веніяминові вороги, що вигнанці будують храма Господеві, Богові Ізраїля.
EZRA|4|2|І прийшли вони до Зоровавеля та до голів батьківських родів, та й сказали їм: І ми будемо будувати з вами, бо ми звертаємось, як ви, до вашого Бога, і ми приносимо Йому жертви від днів Есар-Хаддона, царя асирійського, що привів нас сюди.
EZRA|4|3|І сказав їм Зоровавель і Ісус, та решта голів батьківських родів Ізраїлевих: Не вам і нам разом будувати храм для Бога! Самі бо ми будемо будувати для Господа, Бога Ізраїлевого, як наказав нам цар Кір, цар перський.
EZRA|4|4|І став народ тієї землі ослаблювати руки Юдиного народу та страхати їх при будуванні.
EZRA|4|5|І підкуплювали вони проти них дорадників царських, щоб заламати їхній задум, по всі дні Кіра, царя перського, й аж до царювання Дарія, царя перського.
EZRA|4|6|А за царя Ахашвероша, на початку його царювання, написали вони оскарження на мешканців Юдеї та Єрусалиму.
EZRA|4|7|А за днів Артаксеркса написав Бішлам, Мітредат, Товеїл та решта товаришів його до Артаксеркса, царя перського. А лист був написаний по-арамейськи, а перекладений по-перськи.
EZRA|4|8|Начальник Рехум та писар Шімай написали одного листа проти Єрусалиму до царя Артаксеркса отак.
EZRA|4|9|Тоді начальник Рехум та писар Шімшай та решта товаришів його, судді й урядники, писарчуки, писарі, аркев'яни, вавилоняни, шушаняни, цебто еламіти,
EZRA|4|10|та решта народів, яких повиганяв Аснаппар, великий та славний, й осадив їх у місті Самарії та в решті Заріччя.
EZRA|4|11|Оце відпис листа, що послали до нього: До царя Артаксеркса твої раби, люди Заріччя. І ось
EZRA|4|12|щоб було відоме цареві, що Юдеї, які вийшли від тебе до нас, прибули до Єрусалиму. Вони будують місто бунтівниче та шкідливе, і вдосконалюють мури, а підвалини поліпшили.
EZRA|4|13|А тепер щоб було відоме цареві, що коли тільки це місто буде збудоване, а мури закінчаться, вони не будуть давати ані данини, ані податку, ані мита, а це буде шкодити царському прибуткові.
EZRA|4|14|І ото, беручи на увагу, що сіль царського палацу сіль наша, а царський сором не випадає нам бачити, тому ми посилаємо й завідомляємо царя,
EZRA|4|15|щоб пошукали в книзі споминів батьків твоїх, і ти знайдеш у книзі споминів, і знатимеш, що місто це місто бунтівниче та шкідливе царям та округам, і що в ньому підіймали бунт від правіку, чому місто це було зруйноване.
EZRA|4|16|Ми сповіщаємо царя, що коли тільки місто це буде добудоване, а мури закінчаться, то через те не буде тобі частки в Заріччі.
EZRA|4|17|Цар послав відповідь: Начальникові Рехумові, і писареві Шімшаєві, та решті їхніх товаришів, що сидять у Самарії, і решта Заріччя: Мир вам! А тепер,
EZRA|4|18|лист, якого ви послали до нас, виразно прочитаний передо мною.
EZRA|4|19|І був виданий від мене наказ, і шукали та й знайшли, що місто це з давніх-давен підіймалося на царів, і повстання та бунт робилися в ньому.
EZRA|4|20|І могутні царі були над Єрусалимом, і панували в усьому Заріччі, а данина, податок та мито давалися їм.
EZRA|4|21|А тепер видайте наказа, щоб спинилися ці люди, а місто це не будувалося, поки від мене не буде виданий новий наказ.
EZRA|4|22|І будьте бережні, щоб через це не зробити помилки. Нащо ростиме зло на шкоду царям?
EZRA|4|23|Тоді, як тільки був прочитаний відпис листа царя Артаксеркса перед Рехумом і писарем Шімшаєм та їхніми товаришами, пішли вони поспішно до Єрусалиму, і спинили роботу їх зброєю та насиллям!
EZRA|4|24|Тим спинилася робота Божого дому, що в Єрусалимі, і спинилася вона аж до другого року царювання Дарія, царя перського...
EZRA|5|1|І пророкував пророк Огій та Захарій, син Іддо, пророки, на юдеїв, що в Юдеї та в Єрусалимі, в Ім'я Бога Ізраїля, що над ними.
EZRA|5|2|Тоді встали Зоровавель, син Шеалтіїлів, та Ісус, син Йоцадаків, і зачали будувати Божий дім, що в Єрусалимі, а з ними Божі пророки, що допомагали їм.
EZRA|5|3|Того часу прийшов до них Таттенай, намісник Заріччя, і Шетар-Бозенай та їхні товариші, і сказали їм так: Хто видав вам наказа будувати цей храм і кінчати цю будову?
EZRA|5|4|Тоді ми сказали їм імена тих мужів, що будують цього будинка.
EZRA|5|5|Та око їхнього Бога було на юдейських старших, і вони не спинили їх, аж поки не піде донесення до Дарія, і тоді дадуть писемну відповідь про це.
EZRA|5|6|Ось відпис листа, що послав Таттенай, намісник Заріччя, і Шетар-Бозенай, та товариство його, і перси, що в Заріччі, до царя Дарія,
EZRA|5|7|вони послали йому донесення, а в ньому писано так: Цареві Дарієві усякого миру!
EZRA|5|8|Щоб було відоме цареві, що ми ходили до Юдейської округи, до дому великого Бога, а він будується з великого каменя, і дерево кладеться в стіни. А робота та робиться докладно, і успіх у їхній руці.
EZRA|5|9|Тоді ми питалися тих старших, і сказали їм так: Хто видав вам наказа будувати цей храм і кінчати цю святиню?
EZRA|5|10|А також питалися ми їх про їхні імена, щоб повідомити тебе, що запишемо ім'я тих мужів, які за голову в них.
EZRA|5|11|А вони так відповіли нам та сказали: Ми то раби Бога небес та землі, і будуємо храма, що був збудований за багато літ перед цим, а збудував його й докінчив його великий Ізраїлів цар.
EZRA|5|12|Але згодом, коли наші батьки розгнівили були Бога небес, Він віддав їх у руку Навуходоносора, царя вавилонського, халдея, а храм той він зруйнував його, а народ вигнав до Вавилону.
EZRA|5|13|Але першого року Кіра, царя вавилонського, цар Кір видав наказа будувати цей дім Божий.
EZRA|5|14|А також посуд Божого дому, золотий та срібний, що Навуходоносор був виніс із єрусалимського храму й заніс його до храму вавилонського, виніс його цар Кір із вавилонського храму й дав мужеві, ім'я його Шешбаццар, якого він настановив намісником.
EZRA|5|15|І сказав він йому: Візьми цей посуд, іди, віднеси його до храму, що в Єрусалимі, а дім Божий нехай будується на своєму місці.
EZRA|5|16|Тоді той Шешбаццар прийшов, заклав підвалини Божого дому в Єрусалимі, і відтоді й аж до цього часу він будується, і не скінчений.
EZRA|5|17|І ось, якщо це цареві добре, нехай пошукається в домі царських скарбів там, у Вавилоні, чи справді від царя Кіра виданий був наказ будувати цей Божий дім в Єрусалимі, а царську волю про це нехай пошлють до нас.
EZRA|6|1|Тоді цар Дарій видав наказа, і шукали в домі, де складають скарби книжок у Вавилоні.
EZRA|6|2|І був знайдений один звій в замку Ахметі, що в мідійській окрузі, а в ньому написано так: На пам'ять.
EZRA|6|3|Першого року царя Кіра цар Кір видав наказа: Дім Божий в Єрусалимі дім той нехай будується на місці, де приносять жертви, а його підвалини заложені. Вишина його шістдесят ліктів, ширина його шістдесят ліктів.
EZRA|6|4|Три ряди з великого каменю, й один ряд з дерева, а видатки будуть дані з царського дому.
EZRA|6|5|А посуд Божого дому, золотий та срібний, що Навуходоносор виніс був із храму, що в Єрусалимі, і переніс до Вавилону, нехай повернуть, і нехай він піде до храму, що в Єрусалимі, на своє місце, і покладеш те в Божому домі...
EZRA|6|6|Тепер же ти, Таттенаю, наміснику Заріччя, ти, Шетор-Бозенаю з товаришами своїми, перси, що в Заріччі, віддаліться звідти!
EZRA|6|7|Позоставте працю цього Божого дому, юдейський намісник та юдейські старші збудують той Божий дім на його місці.
EZRA|6|8|А від мене даний наказ про те, що ви будете робити з тими юдейськими старшими, щоб збудувати цей Божий дім, а з царського добра, з данини Заріччя, нехай докладно дається видаток тим людям, щоб не спиняти роботи.
EZRA|6|9|А що буде потрібне, чи телят, чи баранів, чи овечок на принесення Небесному Богові, пшеницю, сіль, вино та оливу, що скажуть священики, які в Єрусалимі, щоб без омани видавалося їм день-у-день,
EZRA|6|10|щоб вони завжди приносили пахощі в жертву Небесному Богові та молилися за життя царя та синів його.
EZRA|6|11|А від мене виданий наказ, що коли який чоловік змінить це моє слово, то буде вирване дерево з дому його, і буде поставлене, а він буде прибитий на ньому, а дім його буде обернений за це в руїну!
EZRA|6|12|А Бог, що вчинив, щоб там пробувало Ім'я Його, знищить кожного царя та народ, що простягне свою руку, щоб змінити це, щоб ушкодити той Божий дім, що в Єрусалимі! Я, Дарій, видав цього наказа, нехай він докладно буде виконаний!
EZRA|6|13|Тоді Таттенай, намісник Заріччя, Шетар-Бозенай та їхні товариші докладно зробили згідно з тим, як послав цар Дарій.
EZRA|6|14|А юдейські старші будували, і щастило їм за пророцтвом пророка Огія та Захарія, сина Іддо. І вони збудували й закінчили з наказу Бога Ізраїлевого та з наказу Кіра, і Дарія, і Артаксеркса, царя перського.
EZRA|6|15|І закінчений був цей храм до третього місяця адара, що він місяць дванадцятий, шостого року царювання царя Дарія.
EZRA|6|16|І справили Ізраїлеві сини, священики й Левити та решта вигнанців свято відновлення того Божого дому з радістю.
EZRA|6|17|І принесли в жертву на свято відновлення того Божого дому: волів сотню, баранів двісті, ягнят чотири сотні, а козлят у жертву за гріх за всього Ізраїля дванадцять, за числом Ізраїлевих племен.
EZRA|6|18|І поставили священиків за їхніми частинами, а Левитів за чергами їхніми на службу Божого дому, що в Єрусалимі, як написано в книзі Мойсея.
EZRA|6|19|А поверненці справили Пасху чотирнадцятого дня першого місяця,
EZRA|6|20|бо очистилися священики та Левити, як один, усі вони чисті. І вони зарізали пасхальне ягня для всіх поверненців, для своїх братів священиків та для себе.
EZRA|6|21|І їли Ізраїлеві сини, що вернулися з вигнання, і також усі, хто відділився до них від нечистости народів землі, щоб звертатися до Господа, Бога Ізраїлевого.
EZRA|6|22|І справляли вони свято Опрісноків сім день у радості, бо Господь їх потішив і обернув до них серце асирійського царя, щоб зміцнити їхні руки при праці дому Бога, Бога Ізраїлевого.
EZRA|7|1|А по цих пригодах, за царювання Артаксеркса, царя перського, Ездра, син Азарії, сина Хійлкійї,
EZRA|7|2|сина Шаллуна, сина Садока, сина Ахітуви,
EZRA|7|3|сина Амарії, сина Азарії, сина Мерайота,
EZRA|7|4|сина Захарія, сина Уззі, сина Буккі,
EZRA|7|5|сина Авішуї, сина Пінхаса, сина Елеазара, сина Аарона, первосвященика,
EZRA|7|6|цей Ездра вийшов із Вавилону, а він був учитель, знавець Мойсеєвого Закону, що його дав Господь, Бог Ізраїлів. І дав йому цар згідно з тим, як була на ньому рука Господа, Бога його, всяке його пожадання.
EZRA|7|7|І пішли з ним дехто з Ізраїлевих синів, і з священиків, і Левитів, і співаків, і придверних, і храмових підданців до Єрусалиму сьомого року царя Артаксеркса.
EZRA|7|8|І прибув він до Єрусалиму п'ятого місяця, а то сьомий рік царювання.
EZRA|7|9|Бо першого дня місяця першого був початок виходу з Вавилону, а першого дня п'ятого місяця він прийшов до Єрусалиму, бо рука його Бога була добра на ньому.
EZRA|7|10|Бо Ездра приготовив своє серце досліджувати Господнього Закона, і виконувати його, і навчати в Ізраїлі устава та права.
EZRA|7|11|А оце відпис писання, що цар Артаксеркс дав священикові Ездрі, учителеві, що пише слова заповідей Господа та Його устави над Ізраїлем:
EZRA|7|12|Артаксеркс, цар над царями, до священика Ездри, досконалого вчителя Закону Бога Небесного, і так далі.
EZRA|7|13|А ось виданий від мене наказ, щоб кожен, хто в моїм царстві з Ізраїлевого народу, і їхніх священиків, і Левитів з доброї волі бажає йти до Єрусалиму з тобою, нехай іде,
EZRA|7|14|через те, що ти посланий від царя та семи його дорадників, щоб дослідити про Юдею та про Єрусалим за правом твого Бога, правом, що в руці твоїй,
EZRA|7|15|і щоб відправити срібло та золото, що цар та дорадники його пожертвували для Бога Ізраїлевого, Якого місце перебування в Єрусалимі,
EZRA|7|16|і все срібло та золото, яке ти знайдеш у всій вавилонській окрузі разом із пожертвами народу та священиків, які жертвують для дому їхнього Бога, що в Єрусалимі.
EZRA|7|17|Тому ти невідкладно купиш за це срібло биків, баранів, овечок, і їх жертви хлібні та їх жертви ливні, і принесеш їх на жертівнику дому вашого Бога, що в Єрусалимі.
EZRA|7|18|А що тобі та браттям твоїм буде добре вчинити з рештою срібла та золота, те зробіть за вподобанням вашого Бога.
EZRA|7|19|А посуд, що даний тобі на служення дому твого Бога, віддай у цілості перед Богом Єрусалиму.
EZRA|7|20|А решта потрібного для дому Бога твого, що випаде тобі дати, буде дана з дому царських скарбів.
EZRA|7|21|А від мене я цар Артаксеркс виданий наказ для всіх скарбників, що в Заріччі, що все, чого зажадає від вас священик Ездра, учитель Закону Бога Небесного, нехай буде докладно зроблене:
EZRA|7|22|срібла аж до сотні талантів, і пшениці аж до сотні корів, і вина аж до сотні батів, і оливи аж до сотні батів, за соли без запису.
EZRA|7|23|Усе, що з наказу Небесного Бога, нехай буде горливо зроблене для дому Небесного Бога, бо нащо був би гнів на царство царя та на синів його?
EZRA|7|24|І вас завідомляємо, що всі священики та Левити, співаки, придверні, храмові підданці та працівники того Божого дому вільні, данини, податку, чи мита не належить накладати на них!
EZRA|7|25|А ти, Ездро, за мудрістю Бога твого, яка в руці твоїй, попризначай суддів та виконавців Закону, щоб судили для всього народу, що в Заріччі, для всіх, хто знає закони твого Бога, а хто не знає, тих навчите.
EZRA|7|26|А кожен, хто не буде виконувати Закона твого Бога та закона царського докладно, щоб чинився над ним суд: чи то на смерть, чи то на вигнання, чи то на кару маєткову, чи то на ув'язнення.
EZRA|7|27|Благословенний Господь, Бог наших батьків, що вклав у цареве серце, щоб оздобити дім Господній, що в Єрусалимі,
EZRA|7|28|а на мене нахилив милість перед царем та його дорадниками, та всіма хоробрими царевими зверхниками! А я зміцнився, бо рука Господа, Бога, була надо мною, і я зібрав провідних людей з Ізраїля, щоб вони пішли зо мною.
EZRA|8|1|А оце голови їхніх батьків та їх родовід, що пішли зо мною, за царювання царя Артаксеркса, з Вавилону:
EZRA|8|2|з Пінхасових синів: Ґершом, з Ітамарових синів: Даніїл, з Давидових синів: Хаттуш.
EZRA|8|3|З Шеханіїних синів, з Пар'ошових синів: Захарій, а з ним за родоводом сто й п'ятдесят мужчин.
EZRA|8|4|З Пахат-Моавових синів: Ел'єгоенай, син Зерахіїн, а з ним двісті мужчин.
EZRA|8|5|З синів Затту: Шеханія, син Яхазіїлів, а з ним три сотні мужчин.
EZRA|8|6|А з Адінових синів: Евед, син Йонатанів, а з ним п'ятдесят мужчин.
EZRA|8|7|А з Еламових синів: Єшая, син Аталіїн, а з ним сімдесят мужчин.
EZRA|8|8|А з Шефатіїних синів: Зевадія, син Михаїлів, а з ним вісімдесят мужчин.
EZRA|8|9|З Йоавових синів: Овадія, син Єгіїлів, а з ним двісті й вісімнадцять мужчин.
EZRA|8|10|А з синів Бані: Шеломіт, син Йосіфіїн, а з ним сотня й шістдесят мужчин.
EZRA|8|11|А з Беваєвих синів: Захарій, син Беваїв, а з ним двадцять і вісім мужчин.
EZRA|8|12|А з Азґадових синів: Йоханан, син Катанів, а з ним сотня й десять мужчин.
EZRA|8|13|А з Адонікамових синів останні, а оце їхні імена: Еліфелет, Єіїл, і Шемая, а з ними шістдесят мужчин.
EZRA|8|14|А з Біґваєвих синів: Утай і Заввуд, а з ними сімдесят мужчин.
EZRA|8|15|І зібрав я їх до річки, що впадає до Агави, і ми таборували там три дні. І переглянув я народ та священиків, і не знайшов там нікого з Левієвих синів.
EZRA|8|16|І послав я по Еліезера, по Аріїла, по Шемаю, по Елнатана, і по Яріва, і по Елнатана, і по Натана, і по Захарія, і по Мешуллама, голів, і по Йойаріва, і по Елнатана, учителів.
EZRA|8|17|І відправив я їх до Іддо, голови в місцевості Касіф'я, і вклав в їхні уста слова, щоб говорити до Іддо та братів його, підданих у місцевості Касіф'я, щоб вони привели нам служителів для дому нашого Бога.
EZRA|8|18|І привели вони нам, бо рука нашого Бога була добра до нас, чоловіка розумного з синів Махлі, сина Левія, Ізраїлевого сина, та Шеревею й синів його та братів його, вісімнадцять,
EZRA|8|19|та Хашавію, а з ним Єшаю, з синів Мерарієвих, братів його та синів його двадцять,
EZRA|8|20|а з підданців храму, яких дав Давид та зверхники на роботу Левитам, двісті й двадцять підданців: усі вони були означені поіменно.
EZRA|8|21|І проголосив я там піст, над річкою Агавою, щоб упокорятися нам перед лицем нашого Бога, щоб просити від Нього щасливої дороги для нас і для дітей наших та для всього нашого маєтку,
EZRA|8|22|бо я соромився просити від царя війська та верхівців, щоб помагали нам у дорозі проти ворога, бо сказали ми цареві, говорячи: Рука нашого Бога на добро для всіх, хто шукає Його, а сила Його та гнів Його на всіх, хто кидає Його!
EZRA|8|23|І постили ми, і просили нашого Бога про це, і Він дав нам ублагати Себе.
EZRA|8|24|І я відділив із священичих зверхників дванадцять до Шеревеї, Хашавії, і до десятьох їхніх братів з ними.
EZRA|8|25|І відважив я їм срібло й золото та посуд принесення нашого Божого дому, що принесли цар, і його дорадники, і його зверхники та ввесь Ізраїль, що знаходився там.
EZRA|8|26|І відважив я на їхню руку шість сотень і п'ятдесят талантів срібла, а срібних речей сто талантів, золота сто талантів,
EZRA|8|27|а золотих чаш двадцять на тисячу дарейків, а посудин з золоченої й доброї міді дві, дорогі, як золото.
EZRA|8|28|І сказав я до них: Ви святість для Господа, і цей посуд святість, а те срібло та золото добровільна жертва для Господа, Бога ваших батьків.
EZRA|8|29|Пильнуйте й бережіть це, аж поки не відважите його перед зверхниками священиків і Левитів та зверхниками батьківських родів Ізраїлевих в Єрусалимі до кімнат Господнього дому.
EZRA|8|30|І прийняли священики та Левити вагу того срібла та золота та того посуду, щоб віднести до Єрусалиму, до дому нашого Бога.
EZRA|8|31|І рушили ми з річки Агави двадцятого дня першого місяця, щоб іти до Єрусалиму. А рука нашого Бога була над нами, і Він урятував нас з руки ворога та чатівника на дорозі.
EZRA|8|32|І прийшли ми до Єрусалиму, і сиділи там три дні.
EZRA|8|33|А четвертого дня відважили ми те срібло й золото та той посуд у домі нашого Бога на руку священика Меремота, сина Урійїного, а з ним був Елеазар, син Пінхасів, а з ними Йозавад, син Єшуїн, та Ноадія, син Біннуїв, Левити,
EZRA|8|34|за числом, за вагою на все. І того часу була записана вся та вага.
EZRA|8|35|Ті, що прийшли з полону, сини вигнання, принесли цілопалення для Бога Ізраїля: дванадцять биків за всього Ізраїля, дев'ятдесят і шість баранів, сімдесят і сім овець, дванадцять козлів на жертву за гріх, це все цілопалення для Господа.
EZRA|8|36|І віддали цареві накази царським сатрапам та намісникам Заріччя, а ті підтримували народ та Божий дім.
EZRA|9|1|А як скінчилося це, підійшли до мене зверхники, говорячи: Цей народ, Ізраїль, і священики та Левити не відділилися від народів цих країв з їхніми гидотами, від хананеян, періззеян, євусеян, аммонеян, моавітян, єгиптян та амореян,
EZRA|9|2|бо побрали з їхніх дочок собі та своїм синам, змішалося святе насіння з народами цих країв, а рука зверхників та представників була перша в цьому спроневіренні.
EZRA|9|3|А коли я почув це слово, то роздер я одежу свою та плаща свого, і рвав волосся з голови своєї та з бороди своєї, і сидів остовпілий...
EZRA|9|4|І зібралися до мене всі тремтячі перед словами Бога Ізраїлевого за спроневірення поверненців, а я сидів остовпілий аж до жертви вечірньої.
EZRA|9|5|А за вечірньої жертви встав я з упокорення свого, і, роздерши шату свою та плаща свого, упав я на коліна свої, і простягнув руки свої до Господа, Бога мого...
EZRA|9|6|І сказав я: Боже мій, соромлюся я та стидаюся піднести, Боже мій, обличчя своє до Тебе, бо беззаконня наші помножилися понад голову, а наша провина виросла аж до неба!...
EZRA|9|7|Від днів наших батьків ми в великій провині аж до дня цього, а за наші беззаконня були віддані ми, наші царі, наші священики в руку царів цих країв на меча, на полон, і на грабіж, і на посоромлення обличчя, як цього дня.
EZRA|9|8|А тепер на малу хвилю сталася нам милість від Господа, Бога нашого, щоб позоставити нам останок, і дати нам затвердитися на місці святині Його, щоб освітити очі наші, Боже наш, і дати нам трохи ожити в нашій неволі!
EZRA|9|9|Бо раби ми, та в нашій неволі не покинув нас Бог наш, і прихилив до нас милість перед перськими царями, щоб дати нам ожити, щоб піднести дім нашого Бога й щоб відбудувати руїни його, та щоб дати нам захист в Юдеї та в Єрусалимі.
EZRA|9|10|А тепер що скажемо, Боже наш, по цьому? Бо ми покинули заповіді Твої,
EZRA|9|11|які Ти наказав через Своїх рабів пророків, говорячи: Цей Край, що ви йдете посісти, він край нечистий через нечистість народу цих країв, через їхні гидоти, що наповнили його від краю до краю своєю нечистістю.
EZRA|9|12|А тепер дочок своїх не давайте їхнім синам, а їхніх дочок не беріть для своїх синів, і не питайте їх про мир та про добро їх аж навіки, щоб ви стали сильні, та споживали добро цієї землі, і віддали на спадок вашим синам аж навіки.
EZRA|9|13|А по тому всьому, що прийшло на нас за наші злі чини та за нашу велику провину, бо Ти, Боже наш, стримав кару більше від гріха нашого, і дав нам таку рештку,
EZRA|9|14|чи знову ми ламатимемо заповіді Твої, і будемо посвоячуватися з оцими мерзотними народами? Чи ж Ти не розгніваєшся на нас аж до вигублення нас, так що ніхто не позостався б і не врятувався?
EZRA|9|15|Господи, Боже Ізраїлів, Ти праведний, бо ми позосталися останком, як цього дня. Ось ми в провині своїй перед лицем Твоїм, бо не встояти нам за це перед лицем Твоїм!...
EZRA|10|1|А коли Ездра молився та сповідався, плакав та припадав перед Божим домом, зібрався до нього з Ізраїля дуже великий збір, чоловіки, і жінки та діти, бо народ плакав ревним плачем...
EZRA|10|2|І відповів Шеханія, Єхіїлів син, з Еламових синів, та й сказав до Ездри: Ми спроневірилися нашому Богові, бо взяли ми чужинок із народів цього краю за жінок. Але є ще надія для Ізраїля в цьому!
EZRA|10|3|А тепер складімо заповіта нашому Богові, що випровадимо від себе всіх жінок та народжене від них, за радою пана нашого, та тих, хто тремтить перед заповіддю нашого Бога, і буде зроблене за Законом.
EZRA|10|4|Устань, бо на тобі ця річ, а ми з тобою. Будь мужній і дій!
EZRA|10|5|І встав Ездра, і заприсяг зверхників, священиків і Левитів та всього Ізраїля, щоб робити за цим словом. І вони заприсягли.
EZRA|10|6|І Ездра встав з-перед Божого дому й пішов до кімнати Єгохонана, Ел'яшівового сина, і ночував там. Хліба він не їв і води не пив, бо був у жалобі за спроневірення поверненців.
EZRA|10|7|І оголосили в Юдеї та в Єрусалимі до всіх поверненців, щоб зібратися до Єрусалиму.
EZRA|10|8|А кожен, хто не прийде до трьох день, за порадою зверхників та старших, увесь маєток того буде зроблений закляттям, а він буде вилучений із громади поверненців.
EZRA|10|9|І зібралися всі люди Юди та Веніямина до Єрусалиму до трьох день, це був дев'ятий місяць, двадцятого дня місяця. І сидів увесь народ на площі Божого дому, тремтячи від цієї справи та від дощу.
EZRA|10|10|І встав священик Ездра та й сказав до них: Ви спроневірилися, і взяли чужинних жінок, щоб побільшити Ізраїлеву провину.
EZRA|10|11|А тепер повиніться Господеві, Богові ваших батьків, і чиніть Його волю! І віддаліться від народів цього Краю та від тих чужих жінок!
EZRA|10|12|І відповіла вся громада, і сказали гучним голосом: Так, за словом твоїм, ми повинні зробити!
EZRA|10|13|Але народ численний, і час дощів, і нема сили стояти на вулиці. Та й праці не на один день і не на два, бо ми багато нагрішили в цій справі.
EZRA|10|14|Нехай же стануть наші зверхники за ввесь збір, а кожен, хто є в наших містах, хто взяв чужинних жінок, нехай прийде на означені часи, а з ними старші кожного міста та судді його, аж поки не відвернеться від нас жар гніву нашого Бога за цю річ.
EZRA|10|15|Особливо стали над цим Йонатан, син Асагелів, та Яхзея, син Тіквин, а Мешуллам та Левит Шеббетай допомагали їм.
EZRA|10|16|І зробили так поверненці. І відділив собі священик Ездра людей, голів батьків за родом їхніх батьків, і всі вони поіменно. І сіли вони першого дня десятого місяця, щоб дослідити цю справу.
EZRA|10|17|І скінчили до першого дня першого місяця справи про всіх тих людей, що взяли були чужинних жінок.
EZRA|10|18|І знайшлися поміж священичими синами, що взяли чужинних жінок, із синів Єшуї, сина Йоцадакового, та братів його: Моасея, і Еліезер, і Ярів, і Ґедалія.
EZRA|10|19|І дали вони руку свою, що повипроваджують жінок своїх, а винні принесли в жертву барана з отари за провину свою.
EZRA|10|20|А з синів Іммерових: Ханані та Зевадія.
EZRA|10|21|І з синів Харімових: Массея, і Елійя, і Шемая, і Єхіїл, і Уззійя.
EZRA|10|22|І з синів Пашхурових: Ел'йоенай, Маасея, Ізмаїл, Натанаїл, Йозавад та Ел'аса.
EZRA|10|23|А з Левитів: Йозавад, і Шім'ї, і Келая, він Келіта, Петахія, Юда та Еліезер.
EZRA|10|24|А з співаків: Ел'яшів. А з придверних: Шаллум, і Телем, та Урі.
EZRA|10|25|А з Ізраїля, з синів Пар'ошових: Рам'я, і Їззійя, і Малкійя, і Мійямін, і Елеазар, і Малкійя та Беная.
EZRA|10|26|А з синів Еламових: Маттанія, Захарій, і Єхіїл, і Авді, і Єремот, і Елійя.
EZRA|10|27|І з синів Затту: Ел'йоенай, Ел'яшів, Маттанія, і Еремот, і Завад та Азіза.
EZRA|10|28|А з синів Беваєвих: Єгоханан, Хананія, Заббай, Атлай.
EZRA|10|29|І з синів Банієвих: Мешуллам, Маллух, і Адая, Яшув, і Шеал та Рамот.
EZRA|10|30|І з синів Пахатових: Моав, Адна, і Хелал, Беная, Маасея, Маттанія, Веселіїл, і Біннуй та Манасія.
EZRA|10|31|І з синів Харімових: Еліезер, Їшшійя, Малкійя, Шемая, Шімон,
EZRA|10|32|Веніямин, Маллух, Шемарія.
EZRA|10|33|З синів Хашумових: Маттенай, Маттатта, Завад, Еліфелет, Єремай, Манасія, Шім'ї.
EZRA|10|34|З синів Банаєвих: Маадай, Амрам, і Уїл,
EZRA|10|35|Беная, Бедея, Келугу,
EZRA|10|36|Ванія, Меремот, Ел'ятів,
EZRA|10|37|Маттанія, Маттенай, і Яасай,
EZRA|10|38|і Бані, і Біннуй, Шім'ї,
EZRA|10|39|і Шелемія, і Натан, і Адая,
EZRA|10|40|Махнадвай, Шашай, Шарай,
EZRA|10|41|Азаріїл, і Шелемія, Шемарія,
EZRA|10|42|Шаллум, Амарія, Йосип.
EZRA|10|43|А з синів Нево: Єіїл, Маттітія, Завад, Зевіна, Яддай, і Йоїл, Беная.
EZRA|10|44|Усі оці взяли були чужинних жінок, а деякі з цих жінок і дітей породили.
