JUDG|1|1|По смерти Иисуса вопрошали сыны Израилевы Господа, говоря: кто из нас прежде пойдет на Хананеев – воевать с ними?
JUDG|1|2|И сказал Господь: Иуда пойдет; вот, Я предаю землю в руки его.
JUDG|1|3|Иуда же сказал Симеону, брату своему: войди со мною в жребий мой, и будем воевать с Хананеями; и я войду с тобою в твой жребий. И пошел с ним Симеон.
JUDG|1|4|И пошел Иуда, и предал Господь Хананеев и Ферезеев в руки их, и побили они из них в Везеке десять тысяч человек.
JUDG|1|5|В Везеке встретились они с Адони–Везеком, сразились с ним и разбили Хананеев и Ферезеев.
JUDG|1|6|Адони–Везек побежал, но они погнались за ним и поймали его и отсекли большие пальцы на руках его и на ногах его.
JUDG|1|7|Тогда сказал Адони–Везек: семьдесят царей с отсеченными на руках и на ногах их большими пальцами собирали [крохи] под столом моим; как делал я, так и мне воздал Бог. И привели его в Иерусалим, и он умер там.
JUDG|1|8|И воевали сыны Иудины против Иерусалима и взяли его, и поразили его мечом и город предали огню.
JUDG|1|9|Потом пошли сыны Иудины воевать с Хананеями, которые жили на горах и на полуденной земле и на низменных местах.
JUDG|1|10|И пошел Иуда на Хананеев, которые жили в Хевроне (имя же Хеврону [было] прежде Кириаф–Арбы), и поразили Шешая, Ахимана и Фалмая.
JUDG|1|11|Оттуда пошел он против жителей Давира; имя Давиру [было] прежде Кириаф–Сефер.
JUDG|1|12|И сказал Халев: кто поразит Кириаф–Сефер и возьмет его, тому отдам Ахсу, дочь мою, в жену.
JUDG|1|13|И взял его Гофониил, сын Кеназа, младшего брата Халевова, и [Халев] отдал в жену ему Ахсу, дочь свою.
JUDG|1|14|Когда надлежало ей идти, [Гофониил] научил ее просить у отца ее поле, и она сошла с осла. Халев сказал ей: что тебе?
JUDG|1|15|[Ахса] сказала ему: дай мне благословение; ты дал мне землю полуденную, дай мне и источники воды. И дал ей [Халев] источники верхние и источники нижние.
JUDG|1|16|И сыны [Иофора] Кенеянина, тестя Моисеева, пошли из города Пальм с сынами Иудиными в пустыню Иудину, которая на юг от Арада, и пришли и поселились среди народа.
JUDG|1|17|И пошел Иуда с Симеоном, братом своим, и поразили Хананеев, живших в Цефафе, и предали его заклятию, и [от того] называется город сей Хорма.
JUDG|1|18|Иуда взял также Газу с пределами ее, Аскалон с пределами его, и Екрон с пределами его.
JUDG|1|19|Господь был с Иудою, и он овладел горою; но жителей долины не мог прогнать, потому что у них были железные колесницы.
JUDG|1|20|И отдали Халеву Хеврон, как говорил Моисей, и изгнал [он] оттуда трех сынов Енаковых.
JUDG|1|21|Но Иевусеев, которые жили в Иерусалиме, не изгнали сыны Вениаминовы, и живут Иевусеи с сынами Вениамина в Иерусалиме до сего дня.
JUDG|1|22|И сыны Иосифа пошли также на Вефиль, и Господь был с ними.
JUDG|1|23|И остановились и высматривали сыны Иосифовы Вефиль (имя же городу [было] прежде Луз).
JUDG|1|24|И увидели стражи человека, идущего из города, и сказали ему: покажи нам вход в город, и сделаем с тобою милость.
JUDG|1|25|Он показал им вход в город, и поразили они город мечом, а человека сего и все родство его отпустили.
JUDG|1|26|Человек сей пошел в землю Хеттеев, и построил город и нарек имя ему Луз. Это имя его до сего дня.
JUDG|1|27|И Манассия не выгнал [жителей] Бефсана и зависящих от него городов, Фаанаха и зависящих от него городов, жителей Дора и зависящих от него городов, жителей Ивлеама и зависящих от него городов, жителей Мегиддона и зависящих от него городов; и остались Хананеи жить в земле сей.
JUDG|1|28|Когда Израиль пришел в силу, тогда сделал он Хананеев данниками, но изгнать не изгнал их.
JUDG|1|29|И Ефрем не изгнал Хананеев, живущих в Газере; и жили Хананеи среди их в Газере.
JUDG|1|30|И Завулон не изгнал жителей Китрона и жителей Наглола, и жили Хананеи среди их и платили им дань.
JUDG|1|31|И Асир не изгнал жителей Акко и жителей Сидона и Ахлава, Ахзива, Хелвы, Афека и Рехова.
JUDG|1|32|И жил Асир среди Хананеев, жителей земли той, ибо не изгнал их.
JUDG|1|33|И Неффалим не изгнал жителей Вефсамиса и жителей Бефанафа и жил среди Хананеев, жителей земли той; жители же Вефсамиса и Бефанафа были его данниками.
JUDG|1|34|И стеснили Аморреи сынов Дановых в горах, ибо не давали им сходить на долину.
JUDG|1|35|И остались Аморреи жить на горе Херес, в Аиалоне и Шаалвиме; но рука сынов Иосифовых одолела [Аморреев], и сделались они данниками им.
JUDG|1|36|Пределы Аморреев от возвышенности Акравим и от Селы простирались и далее.
JUDG|2|1|И пришел Ангел Господень из Галгала в Бохим и сказал: Я вывел вас из Египта и ввел вас в землю, о которой клялся отцам вашим – [дать вам], и сказал Я: "не нарушу завета Моего с вами вовек;
JUDG|2|2|и вы не вступайте в союз с жителями земли сей; жертвенники их разрушьте". Но вы не послушали гласа Моего. Что вы это сделали?
JUDG|2|3|И потому говорю Я: не изгоню их от вас, и будут они вам петлею, и боги их будут для вас сетью.
JUDG|2|4|Когда Ангел Господень сказал слова сии всем сынам Израилевым, то народ поднял громкий вопль и заплакал.
JUDG|2|5|От сего и называют то место Бохим. Там принесли они жертву Господу.
JUDG|2|6|Когда Иисус распустил народ, и пошли сыны Израилевы, каждый в свой удел, чтобы получить в наследие землю,
JUDG|2|7|тогда народ служил Господу во все дни Иисуса и во все дни старейшин, которых жизнь продлилась после Иисуса и которые видели все великие дела Господни, какие Он сделал Израилю.
JUDG|2|8|Но когда умер Иисус, сын Навин, раб Господень, будучи ста десяти лет,
JUDG|2|9|и похоронили его в пределе удела его в Фамнаф–Сараи, на горе Ефремовой, на север от горы Гааша;
JUDG|2|10|и когда весь народ оный отошел к отцам своим, и восстал после них другой род, который не знал Господа и дел Его, какие Он делал Израилю, –
JUDG|2|11|тогда сыны Израилевы стали делать злое пред очами Господа и стали служить Ваалам;
JUDG|2|12|оставили Господа Бога отцов своих, Который вывел их из земли Египетской, и обратились к другим богам, богам народов, окружавших их, и стали поклоняться им, и раздражили Господа;
JUDG|2|13|оставили Господа и стали служить Ваалу и Астартам.
JUDG|2|14|И воспылал гнев Господень на Израиля, и предал их в руки грабителей, и грабили их; и предал их в руки врагов, окружавших их, и не могли уже устоять пред врагами своими.
JUDG|2|15|Куда они ни пойдут, рука Господня везде была им во зло, как говорил им Господь и как клялся им Господь. И им было весьма тесно.
JUDG|2|16|И воздвигал [им] Господь судей, которые спасали их от рук грабителей их;
JUDG|2|17|но и судей они не слушали, а ходили блудно вслед других богов и поклонялись им, скоро уклонялись от пути, коим ходили отцы их, повинуясь заповедям Господним. Они так не делали.
JUDG|2|18|Когда Господь воздвигал им судей, то Сам Господь был с судьею и спасал их от врагов их во все дни судьи: ибо жалел [их] Господь, слыша стон их от угнетавших и притеснявших их.
JUDG|2|19|Но как скоро умирал судья, они опять делали хуже отцов своих, уклоняясь к другим богам, служа им и поклоняясь им. Не отставали от дел своих и от стропотного пути своего.
JUDG|2|20|И воспылал гнев Господень на Израиля, и сказал Он: за то, что народ сей преступает завет Мой, который Я поставил с отцами их, и не слушает гласа Моего,
JUDG|2|21|и Я не стану уже изгонять от них ни одного из тех народов, которых оставил Иисус, когда умирал, –
JUDG|2|22|чтобы искушать ими Израиля: станут ли они держаться пути Господня и ходить по нему, как держались отцы их, или нет?
JUDG|2|23|И оставил Господь народы сии и не изгнал их вскоре и не предал их в руки Иисуса.
JUDG|3|1|Вот те народы, которых оставил Господь, чтобы искушать ими Израильтян, всех, которые не знали о всех войнах Ханаанских, –
JUDG|3|2|для того только, чтобы знали и учились войне последующие роды сынов Израилевых, которые прежде не знали ее:
JUDG|3|3|пять владельцев Филистимских, все Хананеи, Сидоняне и Евеи, живущие на горе Ливане, от горы Ваал–Ермона до входа в Емаф.
JUDG|3|4|Они были [оставлены], чтобы искушать ими Израильтян и узнать, повинуются ли они заповедям Господним, которые Он заповедал отцам их чрез Моисея.
JUDG|3|5|И жили сыны Израилевы среди Хананеев, Хеттеев, Аморреев, Ферезеев, Евеев, и Иевусеев,
JUDG|3|6|и брали дочерей их себе в жены, и своих дочерей отдавали за сыновей их, и служили богам их.
JUDG|3|7|И сделали сыны Израилевы злое пред очами Господа, и забыли Господа Бога своего, и служили Ваалам и Астартам.
JUDG|3|8|И воспылал гнев Господень на Израиля, и предал их в руки Хусарсафема, царя Месопотамского, и служили сыны Израилевы Хусарсафему восемь лет.
JUDG|3|9|Тогда возопили сыны Израилевы к Господу, и воздвигнул Господь спасителя сынам Израилевым, который спас их, Гофониила, сына Кеназа, младшего брата Халевова.
JUDG|3|10|На нем был Дух Господень, и был он судьею Израиля. Он вышел на войну, и предал Господь в руки его Хусарсафема, царя Месопотамского, и преодолела рука его Хусарсафема.
JUDG|3|11|И покоилась земля сорок лет. И умер Гофониил, сын Кеназа.
JUDG|3|12|Сыны Израилевы опять стали делать злое пред очами Господа, и укрепил Господь Еглона, царя Моавитского, против Израильтян, за то, что они делали злое пред очами Господа.
JUDG|3|13|Он собрал к себе Аммонитян и Амаликитян, и пошел и поразил Израиля, и овладели они городом Пальм.
JUDG|3|14|И служили сыны Израилевы Еглону, царю Моавитскому, восемнадцать лет.
JUDG|3|15|Тогда возопили сыны Израилевы к Господу, и Господь воздвигнул им спасителя Аода, сына Геры, сына Иеминиева, который был левша. И послали сыны Израилевы с ним дары Еглону, царю Моавитскому.
JUDG|3|16|Аод сделал себе меч с двумя остриями, длиною в локоть, и припоясал его под плащом своим к правому бедру,
JUDG|3|17|и поднес дары Еглону, царю Моавитскому; Еглон же был человек очень тучный.
JUDG|3|18|Когда поднес [Аод] все дары и проводил людей, принесших дары,
JUDG|3|19|то сам возвратился от истуканов, которые в Галгале, и сказал: у меня есть тайное слово до тебя, царь. Он сказал: тише! И вышли от него все стоявшие при нем.
JUDG|3|20|Аод вошел к нему: он сидел в прохладной горнице, которая была у него отдельно. И сказал Аод: у меня есть до тебя, слово Божие. [Еглон] встал со стула.
JUDG|3|21|Аод простер левую руку свою и взял меч с правого бедра своего и вонзил его в чрево его,
JUDG|3|22|так что вошла за острием и рукоять, и тук закрыл острие, ибо Аод не вынул меча из чрева его, и он прошел в задние части.
JUDG|3|23|И вышел Аод в преддверие, и затворил за собою двери горницы, и замкнул.
JUDG|3|24|Когда он вышел, рабы [Еглона] пришли и видят, вот, двери горницы замкнуты, и говорят: верно он для нужды в прохладной комнате.
JUDG|3|25|Ждали довольно долго, но видя, что никто не отпирает дверей горницы, взяли ключ и отперли, и вот, господин их лежит на земле мертвый.
JUDG|3|26|Пока они недоумевали, Аод между тем ушел, прошел мимо истуканов и спасся в Сеираф.
JUDG|3|27|Придя же вострубил трубою на горе Ефремовой, и сошли с ним сыны Израилевы с горы, и он [шел] впереди их.
JUDG|3|28|И сказал им: идите за мною, ибо предал Господь врагов ваших Моавитян в руки ваши. И пошли за ним, и перехватили переправу через Иордан к Моаву, и не давали никому переходить.
JUDG|3|29|И побили в то время Моавитян около десяти тысяч человек, все здоровых и сильных, и никто не убежал.
JUDG|3|30|Так смирились в тот день Моавитяне пред Израилем, и покоилась земля восемьдесят лет.
JUDG|3|31|После него был Самегар, сын Анафов, который шестьсот человек Филистимлян побил воловьим рожном; и он также спас Израиля.
JUDG|4|1|Когда умер Аод, сыны Израилевы стали опять делать злое пред очами Господа.
JUDG|4|2|И предал их Господь в руки Иавина, царя Ханаанского, который царствовал в Асоре; военачальником у него был Сисара, который жил в Харошеф–Гоиме.
JUDG|4|3|И возопили сыны Израилевы к Господу, ибо у него было девятьсот железных колесниц, и он жестоко угнетал сынов Израилевых двадцать лет.
JUDG|4|4|В то время была судьею Израиля Девора пророчица, жена Лапидофова;
JUDG|4|5|она жила под Пальмою Девориною, между Рамою и Вефилем, на горе Ефремовой; и приходили к ней сыны Израилевы на суд.
JUDG|4|6|[Девора] послала и призвала Варака, сына Авиноамова, из Кедеса Неффалимова, и сказала ему: повелевает [тебе] Господь Бог Израилев: пойди, взойди на гору Фавор и возьми с собою десять тысяч человек из сынов Неффалимовых и сынов Завулоновых;
JUDG|4|7|а Я приведу к тебе, к потоку Киссону, Сисару, военачальника Иавинова, и колесницы его и многолюдное [войско] его, и предам его в руки твои.
JUDG|4|8|Варак сказал ей: если ты пойдешь со мною, пойду; а если не пойдешь со мною, не пойду.
JUDG|4|9|Она сказала [ему]: пойти пойду с тобою; только не тебе уже будет слава на сем пути, в который ты идешь; но в руки женщины предаст Господь Сисару. И встала Девора и пошла с Вараком в Кедес.
JUDG|4|10|Варак созвал Завулонян и Неффалимлян в Кедес, и пошли вслед за ним десять тысяч человек, и Девора пошла с ним.
JUDG|4|11|Хевер Кенеянин отделился [тогда] от Кенеян, сынов Ховава, родственника Моисеева, и раскинул шатер свой у дубравы в Цаанниме близ Кедеса.
JUDG|4|12|И донесли Сисаре, что Варак, сын Авиноамов, взошел на гору Фавор.
JUDG|4|13|Сисара созвал все колесницы свои, девятьсот железных колесниц, и весь народ, который у него, из Харошеф–Гоима к потоку Киссону.
JUDG|4|14|И сказала Девора Вараку: встань, ибо это тот день, в который Господь предаст Сисару в руки твои; Сам Господь пойдет пред тобою. И сошел Варак с горы Фавора, и за ним десять тысяч человек.
JUDG|4|15|Тогда Господь привел в замешательство Сисару и все колесницы его и все ополчение его от меча Варакова, и сошел Сисара с колесницы и побежал пеший.
JUDG|4|16|Варак преследовал колесницы [его] и ополчение до Харошеф–Гоима, и пало все ополчение Сисарино от меча, не осталось никого.
JUDG|4|17|Сисара же убежал пеший в шатер Иаили, жены Хевера Кенеянина; ибо между Иавином, царем Асорским, и домом Хевера Кенеянина был мир.
JUDG|4|18|И вышла Иаиль навстречу Сисаре и сказала ему: зайди, господин мой, зайди ко мне, не бойся. Он зашел к ней в шатер, и она покрыла его ковром.
JUDG|4|19|[Сисара] сказал ей: дай мне немного воды напиться, я пить хочу. Она развязала мех с молоком, и напоила его и [опять] покрыла его.
JUDG|4|20|[Сисара] сказал ей: стань у дверей шатра, и если кто придет и спросит у тебя и скажет: "нет ли здесь кого?", ты скажи: "нет".
JUDG|4|21|Иаиль, жена Хеверова, взяла кол от шатра, и взяла молот в руку свою, и подошла к нему тихонько, и вонзила кол в висок его так, что приколола к земле; а он спал от усталости – и умер.
JUDG|4|22|И вот, Варак гонится за Сисарою. Иаиль вышла навстречу ему и сказала ему: войди, я покажу тебе человека, которого ты ищешь. Он вошел к ней, и вот, Сисара лежит мертвый, и кол в виске его.
JUDG|4|23|И смирил Бог в тот день Иавина, царя Ханаанского, пред сынами Израилевыми.
JUDG|4|24|Рука сынов Израилевых усиливалась более и более над Иавином, царем Ханаанским, доколе не истребили они Иавина, царя Ханаанского.
JUDG|5|1|В тот день воспела Девора и Варак, сын Авиноамов, сими словами:
JUDG|5|2|Израиль отмщен, народ показал рвение; прославьте Господа!
JUDG|5|3|Слушайте, цари, внимайте, вельможи: я Господу, я пою, бряцаю Господу Богу Израилеву.
JUDG|5|4|Когда выходил Ты, Господи, от Сеира, когда шел с поля Едомского, тогда земля тряслась, и небо капало, и облака проливали воду;
JUDG|5|5|горы таяли от лица Господа, даже этот Синай от лица Господа Бога Израилева.
JUDG|5|6|Во дни Самегара, сына Анафова, во дни Иаили, были пусты дороги, и ходившие прежде путями прямыми ходили тогда окольными дорогами.
JUDG|5|7|Не стало обитателей в селениях у Израиля, не стало, доколе не восстала я, Девора, доколе не восстала я, мать в Израиле.
JUDG|5|8|Избрали новых богов, от того война у ворот. Виден ли был щит и копье у сорока тысяч Израиля?
JUDG|5|9|Сердце мое к вам, начальники Израилевы, к ревнителям в народе; прославьте Господа!
JUDG|5|10|Ездящие на ослицах белых, сидящие на коврах и ходящие по дороге, пойте песнь!
JUDG|5|11|Среди голосов собирающих стада при колодезях, там да воспоют хвалу Господу, хвалу вождям Израиля! Тогда выступил ко вратам народ Господень.
JUDG|5|12|Воспряни, воспряни, Девора! воспряни, воспряни! воспой песнь! Восстань, Варак! и веди пленников твоих, сын Авиноамов!
JUDG|5|13|Тогда немногим из сильных подчинил Он народ; Господь подчинил мне храбрых.
JUDG|5|14|От Ефрема пришли укоренившиеся в земле Амалика; за тобою Вениамин, среди народа твоего; от Махира шли начальники, и от Завулона владеющие тростью писца.
JUDG|5|15|И князья Иссахаровы с Деворою, и Иссахар так же, как Варак, бросился в долину пеший. В племенах Рувимовых большое разногласие.
JUDG|5|16|Что сидишь ты между овчарнями, слушая блеяние стад? В племенах Рувимовых большое разногласие.
JUDG|5|17|Галаад живет [спокойно] за Иорданом, и Дану чего бояться с кораблями? Асир сидит на берегу моря и у пристаней своих живет спокойно.
JUDG|5|18|Завулон – народ, обрекший душу свою на смерть, и Неффалим – на высотах поля.
JUDG|5|19|Пришли цари, сразились, тогда сразились цари Ханаанские в Фанаахе у вод Мегиддонских, но не получили нимало серебра.
JUDG|5|20|С неба сражались, звезды с путей своих сражались с Сисарою.
JUDG|5|21|Поток Киссон увлек их, поток Кедумим, поток Киссон. Попирай, душа моя, силу!
JUDG|5|22|Тогда ломались копыта конские от побега, от побега сильных его.
JUDG|5|23|Прокляните Мероз, говорит Ангел Господень, прокляните, прокляните жителей его за то, что не пришли на помощь Господу, на помощь Господу с храбрыми.
JUDG|5|24|Да будет благословенна между женами Иаиль, жена Хевера Кенеянина, между женами в шатрах да будет благословенна!
JUDG|5|25|Воды просил он: молока подала она, в чаше вельможеской принесла молока лучшего.
JUDG|5|26|[Левую] руку свою протянула к колу, а правую свою к молоту работников; ударила Сисару, поразила голову его, разбила и пронзила висок его.
JUDG|5|27|К ногам ее склонился, пал и лежал, к ногам ее склонился, пал; где склонился, там и пал сраженный.
JUDG|5|28|В окно выглядывает и вопит мать Сисарина сквозь решетку: что долго не идет конница его, что медлят колеса колесниц его?
JUDG|5|29|Умные из ее женщин отвечают ей, и сама она отвечает на слова свои:
JUDG|5|30|верно, они нашли, делят добычу, по девице, по две девицы на каждого воина, в добычу полученная разноцветная [одежда] Сисаре, полученная в добычу разноцветная одежда, вышитая с обеих сторон, снятая с плеч пленника.
JUDG|5|31|Так да погибнут все враги Твои, Господи! Любящие же Его [да] [будут] как солнце, восходящее во всей силе своей! – И покоилась земля сорок лет.
JUDG|6|1|Сыны Израилевы стали [опять] делать злое пред очами Господа, и предал их Господь в руки Мадианитян на семь лет.
JUDG|6|2|Тяжела была рука Мадианитян над Израилем, и сыны Израилевы сделали себе от Мадианитян ущелья в горах и пещеры и укрепления.
JUDG|6|3|Когда посеет Израиль, придут Мадианитяне и Амаликитяне и жители востока и ходят у них;
JUDG|6|4|и стоят у них шатрами, и истребляют произведения земли до самой Газы, и не оставляют для пропитания Израилю ни овцы, ни вола, ни осла.
JUDG|6|5|Ибо они приходили со скотом своим и с шатрами своими, приходили в таком множестве, как саранча; им и верблюдам их не было числа, и ходили по земле Израилевой, чтоб опустошать ее.
JUDG|6|6|И весьма обнищал Израиль от Мадианитян, и возопили сыны Израилевы к Господу.
JUDG|6|7|И когда возопили сыны Израилевы к Господу на Мадианитян,
JUDG|6|8|послал Господь пророка к сынам Израилевым, и сказал им: так говорит Господь Бог Израилев: Я вывел вас из Египта, вывел вас из дома рабства;
JUDG|6|9|избавил вас из руки Египтян и из руки всех, угнетавших вас, прогнал их от вас, и дал вам землю их,
JUDG|6|10|и сказал вам: "Я – Господь Бог ваш; не чтите богов Аморрейских, в земле которых вы живете"; но вы не послушали гласа Моего.
JUDG|6|11|И пришел Ангел Господень и сел в Офре под дубом, принадлежащим Иоасу, потомку Авиезерову; сын его Гедеон выколачивал тогда пшеницу в точиле, чтобы скрыться от Мадианитян.
JUDG|6|12|И явился ему Ангел Господень и сказал ему: Господь с тобою, муж сильный!
JUDG|6|13|Гедеон сказал ему: господин мой! если Господь с нами, то отчего постигло нас все это? и где все чудеса Его, о которых рассказывали нам отцы наши, говоря: "из Египта вывел нас Господь"? Ныне оставил нас Господь и предал нас в руки Мадианитян.
JUDG|6|14|Господь, воззрев на него, сказал: иди с этою силою твоею и спаси Израиля от руки Мадианитян; Я посылаю тебя.
JUDG|6|15|[Гедеон] сказал ему: Господи! как спасу я Израиля? вот, и племя мое в [колене] Манассиином самое бедное, и я в доме отца моего младший.
JUDG|6|16|И сказал ему Господь: Я буду с тобою, и ты поразишь Мадианитян, как одного человека.
JUDG|6|17|[Гедеон] сказал Ему: если я обрел благодать пред очами Твоими, то сделай мне знамение, что Ты говоришь со мною:
JUDG|6|18|не уходи отсюда, доколе я не приду к Тебе и не принесу дара моего и не предложу Тебе. Он сказал: Я останусь до возвращения твоего.
JUDG|6|19|Гедеон пошел и приготовил козленка и опресноков из ефы муки; мясо положил в корзину, а похлебку влил в горшок и принес к Нему под дуб и предложил.
JUDG|6|20|И сказал ему Ангел Божий: возьми мясо и опресноки, и положи на сей камень, и вылей похлебку. Он так и сделал.
JUDG|6|21|Ангел Господень простер конец жезла, который был в руке его, прикоснулся к мясу и опреснокам; и вышел огонь из камня и поел мясо и опресноки; и Ангел Господень скрылся от глаз его.
JUDG|6|22|И увидел Гедеон, что это Ангел Господень, и сказал Гедеон: [увы] [мне], Владыка Господи! потому что я видел Ангела Господня лицем к лицу.
JUDG|6|23|Господь сказал ему: мир тебе, не бойся, не умрешь.
JUDG|6|24|И устроил там Гедеон жертвенник Господу и назвал его: Иегова Шалом. Он еще до сего дня в Офре Авиезеровой.
JUDG|6|25|В ту ночь сказал ему Господь: возьми тельца из стада отца твоего и другого тельца семилетнего, и разрушь жертвенник Ваала, который у отца твоего, и сруби священное дерево, которое при нем,
JUDG|6|26|и поставь жертвенник Господу Богу твоему, на вершине скалы сей, в порядке, и возьми второго тельца и принеси во всесожжение на дровах дерева, которое срубишь.
JUDG|6|27|Гедеон взял десять человек из рабов своих и сделал, как говорил ему Господь; но как сделать это днем он боялся домашних отца своего и жителей города, то сделал ночью.
JUDG|6|28|Поутру встали жители города, и вот, жертвенник Ваалов разрушен, и дерево при нем срублено, и второй телец вознесен во всесожжение на новоустроенном жертвеннике.
JUDG|6|29|И говорили друг другу: кто это сделал? Искали, расспрашивали и сказали: Гедеон, сын Иоасов, сделал это.
JUDG|6|30|И сказали жители города Иоасу: выведи сына твоего; он должен умереть за то, что разрушил жертвенник Ваала и срубил дерево, которое было при нем.
JUDG|6|31|Иоас сказал всем приступившим к нему: вам ли вступаться за Ваала, вам ли защищать его? кто вступится за него, тот будет предан смерти в это же утро; если он Бог, то пусть сам вступится за себя, потому что он разрушил его жертвенник.
JUDG|6|32|И стал звать его с того дня Иероваалом, потому что сказал: пусть Ваал сам судится с ним за то, что он разрушил жертвенник его.
JUDG|6|33|Между тем все Мадианитяне и Амаликитяне и жители востока собрались вместе, перешли [реку] и стали станом на долине Изреельской.
JUDG|6|34|И Дух Господень объял Гедеона; он вострубил трубою, и созвано было племя Авиезерово идти за ним.
JUDG|6|35|И послал послов по всему колену Манассиину, и оно вызвалось идти за ним; также послал послов к Асиру, Завулону и Неффалиму, и сии пришли навстречу им.
JUDG|6|36|И сказал Гедеон Богу: если Ты спасешь Израиля рукою моею, как говорил Ты,
JUDG|6|37|то вот, я расстелю [здесь] на гумне стриженую шерсть: если роса будет только на шерсти, а на всей земле сухо, то буду знать, что спасешь рукою моею Израиля, как говорил Ты.
JUDG|6|38|Так и сделалось: на другой день, встав рано, он стал выжимать шерсть и выжал из шерсти росы целую чашу воды.
JUDG|6|39|И сказал Гедеон Богу: не прогневайся на меня, если еще раз скажу и еще только однажды сделаю испытание над шерстью: пусть будет сухо на одной только шерсти, а на всей земле пусть будет роса.
JUDG|6|40|Бог так и сделал в ту ночь: только на шерсти было сухо, а на всей земле была роса.
JUDG|7|1|Иероваал, он же и Гедеон, встал поутру и весь народ, бывший с ним, и расположились станом у источника Харода; Мадиамский же стан был от него к северу у холма Море в долине.
JUDG|7|2|И сказал Господь Гедеону: народа с тобою слишком много, не могу Я предать Мадианитян в руки их, чтобы не возгордился Израиль предо Мною и не сказал: "моя рука спасла меня";
JUDG|7|3|итак провозгласи вслух народа и скажи: "кто боязлив и робок, тот пусть возвратится и пойдет назад с горы Галаада". И возвратилось народа двадцать две тысячи, а десять тысяч осталось.
JUDG|7|4|И сказал Господь Гедеону: все еще много народа; веди их к воде, там Я выберу их тебе; о ком Я скажу: "пусть идет с тобою", тот и пусть идет с тобою; а о ком скажу тебе: "не должен идти с тобою", тот пусть и не идет.
JUDG|7|5|Он привел народ к воде. И сказал Господь Гедеону: кто будет лакать воду языком своим, как лакает пес, того ставь особо, также и тех всех, которые будут наклоняться на колени свои и пить.
JUDG|7|6|И было число лакавших ртом своим с руки триста человек; весь же остальной народ наклонялся на колени свои пить воду.
JUDG|7|7|И сказал Господь Гедеону: тремя стами лакавших Я спасу вас и предам Мадианитян в руки ваши, а весь народ пусть идет, каждый в свое место.
JUDG|7|8|И взяли они съестной запас у народа себе и трубы их, и отпустил Гедеон всех Израильтян по шатрам и удержал у себя триста человек; стан же Мадиамский был у него внизу в долине.
JUDG|7|9|В ту ночь сказал ему Господь: встань, сойди в стан, Я предаю его в руки твои;
JUDG|7|10|если же ты боишься идти [один], то пойди в стан ты и Фура, слуга твой;
JUDG|7|11|и услышишь, что говорят, и тогда укрепятся руки твои, и пойдешь в стан. И сошел он и Фура, слуга его, к самому [полку] вооруженных, которые были в стане.
JUDG|7|12|Мадианитяне же и Амаликитяне и все жители востока расположились на долине в таком множестве, как саранча; верблюдам их не было числа, много было их, как песку на берегу моря.
JUDG|7|13|Гедеон пришел. И вот, один рассказывает другому сон и говорит: снилось мне, будто круглый ячменный хлеб катился по стану Мадиамскому и, прикатившись к шатру, ударил в него так, что он упал, опрокинул его, и шатер распался.
JUDG|7|14|Другой сказал в ответ ему: это не иное что, как меч Гедеона, сына Иоасова, Израильтянина; предал Бог в руки его Мадианитян и весь стан.
JUDG|7|15|Гедеон, услышав рассказ сна и толкование его, поклонился [Господу] и возвратился в стан Израильский и сказал: вставайте! предал Господь в руки ваши стан Мадиамский.
JUDG|7|16|И разделил триста человек на три отряда и дал в руки всем им трубы и пустые кувшины и в кувшины светильники.
JUDG|7|17|И сказал им: смотрите на меня и делайте то же; вот, я подойду к стану, и что буду делать, то и вы делайте;
JUDG|7|18|когда я и находящиеся со мною затрубим трубою, трубите и вы трубами вашими вокруг всего стана и кричите: [меч] Господа и Гедеона!
JUDG|7|19|И подошел Гедеон и сто человек с ним к стану, в начале средней стражи, и разбудили стражей, и затрубили трубами и разбили кувшины, которые были в руках их.
JUDG|7|20|И затрубили [все] три отряда трубами, и разбили кувшины, и держали в левой руке своей светильники, а в правой руке трубы, и трубили, и кричали: меч Господа и Гедеона!
JUDG|7|21|И стоял всякий на своем месте вокруг стана; и стали бегать во всем стане, и кричали, и обратились в бегство.
JUDG|7|22|Между тем как триста человек трубили трубами, обратил Господь меч одного на другого во всем стане, и бежало ополчение до Бефшитты к Царере, до предела Авелмехолы, близ Табафы.
JUDG|7|23|И созваны Израильтяне из колена Неффалимова, Асирова и всего колена Манассиина, и погнались за Мадианитянами.
JUDG|7|24|Гедеон же послал послов на всю гору Ефремову сказать: выйдите навстречу Мадианитянам и перехватите у них [переправу через] воду до Бефвары и Иордан. И созваны все Ефремляне и перехватили [переправы] [через] воду до Бефвары и Иордан;
JUDG|7|25|и поймали двух князей Мадиамских: Орива и Зива, и убили Орива в Цур–Ориве, а Зива в Иекев–Зиве и преследовали Мадианитян; головы же Орива и Зива принесли к Гедеону за Иордан.
JUDG|8|1|И сказали ему Ефремляне: зачем ты это сделал, что не позвал нас, когда шел воевать с Мадианитянами? И сильно ссорились с ним.
JUDG|8|2|[Гедеон] отвечал им: сделал ли я что такое, как вы ныне? Не счастливее ли Ефрем добирал виноград, нежели Авиезер обирал?
JUDG|8|3|В ваши руки предал Бог князей Мадиамских Орива и Зива, и что мог сделать я такое, как вы? Тогда успокоился дух их против него, когда сказал он им такие слова.
JUDG|8|4|И пришел Гедеон к Иордану, и перешел сам и триста человек, бывшие с ним. Они были утомлены, преследуя [врагов].
JUDG|8|5|И сказал он жителям Сокхофа: дайте хлеба народу, который идет за мною; они утомились, а я преследую Зевея и Салмана, царей Мадиамских.
JUDG|8|6|Князья Сокхофа сказали: разве рука Зевея и Салмана уже в твоей руке, чтобы нам войску твоему давать хлеб?
JUDG|8|7|И сказал Гедеон: за это, когда предаст Господь Зевея и Салмана в руки мои, я растерзаю тело ваше терновником пустынным и молотильными зубчатыми досками.
JUDG|8|8|Оттуда пошел он в Пенуэл и то же сказал жителям его, и жители Пенуэла отвечали ему то же, что отвечали жители Сокхофа.
JUDG|8|9|Он сказал и жителям Пенуэла: когда я возвращусь в мире, разрушу башню сию.
JUDG|8|10|Зевей же и Салман были в Каркоре и с ними их ополчение до пятнадцати тысяч, все, что осталось из всего ополчения жителей востока; пало же сто двадцать тысяч человек, обнажающих меч.
JUDG|8|11|Гедеон пошел к живущим в шатрах на восток от Новы и Иогбеги и поразил стан, когда стан стоял беспечно.
JUDG|8|12|Зевей и Салман побежали; он погнался за ними и схватил обоих царей Мадиамских, Зевея и Салмана, и весь стан привел в замешательство.
JUDG|8|13|И возвратился Гедеон, сын Иоаса, с войны от возвышенности Хереса.
JUDG|8|14|И захватил юношу из жителей Сокхофа и выспросил у него; и он написал ему князей и старейшин Сокхофских семьдесят семь человек.
JUDG|8|15|И пришел он к жителям Сокхофским, и сказал: вот Зевей и Салман, за которых вы посмеялись надо мною, говоря: разве рука Зевея и Салмана уже в твоей руке, чтобы нам давать хлеб утомившимся людям твоим?
JUDG|8|16|И взял старейшин города и терновник пустынный и зубчатые молотильные доски и наказал ими жителей Сокхофа;
JUDG|8|17|и башню Пенуэльскую разрушил, и перебил жителей города.
JUDG|8|18|И сказал Зевею и Салману: каковы были те, которых вы убили на Фаворе? Они сказали: они были такие, как ты, каждый имел вид сынов царских.
JUDG|8|19|[Гедеон] сказал: это были братья мои, сыны матери моей. Жив Господь! если бы вы оставили их в живых, я не убил бы вас.
JUDG|8|20|И сказал Иеферу, первенцу своему: встань, убей их. Но юноша не извлек меча своего, потому что боялся, так как был еще молод.
JUDG|8|21|И сказали Зевей и Салман: встань сам и порази нас, потому что по человеку и сила его. И встал Гедеон, и убил Зевея и Салмана, и взял пряжки, бывшие на шеях верблюдов их.
JUDG|8|22|И сказали Израильтяне Гедеону: владей нами ты и сын твой и сын сына твоего, ибо ты спас нас из руки Мадианитян.
JUDG|8|23|Гедеон сказал им: ни я не буду владеть вами, ни мой сын не будет владеть вами; Господь да владеет вами.
JUDG|8|24|И сказал им Гедеон: прошу у вас одного, дайте мне каждый по серьге из добычи своей. (Ибо у [неприятелей] много было золотых серег, потому что они были Измаильтяне.)
JUDG|8|25|Они сказали: дадим. И разостлали одежду и бросали туда каждый по серьге из добычи своей.
JUDG|8|26|Весу в золотых серьгах, которые он выпросил, было тысяча семьсот золотых [сиклей], кроме пряжек, пуговиц и пурпуровых одежд, которые были на царях Мадиамских, и кроме [золотых] цепочек, которые были на шее у верблюдов их.
JUDG|8|27|Из этого сделал Гедеон ефод и положил его в своем городе, в Офре, и стали все Израильтяне блудно ходить туда за ним, и был он сетью Гедеону и всему дому его.
JUDG|8|28|Так смирились Мадианитяне пред сынами Израиля и не стали уже поднимать головы своей, и покоилась земля сорок лет во дни Гедеона.
JUDG|8|29|И пошел Иероваал, сын Иоасов, и жил в доме своем.
JUDG|8|30|У Гедеона было семьдесят сыновей, происшедших от чресл его, потому что у него много было жен.
JUDG|8|31|Также и наложница, жившая в Сихеме, родила ему сына, и он дал ему имя Авимелех.
JUDG|8|32|И умер Гедеон, сын Иоасов, в глубокой старости, и погребен во гробе отца своего Иоаса, в Офре Авиезеровой.
JUDG|8|33|Когда умер Гедеон, сыны Израилевы опять стали блудно ходить вслед Ваалов и поставили себе богом Ваалверифа;
JUDG|8|34|и не вспомнили сыны Израилевы Господа Бога своего, Который избавлял их из руки всех врагов, окружавших их;
JUDG|8|35|и дому Иероваалову, [или] Гедеонову, не сделали милости за все благодеяния, какие он сделал Израилю.
JUDG|9|1|Авимелех, сын Иероваалов, пошел в Сихем к братьям матери своей и говорил им и всему племени отца матери своей, и сказал:
JUDG|9|2|внушите всем жителям Сихемским: что лучше для вас, чтобы владели вами все семьдесят сынов Иеровааловых, или чтобы владел один? и вспомните, что я кость ваша и плоть ваша.
JUDG|9|3|Братья матери его внушили о нем все сии слова жителям Сихемским; и склонилось сердце их к Авимелеху, ибо говорили они: он брат наш.
JUDG|9|4|И дали ему семьдесят [сиклей] серебра из дома Ваалверифа; Авимелех нанял на оные праздных и своевольных людей, которые и пошли за ним.
JUDG|9|5|И пришел он в дом отца своего в Офру и убил братьев своих, семьдесят сынов Иеровааловых, на одном камне. Остался только Иофам, младший сын Иероваалов, потому что скрылся.
JUDG|9|6|И собрались все жители Сихемские и весь дом Милло, и пошли и поставили царем Авимелеха у дуба, что близ Сихема.
JUDG|9|7|Когда рассказали об этом Иофаму, он пошел и стал на вершине горы Гаризима и, возвысив голос свой, кричал и говорил им: послушайте меня, жители Сихема, и послушает вас Бог!
JUDG|9|8|Пошли некогда дерева помазать над собою царя и сказали маслине: царствуй над нами.
JUDG|9|9|Маслина сказала им: оставлю ли я тук мой, которым чествуют богов и людей и пойду ли скитаться по деревам?
JUDG|9|10|И сказали дерева смоковнице: иди ты, царствуй над нами.
JUDG|9|11|Смоковница сказала им: оставлю ли я сладость мою и хороший плод мой и пойду ли скитаться по деревам?
JUDG|9|12|И сказали дерева виноградной лозе: иди ты, царствуй над нами.
JUDG|9|13|Виноградная лоза сказала им: оставлю ли я сок мой, который веселит богов и человеков, и пойду ли скитаться по деревам?
JUDG|9|14|Наконец сказали все дерева терновнику: иди ты, царствуй над нами.
JUDG|9|15|Терновник сказал деревам: если вы по истине поставляете меня царем над собою, то идите, покойтесь под тенью моею; если же нет, то выйдет огонь из терновника и пожжет кедры Ливанские.
JUDG|9|16|Итак смотрите, по истине ли и по правде ли вы поступили, поставив Авимелеха царем? И хорошо ли вы поступили с Иероваалом и домом его, и сообразно ли с его благодеяниями поступили вы?
JUDG|9|17|За вас отец мой сражался, не дорожил жизнью своею и избавил вас от руки Мадианитян;
JUDG|9|18|а вы теперь восстали против дома отца моего, и убили семьдесят сынов отца моего на одном камне, и поставили царем над жителями Сихемскими Авимелеха, сына рабыни его, потому что он брат ваш.
JUDG|9|19|Если вы ныне по истине и по правде поступили с Иероваалом и домом его, то радуйтесь об Авимелехе, и он пусть радуется о вас;
JUDG|9|20|если же нет, то да изыдет огонь от Авимелеха и да пожжет жителей Сихемских и весь дом Милло и да изыдет огонь от жителей Сихемских и от дома Милло, и да пожжет Авимелеха.
JUDG|9|21|И побежал Иофам, и убежал и пошел в Беэр, и жил там, [укрываясь] от брата своего Авимелеха.
JUDG|9|22|Авимелех же царствовал над Израилем три года.
JUDG|9|23|И послал Бог злого духа между Авимелехом и между жителями Сихема, и не стали покоряться жители Сихемские Авимелеху,
JUDG|9|24|дабы таким образом совершилось мщение за семьдесят сынов Иеровааловых, и кровь их обратилась на Авимелеха, брата их, который убил их, и на жителей Сихемских, которые подкрепили руки его, чтоб убить братьев своих.
JUDG|9|25|Жители Сихемские посадили против него в засаду людей на вершинах гор, которые грабили всякого проходящего мимо их по дороге. О сем донесено было Авимелеху.
JUDG|9|26|Пришел же и Гаал, сын Еведов, с братьями своими в Сихем, и ходили они по Сихему, и жители Сихемские положились на него.
JUDG|9|27|И вышли в поле, и собирали виноград свой, и давили в точилах, и делали праздники, ходили в дом бога своего, и ели и пили, и проклинали Авимелеха.
JUDG|9|28|Гаал, сын Еведов, говорил: кто Авимелех и что Сихем, чтобы нам служить ему? Не сын ли он Иероваалов, и не Зевул ли главный начальник его? Служите лучше потомкам Еммора, отца Сихемова, а ему для чего нам служить?
JUDG|9|29|Если бы кто дал народ сей в руки мои, я прогнал бы Авимелеха. И сказано было Авимелеху: умножь войско твое и выходи.
JUDG|9|30|Зевул, начальник города, услышал слова Гаала, сына Еведова, и воспылал гнев его.
JUDG|9|31|Он хитрым образом отправляет послов к Авимелеху, чтобы сказать: вот, Гаал, сын Еведов, и братья его пришли в Сихем, и вот, они возмущают против тебя город;
JUDG|9|32|итак, встань ночью, ты и народ, находящийся с тобою, и поставь засаду в поле;
JUDG|9|33|поутру же, при восхождении солнца, встань рано и приступи к городу; и когда он и народ, который у него, выйдут к тебе, тогда делай с ними, что может рука твоя.
JUDG|9|34|И встал ночью Авимелех и весь народ, находившийся с ним, и поставили в засаду у Сихема четыре отряда.
JUDG|9|35|Гаал, сын Еведов, вышел и стал у ворот городских; и встал Авимелех и народ, бывший с ним, из засады.
JUDG|9|36|Гаал, увидев народ, говорит Зевулу: вот, народ спускается с вершины гор. А Зевул сказал ему: тень гор тебе кажется людьми.
JUDG|9|37|Гаал опять говорил и сказал: вот, народ спускается с возвышенности, и один отряд идет от дуба Меонним.
JUDG|9|38|И сказал ему Зевул: где уста твои, которые говорили: "кто Авимелех, чтобы мы стали служить ему?" Это тот народ, который ты пренебрегал; выходи теперь и сразись с ним.
JUDG|9|39|И пошел Гаал впереди жителей Сихемских и сразился с Авимелехом.
JUDG|9|40|И погнался за ним Авимелех, и побежал он от него, и много пало убитых до самых ворот города.
JUDG|9|41|И остался Авимелех в Аруме, а Гаала и братьев его Зевул выгнал, чтоб они не жили в Сихеме.
JUDG|9|42|На другой день вышел народ в поле, и донесли о сем Авимелеху.
JUDG|9|43|Он взял свой народ и разделил его на три отряда и поставил в засаду в поле. И увидев, что народ вышел из города, восстал на них и побил их.
JUDG|9|44|Между тем как Авимелех и отряды, бывшие с ним, приступили и стали у ворот городских, другие два отряда напали на всех, бывших в поле, и убивали их.
JUDG|9|45|И сражался Авимелех с городом весь тот день, и взял город, и побил народ, бывший в нем, и разрушил город и засеял его солью.
JUDG|9|46|Услышав об этом, все бывшие в башне Сихемской ушли в башню капища [Ваал–Верифа].
JUDG|9|47|Авимелеху донесено, что собрались [туда] все бывшие в башне Сихемской.
JUDG|9|48|И пошел Авимелех на гору Селмон, сам и весь народ, бывший с ним, и взял Авимелех топоры с собою и нарубил сучьев древесных, и положил на плечи свои, и сказал народу, бывшему с ним: вы видели, что я делал; скорее делайте и вы то же, что я.
JUDG|9|49|И нарубил каждый из всего народа сучьев, и пошли за Авимелехом, и положили к башне, и сожгли посредством их башню огнем, и умерли все бывшие в башне Сихемской, около тысячи мужчин и женщин.
JUDG|9|50|Потом пошел Авимелех в Тевец и осадил Тевец и взял его.
JUDG|9|51|Среди города была крепкая башня, и убежали туда все мужчины и женщины и все жители города, и заперлись и взошли на кровлю башни.
JUDG|9|52|Авимелех пришел к башне и окружил ее и подошел к дверям башни, чтобы сжечь ее огнем.
JUDG|9|53|Тогда одна женщина бросила обломок жернова на голову Авимелеху и проломила ему череп.
JUDG|9|54|[Авимелех] тотчас призвал отрока, оруженосца своего, и сказал ему: обнажи меч твой и умертви меня, чтобы не сказали обо мне: женщина убила его. И пронзил его отрок его, и он умер.
JUDG|9|55|Израильтяне, видя, что умер Авимелех, пошли каждый в свое место.
JUDG|9|56|Так воздал Бог Авимелеху за злодеяние, которое он сделал отцу своему, убив семьдесят братьев своих.
JUDG|9|57|И все злодеяния жителей Сихемских обратил Бог на голову их; и постигло их проклятие Иофама, сына Иероваалова.
JUDG|10|1|После Авимелеха восстал для спасения Израиля Фола, сын Фуи, сына Додова, из колена Иссахарова. Он жил в Шамире на горе Ефремовой.
JUDG|10|2|Он был судьею Израиля двадцать три года, и умер, и погребен в Шамире.
JUDG|10|3|После него восстал Иаир из Галаада и был судьею Израиля двадцать два года.
JUDG|10|4|У него было тридцать сыновей, ездивших на тридцати молодых ослах, и тридцать городов было у них; их до сего дня называют селениями Иаира, что в земле Галаадской.
JUDG|10|5|И умер Иаир и погребен в Камоне.
JUDG|10|6|Сыны Израилевы продолжали делать злое пред очами Господа и служили Ваалам и Астартам, и богам Арамейским, и богам Сидонским, и богам Моавитским, и богам Аммонитским, и богам Филистимским; а Господа оставили и не служили Ему.
JUDG|10|7|И воспылал гнев Господа на Израиля, и Он предал их в руки Филистимлян и в руки Аммонитян;
JUDG|10|8|они теснили и мучили сынов Израилевых с того года восемнадцать лет, всех сынов Израилевых по ту сторону Иордана в земле Аморрейской, которая в Галааде.
JUDG|10|9|Наконец Аммонитяне перешли Иордан, чтобы вести войну с Иудою и Вениамином и с домом Ефремовым. И весьма тесно было сынам Израиля.
JUDG|10|10|И возопили сыны Израилевы к Господу, и говорили: согрешили мы пред Тобою, потому что оставили Бога нашего и служили Ваалам.
JUDG|10|11|И сказал Господь сынам Израилевым: не угнетали ли вас Египтяне, и Аморреи, и Аммонитяне, и Филистимляне,
JUDG|10|12|и Сидоняне, и Амаликитяне, и Моавитяне, и когда вы взывали ко Мне, не спасал ли Я вас от рук их?
JUDG|10|13|А вы оставили Меня и стали служить другим богам; за то Я не буду уже спасать вас:
JUDG|10|14|пойдите, взывайте к богам, которых вы избрали, пусть они спасают вас в тесное для вас время.
JUDG|10|15|И сказали сыны Израилевы Господу: согрешили мы; делай с нами все, что Тебе угодно, только избавь нас ныне.
JUDG|10|16|И отвергли от себя чужих богов и стали служить Господу. И не потерпела душа Его страдания Израилева.
JUDG|10|17|Аммонитяне собрались и расположились станом в Галааде; собрались также сыны Израилевы и стали станом в Массифе.
JUDG|10|18|Народ [и] князья Галаадские сказали друг другу: кто начнет войну против Аммонитян, тот будет начальником всех жителей Галаадских.
JUDG|11|1|Иеффай Галаадитянин был человек храбрый. Он был сын блудницы; от Галаада родился Иеффай.
JUDG|11|2|И жена Галаадова родила ему сыновей. Когда возмужали сыновья жены, изгнали они Иеффая, сказав ему: ты не наследник в доме отца нашего, потому что ты сын другой женщины.
JUDG|11|3|И убежал Иеффай от братьев своих и жил в земле Тов; и собрались к Иеффаю праздные люди и выходили с ним.
JUDG|11|4|Чрез несколько времени Аммонитяне пошли войною на Израиля.
JUDG|11|5|Во время войны Аммонитян с Израильтянами пришли старейшины Галаадские взять Иеффая из земли Тов
JUDG|11|6|и сказали Иеффаю: приди, будь у нас вождем, и сразимся с Аммонитянами.
JUDG|11|7|Иеффай сказал старейшинам Галаадским: не вы ли возненавидели меня и выгнали из дома отца моего? зачем же пришли ко мне ныне, когда вы в беде?
JUDG|11|8|Старейшины Галаадские сказали Иеффаю: для того мы теперь пришли к тебе, чтобы ты пошел с нами и сразился с Аммонитянами и был у нас начальником всех жителей Галаадских.
JUDG|11|9|И сказал Иеффай старейшинам Галаадским: если вы возвратите меня, чтобы сразиться с Аммонитянами, и Господь предаст мне их, то останусь ли я у вас начальником?
JUDG|11|10|Старейшины Галаадские сказали Иеффаю: Господь да будет свидетелем между нами, что мы сделаем по слову твоему!
JUDG|11|11|И пошел Иеффай со старейшинами Галаадскими, и народ поставил его над собою начальником и вождем, и Иеффай произнес все слова свои пред лицем Господа в Массифе.
JUDG|11|12|И послал Иеффай послов к царю Аммонитскому сказать: что тебе до меня, что ты пришел ко мне воевать на земле моей?
JUDG|11|13|Царь Аммонитский сказал послам Иеффая: Израиль, когда шел из Египта, взял землю мою от Арнона до Иавока и Иордана; итак возврати мне ее с миром.
JUDG|11|14|Иеффай в другой раз послал послов к царю Аммонитскому,
JUDG|11|15|сказать ему: так говорит Иеффай: Израиль не взял земли Моавитской и земли Аммонитской;
JUDG|11|16|ибо когда шли из Египта, Израиль пошел в пустыню к Чермному морю и пришел в Кадес;
JUDG|11|17|оттуда послал Израиль послов к царю Едомскому сказать: "позволь мне пройти землею твоею"; но царь Едомский не послушал; и к царю Моавитскому он посылал, но и тот не согласился; посему Израиль оставался в Кадесе.
JUDG|11|18|И пошел пустынею, и миновал землю Едомскую и землю Моавитскую, и, придя к восточному пределу земли Моавитской, расположился станом за Арноном; но не входил в пределы Моавитские, ибо Арнон есть предел Моава.
JUDG|11|19|И послал Израиль послов к Сигону, царю Аморрейскому, царю Есевонскому, и сказал ему Израиль: позволь нам пройти землею твоею в свое место.
JUDG|11|20|Но Сигон не согласился пропустить Израиля чрез пределы свои, и собрал Сигон весь народ свой, и расположился станом в Иааце, и сразился с Израилем.
JUDG|11|21|И предал Господь Бог Израилев Сигона и весь народ его в руки Израилю, и он побил их; и получил Израиль в наследие всю землю Аморрея, жившего в земле той;
JUDG|11|22|и получили они в наследие все пределы Аморрея от Арнона до Иавока и от пустыни до Иордана.
JUDG|11|23|Итак Господь Бог Израилев изгнал Аморрея от лица народа Своего Израиля, а ты хочешь взять его наследие?
JUDG|11|24|Не владеешь ли ты тем, что дал тебе Хамос, бог твой? И мы владеем всем тем, что дал нам в наследие Господь Бог наш.
JUDG|11|25|Разве ты лучше Валака, сына Сепфорова, царя Моавитского? Ссорился ли он с Израилем, или воевал ли с ними?
JUDG|11|26|Израиль уже живет триста лет в Есевоне и в зависящих от него [городах], в Ароере и зависящих от него [городах], и во всех городах, которые близ Арнона; для чего вы в то время не отнимали [их]?
JUDG|11|27|А я не виновен пред тобою, и ты делаешь мне зло, выступив против меня войною. Господь Судия да будет ныне судьею между сынами Израиля и между Аммонитянами!
JUDG|11|28|Но царь Аммонитский не послушал слов Иеффая, с которыми он посылал к нему.
JUDG|11|29|И был на Иеффае Дух Господень, и прошел он Галаад и Манассию, и прошел Массифу Галаадскую, и из Массифы Галаадской пошел к Аммонитянам.
JUDG|11|30|И дал Иеффай обет Господу и сказал: если Ты предашь Аммонитян в руки мои,
JUDG|11|31|то по возвращении моем с миром от Аммонитян, что выйдет из ворот дома моего навстречу мне, будет Господу, и вознесу сие на всесожжение.
JUDG|11|32|И пришел Иеффай к Аммонитянам – сразиться с ними, и предал их Господь в руки его;
JUDG|11|33|и поразил их поражением весьма великим, от Ароера до Минифа двадцать городов, и до Авель–Керамима, и смирились Аммонитяне пред сынами Израилевыми.
JUDG|11|34|И пришел Иеффай в Массифу в дом свой, и вот, дочь его выходит навстречу ему с тимпанами и ликами: она была у него только одна, и не было у него еще ни сына, ни дочери.
JUDG|11|35|Когда он увидел ее, разодрал одежду свою и сказал: ах, дочь моя! ты сразила меня; и ты в числе нарушителей покоя моего! я отверз [о тебе] уста мои пред Господом и не могу отречься.
JUDG|11|36|Она сказала ему: отец мой! ты отверз уста твои пред Господом – и делай со мною то, что произнесли уста твои, когда Господь совершил чрез тебя отмщение врагам твоим Аммонитянам.
JUDG|11|37|И сказала отцу своему: сделай мне только вот что: отпусти меня на два месяца; я пойду, взойду на горы и оплачу девство мое с подругами моими.
JUDG|11|38|Он сказал: пойди. И отпустил ее на два месяца. Она пошла с подругами своими и оплакивала девство свое в горах.
JUDG|11|39|По прошествии двух месяцев она возвратилась к отцу своему, и он совершил над нею обет свой, который дал, и она не познала мужа. И вошло в обычай у Израиля,
JUDG|11|40|что ежегодно дочери Израилевы ходили оплакивать дочь Иеффая Галаадитянина, четыре дня в году.
JUDG|12|1|Ефремляне собрались и перешли в Севину и сказали Иеффаю: для чего ты ходил воевать с Аммонитянами, а нас не позвал с собою? мы сожжем дом твой огнем и с тобою вместе.
JUDG|12|2|Иеффай сказал им: я и народ мой имели с Аммонитянами сильную ссору; я звал вас, но вы не спасли меня от руки их;
JUDG|12|3|видя, что ты не спасаешь меня, я подверг опасности жизнь мою и пошел на Аммонитян, и предал их Господь в руки мои; зачем же вы пришли ныне воевать со мною?
JUDG|12|4|И собрал Иеффай всех жителей Галаадских и сразился с Ефремлянами, и побили жители Галаадские Ефремлян, говоря: вы беглецы Ефремовы, Галаад же среди Ефрема и среди Манассии.
JUDG|12|5|И перехватили Галаадитяне переправу чрез Иордан от Ефремлян, и когда кто из уцелевших Ефремлян говорил: "позвольте мне переправиться", то жители Галаадские говорили ему: не Ефремлянин ли ты? Он говорил: нет.
JUDG|12|6|Они говорили ему "скажи: шибболет", а он говорил: "сибболет", и не мог иначе выговорить. Тогда они, взяв его, заколали у переправы чрез Иордан. И пало в то время из Ефремлян сорок две тысячи.
JUDG|12|7|Иеффай был судьею Израиля шесть лет, и умер Иеффай Галаадитянин и погребен в одном из городов Галаадских.
JUDG|12|8|После него был судьею Израиля Есевон из Вифлеема.
JUDG|12|9|У него было тридцать сыновей, и тридцать дочерей отпустил он из дома [в замужество], а тридцать дочерей взял со стороны за сыновей своих, и был судьею Израиля семь лет.
JUDG|12|10|И умер Есевон и погребен в Вифлееме.
JUDG|12|11|После него был судьею Израиля Елон Завулонянин и судил Израиля десять лет.
JUDG|12|12|И умер Елон Завулонянин и погребен в Аиалоне, в земле Завулоновой.
JUDG|12|13|После него был судьею Израиля Авдон, сын Гиллела, Пирафонянин.
JUDG|12|14|У него было сорок сыновей и тридцать внуков, ездивших на семидесяти молодых ослах; он судил Израиля восемь лет.
JUDG|12|15|И умер Авдон, сын Гиллела, Пирафонянин, и погребен в Пирафоне в земле Ефремовой, на горе Амаликовой.
JUDG|13|1|Сыны Израилевы продолжали делать злое пред очами Господа, и предал их Господь в руки Филистимлян на сорок лет.
JUDG|13|2|В то время был человек из Цоры, от племени Данова, именем Маной; жена его была неплодна и не рождала.
JUDG|13|3|И явился Ангел Господень жене и сказал ей: вот, ты неплодна и не рождаешь; но зачнешь, и родишь сына;
JUDG|13|4|итак берегись, не пей вина и сикера, и не ешь ничего нечистого;
JUDG|13|5|ибо вот, ты зачнешь и родишь сына, и бритва не коснется головы его, потому что от самого чрева младенец сей будет назорей Божий, и он начнет спасать Израиля от руки Филистимлян.
JUDG|13|6|Жена пришла и сказала мужу своему: человек Божий приходил ко мне, которого вид, как вид Ангела Божия, весьма почтенный; я не спросила его, откуда он, и он не сказал мне имени своего;
JUDG|13|7|он сказал мне: "вот, ты зачнешь и родишь сына; итак не пей вина и сикера и не ешь ничего нечистого, ибо младенец от самого чрева до смерти своей будет назорей Божий".
JUDG|13|8|Маной помолился Господу и сказал: Господи! пусть придет опять к нам человек Божий, которого посылал Ты, и научит нас, что нам делать с имеющим родиться младенцем.
JUDG|13|9|И услышал Бог голос Маноя, и Ангел Божий опять пришел к жене, когда она была в поле, и Маноя, мужа ее, не было с нею.
JUDG|13|10|Жена тотчас побежала и известила мужа своего и сказала ему: вот, явился мне человек, приходивший ко мне тогда.
JUDG|13|11|Маной встал и пошел с женою своею, и пришел к тому человеку и сказал ему: ты ли тот человек, который говорил с сею женщиною? [Ангел] сказал: я.
JUDG|13|12|И сказал Маной: итак, если исполнится слово твое, как нам поступать с младенцем сим и что делать с ним?
JUDG|13|13|Ангел Господень сказал Маною: пусть он остерегается всего, о чем я сказал жене;
JUDG|13|14|пусть не ест ничего, что производит виноградная лоза; пусть не пьет вина и сикера и не ест ничего нечистого и соблюдает все, что я приказал ей.
JUDG|13|15|И сказал Маной Ангелу Господню: позволь удержать тебя, пока мы изготовим для тебя козленка.
JUDG|13|16|Ангел Господень сказал Маною: хотя бы ты и удержал меня, но я не буду есть хлеба твоего; если же хочешь совершить всесожжение Господу, то вознеси его. Маной же не знал, что это Ангел Господень.
JUDG|13|17|И сказал Маной Ангелу Господню: как тебе имя? чтобы нам прославить тебя, когда исполнится слово твое.
JUDG|13|18|Ангел Господень сказал ему: что ты спрашиваешь об имени моем? оно чудно.
JUDG|13|19|И взял Маной козленка и хлебное приношение и вознес Господу на камне. И сделал Он чудо, которое видели Маной и жена его.
JUDG|13|20|Когда пламень стал подниматься от жертвенника к небу, Ангел Господень поднялся в пламени жертвенника. Видя это, Маной и жена его пали лицем на землю.
JUDG|13|21|И невидим стал Ангел Господень Маною и жене его. Тогда Маной узнал, что это Ангел Господень.
JUDG|13|22|И сказал Маной жене своей: верно мы умрем, ибо видели мы Бога.
JUDG|13|23|Жена его сказала ему: если бы Господь хотел умертвить нас, то не принял бы от рук наших всесожжения и хлебного приношения, и не показал бы нам всего того, и теперь не открыл бы нам сего.
JUDG|13|24|И родила жена сына, и нарекла имя ему: Самсон. И рос младенец, и благословлял его Господь.
JUDG|13|25|И начал Дух Господень действовать в нем в стане Дановом, между Цорою и Естаолом.
JUDG|14|1|И пошел Самсон в Фимнафу и увидел в Фимнафе женщину из дочерей Филистимских.
JUDG|14|2|Он пошел и объявил отцу своему и матери своей и сказал: я видел в Фимнафе женщину из дочерей Филистимских; возьмите ее мне в жену.
JUDG|14|3|Отец и мать его сказали ему: разве нет женщин между дочерями братьев твоих и во всем народе моем, что ты идешь взять жену у Филистимлян необрезанных? И сказал Самсон отцу своему: ее возьми мне, потому что она мне понравилась.
JUDG|14|4|Отец его и мать его не знали, что это от Господа, и что он ищет случая [отмстить] Филистимлянам. А в то время Филистимляне господствовали над Израилем.
JUDG|14|5|И пошел Самсон с отцом своим и с матерью своею в Фимнафу, и когда подходили к виноградникам Фимнафским, вот, молодой лев рыкая [идет] навстречу ему.
JUDG|14|6|И сошел на него Дух Господень, и он растерзал [льва] как козленка; а в руке у него ничего не было. И не сказал отцу своему и матери своей, что он сделал.
JUDG|14|7|И пришел и поговорил с женщиною, и она понравилась Самсону.
JUDG|14|8|Спустя несколько дней, опять пошел он, чтобы взять ее, и зашел посмотреть труп льва, и вот, рой пчел в трупе львином и мед.
JUDG|14|9|Он взял его в руки свои и пошел, и ел дорогою; и когда пришел к отцу своему и матери своей, дал и им, и они ели; но не сказал им, что из львиного трупа взял мед сей.
JUDG|14|10|И пришел отец его к женщине, и сделал там Самсон пир, как обыкновенно делают женихи.
JUDG|14|11|И как там увидели его, выбрали тридцать брачных друзей, которые были бы при нем.
JUDG|14|12|И сказал им Самсон: загадаю я вам загадку; если вы отгадаете мне ее в семь дней пира и отгадаете верно, то я дам вам тридцать синдонов и тридцать перемен одежд;
JUDG|14|13|если же не сможете отгадать мне, то вы дайте мне тридцать синдонов и тридцать перемен одежд. Они сказали ему: загадай загадку твою, послушаем.
JUDG|14|14|И сказал им: из ядущего вышло ядомое, и из сильного вышло сладкое. И не могли отгадать загадку в три дня.
JUDG|14|15|В седьмой день сказали они жене Самсоновой: уговори мужа твоего, чтоб он разгадал нам загадку; иначе сожжем огнем тебя и дом отца твоего; разве вы призвали нас, чтоб обобрать нас?
JUDG|14|16|И плакала жена Самсонова пред ним и говорила: ты ненавидишь меня и не любишь; ты загадал загадку сынам народа моего, а мне не разгадаешь ее. Он сказал ей: отцу моему и матери моей не разгадал ее; и тебе ли разгадаю?
JUDG|14|17|И плакала она пред ним семь дней, в которые продолжался у них пир. Наконец в седьмой день разгадал ей, ибо она усиленно просила его. А она разгадала загадку сынам народа своего.
JUDG|14|18|И в седьмой день до захождения солнечного сказали ему граждане: что слаще меда, и что сильнее льва! Он сказал им: если бы вы не орали на моей телице, то не отгадали бы моей загадки.
JUDG|14|19|И сошел на него Дух Господень, и пошел он в Аскалон, и, убив там тридцать человек, снял с них одежды, и отдал перемены [платья] их разгадавшим загадку. И воспылал гнев его, и ушел он в дом отца своего.
JUDG|14|20|А жена Самсонова вышла за брачного друга его, который был при нем другом.
JUDG|15|1|Чрез несколько дней, во время жатвы пшеницы, пришел Самсон повидаться с женою своею, принеся с собою козленка; и когда сказал: "войду к жене моей в спальню", отец ее не дал ему войти.
JUDG|15|2|И сказал отец ее: я подумал, что ты возненавидел ее, и я отдал ее другу твоему; вот, меньшая сестра красивее ее; пусть она будет тебе вместо ее.
JUDG|15|3|Но Самсон сказал им: теперь я буду прав пред Филистимлянами, если сделаю им зло.
JUDG|15|4|И пошел Самсон, и поймал триста лисиц, и взял факелы, и связал хвост с хвостом, и привязал по факелу между двумя хвостами;
JUDG|15|5|и зажег факелы, и пустил их на жатву Филистимскую, и выжег и копны и нежатый хлеб, и виноградные сады [и] масличные.
JUDG|15|6|И говорили Филистимляне: кто это сделал? И сказали: Самсон, зять Фимнафянина, ибо этот взял жену его и отдал другу его. И пошли Филистимляне и сожгли огнем ее и отца ее.
JUDG|15|7|Самсон сказал им: хотя вы сделали это, но я отмщу вам самим и тогда только успокоюсь.
JUDG|15|8|И перебил он им голени и бедра, и пошел и засел в ущелье скалы Етама.
JUDG|15|9|И пошли Филистимляне, и расположились станом в Иудее, и протянулись до Лехи.
JUDG|15|10|И сказали жители Иудеи: за что вы вышли против нас? Они сказали: мы пришли связать Самсона, чтобы поступить с ним, как он поступил с нами.
JUDG|15|11|И пошли три тысячи человек из Иудеи к ущелью скалы Етама и сказали Самсону: разве ты не знаешь, что Филистимляне господствуют над нами? что ты это сделал нам? Он сказал им: как они со мною поступили, так и я поступил с ними.
JUDG|15|12|И сказали ему: мы пришли связать тебя, чтобы отдать тебя в руки Филистимлянам. И сказал им Самсон: поклянитесь мне, что вы не убьете меня.
JUDG|15|13|И сказали ему: нет, мы только свяжем тебя и отдадим тебя в руки их, а умертвить не умертвим. И связали его двумя новыми веревками и повели его из ущелья.
JUDG|15|14|Когда он подошел к Лехе, Филистимляне с криком встретили его. И сошел на него Дух Господень, и веревки, бывшие на руках его, сделались, как перегоревший лен, и упали узы его с рук его.
JUDG|15|15|Нашел он свежую ослиную челюсть и, протянув руку свою, взял ее, и убил ею тысячу человек.
JUDG|15|16|И сказал Самсон: челюстью ослиною толпу, две толпы, челюстью ослиною убил я тысячу человек.
JUDG|15|17|Сказав это, бросил челюсть из руки своей и назвал то место: Рамаф–Лехи.
JUDG|15|18|И почувствовал сильную жажду и воззвал к Господу и сказал: Ты соделал рукою раба Твоего великое спасение сие; а теперь умру я от жажды, и попаду в руки необрезанных.
JUDG|15|19|И разверз Бог ямину в Лехе, и потекла из нее вода. Он напился, и возвратился дух его, и он ожил; от того и наречено имя месту сему: "Источник взывающего", который в Лехе до сего дня.
JUDG|15|20|И был он судьею Израиля во дни Филистимлян двадцать лет.
JUDG|16|1|Пришел однажды Самсон в Газу и, увидев там блудницу, вошел к ней.
JUDG|16|2|Жителям Газы сказали: Самсон пришел сюда. И ходили они кругом, и подстерегали его всю ночь в воротах города, и таились всю ночь, говоря: до света утреннего [подождем, и] убьем его.
JUDG|16|3|А Самсон спал до полуночи; в полночь же встав, схватил двери городских ворот с обоими косяками, поднял их вместе с запором, положил на плечи свои и отнес их на вершину горы, которая на пути к Хеврону.
JUDG|16|4|После того полюбил он одну женщину, жившую на долине Сорек; имя ей Далида.
JUDG|16|5|К ней пришли владельцы Филистимские и говорят ей: уговори его, и выведай, в чем великая сила его и как нам одолеть его, чтобы связать его и усмирить его; а мы дадим тебе за то каждый тысячу сто [сиклей] серебра.
JUDG|16|6|И сказала Далида Самсону: скажи мне, в чем великая сила твоя и чем связать тебя, чтобы усмирить тебя?
JUDG|16|7|Самсон сказал ей: если свяжут меня семью сырыми тетивами, которые не засушены, то я сделаюсь бессилен и буду как и прочие люди.
JUDG|16|8|И принесли ей владельцы Филистимские семь сырых тетив, которые не засохли, и она связала его ими.
JUDG|16|9|(Между тем один скрытно сидел у нее в спальне.) И сказала ему: Самсон! Филистимляне [идут] на тебя. Он разорвал тетивы, как разрывают нитку из пакли, когда пережжет ее огонь. И не узнана сила его.
JUDG|16|10|И сказала Далида Самсону: вот, ты обманул меня и говорил мне ложь; скажи же теперь мне, чем связать тебя?
JUDG|16|11|Он сказал ей: если свяжут меня новыми веревками, которые не были в деле, то я сделаюсь бессилен и буду, как прочие люди.
JUDG|16|12|Далида взяла новые веревки и связала его и сказала ему: Самсон! Филистимляне [идут] на тебя. (Между тем один скрытно сидел в спальне.) И сорвал он их с рук своих, как нитки.
JUDG|16|13|И сказала Далида Самсону: все ты обманываешь меня и говоришь мне ложь; скажи мне, чем бы связать тебя? Он сказал ей: если ты воткешь семь кос головы моей в ткань [и прибьешь ее гвоздем к ткальной колоде].
JUDG|16|14|и прикрепила их к колоде, и сказала ему: Филистимляне [идут] на тебя, Самсон! Он пробудился от сна своего и выдернул ткальную колоду вместе с тканью.
JUDG|16|15|И сказала ему [Далида]: как же ты говоришь: "люблю тебя", а сердце твое не со мною? вот, ты трижды обманул меня, и не сказал мне, в чем великая сила твоя.
JUDG|16|16|И как она словами своими тяготила его всякий день и мучила его, то душе его тяжело стало до смерти.
JUDG|16|17|И он открыл ей все сердце свое, и сказал ей: бритва не касалась головы моей, ибо я назорей Божий от чрева матери моей; если же остричь меня, то отступит от меня сила моя; я сделаюсь слаб и буду, как прочие люди.
JUDG|16|18|Далида, видя, что он открыл ей все сердце свое, послала и звала владельцев Филистимских, сказав им: идите теперь; он открыл мне все сердце свое. И пришли к ней владельцы Филистимские и принесли серебро в руках своих.
JUDG|16|19|И усыпила его [Далида] на коленях своих, и призвала человека, и велела ему остричь семь кос головы его. И начал он ослабевать, и отступила от него сила его.
JUDG|16|20|Она сказала: Филистимляне [идут] на тебя, Самсон! Он пробудился от сна своего, и сказал: пойду, как и прежде, и освобожусь. А не знал, что Господь отступил от него.
JUDG|16|21|Филистимляне взяли его и выкололи ему глаза, привели его в Газу и оковали его двумя медными цепями, и он молол в доме узников.
JUDG|16|22|Между тем волосы на голове его начали расти, где они были острижены.
JUDG|16|23|Владельцы Филистимские собрались, чтобы принести великую жертву Дагону, богу своему, и повеселиться, и сказали: бог наш предал Самсона, врага нашего, в руки наши.
JUDG|16|24|Также и народ, видя его, прославлял бога своего, говоря: бог наш предал в руки наши врага нашего и опустошителя земли нашей, который побил многих из нас.
JUDG|16|25|И когда развеселилось сердце их, сказали: позовите Самсона, пусть он позабавит нас. И призвали Самсона из дома узников, и он забавлял их, и поставили его между столбами.
JUDG|16|26|И сказал Самсон отроку, который водил его за руку: подведи меня, чтобы ощупать мне столбы, на которых утвержден дом, и прислониться к ним.
JUDG|16|27|Дом же был полон мужчин и женщин; там были все владельцы Филистимские, и на кровле было до трех тысяч мужчин и женщин, смотревших на забавляющего [их] Самсона.
JUDG|16|28|И воззвал Самсон к Господу и сказал: Господи Боже! вспомни меня и укрепи меня только теперь, о Боже! чтобы мне в один раз отмстить Филистимлянам за два глаза мои.
JUDG|16|29|И сдвинул Самсон с места два средних столба, на которых утвержден был дом, упершись в них, в один правою рукою своею, а в другой левою.
JUDG|16|30|И сказал Самсон: умри, душа моя, с Филистимлянами! И уперся [всею] силою, и обрушился дом на владельцев и на весь народ, бывший в нем. И было умерших, которых умертвил [Самсон] при смерти своей, более, нежели сколько умертвил он в жизни своей.
JUDG|16|31|И пришли братья его и весь дом отца его, и взяли его, и пошли и похоронили его между Цорою и Естаолом, во гробе Маноя, отца его. Он был судьею Израиля двадцать лет.
JUDG|17|1|Был некто на горе Ефремовой, именем Миха.
JUDG|17|2|Он сказал матери своей: тысяча сто [сиклей] серебра, которые у тебя взяты и за которые ты при мне изрекла проклятие, это серебро у меня, я взял его. Мать его сказала: благословен сын мой у Господа!
JUDG|17|3|И возвратил он матери своей тысячу сто [сиклей] серебра. И сказала мать его: это серебро я от себя посвятила Господу для сына моего, чтобы сделать из него истукан и литый кумир; итак отдаю оное тебе.
JUDG|17|4|Но он возвратил серебро матери своей. Мать его взяла двести [сиклей] серебра и отдала их плавильщику. Он сделал из них истукан и литый кумир, который и находился в доме Михи.
JUDG|17|5|И был у Михи дом Божий. И сделал он ефод и терафим и посвятил одного из сыновей своих, чтоб он был у него священником.
JUDG|17|6|В те дни не было царя у Израиля; каждый делал то, что ему казалось справедливым.
JUDG|17|7|Один юноша из Вифлеема Иудейского, из колена Иудина, левит, тогда жил там;
JUDG|17|8|этот человек пошел из города Вифлеема Иудейского, чтобы пожить, где случится, и идя дорогою, пришел на гору Ефремову к дому Михи.
JUDG|17|9|И сказал ему Миха: откуда ты идешь? Он сказал ему: я левит из Вифлеема Иудейского и иду пожить, где случится.
JUDG|17|10|И сказал ему Миха: останься у меня и будь у меня отцом и священником; я буду давать тебе по десяти [сиклей] серебра на год, потребное одеяние и пропитание.
JUDG|17|11|Левит пошел к нему и согласился левит остаться у этого человека, и был юноша у него, как один из сыновей его.
JUDG|17|12|Миха посвятил левита, и этот юноша был у него священником и жил в доме у Михи.
JUDG|17|13|И сказал Миха: теперь я знаю, что Господь будет мне благотворить, потому что левит у меня священником.
JUDG|18|1|В те дни не было царя у Израиля; и в те дни колено Даново искало себе удела, где бы поселиться, потому что дотоле не выпало ему [полного] удела между коленами Израилевыми.
JUDG|18|2|И послали сыны Дановы от племени своего пять человек, мужей сильных, из Цоры и Естаола, чтоб осмотреть землю и узнать ее, и сказали им: пойдите, узнайте землю. Они пришли на гору Ефремову к дому Михи и ночевали там.
JUDG|18|3|Находясь у дома Михи, узнали они голос молодого левита и зашли туда и спрашивали его: кто тебя привел сюда? что ты здесь делаешь и зачем ты здесь?
JUDG|18|4|Он сказал им: то и то сделал для меня Миха, нанял меня, и я у него священником.
JUDG|18|5|Они сказали ему: вопроси Бога, чтобы знать нам, успешен ли будет путь наш, в который мы идем.
JUDG|18|6|Священник сказал им: идите с миром; пред Господом путь ваш, в который вы идете.
JUDG|18|7|И пошли те пять мужей, и пришли в Лаис, и увидели народ, который в нем, что он живет покойно, по обычаю Сидонян, тих и беспечен, и что не было в земле той, кто обижал бы в чем, или имел бы власть: от Сидонян они жили далеко, и ни с кем не было у них никакого дела.
JUDG|18|8|И возвратились к братьям своим в Цору и Естаол, и сказали им братья их: с чем вы?
JUDG|18|9|Они сказали: встанем и пойдем на них; мы видели землю, она весьма хороша; а вы задумались: не медлите пойти и взять в наследие ту землю;
JUDG|18|10|когда пойдете вы, придете к народу беспечному, и земля та обширна; Бог предает ее в руки ваши; это такое место, где нет ни в чем недостатка, что [получается] от земли.
JUDG|18|11|И отправились оттуда из колена Данова, из Цоры и Естаола, шестьсот мужей, препоясавшись воинским оружием.
JUDG|18|12|Они пошли и стали станом в Кириаф–Иариме, в Иудее. Посему и называют то место станом Дановым до сего дня. Он позади Кириаф–Иарима.
JUDG|18|13|Оттуда отправились они на гору Ефремову и пришли к дому Михи.
JUDG|18|14|И сказали те пять мужей, которые ходили осматривать землю Лаис, братьям своим: знаете ли, что в одном из домов сих есть ефод, терафим, истукан и литый кумир? итак подумайте, что сделать.
JUDG|18|15|И зашли туда, и вошли в дом молодого левита, в дом Михи, и приветствовали его.
JUDG|18|16|А шестьсот человек из сынов Дановых, перепоясанные воинским оружием, стояли у ворот.
JUDG|18|17|Пять же человек, ходивших осматривать землю, пошли, вошли туда, взяли истукан и ефод и терафим и литый кумир. Священник стоял у ворот с теми шестьюстами человек, препоясанных воинским оружием.
JUDG|18|18|Когда они вошли в дом Михи и взяли истукан, ефод, терафим и литый кумир, священник сказал им: что вы делаете?
JUDG|18|19|Они сказали ему: молчи, положи руку твою на уста твои и иди с нами и будь у нас отцом и священником; лучше ли тебе быть священником в доме одного человека, нежели быть священником в колене или в племени Израилевом?
JUDG|18|20|Священник обрадовался, и взял ефод, терафим и истукан, и пошел с народом.
JUDG|18|21|Они обратились и пошли, и отпустили детей, скот и тяжести вперед.
JUDG|18|22|Когда они удалились от дома Михи, жители домов соседних с домом Михи собрались и погнались за сынами Дана,
JUDG|18|23|и кричали сынам Дана. [Сыны Дановы] оборотились и сказали Михе: что тебе, что ты так кричишь?
JUDG|18|24|(Миха) сказал: вы взяли богов моих, которых я сделал, и священника, и ушли; чего еще более? как же вы говорите: что тебе?
JUDG|18|25|Сыны Дановы сказали ему: [молчи], чтобы мы не слышали голоса твоего; иначе некоторые из нас, рассердившись, нападут на вас, и ты погубишь себя и семейство твое.
JUDG|18|26|И пошли сыны Дановы путем своим; Миха же, видя, что они сильнее его, пошел назад и возвратился в дом свой.
JUDG|18|27|А [сыны Дановы] взяли то, что сделал Миха, и священника, который был у него, и пошли в Лаис, против народа спокойного и беспечного, и побили его мечом, а город сожгли огнем.
JUDG|18|28|Некому было помочь, потому что он был отдален от Сидона и ни с кем не имел дела. [Город сей] находился в долине, что близ Беф–Рехова. И построили [снова] город и поселились в нем,
JUDG|18|29|и нарекли имя городу: Дан, по имени отца своего Дана, сына Израилева; а прежде имя города тому было: Лаис.
JUDG|18|30|И поставили у себя сыны Дановы истукан; Ионафан же, сын Гирсона, сына Манассии, сам и сыновья его были священниками в колене Дановом до дня переселения [жителей той] земли;
JUDG|18|31|и имели у себя истукан, сделанный Михою, во все то время, когда дом Божий находился в Силоме.
JUDG|19|1|В те дни, когда не было царя у Израиля, жил один левит на склоне горы Ефремовой. Он взял себе наложницу из Вифлеема Иудейского.
JUDG|19|2|Наложница его поссорилась с ним и ушла от него в дом отца своего в Вифлеем Иудейский и была там четыре месяца.
JUDG|19|3|Муж ее встал и пошел за нею, чтобы поговорить к сердцу ее и возвратить ее к себе. С ним был слуга его и пара ослов. Она ввела его в дом отца своего.
JUDG|19|4|Отец этой молодой женщины, увидев его, с радостью встретил его, и удержал его тесть его, отец молодой женщины. И пробыл он у него три дня; они ели и пили и ночевали там.
JUDG|19|5|В четвертый день встали они рано, и он встал, чтоб идти. И сказал отец молодой женщины зятю своему: подкрепи сердце твое куском хлеба, и потом пойдете.
JUDG|19|6|Они остались, и оба вместе ели и пили. И сказал отец молодой женщины человеку тому: останься еще на ночь, и пусть повеселится сердце твое.
JUDG|19|7|Человек тот встал, было, чтоб идти, но тесть его упросил его, и он опять ночевал там.
JUDG|19|8|На пятый день встал он поутру, чтоб идти. И сказал отец молодой женщины той: подкрепи сердце твое [хлебом], и помедлите, доколе преклонится день. И ели оба они.
JUDG|19|9|И встал тот человек, чтоб идти, сам он, наложница его и слуга его. И сказал ему тесть его, отец молодой женщины: вот, день преклонился к вечеру, ночуйте, пожалуйте; вот, дню скоро конец, ночуй здесь, пусть повеселится сердце твое; завтра пораньше встанете в путь ваш, и пойдешь в дом твой.
JUDG|19|10|Но муж не согласился ночевать, встал и пошел; и пришел к Иевусу, что [ныне] Иерусалим; с ним пара навьюченных ослов и наложница его с ним.
JUDG|19|11|Когда они были близ Иевуса, день уже очень преклонился. И сказал слуга господину своему: зайдем в этот город Иевусеев и ночуем в нем.
JUDG|19|12|Господин его сказал ему: нет, не пойдем в город иноплеменников, которые не из сынов Израилевых, но дойдем до Гивы.
JUDG|19|13|И сказал слуге своему: дойдем до одного из сих мест и ночуем в Гиве, или в Раме.
JUDG|19|14|И пошли, и шли, и закатилось солнце подле Гивы Вениаминовой.
JUDG|19|15|И повернули они туда, чтобы пойти ночевать в Гиве. И пришел он и сел на улице в городе; но никто не приглашал их в дом для ночлега.
JUDG|19|16|И вот, идет один старик с работы своей с поля вечером; он родом был с горы Ефремовой и жил в Гиве. Жители же места сего были сыны Вениаминовы.
JUDG|19|17|Он, подняв глаза свои, увидел прохожего на улице городской. И сказал старик: куда идешь? и откуда ты пришел?
JUDG|19|18|Он сказал ему: мы идем из Вифлеема Иудейского к горе Ефремовой, откуда я; я ходил в Вифлеем Иудейский, а теперь иду к дому Господа; и никто не приглашает меня в дом;
JUDG|19|19|у нас есть и солома и корм для ослов наших; также хлеб и вино для меня и для рабы твоей и для сего слуги есть у рабов твоих; ни в чем нет недостатка.
JUDG|19|20|Старик сказал ему: будь спокоен: весь недостаток твой на мне, только не ночуй на улице.
JUDG|19|21|И ввел его в дом свой и дал корму ослам [его], а сами они омыли ноги свои и ели и пили.
JUDG|19|22|Тогда как они развеселили сердца свои, вот, жители города, люди развратные, окружили дом, стучались в двери и говорили старику, хозяину дома: выведи человека, вошедшего в дом твой, мы познаем его.
JUDG|19|23|Хозяин дома вышел к ним и сказал им: нет, братья мои, не делайте зла, когда человек сей вошел в дом мой, не делайте этого безумия;
JUDG|19|24|вот у меня дочь девица, и у него наложница, выведу я их, смирите их и делайте с ними, что вам угодно; а с человеком сим не делайте этого безумия.
JUDG|19|25|Но они не хотели слушать его. Тогда муж взял свою наложницу и вывел к ним на улицу. Они познали ее, и ругались над нею всю ночь до утра. И отпустили ее при появлении зари.
JUDG|19|26|И пришла женщина пред появлением зари, и упала у дверей дома того человека, у которого был господин ее, [и лежала] до света.
JUDG|19|27|Господин ее встал поутру, отворил двери дома и вышел, чтоб идти в путь свой: и вот, наложница его лежит у дверей дома, и руки ее на пороге.
JUDG|19|28|Он сказал ей: вставай, пойдем. Но ответа не было, [потому что она умерла]. Он положил ее на осла, встал и пошел в свое место.
JUDG|19|29|Придя в дом свой, взял нож и, взяв наложницу свою, разрезал ее по членам ее на двенадцать частей и послал во все пределы Израилевы.
JUDG|19|30|Всякий, видевший это, говорил: не бывало и не видано было подобного сему от дня исшествия сынов Израилевых из земли Египетской до сего дня. Обратите внимание на это, посоветуйтесь и скажите.
JUDG|20|1|И вышли все сыны Израилевы, и собралось [все] общество, как один человек, от Дана до Вирсавии, и земля Галаадская пред Господа в Массифу.
JUDG|20|2|И собрались начальники всего народа, все колена Израилевы, в собрание народа Божия, четыреста тысяч пеших, обнажающих меч.
JUDG|20|3|И сыны Вениаминовы услышали, что сыны Израилевы пришли в Массифу. И сказали сыны Израилевы: скажите, как происходило это зло?
JUDG|20|4|Левит, муж оной убитой женщины, отвечал и сказал: я с наложницею моею пришел ночевать в Гиву Вениаминову;
JUDG|20|5|и восстали на меня жители Гивы и окружили из–за меня дом ночью; меня намеревались убить, и наложницу мою замучили, так, что она умерла;
JUDG|20|6|я взял наложницу мою, разрезал ее и послал ее во все области владения Израилева, ибо они сделали беззаконное и срамное дело в Израиле;
JUDG|20|7|вот все вы, сыны Израилевы, рассмотрите это дело и решите здесь.
JUDG|20|8|И восстал весь народ, как один человек, и сказал: не пойдем никто в шатер свой и не возвратимся никто в дом свой;
JUDG|20|9|и вот что мы сделаем ныне с Гивою: [пойдем] на нее по жребию;
JUDG|20|10|и возьмем по десяти человек из ста от всех колен Израилевых, по сто от тысячи и по тысяче от тьмы, чтоб они принесли съестных припасов для народа, который пойдет против Гивы Вениаминовой, наказать ее за срамное дело, которое она сделала в Израиле.
JUDG|20|11|И собрались все Израильтяне против города единодушно, как один человек.
JUDG|20|12|И послали колена Израилевы во все колено Вениаминово сказать: какое это гнусное дело сделано у вас!
JUDG|20|13|Выдайте развращенных оных людей, которые в Гиве; мы умертвим их и искореним зло из Израиля. Но сыны Вениаминовы не хотели послушать голоса братьев своих, сынов Израилевых;
JUDG|20|14|а собрались сыны Вениаминовы из городов в Гиву, чтобы пойти войною против сынов Израилевых.
JUDG|20|15|И насчиталось в тот день сынов Вениаминовых, [собравшихся] из городов, двадцать шесть тысяч человек, обнажающих меч; кроме того, из жителей Гивы насчитано семьсот отборных;
JUDG|20|16|из всего народа сего было семьсот человек отборных, которые были левши, и все сии, бросая из пращей камни в волос, не бросали мимо.
JUDG|20|17|Израильтян же, кроме сынов Вениаминовых, насчиталось четыреста тысяч человек, обнажающих меч; все они были способны к войне.
JUDG|20|18|И встали и пошли в дом Божий, и вопрошали Бога и сказали сыны Израилевы: кто из нас прежде пойдет на войну с сынами Вениамина? И сказал Господь: Иуда [пойдет] впереди.
JUDG|20|19|И встали сыны Израилевы поутру и расположились станом подле Гивы;
JUDG|20|20|и выступили Израильтяне на войну против Вениамина, и стали сыны Израилевы в боевой порядок близ Гивы.
JUDG|20|21|И вышли сыны Вениаминовы из Гивы и положили в тот день двадцать две тысячи Израильтян на землю.
JUDG|20|22|Но народ Израильский ободрился, и опять стали в боевой порядок на том месте, где стояли в прежний день.
JUDG|20|23|И пошли сыны Израилевы, и плакали пред Господом до вечера, и вопрошали Господа: вступать ли мне еще в сражение с сынами Вениамина, брата моего? Господь сказал: идите против него.
JUDG|20|24|И подступили сыны Израилевы к сынам Вениамина во второй день.
JUDG|20|25|Вениамин вышел против них из Гивы во второй день, и еще положили на землю из сынов Израилевых восемнадцать тысяч человек, обнажающих меч.
JUDG|20|26|Тогда все сыны Израилевы и весь народ пошли и пришли в дом Божий и, сидя там, плакали пред Господом, и постились в тот день до вечера, и вознесли всесожжения и мирные жертвы пред Господом.
JUDG|20|27|И вопрошали сыны Израилевы Господа (в то время ковчег завета Божия находился там,
JUDG|20|28|и Финеес, сын Елеазара, сына Ааронова, предстоял пред ним): выходить ли мне еще на сражение с сынами Вениамина, брата моего, или нет? Господь сказал: идите; Я завтра предам его в руки ваши.
JUDG|20|29|И поставил Израиль засаду вокруг Гивы.
JUDG|20|30|И пошли сыны Израилевы на сынов Вениамина в третий день и стали в боевой порядок пред Гивою, как прежде.
JUDG|20|31|Сыны Вениаминовы выступили против народа и отдалились от города, и начали, как прежде, убивать из народа на дорогах, из которых одна идет к Вефилю, а другая к Гиве полем, и [убили] до тридцати человек из Израильтян.
JUDG|20|32|И сказали сыны Вениаминовы: они падают пред нами, как и прежде. А сыны Израилевы сказали: побежим от них и отвлечем их от города на дороги.
JUDG|20|33|И все Израильтяне встали с своего места и выстроились в Ваал–Фамаре. И засада Израилева устремилась из своего места, с западной стороны Гивы.
JUDG|20|34|И пришли пред Гиву десять тысяч человек отборных из всего Израиля, и началось жестокое сражение; но [сыны Вениамина] не знали, что предстоит им беда.
JUDG|20|35|И поразил Господь Вениамина пред Израильтянами, и положили в тот день Израильтяне из сынов Вениамина двадцать пять тысяч сто человек, обнажавших меч.
JUDG|20|36|Когда сыны Вениамина увидели, что они поражены, тогда Израильтяне уступили место сынам Вениамина, ибо надеялись на засаду, которую они поставили близ Гивы.
JUDG|20|37|Засада же поспешила и устремилась к Гиве, и вступила и поразила весь город мечом.
JUDG|20|38|Израильтяне поставили с засадою [условленным] знаком к нападению поднимающийся дым из города.
JUDG|20|39|Итак, когда Израильтяне отступили с места сражения, и Вениамин начал поражать и поверг Израильтян до тридцати человек и говорил: "опять падают они пред нами, как и в прежние сражения",
JUDG|20|40|тогда начал подниматься из города дым столбом. Вениамин оглянулся назад, и вот, [дым] от всего города восходит к небу.
JUDG|20|41|Израильтяне воротились, а Вениамин оробел, ибо увидел, что постигла его беда.
JUDG|20|42|И побежали они от Израильтян по дороге к пустыне; но сеча преследовала их, и выходившие из городов побивали их там;
JUDG|20|43|окружили Вениамина, и преследовали его до Менухи и поражали до самой восточной стороны Гивы.
JUDG|20|44|И пало из сынов Вениамина восемнадцать тысяч человек, людей сильных.
JUDG|20|45|[Оставшиеся] оборотились и побежали к пустыне, к скале Риммону, и побили еще [Израильтяне] на дорогах пять тысяч человек; и гнались за ними до Гидома и еще убили из них две тысячи человек.
JUDG|20|46|Всех же сынов Вениаминовых, павших в тот день, было двадцать пять тысяч человек, обнажавших меч, и все они были мужи сильные.
JUDG|20|47|И [обратились оставшиеся] и убежали в пустыню, к скале Риммону, шестьсот человек, и оставались там в каменной горе Риммоне четыре месяца.
JUDG|20|48|Израильтяне же опять пошли к сынам Вениаминовым и поразили их мечом, и людей в городе, и скот, и все, что ни встречалось, и все находившиеся [на пути] города сожгли огнем.
JUDG|21|1|И поклялись Израильтяне в Массифе, говоря: никто из нас не отдаст дочери своей сынам Вениамина в замужество.
JUDG|21|2|И пришел народ в дом Божий, и сидели там до вечера пред Богом, и подняли громкий вопль, и сильно плакали,
JUDG|21|3|и сказали: Господи, Боже Израилев! для чего случилось это в Израиле, что не стало теперь у Израиля одного колена?
JUDG|21|4|На другой день встал народ поутру, и устроили там жертвенник, и вознесли всесожжения и мирные жертвы.
JUDG|21|5|И сказали сыны Израилевы: кто не приходил в собрание пред Господа из всех колен Израилевых? Ибо великое проклятие [произнесено] было на тех, которые не пришли пред Господа в Массифу, и сказано было, что те преданы будут смерти.
JUDG|21|6|И сжалились сыны Израилевы над Вениамином, братом своим, и сказали: ныне отсечено одно колено от Израиля;
JUDG|21|7|как поступить нам с оставшимися из них [касательно] жен, когда мы поклялись Господом не давать им жен из дочерей наших?
JUDG|21|8|И сказали: нет ли кого из колен Израилевых, кто не приходил пред Господа в Массифу? И оказалось, что из Иависа Галаадского никто не приходил пред Господа в стан на собрание.
JUDG|21|9|И осмотрен народ, и вот, не было там ни одного из жителей Иависа Галаадского.
JUDG|21|10|И послало туда общество двенадцать тысяч человек, мужей сильных, и дали им приказание, говоря: идите и поразите жителей Иависа Галаадского мечом, и женщин и детей;
JUDG|21|11|и вот что сделайте: всякого мужчину и всякую женщину, познавшую ложе мужеское, предайте заклятию.
JUDG|21|12|И нашли они между жителями Иависа Галаадского четыреста девиц, не познавших ложа мужеского, и привели их в стан в Силом, что в земле Ханаанской.
JUDG|21|13|И послало все общество переговорить с сынами Вениамина, бывшими в скале Риммоне, и объявило им мир.
JUDG|21|14|Тогда возвратились сыны Вениамина, и дали им (Израильтяне) жен, которых оставили в живых из женщин Иависа Галаадского; но оказалось, что этого было недостаточно.
JUDG|21|15|Народ же сожалел о Вениамине, что Господь не сохранил целости колен Израилевых.
JUDG|21|16|И сказали старейшины общества: что нам делать с оставшимися [касательно] жен, ибо истреблены женщины у Вениамина?
JUDG|21|17|И сказали: наследственная земля пусть остается уцелевшим сынам Вениамина, чтобы не исчезло колено от Израиля;
JUDG|21|18|но мы не можем дать им жен из дочерей наших; ибо сыны Израилевы поклялись, говоря: проклят, кто даст жену Вениамину.
JUDG|21|19|И сказали: вот, каждый год бывает праздник Господень в Силоме, который на север от Вефиля и на восток от дороги, ведущей от Вефиля в Сихем, и на юг от Левоны.
JUDG|21|20|И приказали сынам Вениамина и сказали: подите и засядьте в виноградниках,
JUDG|21|21|и смотрите, когда выйдут девицы Силомские плясать в хороводах, тогда выйдите из виноградников и схватите себе каждый жену из девиц Силомских и идите в землю Вениаминову;
JUDG|21|22|и когда придут отцы их, или братья их с жалобою к нам, мы скажем им: простите нас за них, ибо мы не взяли для каждого из них жены на войне, и вы не дали им; теперь вы виновны.
JUDG|21|23|Сыны Вениамина так и сделали, и взяли жен по числу своему из бывших в хороводе, которых они похитили, и пошли и возвратились в удел свой, и построили города и стали жить в них.
JUDG|21|24|В то же время Израильтяне разошлись оттуда каждый в колено свое и в племя свое, и пошли оттуда каждый в удел свой.
JUDG|21|25|В те дни не было царя у Израиля; каждый делал то, что ему казалось справедливым.
