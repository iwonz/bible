2TIM|1|1|Paul, an apostle of Christ Jesus by the will of God according to the promise of the life that is in Christ Jesus,
2TIM|1|2|To Timothy, my beloved child: Grace, mercy, and peace from God the Father and Christ Jesus our Lord.
2TIM|1|3|I thank God whom I serve, as did my ancestors, with a clear conscience, as I remember you constantly in my prayers night and day.
2TIM|1|4|As I remember your tears, I long to see you, that I may be filled with joy.
2TIM|1|5|I am reminded of your sincere faith, a faith that dwelt first in your grandmother Lois and your mother Eunice and now, I am sure, dwells in you as well.
2TIM|1|6|For this reason I remind you to fan into flame the gift of God, which is in you through the laying on of my hands,
2TIM|1|7|for God gave us a spirit not of fear but of power and love and self-control.
2TIM|1|8|Therefore do not be ashamed of the testimony about our Lord, nor of me his prisoner, but share in suffering for the gospel by the power of God,
2TIM|1|9|who saved us and called us to a holy calling, not because of our works but because of his own purpose and grace, which he gave us in Christ Jesus before the ages began,
2TIM|1|10|and which now has been manifested through the appearing of our Savior Christ Jesus, who abolished death and brought life and immortality to light through the gospel,
2TIM|1|11|for which I was appointed a preacher and apostle and teacher,
2TIM|1|12|which is why I suffer as I do. But I am not ashamed, for I know whom I have believed, and I am convinced that he is able to guard until that Day what has been entrusted to me.
2TIM|1|13|Follow the pattern of the sound words that you have heard from me, in the faith and love that are in Christ Jesus.
2TIM|1|14|By the Holy Spirit who dwells within us, guard the good deposit entrusted to you.
2TIM|1|15|You are aware that all who are in Asia turned away from me, among whom are Phygelus and Hermogenes.
2TIM|1|16|May the Lord grant mercy to the household of Onesiphorus, for he often refreshed me and was not ashamed of my chains,
2TIM|1|17|but when he arrived in Rome he searched for me earnestly and found me-
2TIM|1|18|may the Lord grant him to find mercy from the Lord on that Day!- and you well know all the service he rendered at Ephesus.
2TIM|2|1|You then, my child, be strengthened by the grace that is in Christ Jesus,
2TIM|2|2|and what you have heard from me in the presence of many witnesses entrust to faithful men who will be able to teach others also.
2TIM|2|3|Share in suffering as a good soldier of Christ Jesus.
2TIM|2|4|No soldier gets entangled in civilian pursuits, since his aim is to please the one who enlisted him.
2TIM|2|5|An athlete is not crowned unless he competes according to the rules.
2TIM|2|6|It is the hard-working farmer who ought to have the first share of the crops.
2TIM|2|7|Think over what I say, for the Lord will give you understanding in everything.
2TIM|2|8|Remember Jesus Christ, risen from the dead, the offspring of David, as preached in my gospel,
2TIM|2|9|for which I am suffering, bound with chains as a criminal. But the word of God is not bound!
2TIM|2|10|Therefore I endure everything for the sake of the elect, that they also may obtain the salvation that is in Christ Jesus with eternal glory.
2TIM|2|11|The saying is trustworthy, for: If we have died with him, we will also live with him;
2TIM|2|12|if we endure, we will also reign with him; if we deny him, he also will deny us;
2TIM|2|13|if we are faithless, he remains faithful- for he cannot deny himself.
2TIM|2|14|Remind them of these things, and charge them before God not to quarrel about words, which does no good, but only ruins the hearers.
2TIM|2|15|Do your best to present yourself to God as one approved, a worker who has no need to be ashamed, rightly handling the word of truth.
2TIM|2|16|But avoid irreverent babble, for it will lead people into more and more ungodliness,
2TIM|2|17|and their talk will spread like gangrene. Among them are Hymenaeus and Philetus,
2TIM|2|18|who have swerved from the truth, saying that the resurrection has already happened. They are upsetting the faith of some.
2TIM|2|19|But God's firm foundation stands, bearing this seal: "The Lord knows those who are his," and, "Let everyone who names the name of the Lord depart from iniquity."
2TIM|2|20|Now in a great house there are not only vessels of gold and silver but also of wood and clay, some for honorable use, some for dishonorable.
2TIM|2|21|Therefore, if anyone cleanses himself from what is dishonorable, he will be a vessel for honorable use, set apart as holy, useful to the master of the house, ready for every good work.
2TIM|2|22|So flee youthful passions and pursue righteousness, faith, love, and peace, along with those who call on the Lord from a pure heart.
2TIM|2|23|Have nothing to do with foolish, ignorant controversies; you know that they breed quarrels.
2TIM|2|24|And the Lord's servant must not be quarrelsome but kind to everyone, able to teach, patiently enduring evil,
2TIM|2|25|correcting his opponents with gentleness. God may perhaps grant them repentance leading to a knowledge of the truth,
2TIM|2|26|and they may escape from the snare of the devil, after being captured by him to do his will.
2TIM|3|1|But understand this, that in the last days there will come times of difficulty.
2TIM|3|2|For people will be lovers of self, lovers of money, proud, arrogant, abusive, disobedient to their parents, ungrateful, unholy,
2TIM|3|3|heartless, unappeasable, slanderous, without self-control, brutal, not loving good,
2TIM|3|4|treacherous, reckless, swollen with conceit, lovers of pleasure rather than lovers of God,
2TIM|3|5|having the appearance of godliness, but denying its power. Avoid such people.
2TIM|3|6|For among them are those who creep into households and capture weak women, burdened with sins and led astray by various passions,
2TIM|3|7|always learning and never able to arrive at a knowledge of the truth.
2TIM|3|8|Just as Jannes and Jambres opposed Moses, so these men also oppose the truth, men corrupted in mind and disqualified regarding the faith.
2TIM|3|9|But they will not get very far, for their folly will be plain to all, as was that of those two men.
2TIM|3|10|You, however, have followed my teaching, my conduct, my aim in life, my faith, my patience, my love, my steadfastness,
2TIM|3|11|my persecutions and sufferings that happened to me at Antioch, at Iconium, and at Lystra- which persecutions I endured; yet from them all the Lord rescued me.
2TIM|3|12|Indeed, all who desire to live a godly life in Christ Jesus will be persecuted,
2TIM|3|13|while evil people and impostors will go on from bad to worse, deceiving and being deceived.
2TIM|3|14|But as for you, continue in what you have learned and have firmly believed, knowing from whom you learned it
2TIM|3|15|and how from childhood you have been acquainted with the sacred writings, which are able to make you wise for salvation through faith in Christ Jesus.
2TIM|3|16|All Scripture is breathed out by God and profitable for teaching, for reproof, for correction, and for training in righteousness,
2TIM|3|17|that the man of God may be competent, equipped for every good work.
2TIM|4|1|I charge you in the presence of God and of Christ Jesus, who is to judge the living and the dead, and by his appearing and his kingdom:
2TIM|4|2|preach the word; be ready in season and out of season; reprove, rebuke, and exhort, with complete patience and teaching.
2TIM|4|3|For the time is coming when people will not endure sound teaching, but having itching ears they will accumulate for themselves teachers to suit their own passions,
2TIM|4|4|and will turn away from listening to the truth and wander off into myths.
2TIM|4|5|As for you, always be sober-minded, endure suffering, do the work of an evangelist, fulfill your ministry.
2TIM|4|6|For I am already being poured out as a drink offering, and the time of my departure has come.
2TIM|4|7|I have fought the good fight, I have finished the race, I have kept the faith.
2TIM|4|8|Henceforth there is laid up for me the crown of righteousness, which the Lord, the righteous judge, will award to me on that Day, and not only to me but also to all who have loved his appearing.
2TIM|4|9|Do your best to come to me soon.
2TIM|4|10|For Demas, in love with this present world, has deserted me and gone to Thessalonica. Crescens has gone to Galatia, Titus to Dalmatia.
2TIM|4|11|Luke alone is with me. Get Mark and bring him with you, for he is very useful to me for ministry.
2TIM|4|12|Tychicus I have sent to Ephesus.
2TIM|4|13|When you come, bring the cloak that I left with Carpus at Troas, also the books, and above all the parchments.
2TIM|4|14|Alexander the coppersmith did me great harm; the Lord will repay him according to his deeds.
2TIM|4|15|Beware of him yourself, for he strongly opposed our message.
2TIM|4|16|At my first defense no one came to stand by me, but all deserted me. May it not be charged against them!
2TIM|4|17|But the Lord stood by me and strengthened me, so that through me the message might be fully proclaimed and all the Gentiles might hear it. So I was rescued from the lion's mouth.
2TIM|4|18|The Lord will rescue me from every evil deed and bring me safely into his heavenly kingdom. To him be the glory forever and ever. Amen.
2TIM|4|19|Greet Prisca and Aquila, and the household of Onesiphorus.
2TIM|4|20|Erastus remained at Corinth, and I left Trophimus, who was ill, at Miletus.
2TIM|4|21|Do your best to come before winter. Eubulus sends greetings to you, as do Pudens and Linus and Claudia and all the brothers.
2TIM|4|22|The Lord be with your spirit. Grace be with you.
