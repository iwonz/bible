1SAM|1|1|І був один чоловік із Раматаїм-Цофіму, з Єфремових гір, а ім'я йому Елкана, син Єрохама, сина Ілія, сина Тоху, сина Цуфа, єфремлянин.
1SAM|1|2|А він мав дві жінки, ім'я одній Анна, а ім'я другій Пеніна. І були в Пеніни діти, а в Анни дітей не було.
1SAM|1|3|А той чоловік рік-у-рік ходив із свого міста до Шіло, щоб вклонятися та приносити жертви Господу Саваоту. А там два Ілієві сини, Гофні та Пінхас, були священиками для Господа.
1SAM|1|4|І як бував той день, і Елкана приносив жертви, то він давав своїй жінці Пеніні й усім синам її та дочкам її частини,
1SAM|1|5|а Анні давав частину подвійну, бо любив її. Та Господь замкнув її утробу.
1SAM|1|6|А її суперниця розпалювала їй гнів, щоб докучати їй, бо Господь замкнув її утробу.
1SAM|1|7|І так робив він рік-у-рік, коли вона входила до Господнього дому, а та так гнівила її. І вона плакала й не їла.
1SAM|1|8|І сказав їй чоловік її Елкана: Анно, чого ти плачеш і чому не їси? І чого сумне твоє серце? Чи ж я не ліпший тобі за десятьох синів?
1SAM|1|9|І встала Анна по їді та по питті в Шіло, а священик Ілій сидів на стільці при бічному одвірку Господнього храму.
1SAM|1|10|А вона була скорбна духом, і молилася до Господа та плакала гірко.
1SAM|1|11|І склала вона обітницю, та й сказала: Господи Саваоте, якщо дійсно споглянеш на біду Твоєї невільниці, і згадаєш мене, і не забудеш Своєї невільниці, і даси Своїй невільниці нащадка чоловічої статі, то я дам його Господеві на всі дні життя його, а бритва не торкнеться його голови.
1SAM|1|12|І сталося, коли вона довго молилася перед Господнім лицем, то Ілій пильнував за її устами.
1SAM|1|13|А Анна вона говорила в серці своїм: тільки губи її порушувалися, а голос її не був чутий. І вважав її Ілій за п'яну.
1SAM|1|14|І сказав до неї Ілій: Аж доки ти будеш п'яною? Витверезись зо свого вина!
1SAM|1|15|А Анна відповіла та й сказала: Ні, пане мій, я жінка скорбна духом, а вина та п'янкого напою не пила я. І я вилила душу свою перед Господнім лицем.
1SAM|1|16|Не вважай своєї невільниці за негідницю, бо я говорила аж доти з великої своєї скорботи та з туги своєї.
1SAM|1|17|І відповів Ілій та й сказав: Іди з миром! А Бог Ізраїлів дасть тобі бажання твоє, яке ти від Нього жадала.
1SAM|1|18|А вона сказала: Нехай невільниця твоя знайде милість в очах твоїх! І пішла та жінка своєю дорогою, та й їла, а обличчя її не було вже сумне.
1SAM|1|19|І встала вона рано вранці, і вклонилася перед Господнім лицем. І вернулися вони, і ввійшли до свого дому до Рами. І Елкана пізнав свою жінку Анну, а Господь згадав про неї.
1SAM|1|20|І сталося по році, і завагітніла Анна, та й сина породила. І назвала вона ім'я йому: Самуїл, бо від Господа жадала його.
1SAM|1|21|І пішов той чоловік Елкана та ввесь дім його вчинити для Господа річну жертву та обітниці свої.
1SAM|1|22|А Анна не пішла, бо сказала до чоловіка свого: Аж коли буде відлучений цей хлопчик, то відведу його, і він з'явиться перед Господнім лицем, і назавжди позостанеться там!
1SAM|1|23|І сказав їй чоловік її Елкана: Роби те, що добре в очах твоїх! Залишайся, аж поки відлучиш його, тільки нехай виконає Господь Своє слово. І залишалась та жінка, і годувала свого сина, аж поки вона відлучила його.
1SAM|1|24|А коли відлучила, то повела його з собою та з трьома бичками й одною ефою муки, і бурдюком вина, і привела його до Господнього дому до Шіло. А той хлопчик був ще малий.
1SAM|1|25|І зарізали бичка, і привели того хлопчика до Ілія.
1SAM|1|26|І вона сказала: О, пане мій, як жива душа твоя, мій пане, я та жінка, що стояла з тобою отут, щоб молитися Господеві.
1SAM|1|27|Я молилася за дитину цю, і Господь дав мені жадання моє, що я просила від Нього.
1SAM|1|28|А тепер я віддаю його Господеві на всі дні, скільки він жаданий для Господа. І вклонилася там Господеві.
1SAM|2|1|І молилася Анна та й проказала: Звеселилося Господом серце моє, мій ріг став високим у Господі! Розкрилися уста мої на моїх ворогів, бо радію з спасіння Твого!
1SAM|2|2|Немає святого, подібного Господу, немає нікого, крім Тебе, і скелі немає, як Бог наш!
1SAM|2|3|Більше не говоріть зарозуміло, нехай з ваших уст не виходить зухвальство, бо Господь Бог знання, і Він упляновує вчинки!
1SAM|2|4|Лук сильних поламаний, а немічні оперезалися силою!
1SAM|2|5|Наймаються ситі за хліб, а голодні відпочивають, аж неплідна сімох породила, а многодітна знесиліла.
1SAM|2|6|Господь побиває й оживлює, до шеолу знижає й підносить до неба.
1SAM|2|7|Господь зубожує та збагачує, понижує Він та звеличує.
1SAM|2|8|Підіймає нужденного з пороху, підносить убогого зо смітників, щоб посадити з вельможами й престол слави їм дать на спадщину, бо Господні основи землі, і на них Він поставив вселенну.
1SAM|2|9|Він ноги святих Своїх стереже, нечестиві ж погинуть у темряві, бо сильним не з сили стає чоловік.
1SAM|2|10|Господь хай поламані будуть Його супротивники! У небі Господь загримить, і розсудить Він кінці землі! І Він подасть силу Своєму цареві, і рога повищить Свого помазанця!
1SAM|2|11|І пішов Елкана до Рами, до дому свого. А той отрок служив Господеві при священикові Ілії.
1SAM|2|12|А сини Ілія були люди негідні, вони не знали Господа,
1SAM|2|13|ані звичаю священичого з народом. Коли хто приносив жертву, то, як варилося м'ясо, приходив священиків слуга, а в його руці тризубе видельце.
1SAM|2|14|І він із грюкотом стромляв до мідниці, або до кітла, або до горшка, або до горняти, і все, що витягне видельце, священик собі брав. Так вони робили всьому Ізраїлеві, що приходив туди до Шіло.
1SAM|2|15|Також поки палили лій, то приходив священиків слуга, та й говорив до чоловіка, що приносив жертву: Дай м'яса на печеню для священика, бо він не візьме від тебе м'яса вареного, а тільки сире!
1SAM|2|16|А як той чоловік відповідав йому: Нехай перше спалять і той лій, а ти потім візьми собі, скільки буде жадати душа твоя! А той говорив: Ні, таки зараз давай! А коли ні, візьму силою!
1SAM|2|17|І був гріх тих юнаків дуже великий перед Господнім лицем, бо ті люди безчестили Господню жертву.
1SAM|2|18|А Самуїл служив перед Господнім лицем. Отрок був оперезаний лляним ефодом.
1SAM|2|19|А малу верхню одежину робила йому його мати, і приносила йому з року на рік, коли приходила з своїм мужем приносити річну жертву.
1SAM|2|20|А Ілій поблагословив Елкану й його жінку та й сказав: Нехай Господь дасть тобі нащадків від цієї жінки, за відданого, що Господь узяв. І пішли вони на місце своє.
1SAM|2|21|І Господь згадав про Анну, і вона завагітніла, та й породила трьох синів та дві дочки. А отрок Самуїл ріс із Господом.
1SAM|2|22|А Ілій був дуже старий. І почув він усе, що сини його роблять усьому Ізраїлеві, і що вони злягаються з жінками, які відбувають службу при вході скинії заповіту.
1SAM|2|23|І він сказав їм: Нащо ви робите такі речі, про які я чую? Про ваші злі вчинки я чую від усього цього народу.
1SAM|2|24|Ні, сини мої, недобра та чутка, що я чую, ви відхиляєте Господній народ від Закону!
1SAM|2|25|Якщо хто згрішить супроти людини, то помоляться за неї перед Богом. А якщо людина згрішить супроти Господа, хто заступиться за неї? Та вони не слухали голосу батька свого, бо Господь постановив погубити їх.
1SAM|2|26|А отрок Самуїл усе ріс, та здобував ласку як у Господа, так і в людей.
1SAM|2|27|І прийшов Божий чоловік до Ілія, та й сказав йому: Так сказав Господь: Чи ж Я справді не об'явився домові твого батька, як були вони в Єгипті, у фараоновім домі?
1SAM|2|28|Я вибрав його Собі зо всіх Ізраїлевих племен за священика, щоб він входив до Мого жертівника, щоб кадив кадило, щоб носив ефода перед Моїм лицем. І дав Я домові твого батька всі жертви Ізраїлевих синів.
1SAM|2|29|Чого ж ви берете під ноги Мою жертву та Мою жертву хлібну, що Я заповів для скинії? І ти вшанував синів своїх більш, як Мене, щоб ви потовстіли від найкращих частин усякого Ізраїлевого дару перед лицем Моїм.
1SAM|2|30|Тому то слово Господа, Бога Ізраїлевого, таке: Говорячи, сказав Я: Дім твій та дім батька твого будуть ходити перед Моїм лицем аж навіки. А тепер слово Господнє: Не буде в Мене такого, бо Я шаную тих, хто шанує Мене, а ті, хто зневажає Мене, будуть зневажені!
1SAM|2|31|Ось приходять дні, і Я відітну рамено твоє та рамено дому батька твого, щоб не було старого в домі твоєму.
1SAM|2|32|І побачиш біду Мого мешкання, хоч у всьому Я добре чинив Ізраїлеві, і не буде старого в домі твоїм по всі дні.
1SAM|2|33|Я не витну в тебе всіх від Мого жертівника, щоб вибрати очі твої, і щоб зробити біль душі твоїй, та ввесь доріст твого дому повмирає в силі віку.
1SAM|2|34|А оце тобі ознака, що прийде на обох синів твоїх, на Хофні та Пінхаса, обидва вони помруть одного дня.
1SAM|2|35|А Я поставлю Собі священика вірного, він буде робити згідно з серцем Моїм та з Моєю душею. І Я збудую йому тривалий дім, і він буде ходити перед Моїм помазанцем по всі дні.
1SAM|2|36|І станеться, кожен, хто полишиться в домі твоїм, прийде вклонятися йому за аґору срібла та за буханець хліба, і скаже: Долучи мене до одного з священицтв, щоб їсти кавалок хліба.
1SAM|3|1|А отрок Самуїл служив Господеві при Ілії. А Господнє слово було рідке за тих днів, видіння не було часте.
1SAM|3|2|І сталося того дня, коли Ілій лежав на своєму місці, а очі його стали затемнятися, він не міг бачити,
1SAM|3|3|і поки Божий світильник ще не погас, а Самуїл лежав у Господньому храмі, там, де Божий ковчег,
1SAM|3|4|то покликав Господь до Самуїла: Самуїле, Самуїле! А він відказав: Ось я!
1SAM|3|5|І побіг він до Ілія та й сказав: Ось я, бо ти кликав мене. А той відказав: Я не кликав. Вернися, лягай. І він пішов і ліг.
1SAM|3|6|А Господь далі покликав: Самуїле, Самуїле! І встав Самуїл, і пішов до Ілія та й сказав: Ось я, бо ти кликав мене. А той відказав: Не кликав я, сину мій. Вернися, лягай.
1SAM|3|7|А Самуїл ще не пізнав голосу Господа, і ще не відкрилося йому Господнє слово.
1SAM|3|8|А Господь далі покликав Самуїла третій раз. І він устав, і пішов до Ілія та й сказав: Ось я, бо ти кликав мене. І зрозумів Ілій, що то Господь кличе отрока.
1SAM|3|9|І сказав Ілій до Самуїла: Іди, лягай. І якщо знову покличе тебе, то скажеш: Говори, Господи, бо раб Твій слухає Тебе! І пішов Самуїл, та й ліг на своє місце.
1SAM|3|10|І ввійшов Господь, і став, і покликав, як перед тим: Самуїле, Самуїле! А Самуїл відказав: Говори, Господи, бо раб Твій слухає!
1SAM|3|11|І сказав Господь до Самуїла: Ось Я зроблю таку річ серед Ізраїля, що в кожного, хто почує про неї, задзвенить в обох вухах його.
1SAM|3|12|Того дня Я виконаю над Ілієм все, що Я говорив про дім його, від початку й до кінця.
1SAM|3|13|І розповім йому, що Я суджу дім його навіки за гріх, про який він знав, що сини його богозневажають, та не спиняв їх.
1SAM|3|14|Тому присягнув Я домом Ілія, що не очиститься гріх Ілієвого дому жертвою та жертвою хлібною навіки.
1SAM|3|15|І лежав Самуїл аж до ранку, і відчинив двері Господнього дому. А Самуїл боявся розповісти Ілієві про те видіння.
1SAM|3|16|І покликав Ілій Самуїла, та й сказав: Самуїле, сину мій! А той сказав: Ось я!
1SAM|3|17|І сказав він: Що то за річ, про яку Він говорив до тебе? Не крий правди передо мною. Нехай Господь зробить тобі так, і нехай додасть, якщо ти скажеш неправду передо мною про щось зо всього того, що говорив Він до тебе!
1SAM|3|18|І розповів йому Самуїл усе те, і не сказав неправди перед ним. А той сказав: Він Господь, нехай зробить те, що добре в очах Його!
1SAM|3|19|І виростав Самуїл, а Господь був із ним, і не опустив ані жодного зо всіх Його слів.
1SAM|3|20|І ввесь Ізраїль, від Дана аж до Беер-Шеви, пізнав, що Самуїл вірний, як пророк Господній.
1SAM|3|21|А Господь далі показувався в Шіло, бо Господь явився був у Шіло Самуїлові в слові Господньому.
1SAM|4|1|І було Самуїлове слово для всього Ізраїля. І вийшов Ізраїль на війну проти филистимлян, та й таборував при Евен-Гаезері, а филистимляни таборували в Афеку.
1SAM|4|2|І вишикувались филистимляни навпроти Ізраїля, а коли бій став тяжкий, то Ізраїль був побитий перед филистимлянами. І вони побили в боєвому шикові на полі близько чотирьох тисяч чоловіка.
1SAM|4|3|І прийшов народ до табору, а Ізраїлеві старші сказали: Чому вдарив нас Господь сьогодні перед филистимлянами? Візьмімо собі з Шіло ковчега Господнього заповіту, і нехай ввійде поміж нас, і нехай спасе нас із рук наших ворогів.
1SAM|4|4|І послав народ до Шіло, і понесли звідти ковчега заповіту Господа Саваота, що сидить на херувимах. А там були двоє Ілієвих синів, Хофні та Пінхас, із ковчегом Божого заповіту.
1SAM|4|5|І сталося, як ковчег заповіту Господнього прибув до табору, то ввесь Ізраїль скрикнув великим окриком, аж застогнала земля!
1SAM|4|6|А филистимляни почули голос окрику, та й сказали: Що це за голос цього великого окрику в єврейському таборі? І довідалися вони, що Господній ковчег прибув до табору.
1SAM|4|7|І полякалися филистимляни, і говорили: Бог прибув до табору! І сказали вони: Біда нам, бо такого, як це, не було ще ніколи!
1SAM|4|8|Біда нам! Хто нас урятує від руки цих потужних богів? Оце вони, ті боги, що вдарили були Єгипет усякою поразою у пустині!
1SAM|4|9|Зміцніться та будьте мужні, филистимляни, щоб ви не служили євреям, як вони служили вам. І будьте мужні, і воюйте!
1SAM|4|10|І воювали филистимляни. І був побитий Ізраїль, і кожен утікав до свого намету. І та поразка була дуже велика. І впало з Ізраїля тридцять тисяч піхоти.
1SAM|4|11|А Божий ковчег був узятий, і два Ілієві сини, Хофні та Пінхас, полягли...
1SAM|4|12|І побіг один веніяминівець із бою, і прибув того дня до Шіло; а одежа його була подерта, і порох на голові його.
1SAM|4|13|І прибув він, аж ось Ілій сидить на стільці при дорозі й виглядає, бо серце йому тремтіло за Божого ковчега. А той чоловік прийшов, і розповів у місті, і закричало все місто!
1SAM|4|14|А Ілій почув голос того крику та й сказав: Що це за голос того натовпу? А той чоловік поспішив і прийшов, та й розповів Ілієві.
1SAM|4|15|А Ілій був віку дев'ятидесяти й восьми літ, а очі його померкли, і він не міг бачити.
1SAM|4|16|І сказав той чоловік до Ілія: Я той, що прибіг із бою, і я втік сьогодні з бойових лав. І сказав Ілій: Що то сталося, мій сину?
1SAM|4|17|І відповів вісник і сказав: Ізраїль побіг перед филистимлянами, і сталась велика поразка в народі. І обидва сини твої, Хофні та Пінхас, полягли. А ковчег Божий узятий!
1SAM|4|18|І сталося, як згадав він про Божого ковчега, то впав Ілій зо стільця навзнак при брамі, зламався карк йому, і він помер, бо той муж був старий та тяжкий. А він судив Ізраїля сорок літ.
1SAM|4|19|А невістка його, Пінхасова жінка, була важка, близька до родів. І як зачула вона ту звістку, що взятий Божий ковчег і помер тесть її та чоловік її, то впала на коліна, та й породила, бо прийшли на неї породільні болі її.
1SAM|4|20|А як настав час смерти її, то казали ті, що стояли при ній: Не бійся, бо ти породила сина! Та вона не відповіла, і не взяла цього до серця свого.
1SAM|4|21|І вона назвала ім'я тому хлопцеві: Іхавод, кажучи: Відійшла Ізраїлева слава! Бо почула про взяття Божого ковчегу, і про тестя свого та про мужа свого,
1SAM|4|22|та й сказала: Відійшла слава від Ізраїля, бо взятий Божий ковчег.
1SAM|5|1|А филистимляни взяли Божого ковчега, і принесли його з Евен-Гаезеру до Ашдоду.
1SAM|5|2|І взяли филистимляни Божого ковчега, і принесли його до Даґонового дому, і поставили його біля Даґона.
1SAM|5|3|А другого дня вранці повставали ашдодяни, аж ось Даґон лежить ницьма на землі перед Господнім ковчегом! І взяли вони Даґона, і поставили його на його місце.
1SAM|5|4|А наступного дня повставали вони рано, аж ось Даґон лежить ницьма на землі перед Господнім ковчегом! А Даґонова голова та обидві долоні рук його лежать відтяті на порозі, тільки тулуб Даґонів позостав при ньому.
1SAM|5|5|Тому то жерці та всі, хто входить до Даґонового дому, не ступають на Даґонів поріг у Ашдоді аж до цього дня.
1SAM|5|6|І стала тяжка Господня рука на ашдодян, і Він їх пустошив та бив їх болячками, Ашдод та довкілля його.
1SAM|5|7|І побачили ашдодяни, що так, та й сказали: Нехай не зостається з нами ковчег Ізраїлевого Бога, бо стала тяжкою Його рука на нас та на Даґона, бога нашого!
1SAM|5|8|І послали вони, і зібрали до себе всіх филистимських володарів, та й сказали: Що ми зробимо з ковчегом Ізраїлевого Бога? А ті відказали: Нехай ковчег Ізраїлевого Бога перейде до Ґату. І вони перенесли ковчега Ізраїлевого Бога.
1SAM|5|9|І сталося по тому, як вони перенесли його, то Господня рука була проти міста, сталося дуже велике замішання. І вдарив Він людей того міста від малого й аж до великого, і появилися на них болячки.
1SAM|5|10|І вони вислали Божого ковчега до Екрону. І сталося, як Божий ковчег прибув до Екрону, то екроняни стали кричати, говорячи: Перенесли до нас ковчега Ізраїлевого Бога, щоб вигубив нас та народ наш!
1SAM|5|11|І послали вони, і зібрали всіх филистимських володарів, та й говорили: Відішліть ковчега Ізраїлевого Бога, нехай вернеться на місце своє, і нехай не поб'є нас та народа нашого, бо було смертельне замішання в усьому місті. І Божа рука стала там дуже тяжка.
1SAM|5|12|А ті люди, хто не повмирав, були вдарені болячками, і зойк міста піднявся до неба!
1SAM|6|1|І був Божий ковчег у филистимській землі сім місяців.
1SAM|6|2|І покликали филистимляни жерців та ворожбитів, говорячи: Що робити з Господнім ковчегом? Скажіть нам, як відіслати його на його місце?
1SAM|6|3|А ті сказали: Якщо ви відсилаєте ковчега Ізраїлевого Бога, то не відсилайте його порожньо, але конче принесіть Йому жертву за провину, тоді будете вилікувані, і ви пізнаєте, чому не відступає Його рука від вас.
1SAM|6|4|І ті спитали: Яка ж та жертва за провину, що ми принесемо Йому? А ті відказали: За числом филистимських володарів п'ять золотих болячок та п'ять золотих мишей. Бо одна пораза для всіх вас та для ваших володарів.
1SAM|6|5|І зробіть подоби ваших болячок та подоби ваших мишей, що вигублюють землю, і воздайте славу Ізраїлевому Богові, може Він полегчить Свою руку з-над вас і з-над ваших богів та з-над вашого краю.
1SAM|6|6|І чого ви будете робити запеклими свої серця, як робили запеклим серце своє Єгипет та фараон? Чи ж не тоді, як Він чинив дивні речі з ними, не відпустили їх, і вони пішли?
1SAM|6|7|А тепер візьміть, і зробіть одного нового воза, і візьміть дві дійні корові, що на них не накладалося ярма, і запряжіть ті корови до воза, а їхні телята відведете від них додому.
1SAM|6|8|І візьмете Господнього ковчега, та й поставите його на воза, а золоті речі, що ви принесете Йому жертвою за провину, покладете в скрині збоку її. І відпустите його, і він піде.
1SAM|6|9|І побачите: Якщо він увійде до Бет-Шемешу дорогою до своєї границі, він зробив нам це велике зло. А якщо ні, то пізнаємо, що не його рука доторкнулася нас, випадок то був нам.
1SAM|6|10|І зробили ті люди так. І взяли вони дві дійні корові, і запрягли їх до воза, а їхніх телят замкнули вдома.
1SAM|6|11|І поставили вони Господнього ковчега на воза, і скриню, і золоті миші, і подоби їхніх болячок.
1SAM|6|12|І корови пішли просто дорогою до Бет-Шемешу. Ішли вони однією битою дорогою та все ревли, і не відхилялися ні праворуч, ні ліворуч. А филистимські володарі йшли за ними аж до границі Бет-Шемешу.
1SAM|6|13|А люди Бет-Шемешу жали пшеницю в долині. І звели вони очі свої та й побачили ковчега, і зраділи, що побачили!
1SAM|6|14|А віз увійшов на поле бетшемешанина Ісуса, та й став там, а там був великий камінь. І вони накололи дров із воза, а корів принесли цілопаленням для Господа.
1SAM|6|15|А Левити зняли Господнього ковчега та скриню, що була з ним, що в нім були золоті речі, та й поставили при великому камені. А люди Бет-Шемешу принесли цілопалення, і приносили того дня жертви для Господа.
1SAM|6|16|А п'ять филистимських володарів бачили це, і вернулися того дня до Екрону.
1SAM|6|17|А оце ті золоті болячки, що филистимляни звернули Господеві жертвою за провину: одна за Ашдод, одна за Газу, одна за Ашкелон, одна за Ґат, одна за Екрон.
1SAM|6|18|А золоті миші були за числом усіх филистимських міст п'ятьох володарів, від міста твердинного й аж до безмурного села, і аж до великого каменя, що на ньому поставили Господнього ковчега, і він знаходиться аж до цього дня на полі бет-шемешанина Ісуса.
1SAM|6|19|І вдарив Господь людей Бет-Шемешу, бо вони заглядали в Господній ковчег. І вибив Він між народом п'ятдесят тисяч чоловіка та сімдесят чоловіка. І був народ у жалобі, бо Господь ударив народ великою поразкою.
1SAM|6|20|І сказали люди Бет-Шемешу: Хто зможе стати перед лицем Господа, Того Бога Святого? І до кого Він піде від нас?
1SAM|6|21|І вони послали послів до мешканців Кір'ят-Єаріму, говорячи: Филистимляни вернули Господнього ковчега. Зійдіть, знесіть його до себе.
1SAM|7|1|І поприходили люди Кір'ят-Єаріму, та й підняли Господнього ковчега, і внесли його до Авінадавого дому на узгір'ї в Ґів'ї, а сина його Елеазара посвятили стерегти Господнього ковчега.
1SAM|7|2|І сталося, від дня, коли ковчег полишився у Кір'ят-Єарімі, минуло багато часу, а було його двадцять літ. А ввесь Ізраїлів дім плакав за Господом.
1SAM|7|3|І сказав Самуїл до всього Ізраїлевого дому, говорячи: Якщо ви цілим вашим серцем вертаєтеся до Господа, повикидайте з-поміж себе чужих богів та Астарт, і міцно прихиліть свої серця до Господа, і служіть Самому Йому, і Він спасе вас із руки филистимлян.
1SAM|7|4|І повикидали Ізраїлеві сини Ваалів та Астарт, та й служили Господеві, Самому Йому.
1SAM|7|5|І сказав Самуїл: Зберіть усього Ізраїля до Міцпи, а я буду молитися за вас до Господа!
1SAM|7|6|І зібралися до Міцпи, і черпали воду та лили перед Господнім лицем, і постили того дня, та й казали там: Ми згрішили перед Господом! І судив Самуїл Ізраїлевих синів у Міцпі.
1SAM|7|7|І почули филистимляни, що Ізраїлеві сини зібралися до Міцпи, і піднялися филистимські володарі на Ізраїля. І почули про це Ізраїлеві сини, та й злякалися филистимлян.
1SAM|7|8|І сказали Ізраїлеві сини до Самуїла: Не переставай кликати за нас до Господа, нашого Бога, і нехай Він спасе нас від руки филистимлян.
1SAM|7|9|І взяв Самуїл одне молочне ягня, і приніс його повним цілопаленням для Господа. І кликав Самуїл до Господа за Ізраїля, а Господь відповів йому.
1SAM|7|10|І приносив Самуїл цілопалення, а филистимляни приступили до бою проти Ізраїля. І загримів Господь того дня сильним громом на филистимлян, та й привів їх у замішання, і були вони побиті перед Ізраїлем.
1SAM|7|11|І повиходили Ізраїлеві люди з Міцпи, та й гнали филистимлян, і били їх аж під Бет-Кар.
1SAM|7|12|І взяв Самуїл одного каменя, і поклав між Міцпою та між Шенам, та й назвав ім'я йому: Евен-Єзер. І він сказав: Аж доти допоміг нам Господь.
1SAM|7|13|І були филистимляни переможені, і далі вже не входили в Ізраїлеві границі. І була Господня рука на филистимлянах за всі дні Самуїлові.
1SAM|7|14|І вернулися до Ізраїля ті міста, що филистимляни забрали були від Ізраїля, від Екрону й аж до Ґату, а їхню границю Ізраїль урятував від руки филистимлян. І був мир між Ізраїлем та між Амореянином.
1SAM|7|15|І судив Самуїл Ізраїля всі дні життя свого.
1SAM|7|16|І ходив він рік-річно, і обходив Бет-Ел, і Ґілґал, і Міцпу, і судив Ізраїля по всіх тих місцях.
1SAM|7|17|І вертався до Рами, бо там був дім його, і там судив Ізраїля. І він збудував там жертівника для Господа.
1SAM|8|1|І сталося, як Самуїл постарівся, то поставив синів своїх за суддів для Ізраїля.
1SAM|8|2|І було ім'я перворідного сина його Йоїл, а ім'я другого його Авійя, судді в Беер-Шеві.
1SAM|8|3|А сини його не йшли його дорогою, і вхилялись до зиску, і брали підкупа, і ламали Закона.
1SAM|8|4|І зібралися всі Ізраїлеві старші, і прийшли до Самуїла до Рами,
1SAM|8|5|та й сказали до нього: Ось ти постарівся, а сини твої не йдуть дорогами твоїми. Тепер настанови нам царя, щоб судив нас, як у всіх народів.
1SAM|8|6|І була та річ зла в Самуїлових очах, як вони сказали: Настанови нам царя, щоб судив нас. І молився Самуїл до Господа.
1SAM|8|7|І сказав Господь до Самуїла: Послухай голосу того народу щодо всього, про що він сказав тобі, бо не тобою вони погордували, але Мною погордували, щоб Я не царював над ними.
1SAM|8|8|Як усі ті діла, що вони чинили від дня, коли Я вивів їх з Єгипту, і аж до цього дня, і як вони кидали Мене й служили іншим богам, так вони чинять і тобі.
1SAM|8|9|А тепер послухай їхнього голосу, тільки конче остережеш їх, і розповіси їм право того царя, що буде царювати над ними.
1SAM|8|10|І переказав Самуїл всі Господні слова до народу, що жадав від нього царя,
1SAM|8|11|і сказав: Оце буде право царя, що царюватиме над вами: він візьме синів ваших і поставить собі в колесниці свої та серед їздців своїх, і вони будуть бігати перед колесницею його;
1SAM|8|12|і щоб поставити собі тисячників та п'ятдесятників, і щоб орати орку його, і щоб жати жниво його, і щоб робити зброю військову його та колесничні приладдя його.
1SAM|8|13|А дочок ваших забере за мироварниць, і за кухарок, і за пекарок.
1SAM|8|14|І він позабирає поля ваші, і виноградники ваші, та кращі ваші оливки, і пороздає своїм слугам.
1SAM|8|15|А з вашого посіву та з ваших виноградників братиме десятину, і даватиме своїм евнухам та своїм слугам.
1SAM|8|16|І він забере рабів ваших, і ваших невільниць, і найліпших ваших юнаків, і ваших ослів, і буде вживати їх на роботу свою.
1SAM|8|17|Він братиме десятину з вашої отари, а ви станете йому за рабів.
1SAM|8|18|І ви будете кликати того дня проти вашого царя, якого собі вибрали, та не відповість вам Господь того дня!
1SAM|8|19|Та народ відмовився слухати Самуїлового голосу, та й сказав: Ні, нехай тільки цар буде над нами!
1SAM|8|20|І будемо ми, як усі люди, і буде нас судити наш цар. І він ходитиме перед нами, і провадитиме наші війни.
1SAM|8|21|І вислухав Самуїл усі слова народу, і переказав їх голосно Господеві.
1SAM|8|22|А Господь сказав до Самуїла: Послухайся їхнього голосу, і постав їм царя! І сказав Самуїл до Ізраїлевих людей: Ідіть кожен до міста свого!
1SAM|9|1|І був чоловік із Веніяминового племени, а ім'я йому Кіш, син Авіїла, сина Церорового, сина Бехоратового, сина Афіяхового, веніяминівець, людина заможна.
1SAM|9|2|І був у нього син, а ім'я йому Саул, молодий та гарний. І з Ізраїлевих синів не було нікого вродливішого за нього, цілою головою він був вищий від кожного з усього народу.
1SAM|9|3|І пропали були Кішові, Сауловому батькові, ослиці. І сказав Кіш до свого сина Саула: Візьми з собою одного із слуг, і встань, іди, пошукай ослиці!
1SAM|9|4|І він перейшов Єфремові гори, і перейшов край Шаліша, та не знайшли. І перейшли вони край Шеаліму, та нема. І перейшов він край Веніяминів, та не знайшли.
1SAM|9|5|Увійшли вони до краю Цуф, і Саул сказав до свого слуги, що з ним: Давай вернімося, щоб не занехав батько ослиць, та не став журитися за нами!
1SAM|9|6|А той відказав йому: Ось у цьому місті є чоловік Божий, а той чоловік шанований. Усе, що він говорить, конче справджується. Тепер сходімо туди, може він покаже нам нашу дорогу, що нею ми пішли б.
1SAM|9|7|І сказав Саул до свого слуги: Ось ми підемо, та що ми принесемо цьому чоловікові? Бо хліб вийшов із наших торб, а подарунка нема, щоб принести Божому чоловікові. Що ми маємо?
1SAM|9|8|А той слуга далі відповідав Саулові та й сказав: Ось у руці моїй знаходиться чверть шекля срібла, і я дам Божому чоловікові, а він розповість нам про нашу дорогу.
1SAM|9|9|Колись в Ізраїлі, коли хто ходив питатися Бога, то так говорив: Давайте підемо до провидця. Бо що сьогодні, пророк, колись звалося провидець.
1SAM|9|10|І сказав Саул до свого слуги: Добре твоє слово. Давай підемо! І пішли вони до того міста, де був чоловік Божий.
1SAM|9|11|Коли вони підіймалися по узбіччях до міста, то знайшли дівчат, що вийшли були набрати води. І сказали вони до них: Чи є тут провидець?
1SAM|9|12|А ті відповіли їм та й сказали: Є, ось перед тобою! Поспіши тепер, бо сьогодні він прийшов до міста, бо сьогодні в народа жертва на пагірку.
1SAM|9|13|Як увійдете до міста, так знайдете його, поки він не вийде на пагірок їсти, бо народ не їсть аж до його приходу, бо він благословляє жертву, потім їдять покликані. А тепер увійдіть, бо зараз ви знайдете його.
1SAM|9|14|І піднялися вони до міста. Як вони входили до середини того міста, аж ось Самуїл виходить навпроти них, щоб іти на пагірок.
1SAM|9|15|А Господь, за день перед Сауловим приходом, виявив був Самуїлові, говорячи:
1SAM|9|16|Цього часу взавтра пошлю до тебе чоловіка з Веніяминового краю, і ти помажеш його на володаря над Моїм Ізраїлевим народом, і він спасе народ Мій від руки филистимлян. Я бо зглянувся на народ Мій, бо голосіння його дійшло до Мене!
1SAM|9|17|А коли Самуїл побачив Саула, то Господь сказав йому: Оце той чоловік, що Я казав тобі, він володітиме народом Моїм.
1SAM|9|18|І підійшов Саул до Самуїла в середині брами та й сказав: Скажи мені, де тут дім провидця?
1SAM|9|19|І відповів Самуїл Саулові та й сказав: Я той провидець. Вийди перед мене на пагірок, і ви будете їсти зо мною сьогодні. А рано я відпущу тебе, і про все, що в серці твоїм, я розповім тобі.
1SAM|9|20|А щодо ослиць, що пропали тобі, сьогодні вже три дні, не журися за них, бо знайшлися вони. Та для кого все пожадане в Ізраїлі? Хіба ж не для тебе та для всього дому батька твого?
1SAM|9|21|І відповів Саул та й сказав: Чи ж я не веніяминівець, із найменших Ізраїлевих племен? А рід мій найменший з усіх родів Веніяминового племени. І чого ти говориш мені отаке слово?
1SAM|9|22|І взяв Самуїл Саула та слугу його, і ввів їх до кімнати, і дав їм місце на чолі покликаних, а тих було близько тридцяти чоловіка.
1SAM|9|23|І сказав Самуїл до кухаря: Дай же ту частку, що дав я тобі, що про неї я сказав тобі: Відклади її в себе!
1SAM|9|24|І подав кухар стегно та те, що на ньому, і поклав перед Саулом. А Самуїл сказав: Оце позоставлене! Поклади перед собою та їж, бо воно сховане для тебе на умовлений час, коли я сказав: Покликав я народ. І Саул їв із Самуїлом того дня.
1SAM|9|25|І зійшли вони з пагірка до міста, і він розмовляв із Саулом на даху свого дому.
1SAM|9|26|І повставали вони рано вранці. І сталося, як зійшла рання зоря, то Самуїл кликнув до Саула на дах, говорячи: Уставай же, і я відпушу тебе! І встав Саул, і вони вийшли обоє, він та Саул, на вулицю.
1SAM|9|27|Коли вони підходили на край міста, то Самуїл сказав до Саула: Скажи тому слузі, і нехай він іде перед нами. І той пішов. А ти зараз спинися, я оголошу тобі Боже слово!
1SAM|10|1|І взяв Самуїл посудинку оливи, та й вилляв на його голову, і поцілував його та й сказав: Чи це не помазав тебе Господь над спадком Своїм на володаря? (І будеш ти царювати над народом Господнім, і ти визволиш його від руки ворогів його навколо. І ось тобі ознака, що Господь помазав тебе над спадком Своїм на володаря.)
1SAM|10|2|Як підеш ти сьогодні від мене, то при Рахилинім гробі, у Веніяминовій країні в Целцаху, знайдеш двох людей, і вони скажуть тобі: Знайдені ті ослиці, яких ти шукати ходив. А оце батько твій занехаяв справи тих ослиць, та й зажурився за вас, говорячи: Що я зроблю для свого сина?
1SAM|10|3|І перейдеш ти звідти й далі, і підеш аж до діброви Фаворської, а там знайдуть тебе три чоловіки, що йдуть до Бога до Бет-Елу, один несе трьох ягнят, а один несе три буханці хліба, а один несе бурдюка вина.
1SAM|10|4|І запитають вони тебе про мир, та дадуть тобі два хліби, і ти візьмеш із їхньої руки.
1SAM|10|5|Потому вийдеш ти на Божий горбок, де намісники филистимські. І станеться, як ти ввійдеш там до міста, то стрінеш громаду пророків, що сходять з пагірка, а перед ними арфа, та бубон, та сопілка, та цитра, і вони пророкують.
1SAM|10|6|І злине на тебе Дух Господній, і ти будеш з ними пророкувати, і станеш іншою людиною.
1SAM|10|7|І станеться, коли збудуться тобі ці ознаки, роби собі, що знайде рука твоя, бо Бог з тобою.
1SAM|10|8|І зійдеш ти передо мною до Ґілґалу, а я зійду до тебе, щоб принести цілопалення, щоб приносити мирні жертви. Сім день будеш чекати, аж поки прийду я до тебе, і завідомлю тебе, що будеш робити.
1SAM|10|9|І сталося, як повернувся він, щоб іти від Самуїла, то Бог змінив йому серце на інше, а всі ті ознаки прийшли того дня.
1SAM|10|10|І прийшли вони туди до Ґів'ї, аж ось громада пророків назустріч йому. І злинув на нього Дух Божий, і він пророкував серед них.
1SAM|10|11|І сталося, кожен, хто знав його віддавна, а тепер побачили, ось він пророкує разом із пророками, то казали один до одного: Що то сталося Кішовому синові? Чи й Саул між пророками?
1SAM|10|12|І відповів чоловік звідти й сказав: А хто їній батько? Тому то стало за приказку: Чи й Саул між пророками?
1SAM|10|13|І перестав він пророкувати, і прийшов на пагірок.
1SAM|10|14|І сказав Саулів дядько до нього та до слуги його: Куди ви ходили? А той відказав: Шукати ослиць. І побачили ми, що нема, і прийшли до Самуїла.
1SAM|10|15|А дядько Саулів сказав: Скажи ж мені, що сказав вам Самуїл?
1SAM|10|16|І сказав Саул до дядька свого: Справді розповів нам, що знайдені ті ослиці. А про справу царства, що говорив Самуїл, не розповів йому.
1SAM|10|17|І скликав Самуїл народ до Господа, до Міцпи,
1SAM|10|18|та й сказав до Ізраїлевих синів: Так сказав Господь, Бог Ізраїлів: Я вивів Ізраїля з Єгипту, і спас вас із руки Єгипту та з руки всіх царств, що гнобили вас.
1SAM|10|19|А ви сьогодні погордували своїм Богом, що Він спасає вас з усіх нещасть ваших та утисків ваших. І ви сказали йому: Ні, таки царя постав над нами. А тепер ставайте перед Господнім лицем за вашими племенами та за вашими тисячами.
1SAM|10|20|І привів Самуїл усі Ізраїлеві племена, і було виявлене Веніяминове плем'я.
1SAM|10|21|І привів він Веніяминове плем'я за родами його, і був виявлений рід Матріїв. І привів він рід Матріїв за їхніми мужчинами, і був виявлений Саул, син Кішів. І шукали його, та не знаходили.
1SAM|10|22|І питалися Господа ще: Чи прийде він ще сюди? А Господь відповів: Он він заховався між речами!
1SAM|10|23|І вони побігли, і взяли його звідти. І він став серед народу, і був вищий від усього народу на цілу голову.
1SAM|10|24|І сказав Самуїл до всього народу: Чи бачите, кого вибрав Господь? Бо нема такого, як він, серед усього народу. І ввесь народ ізняв крик та й сказав: Хай живе цар!
1SAM|10|25|А Самуїл промовляв до народу про права царства, і записав те до книги, та й поклав перед Господнім лицем. І відпустив Самуїл увесь народ, кожного до дому свого.
1SAM|10|26|І також Саул пішов до дому свого до Ґів'ї, а з ним пішли ті вояки, що Господь діткнувся їхніх сердець.
1SAM|10|27|А негідні сини говорили: Що, нас спасе отакий? І гордували ним, і не принесли йому дара. Та він мовчав.
1SAM|11|1|І вийшов аммонітянин Нахаш, і таборував при ґілеадському Явешу. І сказали всі явеські люди до Нахаша: Склади з нами умову, і ми будемо служити тобі!
1SAM|11|2|І сказав до них аммонітянин Нахаш: Про це складу з вами умову, щоб кожному з вас вибрати праве око, і я вчиню це на ганьбу для всього Ізраїля.
1SAM|11|3|І сказали до нього явеські старші: Зачекай нам сім день, і нехай ми пошлемо послів у всі Ізраїлеві краї. І якщо нема нам порятунку, то вийдемо до тебе.
1SAM|11|4|І прийшли ті посли до Саулової Ґів'ї, і говорили ті слова до ушей народу. І ввесь народ підніс свій голос, та й заплакав.
1SAM|11|5|Аж ось Саул іде худобою з поля. І сказав Саул: Що народові, що плачуть? І розповіли йому слова явеських людей.
1SAM|11|6|І злинув Божий Дух на Саула, як слухав він ті слова, і дуже запалав його гнів!
1SAM|11|7|І взяв він пару худобин, і порізав її, і порозсилав по всім Ізраїлевім Краї через послів, говорячи: Хто не вийде за Саулом та за Самуїлом, отак буде зроблено худобі його! І великий страх спав на людей, і вони повиходили, як один чоловік.
1SAM|11|8|І він перелічив їх у Безеку, і було Ізраїлевих синів триста тисяч, а Юдиних людей тридцять тисяч.
1SAM|11|9|І сказали вони до послів, що прийшли: Так скажете мешканцям ґілеадського Явешу: Узавтра, як пригріє сонце, буде вам порятунок. І прийшли ті посли, і розповіли явеським людям, і вони зраділи.
1SAM|11|10|І сказали явеські люди: Узавтра ми вийдемо до вас, а ви зробите нам усе, що добре в очах ваших.
1SAM|11|11|І сталося назавтра, і склав Саул із народу три відділи, і вони пройшли в середину табору за ранньої сторожі, та й били Аммона аж до спекоти дня. І сталося, позосталі розбіглися, і не позосталося між ними двох разом.
1SAM|11|12|І сказав народ до Самуїла: Хто той, що запитував: Саул буде царювати над нами? Дайте тих людей, а ми їх повбиваємо!
1SAM|11|13|Та Саул сказав: Ніхто не буде забитий цього дня, бо Господь сьогодні зробив спасіння серед Ізраїля.
1SAM|11|14|А Самуїл сказав до народу: Ходіть, і підемо в Ґілґал, та й відновимо там царство!
1SAM|11|15|І пішов увесь народ до Ґілґалу, і настановили царем там Саула перед Господнім лицем у Ґілґалі, і приносили мирні жертви перед Господнім лицем. І дуже радів там Саул та всі Ізраїлеві мужі!
1SAM|12|1|І сказав Самуїл до всього Ізраїля: Ось я послухався вашого голосу в усьому, що ви говорили мені, і поставив над вами царя.
1SAM|12|2|А тепер той цар ось ходить перед вами. А я постарів та посивів, а сини мої ось вони з вами. І я ходив перед вами від своєї молодости аж до до цього дня.
1SAM|12|3|Ось! Свідкуйте проти мене перед Господом та перед Його помазанцем: чийого вола я взяв, чи осла чийого взяв я? А кого я гнобив, кому чинив насильство? І з чиєї руки взяв я підкупа, і відвернув свої очі від нього? І все це я поверну вам.
1SAM|12|4|А вони сказали: Не гнобив ти нас, і не чинив нам насильства, і ні від кого нічого не брав.
1SAM|12|5|І він сказав: Господь свідок на вас, і свідок Його помазанець цього дня, що ви нічого не знайшли в моїй руці. А народ сказав: Свідок!
1SAM|12|6|І сказав Самуїл до народу: Свідок Господь, що поставив Мойсея та Аарона, і що вивів наших батьків із єгипетського краю.
1SAM|12|7|А тепер станьте, і я буду судитися з вами перед Господнім лицем про всі добродійства Господні, які Він учинив із вами та з вашими батьками.
1SAM|12|8|Як Яків прийшов був до Єгипту, і батьки ваші кликали до Господа, то Господь послав Мойсея та Аарона, і вони вивели ваших батьків із Єгипту, і осадили їх у цьому місці.
1SAM|12|9|Та вони забули Господа, Бога свого, і Він передав їх у руку Сісери, начальника хацорського війська, і в руку филистимлян та в руку моавського царя, і вони воювали проти них.
1SAM|12|10|І кликали вони до Господа та говорили: Згрішили ми, бо покинули Господа та й служили Ваалам та Астартам. А тепер урятуй нас із руки наших ворогів, і ми будемо служити Тобі.
1SAM|12|11|І послав Господь Єруббаала, і Бедана, і Їфтаха, і Самуїла, і врятував вас із руки довколишніх ваших ворогів, і ви сиділи безпечно.
1SAM|12|12|А коли ви побачили, що Нахаш, цар аммонських синів, прийшов на вас, то сказали мені: Ні, нехай царює над нами цар! А Цар ваш Господь, Бог ваш.
1SAM|12|13|А тепер ось той цар, якого ви вибрали, якого жадали, і ось дав Господь над вами царя.
1SAM|12|14|Якщо ви будете боятися Господа, і будете служити Йому, і будете слухатися Його голосу, і не будете непокірні до Господніх заповідей, то будете й ви, і цар, що царює над вами, ходити за Господом, Богом вашим.
1SAM|12|15|А якщо ви не будете слухатися Господнього голосу, і будете непокірні до Господніх заповідей, то Господня рука буде проти вас та проти ваших батьків!
1SAM|12|16|І ось тепер станьте, і побачте ту велику річ, що Господь зробить на ваших очах.
1SAM|12|17|Чи ж сьогодні не жнива на пшеницю? Я покличу до Господа, і Він пошле грім та дощ, а ви пізнаєте й побачите, що велике ваше зло, яке ви зробили в Господніх очах жаданням для себе царя.
1SAM|12|18|І кликнув Самуїл до Господа, а Господь послав того дня грім та дощ. І ввесь народ сильно злякався Господа та Самуїла!
1SAM|12|19|І сказав увесь народ до Самуїла: Помолися за своїх рабів до Господа, Бога твого, щоб нам не померти, бо понад усі наші гріхи додали ми ще й оце зло, що жадали для себе царя.
1SAM|12|20|І сказав Самуїл до народу: Не бійтеся! Ви зробили все те зло, тільки не відступіть від Господа, і служіть Господеві всім серцем своїм!
1SAM|12|21|І не відступайте, і не йдіть за марнотами, які не допоможуть і які не врятують, бо марнота вони.
1SAM|12|22|Бо Господь не полишить народу Свого ради Свого великого Ймення, бо зволив Господь зробити вас народом Своїм.
1SAM|12|23|Також я, не дай мені, Боже, грішити проти Господа, щоб перестав я молитися за вас! І я буду наставляти вас на дорогу добру та просту.
1SAM|12|24|Тільки бійтеся Господа, і служіть Йому правдиво всім вашим серцем, бо ви бачили, які великі діла вчинив Він із вами!
1SAM|12|25|А якщо справді будете чинити зло, погинете й ви, і цар ваш!
1SAM|13|1|Рік був, як Саул зацарював, і два роки царював над Ізраїлем.
1SAM|13|2|І вибрав собі Саул три тисячі з Ізраїля, дві тисячі були з Саулом у Міхмаші та на горі Бет-Елу, а тисяча були з Йонатаном у Веніяминовій Ґів'ї. А решту народу відпустив він кожного до наметів своїх.
1SAM|13|3|І побив Йонатан филистимського намісника, що в Ґеві. І почули це филистимляни, а Саул засурмив у сурму по всьому Краю, говорячи: Нехай почують євреї!
1SAM|13|4|А ввесь Ізраїль чув, говорячи: Саул побив филистимського намісника, і тим Ізраїль став ненависним серед филистимлян. І скликаний був народ за Саулом до Ґілґалу.
1SAM|13|5|А филистимляни були зібрані воювати з Ізраїлем, тридцять тисяч возів і шість тисяч верхівців, а народу, щодо численности, як піску на морському березі. І вийшли вони, і таборували в Міхмаші, на схід Бет-Авену.
1SAM|13|6|А Ізраїльтянин побачив, що скрутно йому, що народ був пригноблений, і народ ховався по печерах, і по щілинах, і по скелях, і по льохах та по ямах.
1SAM|13|7|А інші євреї перейшли Йордан до краю Ґада та до Ґілеаду. А Саул був ще у Ґілґалі, а ввесь народ із тривогою поспішав за ним.
1SAM|13|8|І чекав він сім день умовленого часу, що призначив Самуїл, та Самуїл не прийшов до Ґілґалу, і народ став розбігатися від нього.
1SAM|13|9|І сказав Саул: Приведіть до мене призначене на цілопалення та мирні жертви. І він приніс цілопалення.
1SAM|13|10|І сталося, як скінчив він приносити цілопалення, то ось приходить Самуїл. І вийшов Саул, щоб зустріти його, щоб привітати його.
1SAM|13|11|І сказав Самуїл: Що ти зробив? А Саул відказав: Бо я бачив, що народ розбігається від мене, а ти не прийшов на умовлений час тих днів. А филистимляни зібралися в Міхмаші.
1SAM|13|12|І я сказав: Тепер филистимляни зійдуть до мене до Ґілґалу, а Господнього лиця я ще не вблагав. І я вирішив, і приніс цілопалення!
1SAM|13|13|І сказав Самуїл до Саула: Ти зробив нерозумне! Не послухав ти наказів Господа, Бога свого, що наказав був тобі, бо тепер Господь міцно поставив би аж навіки твоє царство над Ізраїлем.
1SAM|13|14|А тепер царство твоє не буде стояти, Господь пошукав Собі мужа за серцем Своїм, і Господь наказав йому бути володарем над народом Своїм, бо ти не виконав, що наказав був тобі Господь.
1SAM|13|15|І встав Самуїл, і зійшов із Ґілґалу до Веніяминової Ґів'ї. А Саул перелічив народ, що знаходився з ним, близько шости сотень чоловіка.
1SAM|13|16|І Саул і син його Йонатан та народ, що знаходився з ним, сиділи в Веніяминовій Ґеві, филистимляни ж таборували в Міхмаші.
1SAM|13|17|І вийшли руїнники з филистимського табору трьома відділами: один відділ звертається на офрійську дорогу до краю Шуал,
1SAM|13|18|і один відділ звертається на дорогу до Бет-Хорону, а один відділ звертається на дорогу до границі, що провадить від Ґе-Цевоїму до пустині.
1SAM|13|19|А коваля не було по всім Ізраїлевім Краї, бо филистимляни сказали: Щоб не робили євреї меча чи списа!
1SAM|13|20|І сходив увесь Ізраїль до филистимлян гострити кожен свого плуга, і заступа свого, і сокиру свою, і серпа свого,
1SAM|13|21|коли тупилися вістря плугів, і заступів, і вил, і сокир, і мусіли сходити, щоб направити вістря рожна.
1SAM|13|22|І сталося за днів війни, і не знайшлося ані меча, ані списа в руці всього народу, що був з Саулом та з Йонатаном, та був знайдений тільки для Саула та для сина його Йонатана.
1SAM|13|23|І вийшла филистимська залога до переходу Міхмашу.
1SAM|14|1|Одного дня сказав Йонатан, син Саулів, до слуги, свого зброєноші: Ходім, і перейдімо до филистимської залоги, що з того боку. А батькові своєму він цього не розповів.
1SAM|14|2|А Саул сидів на кінці згір'я під гранатовим деревом, що в Міґроні. А народу, що з ним, було близько шости сотень чоловіка.
1SAM|14|3|А Ахійя, син Ахітува, брата Іхавода, сина Пінхаса, сина Ілія, священика в Шіло, носив ефода. А народ не знав, що пішов Йонатан.
1SAM|14|4|А між тими переходами, що Йонатан хотів перейти до филистимської залоги, була зубчаста скеля з цього боку переходу й зубчаста скеля з того боку переходу. А ім'я одній Боцец, а ім'я другій Сенне.
1SAM|14|5|Один зуб скеля стовп із півночі, навпроти Міхмашу, а один із півдня, навпроти Ґеви.
1SAM|14|6|І сказав Йонатан до слуги, свого зброєноші: Ходім, і перейдімо до сторожі тих необрізаних, може Господь зробить поміч для нас, бо Господеві нема перешкоди спасати через багатьох чи через небагатьох.
1SAM|14|7|І сказав йому його зброєноша: Роби все, що на серці твоїм! Звертай собі, ось я з тобою, куди хоче серце твоє.
1SAM|14|8|І сказав Йонатан: Ось ми приходимо до тих людей, і покажемось їм.
1SAM|14|9|Якщо вони скажуть до нас так: Стійте тихо, аж ми прийдемо до вас, то ми станемо на своєму місці, і не підіймемося до них.
1SAM|14|10|А якщо вони скажуть так: Підійміться до нас, то підіймемося, бо Господь дав їх у нашу руку. Це для нас буде знаком.
1SAM|14|11|І вони обидва показалися филистимській сторожі. І сказали филистимляни: Ось виходять із щілин євреї, що поховалися там.
1SAM|14|12|І люди залоги відповіли Йонатанові та його зброєноші та й сказали: Підіймися до нас, і ми вам щось скажемо! І сказав Йонатан зброєноші своєму: Підіймайся за мною, бо Господь дав їх у Ізраїлеву руку!
1SAM|14|13|І піднявся Йонатан на руках своїх та на ногах своїх, а за ним його зброєноша. І падали филистимляни перед Йонатаном, а його зброєноша добивав за ним.
1SAM|14|14|І була перша поразка, що вдарив Йонатан та його зброєноша, близько двадцяти чоловіка, на половині скиби оброблюваного парою волів поля на день.
1SAM|14|15|І стався сполох у таборі, на полі, та в усьому народі. Залога та нищителі затремтіли й вони. І задрижала земля, і знявся великий сполох!
1SAM|14|16|І побачили Саулові вартівники в Веніяминовій Ґів'ї, аж ось натовп розпливається, і біжить сюди та туди.
1SAM|14|17|І сказав Саул до народу, що був з ним: Перегляньте й побачте, хто пішов від нас? І переглянули, аж ось нема Йонатана та його зброєноші.
1SAM|14|18|І сказав Саул до Ахійї: Принеси Божого ковчега! Бо Божий ковчег був того дня з Ізраїлевими синами.
1SAM|14|19|І сталося, коли Саул говорив до священика, то замішання в филистимському таборі все більшало та ширилось. І сказав Саул до священика: Спини свою руку!
1SAM|14|20|І зібралися Саул та ввесь народ, що був із ним, і вони пішли аж до місця бою, аж ось меч кожного на його ближнього, замішання дуже велике!
1SAM|14|21|А між филистимлянами, як і давніш, були євреї, що поприходили з ними з табором, і вони теж перейшли, щоб бути з Ізраїлем, що був із Саулом та Йонатаном.
1SAM|14|22|А всі ізраїльтяни, що ховалися в Єфремових горах, почули, що филистимляни втікають, і погналися за ними й вони до бою.
1SAM|14|23|І спас Господь Ізраїля того дня. А бій перейшов аж за Бет-Евен.
1SAM|14|24|Та ізраїльтянин був пригноблений того дня. А Саул наклав клятву на народ, говорячи: Проклятий той чоловік, що буде їсти хліб до вечора, поки я пімщуся на своїх ворогах. І ввесь той народ не їв хліба.
1SAM|14|25|І ввесь народ пішов до лісу, а там був мед на галявині.
1SAM|14|26|І ввійшов народ до того лісу, аж ось струмок меду! Та ніхто не простяг своєї руки до уст своїх, бо народ боявся присяги.
1SAM|14|27|А Йонатан не чув, коли батько його заприсягнув був народ. І простягнув він кінець кия, що був у руці його, і вмочив його в стільник меду, та й підніс руку свою до уст своїх. І роз'яснилися очі йому!
1SAM|14|28|А на це один із народу промовив і сказав: Заприсягаючи, заприсяг твій батько народ, говорячи: Проклятий той чоловік, що буде їсти хліб сьогодні! І змучився від цього народ.
1SAM|14|29|І сказав Йонатан: Знещасливив мій батько цю землю! Подивіться но, як роз'яснилися очі мої, коли я скуштував трохи цього меду.
1SAM|14|30|А що, коли б народ сьогодні справді був їв зо здобичі своїх ворогів, що знайшов? Чи тепер не збільшилася б поразка филистимлян?
1SAM|14|31|І били вони того дня між филистимлянами від Міхмашу аж до Айялону. А народ дуже змучився.
1SAM|14|32|І кинувся народ на здобич, і позабирали худобу дрібну й худобу велику та телят, та й різали на землю. І їв народ із кров'ю!
1SAM|14|33|І розповіли Саулові, кажучи: Ось народ грішить проти Господа, їсть із кров'ю! А той відказав: Зрадили ви! Прикотіть до мене сьогодні великого каменя.
1SAM|14|34|І сказав Саул: Розійдіться між людьми, та й скажіть їм: Приведіть до нас кожен вола свого, і кожен штуку дрібної худобини, і заріжте тут. І будете їсти, і не згрішите проти Господа, якщо не будете їсти з кров'ю. І поприводив увесь народ тієї ночі кожен вола свого своєю рукою, і порізали там.
1SAM|14|35|І збудував Саул жертівника для Господа; його першого зачав він будувати, як жертівника для Господа.
1SAM|14|36|І сказав Саул: Зійдімо вночі за филистимлянами, та й винищуймо їх аж до ранкового світла, і не полишімо між ними нікого. А вони сказали: Роби все, що добре в очах твоїх. А священик сказав: Приступімо тут до Бога!
1SAM|14|37|І запитався Саул Бога: Чи зійти за филистимлянами? Чи даси їх в Ізраїлеву руку? Та Він не відповів йому того дня.
1SAM|14|38|І сказав Саул: Зійдіться сюди всі видатні народу, і пізнайте та побачте, у чому стався той гріх сьогодні.
1SAM|14|39|Бо як живий Господь, що допоміг Ізраїлеві, якщо він був хоча б на сині моїм Йонатані, то конче помре він! Та ніхто не відповів йому з усього народу.
1SAM|14|40|І сказав він до всього Ізраїля: Ви станете на один бік, а я та син мій Йонатан на другий бік. І сказав той народ до Саула: Зроби, що добре в очах твоїх!
1SAM|14|41|І сказав Саул до Господа, Бога Ізраїля: Дай же тумім! І був виявлений жеребком Йонатан та Саул, а народ повиходив оправданим.
1SAM|14|42|І сказав Саул: Киньте поміж мною та поміж сином моїм Йонатаном. І був виявлений Йонатан.
1SAM|14|43|І сказав Саул до Йонатана: Розкажи мені, що ти зробив? І розповів йому Йонатан і сказав: Я справді скуштував кінцем кия, що був у руці моїй, трохи меду. Ось я помру за це!
1SAM|14|44|І сказав Саул: Так нехай зробить Бог, і так нехай додасть, що конче помреш, Йонатане!
1SAM|14|45|А народ сказав до Саула: Чи помирати Йонатанові, що зробив оце велике спасіння в Ізраїлі? Борони Боже! Як живий Господь, не спаде волосина з голови його на землю, бо з Богом робив він цього дня! І визволив народ Йонатана, і він не помер.
1SAM|14|46|І відійшов Саул від филистимлян, а филистимляни пішли на своє місце.
1SAM|14|47|І здобув Саул царювання над Ізраїлем, і воював навколо зо всіма своїми ворогами: з Моавом, і з синами Аммона, і з Едомом, і з царями Цови, і з филистимлянами. І скрізь, проти кого він обертався, мав успіх.
1SAM|14|48|І склав він військо, та й побив Амалика, і врятував Ізраїля з руки грабіжника.
1SAM|14|49|І були в Саула сини: Йонатан, і Їшві, і Малкішуя; а ім'я двох дочок його: ім'я старшій Мерав, а ім'я молодшій Мелхола.
1SAM|14|50|А ім'я Саулової жінки: Ахіноам, дочка Ахімааца. А ім'я провідника його війська: Авнер, син Нера, Саулового дядька.
1SAM|14|51|А Кіш батько Саулів, а Нер батько Авнера, син Авіїлів.
1SAM|14|52|І була сильна війна на филистимлян за всіх Саулових днів. І коли Саул бачив якого чоловіка хороброго та якого сильного, то брав його до себе.
1SAM|15|1|І сказав Самуїл до Саула: Господь послав був мене помазати тебе на царя над народом Його, над Ізраїлем. А тепер послухайся голосу Господніх слів.
1SAM|15|2|Так сказав Господь Саваот: Я згадаю, що зробив був Амалик Ізраїлеві, що клав йому перешкоду на дорозі, коли він виходив із Єгипту.
1SAM|15|3|Тепер іди, і поб'єш Амалика, і вчиниш закляттям усе, що його, і не змилосердишся над ним. І позабиваєш усе, від чоловіка аж до жінки, від дитини й аж до немовляти, від вола й аж до штуки дрібної худобини, від верблюда й аж до осла.
1SAM|15|4|І Саул оповістив народ, і перелічив їх у Телаїмі, і двісті тисяч піхоти та десять тисяч мужа Юди.
1SAM|15|5|І прийшов Саул аж до Амаликового міста, та й засів у долині.
1SAM|15|6|І сказав Саул кенеянам: Ідіть, відокремтесь, вийдіть з-поміж Амаликитянина, щоб я не долучив вас до них, бо ви зробили були милість усім ізраїльтянам, коли вони виходили з Єгипту. І відокремився Кенеянин з-поміж Амалика.
1SAM|15|7|А Саул побив Амалика від Хавіли аж до місця, де йдеш до Шуру, що навпроти Єгипту.
1SAM|15|8|І зловив він Аґаґа, амаликського царя, живого, а ввесь народ зробив закляттям, та й побив вістрям меча.
1SAM|15|9|Та змилосердився Саул і народ над Аґаґом, і над найліпшим з його худоби дрібної й з худоби його великої та з товару вгодованого, і над вівцями, та над усім добром, і не хотіли зробити їх закляттям. А все маловарте й худе його зробили закляттям.
1SAM|15|10|І було Господнє слово до Самуїла й казало:
1SAM|15|11|Жалкую, що Я настановив Саула за царя, бо він відвернувся від Мене, а слів Моїх не виконав. І запалився гнів Самуїлів, і він кликав до Господа цілу ніч.
1SAM|15|12|А рано вранці Самуїл устав, і пішов назустріч Саулові. І Самуїлові донесли, говорячи: Саул прийшов до Кармелу, і ось ставить собі пам'ятника, а потому повернувся й пішов, і зійшов до Ґілґалу.
1SAM|15|13|І прийшов Самуїл до Саула, а Саул сказав йому: Благословенний ти в Господа! Я виконав слово Господнє.
1SAM|15|14|А Самуїл сказав: А що це за мекання цієї отари в ушах моїх, та рик великої худоби, що я чую?
1SAM|15|15|І сказав Саул: Від Амаликитянина привели їх, бо народ змилосердився над найліпшим із худоби дрібної та з худоби великої, щоб зарізати в жертву для Господа, Бога твого, а позостале вчинили закляттям.
1SAM|15|16|А Самуїл сказав до Саула: Покинь, а я розповім тобі, що Господь говорив мені цієї ночі. А той сказав йому: Говори.
1SAM|15|17|І сказав Самуїл: Хоч ти малий був в очах своїх, чи ж ти не голова Ізраїлевих племен? Чи ж не помазав тебе Господь на царя над Ізраїлем?
1SAM|15|18|І послав тебе Господь дорогою, і сказав: Іди, і вчиниш закляттям нечестивих амаликитян, і будеш воювати з ними, аж поки ти не вигубиш їх.
1SAM|15|19|І чому ти не послухався Господнього голосу, але кинувся на здобич, і зробив оце зло в Господніх очах?
1SAM|15|20|І сказав Саул до Самуїла: Та я послухався Господнього голосу, і пішов дорогою, якою послав був мене Господь, і привів я Аґаґа, царя амаликського, а Амалика зробив закляттям.
1SAM|15|21|А народ узяв зо здобичі худобу дрібну та худобу велику, як початок закляття, щоб приносити в жертву Господеві, Богові твоєму, в Ґілґалі.
1SAM|15|22|І сказав Самуїл: Чи жадання Господа цілопалень та жертов таке, як послух Господньому голосу? Таж послух ліпший від жертви, покірливість краща від баранячого лою!
1SAM|15|23|Бо непокірливість як гріх ворожбитства, а свавільство як провина та служба бовванам. Через те, що ти відкинув Господні слова, то Він відкинув тебе, щоб не був ти царем.
1SAM|15|24|І сказав Саул до Самуїла: Прогрішився я, бо переступив накази Господні та слова твої, бо я боявся народу, та послухався його голосу.
1SAM|15|25|А тепер прости ж мій гріх, і вернися зо мною, і я поклонюсь Господеві.
1SAM|15|26|Та Самуїл сказав до Саула: Не вернуся з тобою, бо ти погордив Господнім словом, а Господь погордив тобою, щоб не був ти царем над Ізраїлем.
1SAM|15|27|І повернувся Самуїл, щоб піти, а Саул схопив полу плаща його, та й відірвав.
1SAM|15|28|І сказав до нього Самуїл: Господь відірвав сьогодні від тебе Ізраїлеве царство, та й передав його твоєму ближньому, ліпшому від тебе!
1SAM|15|29|І також Ізраїлева Слава не скаже неправди та не буде каятися, бо Він не людина, щоб каятись.
1SAM|15|30|А Саул сказав: Прогрішився я! Але вшануй й мене перед старшими мого народу та перед Ізраїлем, і вернися зо мною, а я поклонюся Господеві, Богові твоєму.
1SAM|15|31|І вернувся Самуїл за Саулом, і Саул поклонився Господеві.
1SAM|15|32|І сказав Самуїл: Підведіть до мене Аґаґа, царя амаликського. І пішов до нього Аґаґ весело. І сказав Аґаґ: Справді, відступилася гіркота смерти!
1SAM|15|33|А Самуїл сказав: Як твій меч позбавляв жінок дітей, так позбавиться дітей твоя мати між жінками. І посік Самуїл Аґаґа перед Господнім лицем у Ґілґалі.
1SAM|15|34|І пішов Самуїл до Рами, а Саул зійшов до дому свого, до Саулової Ґів'ї.
1SAM|15|35|І більше не бачив Самуїл Саула аж до дня його смерти, та Самуїл сумував за Саулом. А Господь жалкував, що настановив був Саула царем над Ізраїлем.
1SAM|16|1|І сказав Господь до Самуїла: Аж доки ти сумуватимеш за Саулом? Таж Я відкинув його, щоб не царював над Ізраїлем. Наповни рога свого оливою, та й іди, пошлю тебе до віфлеємлянина Єссея, бо Я наглянув Собі царя між синами його.
1SAM|16|2|І сказав Самуїл: Як я піду? А почує Саул, то вб'є мене. А Господь сказав: Візьми в свою руку теля з великої худоби, та й скажеш: Я прийшов, щоб принести жертву для Господа.
1SAM|16|3|І закличеш Єссея на жертву, а Я тобі дам знати, що маєш робити, і помажеш Мені того, кого скажу тобі.
1SAM|16|4|І зробив Самуїл, що Господь говорив. І прийшов він до Віфлеєму, а старші міста вийшли йому назустріч із тремтінням. І сказали вони: Чи твій прихід то мир?
1SAM|16|5|А він відказав: Мир! Я прийшов, щоб принести жертву Господеві. Освятіться, і прийдете зо мною до жертви. І освятив він Єссея та синів його, і покликав їх на жертву.
1SAM|16|6|І сталося, як вони поприходили, то побачив він Еліява, та й сказав: Справді перед Господом помазанець Його!
1SAM|16|7|Та Господь сказав Самуїлові: Не дивись на обличчя його та на високість зросту його, бо Я відкинув його Собі! Бо Бог бачить не те, що бачить людина: чоловік бо дивиться на лице, а Господь дивиться на серце.
1SAM|16|8|І покликав Єссей Авінадава, і привів його перед Самуїла, та той сказав: Також цього не вибрав Господь!
1SAM|16|9|І привів Єссей Шамму, та Самуїл сказав: Також цього не вибрав Господь.
1SAM|16|10|І привів Єссей сімох своїх синів перед Самуїла. І сказав Самуїл до Єссея: Цих не вибрав Господь.
1SAM|16|11|І сказав Самуїл до Єссея: Чи то всі твої діти? А той відказав: Ще позостався найменший, він пасе отару. І сказав Самуїл до Єссея: Пошли ж привести його, бо не сядемо за стіл, аж поки він не прийде сюди.
1SAM|16|12|І послав він, і привів його, а він рум'яний, із гарними очима та хорошого стану. А Господь сказав Самуїлові: Устань, помаж його, бо це він!
1SAM|16|13|І взяв Самуїл рога оливи, та й помазав його серед братів його. І Дух Господній злинув на Давида, і був на ньому від того дня й далі. А Самуїл устав, і пішов до Рами.
1SAM|16|14|І Дух Господній відступився від Саула, а напав його дух злий, посланий від Господа.
1SAM|16|15|І сказали раби Саула до нього: Оце злий дух від Бога нападає на тебе.
1SAM|16|16|Нехай скаже пан наш, раби твої пошукають тобі кого, хто вміє грати на гуслах. І станеться, коли буде на тебе злий дух від Бога, то заграє той рукою своєю, і буде тобі добре.
1SAM|16|17|І сказав Саул до рабів своїх: Нагляньте мені кого, хто добре грає, і приведіть до мене.
1SAM|16|18|І відповів один із слуг, і сказав: Ось бачив я сина віфлеємлянина Єссея, що вміє грати, лицар та вояка, і розуміється на речах, і чоловік хорошої постави. І Господь із ним.
1SAM|16|19|І послав Саул послів до Єссея й сказав: Пошли до мене Давида, сина свого, що при отарі.
1SAM|16|20|І взяв Єссей осла, наладованого хлібом, та бурдюка вина, та одне козля, і послав через сина свого Давида до Саула.
1SAM|16|21|І прийшов Давид до Саула, та й став перед ним. І той сильно полюбив його, і він став йому зброєношею.
1SAM|16|22|І послав Саул до Єссея, говорячи: Нехай остається Давид при мені, бо він знайшов ласку в очах моїх.
1SAM|16|23|І бувало, коли злий дух від Бога нападав на Саула, то Давид брав гусла, та й грав своєю рукою. І легшало Саулові, і ставало йому добре, і відступав від нього той злий дух.
1SAM|17|1|І зібрали филистимляни свої війська на війну. І зібралися вони до Сохо, що Юдине, і таборували між Сохо та між Азекою в Ефес-Даммімі.
1SAM|17|2|І зібралися Саул та ізраїльтяни, і таборували в долині Елі, і вставилися до бою проти филистимлян.
1SAM|17|3|І стояли филистимляни на горі з того боку, а Ізраїль стояв на горі з цього боку, а поміж ними долина.
1SAM|17|4|І вийшов із филистимських таборів одноборець, ім'я йому Ґоліят із Ґату. Високий був шість ліктів і п'ядь.
1SAM|17|5|А на голові його мідяний шолом, і він одягнений був у панцера з луски; а вага того панцера п'ять тисяч шеклів міді.
1SAM|17|6|А на ногах його мідяні наголінники, а за плечима його мідяний спис.
1SAM|17|7|А держак списа його як ткацький вал, а вістря спису його шістсот шеклів заліза. А перед ним ходив щитоноша.
1SAM|17|8|І став він, і кликнув до Ізраїлевих полків, та й сказав до них: Чого ви вийшли ставати до бою? Чи ж я не филистимлянин, а ви не раби Саулові? Оберіть собі кого, і нехай він зійде до мене.
1SAM|17|9|Якщо він зможе воювати зо мною, і вб'є мене, то ми станемо вам за рабів. А якщо я переможу його, і вб'ю його, то ви станете нам за рабів, і будете служити нам.
1SAM|17|10|І сказав филистимлянин: Я цього дня зневажив Ізраїлеві полки. Дайте мені чоловіка, і будемо битися вдвох.
1SAM|17|11|І чув Саул та ввесь Ізраїль ці слова филистимлянина, і вони перестрашилися та сильно налякалися.
1SAM|17|12|А Давид син того мужа ефратянина, з Юдиного Віфлеєму, а ім'я йому Єссей, що мав восьмеро синів. І цей чоловік за Саулових днів був старий, увійшов у літа.
1SAM|17|13|І пішли троє найстарших Єссеєвих синів, пішли за Саулом на війну. А імена трьох синів його, що пішли на війну: перворідний Еліяв, а другий його Авінадав, а третій Шамма.
1SAM|17|14|А Давид він найменший, а три найстарші пішли за Саулом.
1SAM|17|15|А Давид ходив до Саула, та вертався пасти отару свого батька в Віфлеємі.
1SAM|17|16|А той филистимлянин підходив ранком та ввечорі, і виступав сорок день.
1SAM|17|17|І сказав Єссей до сина свого Давида: Візьми но для братів своїх ефу цього праженого зерна, і десять цих хлібів, та й віднеси скоренько до табору до своїх братів.
1SAM|17|18|А цих десять кусків сиру віднесеш для тисячника, і розізнаєш про поводження братів своїх, і вивідай про їхні потреби.
1SAM|17|19|А Саул і вони, та всі ізраїльтяни були в долині Елі, воювали з филистимлянами.
1SAM|17|20|І встав Давид рано вранці, і полишив отару свою на сторожа; і взяв та й пішов, як наказав йому Єссей. І ввійшов він до обозу, а військо виходило до бойового строю, і підняли вони окрик у бою.
1SAM|17|21|І вишикувалися Ізраїль та Филистимлянин лава проти лави.
1SAM|17|22|І Давид позоставив свою ношу в сторожа речей, та й побіг до полку. І ввійшов він, і запитав своїх братів про поводження.
1SAM|17|23|А коли він розмовляв із ними, аж ось виходить із филистимських полків одноборець, филистимлянин Ґоліят ім'я йому, із Ґату. І промовляв він ті самі слова, а Давид почув.
1SAM|17|24|А всі ізраїльтяни, коли бачили того чоловіка, то втікали перед ним та дуже лякалися.
1SAM|17|25|І говорив Ізраїльтянин: Чи бачите ви цього чоловіка, що виходить? А виходить він, щоб зневажати Ізраїля. І буде, того чоловіка, що вб'є його, збагатить його цар великим багатством, і дочку свою віддасть йому, а дім його батька зробить вільним в Ізраїлі.
1SAM|17|26|І спитався Давид тих людей, хто стояв з ним, говорячи: Що буде зроблене тому, хто вб'є цього филистимлянина й здійме образу з Ізраїля? Бо хто цей необрізаний филистимлянин, що так зневажає полки Живого Бога?
1SAM|17|27|А народ сказав йому те саме слово, говорячи: Отак буде зроблено чоловікові, хто вб'є його.
1SAM|17|28|І почув Еліяв, його найстарший брат, як він говорив до людей. І запалився Еліявів гнів на Давида, і він сказав: Чого то зійшов ти? І на кого ти позоставив трохи тієї отари в пустині? Я знаю зарозумілість твою та порожнечу твого серця, бо ти зійшов, щоб подивитися на війну!
1SAM|17|29|А Давид відказав: Та що я зробив тепер? Чи не на наказ батька?
1SAM|17|30|І він відвернувся від нього до іншого, і запитував про те саме. А народ відповів йому те саме, як перше.
1SAM|17|31|І були почуті слова ті, що говорив Давид, і донесли їх Саулові, і він покликав його.
1SAM|17|32|І сказав Давид до Саула: Хай не лякається нічиє серце через нього. Раб твій піде, і буде битися з отим филистимлянином.
1SAM|17|33|І сказав Саул до Давида: Ти не можеш піти на того филистимлянина битися з ним, бо ти малий, а він вояк від своєї молодости.
1SAM|17|34|І сказав Давид до Саула: Твій раб був пастухом свого батька при отарі, і приходив лев, а також ведмідь, та й тягнув штуку дрібної худоби зо стада,
1SAM|17|35|а я виходив за ним, і побивав його, і виривав те з пащі його. А як він ставав на мене, то я хапав його за його гриву, та й побивав його.
1SAM|17|36|І лева, і ведмедя побивав твій раб. І цей необрізаний филистимлянин буде, як один із них, бо він зневажив полки Живого Бога!
1SAM|17|37|І сказав Давид: Господь, що врятував мене з лапи лева та з лапи ведмедя, Він урятує мене з руки цього филистимлянина. І сказав Саул: Іди, і нехай Господь буде з тобою!
1SAM|17|38|І зодягнув Саул Давида в свою одіж, і дав мідяного шолома на його голову, і надів на нього панцера.
1SAM|17|39|І прип'яв Давид меча його на одежу свою, та й силкувався йти, бо він не звик був до того. І сказав Давид до Саула: Не можу в цьому ходити, бо я не звик! І поскидав Давид їх із себе.
1SAM|17|40|І взяв він кия свого в свою руку, і вибрав собі п'ять вигладжених камінців із потоку, і поклав їх у пастушу торбу, яку мав, та в торбину, а його праща у руці його. І він пішов до филистимлянина.
1SAM|17|41|А филистимлянин підходив усе ближче до Давида, і чоловік ніс щита перед ним.
1SAM|17|42|І подивився филистимлянин, та й побачив Давида, і злегковажив його, бо той був ще хлопець, рум'яний юнак стрункої постави.
1SAM|17|43|І сказав филистимлянин до Давида: Чи я пес, що ти вийшов на мене з києм? І филистимлянин прокляв Давида своїми богами.
1SAM|17|44|І сказав филистимлянин до Давида: Ходи ж до мене, а я твоє тіло віддам птаству небесному та звірині польовій.
1SAM|17|45|І сказав Давид до филистимлянина: Ти йдеш на мене з мечем і списом та ратищем, а я йду на тебе в Ім'я Господа Саваота, Бога військ Ізраїлевих, які ти зневажив.
1SAM|17|46|Сьогодні віддасть тебе Господь у мою руку, і я поб'ю тебе, і відітну голову твою з тебе, і дня цього я дам падло филистимського табору птаству небесному та земній звірині. І пізнає вся земля, що є Бог Ізраїлів!
1SAM|17|47|І пізнає вся громада те, що Господь спасає не мечем та списом, бо це війна Господа, і Він віддасть вас у нашу руку.
1SAM|17|48|І сталося, коли филистимлянин устав і пішов, і зблизився до Давида, то Давид поспішив і побіг до лави навпроти филистимлянина.
1SAM|17|49|І простяг Давид руку свою до торби, і взяв звідти каменя, та й кинув із пращі, і вдарив филистимлянина в чоло його. І той камінь втявся йому в чоло, і він упав на обличчя своє на землю.
1SAM|17|50|І отак переміг Давид филистимлянина пращею та каменем, і вдарив він филистимлянина, та й убив його, а меча не було в Давидовій руці.
1SAM|17|51|І підбіг Давид, і став на филистимлянина, і вихопив його меча, і витяг його з його піхви, та й убив його, відтяв ним йому голову! І побачили филистимляни, що помер їх силач, і стали втікати!
1SAM|17|52|А люди Ізраїлеві та Юдині схопилися, і зняли крик, та й погнали филистимлян аж доти, де йдеться до Ґаю, і аж до брами Екрону. І падали трупи филистимлян по дорозі аж до Шаараїму, і аж до Ґату, і аж до Екрону.
1SAM|17|53|І вернулися Ізраїлеві сини з погоні за филистимлянами, та й розграбували їхні табори.
1SAM|17|54|А Давид узяв голову того филистимлянина, і приніс її до Єрусалиму, а зброю його склав у своєму наметі.
1SAM|17|55|А як Саул побачив Давида, що виходив навпроти филистимлянина, то сказав до Авнера, провідника війська: Чий син оцей хлопець, Авнере? А Авнер відказав: Присягаю життям твоїм, о царю, що не знаю!
1SAM|17|56|І сказав цар: Запитай, чий син цей юнак?
1SAM|17|57|А коли Давид вертався, побивши филистимлянина, то Авнер узяв його й привів його перед Саула, а голова филистимлянина у руці його.
1SAM|17|58|І сказав до нього Саул: Чий ти син, хлопче? А Давид відказав: Я син раба твого віфлеємлянина Єссея.
1SAM|18|1|І сталося, як скінчив він говорити до Саула, то Йонатанова душа зв'язалася з душею Давидовою, і полюбив його Йонатан, як душу свою.
1SAM|18|2|І того дня взяв його Саул, і не пустив його вернутися до дому його батька.
1SAM|18|3|І склав Йонатан із Давидом умову, бо полюбив його, як душу свою.
1SAM|18|4|І зняв Йонатан із себе плаща, що був на ньому, та й дав його Давидові, і вбрання своє, і все аж до меча свого, і аж до лука свого, і аж до пояса свого.
1SAM|18|5|І ходив Давид скрізь, куди посилав його Саул, і робив мудро. І настановив його Саул над вояками, і він подобався усьому народові, а також Сауловим рабам.
1SAM|18|6|І сталося, як вони йшли, коли Давид вертався, побивши филистимлянина, то повиходили жінки зо всіх Ізраїлевих міст, щоб співати та танцювати назустріч царя Саула, із бубнами, із радістю, та з цимбалами.
1SAM|18|7|І викрикували ті жінки, що грали, та й казали: Саул повбивав свої тисячі, а Давид десятки тисяч свої!
1SAM|18|8|І дуже запалився Саулів гнів, і та річ була неприємна йому, і він сказав: Давидові дали десятки тисяч, а мені дали тисячі, йому бракує ще тільки царювання!
1SAM|18|9|І від того дня й далі Саул дивився заздрісним оком на Давида.
1SAM|18|10|І сталося другого дня, і напав злий дух від Бога на Саула, і він став несамовитий в себе вдома, а Давид грав своєю рукою, як щоденно, а в Сауловій руці був спис.
1SAM|18|11|І кинув Саул списа, кажучи про себе: Ударю в Давида, і приб'ю його до стіни! Та Давид два рази ухилився від нього.
1SAM|18|12|І боявся Саул Давида, бо з ним був Господь, а від Саула Він відступив.
1SAM|18|13|І віддалив його Саул від себе, і настановив його собі тисячником, і він виходив на війни, і вертався перед народом.
1SAM|18|14|І мав Давид поводження в усіх дорогах своїх, і з ним був Господь.
1SAM|18|15|І побачив Саул, що той має велике поводження, і налякався його.
1SAM|18|16|А ввесь Ізраїль та Юда любили Давида, бо він виходив на війни, і вертався перед ними.
1SAM|18|17|І сказав Саул до Давида: Ось моя найстарша дочка Мерав, її я дам тобі за жінку. Тільки будь мені хоробрим та воюй Господні війни! А про себе Саул сказав: Нехай не буде на ньому моя рука, а нехай буде на ньому рука филистимлян!
1SAM|18|18|А Давид сказав до Саула: Хто я, і яке життя моє та рід мого батька в Ізраїлі, що я стану зятем цареві?
1SAM|18|19|І сталося, коли настав час дати Давидові Мерав, Саулову дочку, то вона була видана за жінку мехолатитянинові Адріїлові,
1SAM|18|20|а Давида покохала Мелхола, друга Саулова дочка. І розповіли про це Саулові, і ця річ була слушна в очах його.
1SAM|18|21|І сказав Саул про себе: Дам я її йому, і нехай вона стане йому за пастку, і нехай буде на ньому рука филистимлян! А до Давида Саул сказав удруге: Посвоячишся сьогодні зо мною.
1SAM|18|22|І наказав Саул своїм рабам: Промовляйте до Давида потиху, говорячи: Ось цар уподобав тебе собі, а всі його раби полюбили тебе, а тепер ти посвоячишся з царем.
1SAM|18|23|І Саулові раби говорили ці слова до Давидових ушей. А Давид сказав: Чи то легко в ваших очах посвоячитися з царем? Таж я людина вбога та маловажна!
1SAM|18|24|І розповіли це раби Саула йому, говорячи: Отак говорив Давид.
1SAM|18|25|І сказав Саул: Так скажете Давидові: Не бажає цар заплати за молоду, а бажає тільки сто крайніх плотів филистимських, щоб пімститися на неприятелях царя. А Саул думав тим зробити, щоб Давид попав до руки филистимлян.
1SAM|18|26|І його раби переказали ці слова Давидові, і ця річ була мила в Давидових очах, щоб посвоячитися з царем. І в недовгому часі
1SAM|18|27|встав Давид, та й пішов він та його люди, і забив серед филистимлян двісті чоловіка. І Давид приніс їхні крайні плоті, і дав їх у повному числі цареві, щоб посвоячитися з царем. І Саул дав йому за жінку дочку свою Мелхолу.
1SAM|18|28|І побачив Саул, і пізнав, що Господь із Давидом, а Мелхола, Саулова дочка, полюбила його.
1SAM|18|29|А Саул ще й далі боявся Давида. І Саул ненавидів Давида по всі дні.
1SAM|18|30|І виходили воювати филистимські провідники, і бувало скільки вони виходили, то Давид мав найбільше поводження від усіх Саулових рабів. І стало ім'я його дуже шановане.
1SAM|19|1|І говорив Саул до свого сина Йонатана та до всіх своїх рабів, щоб убити Давида. Та Йонатан, син Саулів, дуже кохав Давида.
1SAM|19|2|І розповів Йонатан Давидові, говорячи: Батько мій Саул хоче вбити тебе. А тепер уранці стережися, сиди в укритті, і сховайся.
1SAM|19|3|А я вийду, і стану при своєму батькові на полі, де ти будеш, і я буду говорити про тебе до свого батька. І що побачу, те розповім тобі.
1SAM|19|4|І говорив Йонатан своєму батькові Саулові добре про Давида, і сказав йому: Нехай не згрішить цар проти раба свого, проти Давида, бо не згрішив він проти тебе, а вчинки його дуже добрі для тебе.
1SAM|19|5|І наражав він на небезпеку життя своє, і вбив филистимлянина, і Господь учинив велике спасіння для всього Ізраїля. Ти це бачив та радів. І для чого згрішиш ти проти невинної крови, бажаючи вбити Давида безпричинно?
1SAM|19|6|І послухався Саул Йонатанового голосу. І Саул присягнув: Як живий Господь, не буде той убитий!
1SAM|19|7|І покликав Йонатан Давида, і переказав йому Йонатан усі ті слова. І привів Йонатан Давида до Саула, і він був перед ним, як давніше.
1SAM|19|8|А війна була далі. І вийшов Давид, воював з филистимлянами, та й завдав їм велику поразку, і вони повтікали перед ним.
1SAM|19|9|А злий дух від Господа був на Саулі, і він сидів у своїм домі, і спис його в руці його, а Давид грав рукою.
1SAM|19|10|А Саул хотів ударити списом у Давида, прибити його до стіни, та відхилився той перед Саулом, і він увігнав списа в стіну, а Давид утік, і був урятований тієї ночі.
1SAM|19|11|І послав Саул посланців до Давидового дому, щоб стерегли його й щоб убили його вранці. І розповіла Давидові його жінка Мелхола, говорячи: Якщо ти не врятуєш свого життя цієї ночі, то взавтра ти будеш забитий.
1SAM|19|12|І Мелхола спустила Давида через вікно, і він пішов і втік, і врятувався.
1SAM|19|13|І взяла Мелхола домашнього божка, і поклала до ліжка, а подушку з козячого волосу поклала в головах його, та й прикрила плащем.
1SAM|19|14|І послав Саул посланців, щоб узяти Давида, а вона сказала: Він хворий!
1SAM|19|15|І послав Саул тих посланців побачити Давида, говорячи: Принесіть його в ліжку до мене, щоб забити його!
1SAM|19|16|І ввійшли ті посланці, аж ось у ліжку домашній божок, а в головах його подушка з козячого волосу!
1SAM|19|17|І сказав Саул до Мелхоли: Нащо ти так обманила мене, і відпустила мого ворога, і він урятувався? А Мелхола відказала Саулові: Він сказав мені: Відпусти мене, бо інакше вб'ю тебе!
1SAM|19|18|А Давид утік і врятувався. І прийшов він до Самуїла до Рами, і розповів йому все, що зробив йому Саул. І пішов він та Самуїл, та й осілися в Найоті.
1SAM|19|19|І розповіджено Саулові, говорячи: Ось Давид у Найоті в Рамі.
1SAM|19|20|І послав Саул посланців, щоб узяли Давида. І вони побачили громаду пророків, що пророкувала, а Самуїл стояв над ними. І на Саулових посланців злинув Дух Божий, і пророкували й вони.
1SAM|19|21|І розповіли про це Саулові. І послав він інших посланців, та пророкували також і вони. А Саул послав посланців ще третіх, та пророкували й вони.
1SAM|19|22|І пішов і він до Рами, і прийшов аж до великої ями, що в Сеху, і запитав, і сказав: Де Самуїл та Давид? А запитаний відказав: Ось у Найоті в Рамі.
1SAM|19|23|І пішов він туди до Найоту в Рамі. І злинув Божий Дух також на нього, і він усе пророкував, аж поки не прийшов у Найот у Рамі.
1SAM|19|24|І зняв і він одежу свою, і пророкував і він перед Самуїлом, і лежав нагий цілий той день та цілу ніч. Тому то й говорять: Чи й Саул між пророками?
1SAM|20|1|І втік Давид з Найоту в Рамі, і прийшов та й сказав перед Йонатаном: Що я зробив, яка провина моя й який мій гріх перед батьком твоїм, що він шукає моєї душі?
1SAM|20|2|А той відказав: Борони Боже, ти не помреш! Таж батько мій не робить жодної справи, великої чи справи малої, коли не відкриває на вухо мені, то чому мій батько заховає від мене цю справу? Цього не буде!
1SAM|20|3|А Давид іще присягнув та й сказав: Добре пізнав твій батько, що я знайшов милість в очах твоїх. І сказав він: Нехай не довідається про те Йонатан, щоб не був він засмучений. Але як живий Господь і як жива душа твоя, між мною та смертю не більше кроку!
1SAM|20|4|І сказав Йонатан до Давида: Що підкаже душа твоя, те зроблю тобі!
1SAM|20|5|І сказав Давид до Йонатана: Ось узавтра новомісяччя, коли звичайно сиджу я з царем, щоб їсти з ним. Але ти відпусти мене, а я сховаюся в полі аж до третього вечора.
1SAM|20|6|Якщо дійсно згадає про мене твій батько, то скажеш, що конче жадав від мене Давид, щоб йому забігти до свого міста Віфлеєму, бо там річна жертва для всього роду його.
1SAM|20|7|Якщо він скаже так: Добре! то мир твоєму рабові. А якщо дійсно запалає йому гнів, то знай, що постановлене те зло від нього.
1SAM|20|8|І зробиш милість своєму рабові, бо ти ввів свого раба в Господній заповіт із собою. А якщо є на мені провина, убий мене ти, а до батька твого пощо мене вести?
1SAM|20|9|І відказав Йонатан: Борони тебе, Боже! Бо якщо справді пізнаю, що в мого батька постановлене зло, щоб прийшло на тебе, чи ж того я не розкажу тобі?
1SAM|20|10|І сказав Давид до Йонатана: Хто повідомить мене, якщо батько твій відповість тобі жорстоке?
1SAM|20|11|А Йонатан сказав до Давида: Ходи ж, і вийдемо на поле. І вийшли вони обидва на поле.
1SAM|20|12|І сказав Йонатан до Давида: Свідок Господь, Бог Ізраїлів, що післязавтра цього часу вивідаю я батька свого. Нехай скарає мене Бог, якщо тоді не пошлю до тебе, і не сповіщу тебе,
1SAM|20|13|так нехай зробить Господь Йонатану, і так нехай додасть! А якщо моєму батькові вгодно зробити зло тобі, то сповіщу тебе, і відішлю тебе, і ти підеш у мирі, а Господь буде з тобою, як Він був із моїм батьком.
1SAM|20|14|І ти, якщо я буду ще живий, хіба не зробиш зо мною Господньої милости? Коли ж я помру,
1SAM|20|15|то не відбирай своєї милости від дому мого навіки, а навіть тоді, як Господь понищить усіх Давидових ворогів із поверхні землі.
1SAM|20|16|І нехай пошукає Господь душі від Давидових ворогів! І склав Йонатан умову з Давидовим домом.
1SAM|20|17|І Йонатан далі присягався Давидові в своїй любові до нього, бо він покохав його, як свою душу.
1SAM|20|18|І сказав йому Йонатан: Узавтра новомісяччя, і ти будеш згаданий, бо буде порожнє твоє місце.
1SAM|20|19|А третього дня скоро зійдеш, і прийдеш до місця, де ти ховався у день твого чину, і сядеш при камені Азел.
1SAM|20|20|А я пущу три стрілі набік, ніби стріляючи собі до мети.
1SAM|20|21|І ось пошлю я слугу: Іди, знайди ті стріли! Якщо, говорячи, скажу я до хлопця: Он ті стріли тут перед тобою, візьми їх, то приходь, бо мир тобі, і нема нічого злого, як живий Господь!
1SAM|20|22|А якщо я скажу до того юнака так: Он ті стріли з а тобою далі, то втікай, бо Господь відпускає тебе.
1SAM|20|23|А та річ, що про неї говорили ми, я та ти, ось Господь буде свідком між мною та між тобою аж навіки!
1SAM|20|24|І сховався Давид у полі. І було новомісяччя, а цар засів до їжі.
1SAM|20|25|І сів цар на стільці своїм, як раз-у-раз, на стільці при стіні. І встав Йонатан, а Авнер сів збоку Саула, а Давидове місце було порожнє.
1SAM|20|26|Та Саул нічого не говорив того дня, бо сказав собі: Це випадок, Давид не чистий, бо не очистився.
1SAM|20|27|І сталося другого дня, на другий день новомісяччя, було порожнє Давидове місце. І сказав Саул до сина свого Йонатана: Чому не прийшов на хліб Єссеїв син і вчора, і сьогодні?
1SAM|20|28|І відповів Йонатан Саулові: Дійсно просився Давид у мене до Віфлеєму.
1SAM|20|29|І він говорив: Пусти мене, бо в тому місті для нас родова жертва, і запросив мене брат мій. А тепер, якщо знайшов я милість в очах твоїх, нехай я побіжу та побачу братів моїх. Тому не прийшов він до царського столу.
1SAM|20|30|І запалав Саулів гнів на Йонатана, і він сказав йому: Негідний і неслухняний сину! Чи ж не знаю я, що ти вибрав Єссеєвого сина на свій сором та на сором і неславу своєї матері?
1SAM|20|31|Бо всі дні, поки Єссеїв син живий на землі, не будеш міцно стояти ані ти, ані царство твоє. А тепер пошли, і приведи його до мене, бо він призначений на смерть.
1SAM|20|32|І відповів Йонатан своєму батькові Саулові та й сказав йому: Чому він буде забитий? Що він зробив?
1SAM|20|33|Тоді Саул кинув списа на нього, щоб убити його. І пізнав Йонатан, що то постановлене від батька, щоб убити Давида.
1SAM|20|34|І встав Йонатан від столу, розпалений гнівом, і не їв хліба і другого дня новомісяччя, бо був засмучений за Давида, бо його образив його батько.
1SAM|20|35|І сталося вранці, і вийшов Йонатан на поле, на умовлений з Давидом час, а з ним був малий хлопець.
1SAM|20|36|І сказав він до хлопця свого: Побіжи, знайди ті стріли, що я вистріляю. Хлопець побіг, а він пустив стрілу поза нього.
1SAM|20|37|І прийшов хлопець до місця стріли, що пустив Йонатан, а Йонатан кликнув за хлопцем і сказав: Он та стріла за тобою далі!
1SAM|20|38|І кликнув Йонатан за хлопцем: Скоро, поспіши, не ставай! І зібрав Йонатанів хлопець стріли, та й прийшов до свого пана.
1SAM|20|39|А той хлопець нічого не знав, тільки Йонатан та Давид знали ту справу.
1SAM|20|40|І віддав Йонатан свою зброю юнакові, якого мав, та й сказав йому: Іди, занеси це до міста!
1SAM|20|41|Той юнак пішов, а Давид устав із південного боку, і впав на обличчя своє на землю, та й поклонився три рази. І поцілували вони один одного, і оплакували один одного, а Давид гірко плакав.
1SAM|20|42|І сказав Йонатан до Давида: Іди з миром! А що присягнули ми двоє в Господнє Ім'я, говорячи: Господь нехай буде свідком між мною та між тобою, і між насінням моїм та насінням твоїм, нехай буде аж навіки! (21-1) І встав Давид і пішов, а Йонатан пішов до міста.
1SAM|21|1|(21-2) І прийшов Давид до Нова, до священика Ахімелеха. А Ахімелех із тремтінням стрів Давида й сказав йому: Чому ти сам, і нікого немає з тобою?
1SAM|21|2|(21-3) І сказав Давид до священика Ахімелеха: Цар наказав мені справу, і до мене сказав: Нехай ніхто не знає цього, тієї справи, за якою я посилаю тебе, і яку наказав тобі. А слуг я умовив на означене місце.
1SAM|21|3|(21-4) А тепер, що є в тебе під рукою? П'ять хлібів дай у мою руку, або що знайдеться.
1SAM|21|4|(21-5) А священик відповів Давидові та й сказав: Нема в мене звичайного хліба під рукою, а є тільки хліб святий, якщо твої слуги здержалися від жінки.
1SAM|21|5|(21-6) І відповів Давид священикові, та й сказав йому: Так, бо жінок не було при нас як учора, так і позавчора, відколи я вийшов, і тіла слуг були чисті. А то хліб звичайний, особливо коли сьогодні замість цього інший хліб у посудині стане святим.
1SAM|21|6|(21-7) І дав йому священик святе, бо не було там іншого хліба, крім хлібів показних, що були зняті з-перед Господнього лиця, щоб покласти теплий хліб того дня, коли його забирають.
1SAM|21|7|(21-8) А там того дня знаходився один із Саулових рабів перед Господнім лицем, а ім'я йому Доеґ, ідумеянин, провідник пастухів, яких мав Саул.
1SAM|21|8|(21-9) І сказав Давид до Ахімелеха: Чи нема тут у тебе під рукою списа або меча? Бо я не взяв до своєї руки ані меча свого, ані іншої зброї своєї, бо царська справа була нагла.
1SAM|21|9|(21-10) А священик сказав: Є меч филистимлянина Ґоліята, що ти вбив його в долині Ела, ось він за ефодом, загорнений одежею. Якщо візьмеш його собі, візьми, бо тут нема іншого, окрім нього. І сказав Давид: Нема іншого такого, як він, дай його мені!
1SAM|21|10|(21-11) І встав Давид, і втікав того дня перед Саулом, і прибув до Ахіша, царя ґатського.
1SAM|21|11|(21-12) І сказали до нього Ахішеві раби: Чи ж не цей Давид цар Краю? Хіба ж не про нього співають у танцях, говорячи: Саул повбивав свої тисячі, а Давид десятки тисяч свої.
1SAM|21|12|(21-13) І заховав Давид ті слова в своєму серці, і сильно боявся Ахіша, царя ґатського.
1SAM|21|13|(21-14) І змінив він свій розум на їхніх очах, і шалів при них, і бив по дверях брами, і пускав слину свою на свою бороду.
1SAM|21|14|(21-15) І сказав Ахіш до своїх рабів: Ось бачите чоловіка, що сходить із розуму. Нащо привели його до мене?
1SAM|21|15|(21-16) Чи мені бракує безумних, що ви привели його, щоб сходив із розуму передо мною? Чи такий може входити до мого дому?
1SAM|22|1|І пішов Давид звідти, і втік до печери Адуллам. А брати його та ввесь дім батька його почули про це, та й посходилися до нього туди.
1SAM|22|2|І позбиралися до нього кожен пригноблений, і кожен, хто був задовжений, і кожен огірчений в душі, і він став над ними провідником. І було їх із ним близько чотирьох сотень люда.
1SAM|22|3|І пішов Давид ізвідти до Моавської Міцпи, та й сказав до моавського царя: Нехай прийде батько мій та мати моя, і будуть із вами, аж поки я буду знати, що зробить мені Бог.
1SAM|22|4|І він привів їх до моавського царя, і вони осілися з ним на всі дні Давидового перебування в твердині.
1SAM|22|5|А пророк Ґад сказав до Давида: Ти не будеш сидіти в твердині, іди, і перейдеш собі до Юдиного краю! І пішов Давид, і прийшов до лісу Херет.
1SAM|22|6|І почув Саул, що пізнаний Давид та люди, хто з ним. А Саул сидів у Ґів'ї під тамариском на узгір'ї, а спис його був у руці його, і всі його раби стояли при ньому.
1SAM|22|7|І сказав Саул до слуг своїх, що стояли при ньому: Послухайте, веніяминівці! Чи вже ж Єссеїв син дасть усім вам поля та виноградники? Чи вже ж настановить усіх вас тисячниками та сотниками,
1SAM|22|8|що всі ви змовилися на мене, і не донесли до вуха мого, що син мій склав умову з Єссеєвим сином, і ніхто з вас не змилосердився надо мною, і не відкрив мені, що син мій поставив мого раба чатувати на мене, і те діється і цього дня?
1SAM|22|9|І відповів ідумеянин Доеґ, а він стояв при Саулових слугах, і сказав: Я бачив Єссеєвого сина, що приходив до Нова, до Ахімелеха, Ахітувового сина,
1SAM|22|10|і він питав для нього Господа, і дав йому поживи на дорогу, і дав йому меча филистимлянина Ґоліята.
1SAM|22|11|І послав цар покликати священика Ахімелеха, сина Ахітувового, та ввесь дім його батька, священиків, що в Нові. І всі вони прибули до царя.
1SAM|22|12|А Саул сказав: Слухай но, сину Ахітувів! А той відказав: Ось я, мій пане!
1SAM|22|13|І сказав до нього Саул: Нащо ви змовилися на мене, ти та Єссеїв син, коли ти дав йому хліба та меча, і питав для нього Бога, щоб повстав він на мене й чигав, як цього дня?
1SAM|22|14|І відповів Ахімелех цареві та й сказав: А хто серед усіх рабів твоїх вірний, як Давид, царів зять, і має приступ до тайної ради, і шанований у твоєму домі?
1SAM|22|15|Хіба сьогодні зачав я питати для нього Бога? Борони мене Боже! Нехай цар не кладе закиду на раба свого та на ввесь дім батька мого, бо в усьому тому твій раб не знає нічого, ані малого, ані великого.
1SAM|22|16|А цар сказав: Конче помреш, Ахімелеху, ти та ввесь дім батька твого!
1SAM|22|17|І сказав цар слугам, що стояли при ньому: Підійдіть, і повбивайте Господніх священиків, бо й їхня рука разом із Давидом, бо вони знали, що втікає він, та не донесли до вуха мого. Та не хотіли цареві раби простягнути своєї руки, щоб діткнутися до Господніх священиків.
1SAM|22|18|Тоді цар сказав до Доеґа: Підійди ти, і вдар священиків! І підійшов ідумеянин Доеґ, та й ударив священиків, і вбив того дня вісімдесят і п'ять чоловіка, що носять лляного ефода.
1SAM|22|19|А Нов, священиче місто, цар побив вістрям меча все, від чоловіка й аж до жінки, від дитини й аж до немовляти, і вола, і осла, і дрібну худобину, усе побив вістрям меча.
1SAM|22|20|Та втік один син Ахімелеха, Ахітувового сина, а ім'я йому: Евіятар. І втік він до Давида.
1SAM|22|21|І Евіятар доніс Давидові, що Саул повбивав Господніх священиків.
1SAM|22|22|А Давид сказав до Евіятара: Я знав того дня, що там ідумеянин Доеґ, який конче розповість Саулові. Я став причиною загибелі всіх душ дому твого батька!
1SAM|22|23|Зостанься ж зо мною, не бійся, бо той, хто шукатиме моєї душі, шукатиме й душі твоєї, та ти будеш стережений у мене.
1SAM|23|1|І донесли Давидові, говорячи: Ось филистимляни облягли Кеїлу, і грабують клуні.
1SAM|23|2|І запитав Давид Господа, говорячи: Чи піду й переможу тих филистимлян? А Господь сказав до Давида: Іди, і поб'єш филистимлян та спасеш Кеїлу.
1SAM|23|3|А Давидові люди сказали до нього: Ось ми боїмося тут у Юді, а що ж буде, коли підемо в Кеїлу, проти филистимських лав?
1SAM|23|4|А Давид ще далі питався Господа, і Господь відповів та сказав йому: Устань, зійди до Кеїли, бо Я даю филистимлян у твою руку.
1SAM|23|5|І пішов Давид та люди його до Кеїли, та й воював із филистимлянами, і зайняв їхню худобу, і наніс їм велику поразку. І спас Давид мешканців Кеїли.
1SAM|23|6|І сталося, коли втікав Евіятар, син Ахімелеха, до Давида в Кеїлу, то ефод був у його руці.
1SAM|23|7|А Саулові донесено, що Давид увійшов у Кеїлу. І сказав Саул: Бог віддав його в мою руку, бо він замкнув себе, коли ввійшов до міста з воротами та засувом.
1SAM|23|8|І скликав Саул увесь народ на війну, щоб зійти до Кеїли облягти Давида та людей його.
1SAM|23|9|І дізнався Давид, що Саул задумує лихо на нього, і сказав до священика Евіятара: Принеси ефода!
1SAM|23|10|І Давид сказав: Господи, Боже Ізраїлів! Дослухуючися, чув Твій раб, що Саул хоче ввійти до Кеїли, щоб вигубити місто через мене.
1SAM|23|11|Чи видадуть мене громадяни Кеїли в його руку? Чи зійде Саул, як чув твій раб? Господи, Боже Ізраїлів, розповіж же Своєму рабові! І сказав Господь: Зійде.
1SAM|23|12|І запитався Давид: Чи видадуть громадяни Кеїли мене та людей моїх у Саулову руку? А Господь сказав: Видадуть.
1SAM|23|13|І встав Давид та його люди, близько шости сотень чоловіка, та й вийшли з Кеїли, і ходили, де можна було ходити. А Саулові донесено, що Давид утік із Кеїли, і він занехаяв похід.
1SAM|23|14|І осівся Давид у пустині в твердинях, і осівся на горі в пустині Зіф. А Саул шукав його повсякденно, та Бог не дав його в руку йому.
1SAM|23|15|І побачив Давид, що Саул вийшов шукати душі його, а Давид пробував у пустині Зіф у Хореші.
1SAM|23|16|І встав Йонатан, Саулів син, і пішов до Давида до Хорешу, і зміцнив його на дусі в Бозі,
1SAM|23|17|та й сказав до нього: Не бійся, бо не знайде тебе рука мого батька Саула! І ти будеш царювати над Ізраїлем, а я буду тобі заступником. І це знає й батько мій Саул.
1SAM|23|18|І вони обидва склали умову перед Господнім лицем. І осівся Давид у Хорешу, а Йонатан пішов до свого дому.
1SAM|23|19|А зіфеяни прийшли до Саула до Ґів'ї, говорячи: Ось Давид ховається в нас у твердинях у Хорешу, на взгір'ї Хахіла, що з півдня від Єшімону.
1SAM|23|20|А тепер, за всім жаданням своєї душі, о царю, конче зійди, а нам хіба видати його в цареву руку.
1SAM|23|21|І сказав Саул: Благословенні ви в Господа, бо змилосердилися надо мною!
1SAM|23|22|Ідіть же, приготуйте ще, і розпізнайте, і побачте місце його, де буде нога його, хто його там бачив, бо казали мені: сильно хитрує він!
1SAM|23|23|І подивіться, і розізнайте всі схованки, де він ховається, і вернетесь до мене з певною звісткою, і я піду з вами. І буде, якщо він є в Краю, то пошукаю його по всіх Юдиних тисячах.
1SAM|23|24|І встали вони, і пішли в Зіф перед Саулом. А Давид та його люди були в Маонській пустині в Араві, на південь від Єшімону.
1SAM|23|25|А Саул та його люди пішли шукати. І донесли про це Давидові, і він зійшов до Сели, і спинився в Маонській пустині. А Саул прочув, та й гнався за Давидом до Маонської пустині.
1SAM|23|26|І пішов Саул з цього боку гори, а Давид та його люди з того боку гори. І поспішав Давид відійти перед Саулом, а Саул та люди його оточували Давида та людей його, щоб схопити їх.
1SAM|23|27|І прийшов посланець до Саула, говорячи: Іди поспішно, бо филистимляни кинулися на Край!
1SAM|23|28|І вернувся Саул з погоні за Давидом, і пішов навперейми филистимлян. Тому то назвали ім'я тому місцю: Села-Гаммахлекот.
1SAM|23|29|(24-1) А Давид вийшов звідти, і осівся в твердинях Ен-Ґеді.
1SAM|24|1|(24-2) І сталося, як вернувся Саул із погоні за филистимлянами, то донесли йому, говорячи: Ось Давид у пустині Ен-Ґеді.
1SAM|24|2|(24-3) І взяв Саул три тисячі війська, вибраних з усього Ізраїля, і пішов шукати Давида та людей його на поверхні газельських скель.
1SAM|24|3|(24-4) І прийшов він до кошар на отари при дорозі, а там печера. І Саул увійшов туди для потреби, а по боках печери сиділи Давид та люди його.
1SAM|24|4|(24-5) І сказали люди Давида до нього: Оце той день, що Господь говорив до тебе: Ось Я даю ворога твого в твою руку, і ти зробиш йому, як буде добре в твоїх очах. А Давид устав, і тихо відтяв полу Саулового плаща.
1SAM|24|5|(24-6) І сталося потім, і серце Давидове все докоряло йому, що він відтяв полу Саулового плаща.
1SAM|24|6|(24-7) І сказав він до своїх людей: Борони мене, Господи, щоб зробити ту річ моєму панові, Господньому помазанцеві, щоб простягнути руку свою на нього, бо він помазанець Господній!
1SAM|24|7|(24-8) І Давид стримав цими словами людей своїх, і не дав їм повстати на Саула. А Саул устав із печери, і пішов дорогою.
1SAM|24|8|(24-9) А потому Давид устав, і вийшов із печери, та й закричав за Саулом, говорячи: Пане мій, о царю! А Саул озирнувся назад, а Давид схилився обличчям до землі та й поклонився.
1SAM|24|9|(24-10) І сказав Давид до Саула: Нащо ти слухаєш слів того, хто каже: Давид хоче тобі зла?
1SAM|24|10|(24-11) Ось цього дня очі твої бачать те, що Господь дав був тебе сьогодні в мою руку в печері. І радили мені забити тебе, та я змилосердився над тобою й сказав: Не простягну своєї руки на свого пана, бо він помазанець Господній!
1SAM|24|11|(24-12) І подивися, батьку мій, і поглянь на полу плаща свого в моїй руці, бо коли я відрізував цю полу плаща твого, то я не забив тебе. Пізнай та побач, що в моїй руці нема зла та гріха, і не згрішив я проти тебе, а ти чигаєш на душу мою, щоб забрати її!
1SAM|24|12|(24-13) Нехай розсудить Господь між мною та між тобою, і нехай пімститься Господь тобі за мене, а моя рука не буде на тобі!
1SAM|24|13|(24-14) Як говорить стародавня приказка: Від безбожних виходить безбожність, а моя рука не буде на тобі!
1SAM|24|14|(24-15) За ким вийшов Ізраїлів цар? За ким ти ганяєшся? За мертвим псом, за однією блохою?
1SAM|24|15|(24-16) І нехай буде Господь за суддю, і нехай Він розсудить між мною та між тобою. І побачить Він, і заступиться за мою справу, і висудить мене з твоєї руки.
1SAM|24|16|(24-17) І сталося, як Давид скінчив говорити ці слова до Саула, то Саул сказав: Чи це твій голос, сину мій Давиде? І підняв Саул голос свій, та й заплакав.
1SAM|24|17|(24-18) І сказав він до Давида: Справедливіший ти від мене, бо ти робив мені добро, а я робив тобі лихо.
1SAM|24|18|(24-19) Бо ти сьогодні засвідчив, що зробив зо мною добро тим, що Господь видав мене в твою руку, а ти не вбив.
1SAM|24|19|(24-20) Як чоловік знайде свого ворога, то хіба відпускає його доброю дорогою? І Господь відплатить тобі добром за те, що ти зробив мені цього дня.
1SAM|24|20|(24-21) А тепер я ось пізнав, що дійсно будеш ти царювати, і стане в руці твоїй Ізраїлеве царство.
1SAM|24|21|(24-22) А тепер присягни мені Господом, що не вигубиш насіння мого по мені, і що не вигубиш імени мого з дому батька мого.
1SAM|24|22|(24-23) І Давид заприсягнув Саулові. І пішов Саул до дому свого, а Давид та люди його ввійшли до твердині.
1SAM|25|1|І вмер Самуїл, і зібрався ввесь Ізраїль, та й оплакував його, і поховали його в його домі в Рамі. А Давид устав, і пішов у пустиню Паран.
1SAM|25|2|І був чоловік у Маоні, а оселя його на Кармелі, і цей чоловік був дуже багатий, і мав три тисячі дрібної худоби та тисячу кіз. І був він на Кармелі, коли стригли отару його.
1SAM|25|3|А ім'я тому чоловікові Навал, а ім'я жінці його Авіґаїл. А жінка та була доброго розуму та вродлива, чоловік же той був жорстокий та злочинний, із роду Калева.
1SAM|25|4|А Давид почув у пустині, що Навал стриже свою отару.
1SAM|25|5|І послав Давид десять хлопців. І сказав Давид до тих хлопців: Вийдіть на Кармел, і прийдете до Навала й запитаєте його в моєму йменні про мир,
1SAM|25|6|та й скажете так братові моєму: І тобі мир, і дому твоєму мир, і всьому, що твоє, мир!
1SAM|25|7|А тепер почув я, що в тебе стрижуть. Пастухи твої були з нами, ми не кривдили їх, і нічого не пропало їм по всі дні перебування їх на Кармелі.
1SAM|25|8|Запитай своїх слуг, і вони розповідять тобі. І нехай знайдуть в очах твоїх милість мої хлопці, бо доброго дня ми прийшли. Дай же рабам своїм та синові своєму Давидові, що знайде рука твоя!
1SAM|25|9|І прийшли Давидові хлопці, і промовили до Навала, в імені Давида, усі ці слова. І спинилися.
1SAM|25|10|І відповів Навал Давидовим рабам, і сказав: Хто такий Давид та хто Єссеїв син? Сьогодні намножилося рабів, що вириваються кожен від пана свого!
1SAM|25|11|І я візьму хліб свій і воду свою та зарізане, що нарізав я для своїх стрижіїв, та й дам людям, яких не знаю, звідки то вони?
1SAM|25|12|І Давидові хлопці пішли назад на свою дорогу, і вернулися, і прийшли, і розповіли йому всі ці слова.
1SAM|25|13|А Давид сказав до людей своїх: Припережіть кожен меча свого! І приперезали кожен меча свого, і приперезав і Давид свого меча. І вийшло за Давидом близько чотирьох сотень чоловіка, а дві сотні остались при речах.
1SAM|25|14|А один хлопець із Навалових слуг доніс Авіґаїл, Наваловій жінці, говорячи: Ось Давид послав був із пустині посланців, щоб привітати нашого пана, а він кинувся на них.
1SAM|25|15|А ті люди дуже добрі для нас, і не були ми покривджені, і нічого нам не пропало за всі дні, коли ми ходили з ними, як були ми на полі.
1SAM|25|16|Муром були вони над нами і вночі, і вдень повсякчас, коли ми були з ними, як ми пасли отари.
1SAM|25|17|А тепер пізнай та побач, що зробиш, бо дозріло зло на нашого пана та на ввесь дім його. А він негідний, із ним не можна говорити.
1SAM|25|18|Тоді Авіґаїл поспішно взяла двісті хлібів, і два бурдюки вина, і п'ятеро приготовлених з отари, і п'ять сеїв пряженого зерна, а сто родзинок, та двісті сушених фіґ. І склала це на ослів.
1SAM|25|19|І сказала вона до своїх слуг: Ідіть передо мною, а я ось піду за вами.
1SAM|25|20|І сталося, як вона їхала на ослі й спускалася в гірському укритті, аж ось Давид та люди його сходять навперейми їй. І вона стрінула їх.
1SAM|25|21|А Давид сказав: Надармо ж пильнував я все, що належить тому чоловікові в пустині, і зо всього його нічого не пропало. Та він вернув мені злом за добро!
1SAM|25|22|Так нехай зробить Бог Давидовим ворогам, і так нехай додасть, якщо я позоставлю до ранку зо всього належного йому бодай те, що мочиться до стіни!
1SAM|25|23|А Авіґаїл побачила Давида, і поспішно зійшла з осла, і впала перед Давидом на обличчя своє, та й вклонилася до землі.
1SAM|25|24|І впала вона до ніг йому та й сказала: На мені самій, пане мій, ця провина! І дозволь говорити твоїй невільниці до ушей твоїх, а ти послухай слів своєї невільниці.
1SAM|25|25|Нехай же пан мій не кладе свого серця на цього негідного чоловіка, на Навала, бо яке ім'я його, такий він: Навал ім'я йому, і глупота з ним! А я, невільниця твоя, не бачила хлопців мого пана, що ти посилав.
1SAM|25|26|А тепер, мій пане, як живий Господь і як жива душа твоя! Господь стримає тебе, щоб ти не ввійшов до пролиття крови, і щоб рука твоя не допомогла в цьому тобі! А тепер нехай стануть, як Навал, вороги твої та ті, що шукають зла на пана мого!
1SAM|25|27|А оце дарунок, якого принесла твоя невільниця своєму панові, буде даний хлопцям, що служать моєму панові.
1SAM|25|28|Прости ж провину невільниці своєї, бо конче зробить Господь моєму панові вірний дім, бо пан мій провадить війни Господні, і зло не буде знайдене в тобі за твоїх днів.
1SAM|25|29|І хоч повстане хто гнати тебе, і шукати твоєї душі, то буде душа мого пана зв'язана у в'язці живих із Господом, Богом твоїм, а душу ворогів твоїх нехай Він її кине, як із пращі!
1SAM|25|30|І станеться, коли Господь зробить моєму панові все добре, що говорив про тебе, і настановить тебе володарем над Ізраїлем,
1SAM|25|31|то це не буде тобі на спотикання та на спокусу серця мого пана, як коли б пролив ти надармо кров, і пан мій пімстився сам. А коли Господь зробить добро моєму панові, то ти згадаєш про свою невільницю!
1SAM|25|32|І сказав Давид до Авіґаїл: Благословенний Господь, Бог Ізраїлів, що послав тебе на це навпроти мене!
1SAM|25|33|І благословенний розум твій, і благословенна ти, що стримала мене цього дня, щоб я не пішов на пролиття крови, і щоб рука моя не відімстила за мене.
1SAM|25|34|Але живий Господь, Бог Ізраїлів, що стримав мене зробити тобі зло, бо коли б ти була не поспішила, і не прийшла назустріч мені, то до світла ранку Навалові не зоставлено б навіть те, що мочиться до стіни!
1SAM|25|35|І взяв Давид із руки її те, що вона принесла йому, а їй сказав: Іди з миром до свого дому! Бачиш, я послухався голосу твого, і простив тобі!
1SAM|25|36|І прийшла Авіґаїл до Навала, аж ось у нього прийняття в його домі, немов прийняття царське! А Навалове серце було веселе в ньому, і він був дуже п'яний. І вона не розповіла йому нічого, ані малого, ані великого аж до світла ранку.
1SAM|25|37|І сталося, вранці, коли Навал витверезився, то жінка його розповіла йому про цю справу. І завмерло йому серце в його середині, і він став, як камінь.
1SAM|25|38|І сталося днів через десять, і вразив Господь Навала, і той помер.
1SAM|25|39|І почув Давид, що Навал помер, і сказав: Благословенний Господь, що розсудив справу образи моєї від Навала, а раба Свого стримав від зла, зло Навала звернув Господь на його голову! І Давид послав, і говорив про Авіґаїл, щоб узяти її собі за жінку.
1SAM|25|40|І прийшли Давидові раби до Авіґаїл на Кармел, і промовляли до неї, говорячи: Давид послав нас до тебе, щоб узяти тебе йому за жінку.
1SAM|25|41|А вона встала, і вклонилася лицем до землі, та й сказала: Ось твоя служниця готова стати невільницею, щоб мити ноги рабів пана мого!
1SAM|25|42|І Авіґаїл поспішно встала, і сіла на осла, а п'ятеро служанок її йшли при ногах її. І пішла вона за Давидовими посланцями, та й стала йому за жінку.
1SAM|25|43|А Ахіноам узяв Давида з Їзреелу, і вони обидві стали йому за жінок.
1SAM|25|44|А Саул віддав дочку свою Мелхолу, Давидову жінку, Палтієві, Лаїшевому синові, що з Ґалліму.
1SAM|26|1|І прийшли зіфеяни до Саула до Ґів'ї, говорячи: Он Давид ховається на взгір'ях Гахіли навпроти Єшімону!
1SAM|26|2|І встав Саул, і зійшов у пустиню Зіф, а з ним три тисячі чоловіка, вибраних із Ізраїля, щоб шукати Давида в пустині Зіф.
1SAM|26|3|І таборував Саул на згір'ї Гахіли, що навпроти Єшімону, на дорозі. А Давид пробував у пустині, і побачив, що Саул вийшов за ним до пустині.
1SAM|26|4|І послав Давид підглядачів, і довідався, що Саул дійсно прийшов.
1SAM|26|5|А Давид устав, і прийшов до місця, де таборував Саул. І Давид побачив те місце, де лежав Саул та Авнер, син Нерів, керівник його війська. А Саул лежав у таборі, а народ таборував навколо нього.
1SAM|26|6|І звернувся Давид, і сказав до хіттеянина Ахімелеха та до Авішая, Церуєвого сина, Йоавого брата, говорячи: Хто зійде зо мною до Саула до табору? І сказав Авішай: Я зійду з тобою!
1SAM|26|7|І прийшов Давид та Авішай до Саулового народу вночі, аж ось Саул лежить, спить у таборі, а спис його встромлений у землю в приголів'ї його, а Авнер та народ лежать навколо нього.
1SAM|26|8|І сказав Авішай до Давида: Сьогодні Бог видав твого ворога в руку твою, а тепер проколю я його списом аж до землі одним ударом, і не повторю йому!
1SAM|26|9|І сказав Давид до Авішая: Не губи його, бо хто простягав руку свою на Господнього помазанця, і був невинний?
1SAM|26|10|І сказав Давид: Як живий Господь, тільки Господь уразить його: або прийде день його і він помре, або він піде на війну і загине.
1SAM|26|11|Борони мене, Господи, простягнути свою руку на Господнього помазанця! А тепер візьми цього списа, що в приголів'ї його, та горня води, і ходімо собі!
1SAM|26|12|І взяв Давид списа та горня води з Саулового приголів'я, та й пішли собі. І ніхто не бачив, і не знав, і не збудився, бо всі вони спали, бо на них упав сон від Господа.
1SAM|26|13|І перейшов Давид на той бік, і став здалека на верховині гори, а між ними велика просторінь.
1SAM|26|14|І крикнув Давид до народу та до Авнера, Нерового сина, говорячи: Чи ж не відповіси, Авнере? А Авнер відповів та сказав: Хто ти, що кликав до царя?
1SAM|26|15|І сказав Давид до Авнера: Чи ти не муж? І хто рівний тобі в Ізраїлі? І чому не пильнував ти свого пана, царя? Бо приходив один із народу, щоб погубити царя, твого пана.
1SAM|26|16|Не добра це річ, що ти зробив! Як живий Господь, ви повинні померти, бо не пильнували ви пана свого, Господнього помазанця! А тепер побач, де царів спис, та де горня води, що були в приголів'ї його?
1SAM|26|17|І пізнав Саул Давидів голос, та й сказав: Чи це твій голос, сину мій Давиде? А Давид сказав: Мій голос, пане мій, царю!
1SAM|26|18|І далі сказав: Нащо то пан мій ганяється за своїм рабом? Бо що я зробив, і яке зло в моїй руці?
1SAM|26|19|А тепер нехай пан мій, цар, послухає слів свого раба. Якщо Господь намовив тебе проти мене, то нехай це станеться запашною жертвою, а якщо людські сини, прокляті вони перед Господнім лицем, бо вони відігнали мене сьогодні, щоб я не належав до Господнього спадку, говорячи: Іди, служи іншим богам!
1SAM|26|20|А тепер нехай не проллється моя кров на землю перед Господнім лицем, бо вийшов Ізраїлів цар шукати однієї блохи, як женуть куропатву в горах!
1SAM|26|21|І сказав Саул: Прогрішив я! Вернися, сину мій, Давиде, бо не вчиню вже тобі зла за те, що дороге було моє життя в очах твоїх цього дня. Оце був я нерозумний, і дуже багато помилявся.
1SAM|26|22|А Давид відповів та й сказав: Ось царів спис, і нехай прийде один із слуг, і нехай його візьме.
1SAM|26|23|А Господь відплатить кожному за його справедливість та правду його, що Господь дав тебе сьогодні в руку мою, та я не хотів підіймати своєї руки на Господнього помазанця.
1SAM|26|24|І ось, яке велике було життя твоє цього дня в очах моїх, таке велике нехай буде моє життя в очах Господа, і нехай Він урятує мене від усякого утиску!
1SAM|26|25|І сказав Саул до Давида: Благословенний ти, сину мій Давиде! І ти дійсно зробиш, і дійсно зможеш ти! І пішов Давид на свою дорогу, а Саул вернувся на своє місце.
1SAM|27|1|І сказав Давид у серці своїм: Колись я попадуся в Саулову руку. Нема мені ліпшого, як, утікаючи, утечу до филистимського краю, і відмовиться від мене Саул, щоб шукати мене вже по всій Ізраїлевій країні, і я втечу від руки його.
1SAM|27|2|І встав Давид, і перейшов він та шість сотень чоловіка, що з ним, до Ахіша, Маохового сина, ґатського царя.
1SAM|27|3|І осівся Давид з Ахішем у Ґаті, він та люди його, кожен із домом своїм, Давид та дві жінки його: ізреелітка Ахіноан та Авіґаїл, колишня жінка Навалова, кармелітка.
1SAM|27|4|І донесено Саулові, що Давид утік до Ґату, і він більш уже не шукав його.
1SAM|27|5|А Давид сказав до Ахіша: Якщо я знайшов милість в очах твоїх, нехай дадуть мені місце в одному з міст цієї землі, і нехай я осяду там. І чого сидітиме раб твій у місті твого царства разом із тобою?
1SAM|27|6|І дав йому Ахіш того дня Ціклаґ, чому належить Ціклаґ Юдиним царям аж до цього дня.
1SAM|27|7|А число днів, що Давид сидів на филистимській землі, було рік та чотири місяці.
1SAM|27|8|І сходив Давид та люди його, і нападали на Ґешуреянина, і на Ґірзеянина, і на Амаликитянина, бо вони мешканці цього краю відвіку, аж доти, як іти до Шуру, і аж до єгипетського краю.
1SAM|27|9|І побивав Давид той край, і не лишав при житті ані чоловіка, ані жінки, і забирав худобу дрібну та худобу велику, і осли, і верблюди, і одежу, і вертався, і приходив до Ахіша.
1SAM|27|10|І питався Ахіш: На кого нападали ви сьогодні? А Давид казав: На південь Юдин, і на південь Єрахмеелеянина, і на південь Кенеянина.
1SAM|27|11|А Давид не лишав при житті ані чоловіка, ані жінки, щоб привести до Ґату, говорячи: Щоб не донесли на нас, кажучи: Так зробив Давид, і такий його звичай по всі дні, коли сидів на филистимській землі.
1SAM|27|12|І вірив Ахіш Давидові, говорячи: Справді обриднув він своєму народові в Ізраїлі, і буде мені за вічного раба!
1SAM|28|1|І сталося тими днями, і зібрали филистимляни свої військові табори, щоб воювати з Ізраїлем. І сказав Ахіш до Давида: Щоб ти певно знав, що вийдеш зо мною в таборі, ти та люди твої.
1SAM|28|2|І сказав Давид до Ахіша: Тому тепер ти пізнаєш, що зробить твій раб. А Ахіш сказав до Давида: Тому то зроблю тебе сторожем моєї голови по всі дні.
1SAM|28|3|А Самуїл тоді помер, і оплакував його ввесь Ізраїль, і поховали його в Рамі, у його місті. А Саул повиганяв із Краю ворожбитів та віщунів.
1SAM|28|4|І зібралися филистимляни, і прийшли, і таборували в Шунемі. А Саул зібрав усього Ізраїля, і таборували в Ґілбоа.
1SAM|28|5|І побачив Саул филистимський табір та й злякався, і сильно затремтіло йому серце.
1SAM|28|6|І питався Саул Господа, та не відповів йому Господь ані в снах, ані урімом, ані пророками.
1SAM|28|7|І сказав Саул до своїх рабів: Пошукайте мені жінку ворожку, і я піду до неї, і запитаю її. І відповіли йому раби його: Ось жінка ворожка, в Ен-Дорі.
1SAM|28|8|І перебрався Саул, і надів іншу одежу, і пішов він та двоє людей з ним, і прийшли до тієї жінки вночі. А він сказав: Поворожи мені, і виклич мені того, кого скажу тобі.
1SAM|28|9|А та жінка відповіла йому: Ти ж знаєш, що зробив Саул, що в Краю він вигубив ворожбитів та віщунів. І нащо ти важиш на мою душу, щоб забити її?
1SAM|28|10|І Саул присягнув їй Господом, говорячи: Як живий Господь, не спіткає тебе вина за цю річ!
1SAM|28|11|І сказала та жінка: Кого я викличу тобі? А він відказав: Самуїла виклич мені.
1SAM|28|12|І побачила та жінка Самуїла, та й крикнула сильним голосом! І сказала та жінка до Саула, говорячи: Нащо ти обманив мене, таж ти Саул!
1SAM|28|13|І сказав їй цар; Не бійся! Але що ти бачиш? А та жінка відказала Саулові: Я бачу ніби богів, що виходять із землі!
1SAM|28|14|І він їй сказав: Який його вид? А та відказала: Виходить старий чоловік, зодягнений у довгу одежу. І Саул пізнав, що то Самуїл, і схилив своє обличчя до землі, та й уклонився.
1SAM|28|15|І сказав Самуїл до Саула: Нащо ти непокоїш мене, мене викликаючи? А Саул сказав: Дуже тяжко мені, филистимляни воюють зо мною, а Бог відступився від мене, і не відповідає мені вже ані через пророків, ані в снах. І покликав я тебе, щоб ти навчив мене, що я маю робити.
1SAM|28|16|І сказав Самуїл: І нащо ти питаєш мене, коли Господь відступився від тебе, і став із твоїм ворогом?
1SAM|28|17|І Господь зробив йому, як говорив був через мене, Господь узяв царство з твоєї руки, і дав його твоєму ближньому, Давидові.
1SAM|28|18|Як ти не слухався Господнього голосу, і не виконав полум'яного гніву Його на Амалика, тому Господь зробив тобі цю річ цього дня.
1SAM|28|19|І Господь віддав із тобою також Ізраїля до руки филистимлян. А взавтра ти та сини твої будете разом зо мною; також Ізраїлевого табора віддасть Господь до руки филистимлян.
1SAM|28|20|І Саул відразу повалився на землю всім своїм зростом, сильно він злякався Самуїлових слів, та й сили не було в ньому, бо не їв він хліба цілий той день та цілу ту ніч.
1SAM|28|21|І підійшла та жінка до Саула й побачила, що він дуже пригнічений. І сказала до нього: Ось невільниця твоя послухалася твого голосу, і наразила життя своє на небезпеку, бо я послухалася слів твоїх, що ти говорив мені.
1SAM|28|22|А тепер ти послухай також голосу своєї невільниці, я покладу перед тобою шматок хліба, а ти з'їж і буде в тобі сила, коли підеш дорогою.
1SAM|28|23|А він відмовився й сказав: Не буду їсти! Та сильно просили його слуги його та тая жінка, і він послухався їхнього голосу. І звівся він із землі, і всівся на ліжку.
1SAM|28|24|А та жінка мала в домі годоване теля, і поспішно зарізала його. І взяла вона муки й замісила, і спекла з того прісне.
1SAM|28|25|І принесла те перед Саула та перед слуг його, і вони їли. Потім устали й пішли тієї ночі.
1SAM|29|1|І зібрали филистимляни всі свої війська до Афеку, а Ізраїль таборував в Аїні, що в Їзреелі.
1SAM|29|2|А филистимські князі переходили за сотнями та за тисячами, Давид же та люди його ішли накінці разом з Ахішем.
1SAM|29|3|І казали филистимські князі: Що це за євреї? А Ахіш відказав филистимським князям: Таж це Давид, раб Саула, Ізраїлевого царя, що був зо мною певний час, чи то роки, а я не знайшов у ньому нічого злого від дня його приходу аж до дня цього.
1SAM|29|4|І гнівалися на нього филистимські князі. І сказали йому филистимські князі: Заверни того чоловіка, і нехай він вернеться до свого місця, де ти призначив йому, і нехай він не йде з нами на війну, і не стане нам противником на війні. І чим він може подобатися своєму панові? Хіба головами цих людей?
1SAM|29|5|Чи ж це не той Давид, що про нього співали в танцях, говорячи: Саул повбивав свої тисячі, а Давид десятки тисяч свої!
1SAM|29|6|І покликав Ахіш Давида, і сказав до нього: Як живий Господь, ти правдивий, і в моїх очах добрий твій вихід та вхід твій зо мною в таборі, бо я не знайшов у тобі зла від дня приходу твого до мене аж до цього дня. Та в очах князів ти не добрий.
1SAM|29|7|А тепер вернися та йди в мирі, і не зробиш зла в очах филистимських князів.
1SAM|29|8|А Давид сказав до Ахіша: Що ж зробив я? І що ти знайшов у своєму рабові від дня, коли став я перед твоїм обличчям, аж до цього дня, що я не вийду й не буду воювати з ворогами мого пана, царя?
1SAM|29|9|І відповів Ахіш і сказав до Давида: Знаю я, що ти добрий в очах моїх, немов Ангол Божий. Та филистимські князі сказали: Нехай не йде він із нами на війну!
1SAM|29|10|А тепер устань рано вранці ти та раби пана твого, що прийшли з тобою. І повставайте рано вранці, і як вам розсвіне, ідіть!
1SAM|29|11|І встав рано вранці Давид та люди його, щоб піти ранком і вернутися до филистимського краю. А филистимляни пішли до Ізраїля.
1SAM|30|1|І сталося, коли Давид та люди його йшли до Ціклаґу, третього дня, то амаликитяни вдерлися до півдня та до Ціклаґу, і побили Ціклаґ та спалили його огнем.
1SAM|30|2|І позабирали вони до неволі жінок, що були в ньому, від малого аж до великого, нікого не забили, але забрали, та й пішли своєю дорогою.
1SAM|30|3|І прийшов Давид та його люди до того міста, а воно спалене огнем! А їхні жінки, та сини їхні, та їхні дочки забрані в неволю.
1SAM|30|4|І підніс Давид та народ, що з ним, свій голос, та й плакали, аж поки не стало їм сили плакати.
1SAM|30|5|І були взяті до неволі обидві Давидові жінки: їзреелітка Ахіноам та Авіґаїл, колишня жінка кармелітянина Навала.
1SAM|30|6|І було Давидові дуже гірко, бо народ говорив, щоб його вкаменувати, бо засмутилася душа всього народу, кожен обурився за синів своїх та за дочок своїх. Та Давид зміцнився Господом, Богом, своїм.
1SAM|30|7|І сказав Давид до священика Евіятара, Ахімелехового сина: Принеси до мене ефода! І Евіятар приніс ефода до Давида.
1SAM|30|8|І запитав Давид Господа, говорячи: Чи мені гнатися за тією ордою, чи дожену її? А Він відказав йому: Женися, бо конче доженеш, і конче визволиш.
1SAM|30|9|І пішов Давид, він та шість сотень люда, що з ним, і вони прийшли аж до потоку Бесор; а відсталі спинилися.
1SAM|30|10|І гнався Давид, він та чотири сотні чоловіка. А двісті люда спинилися, бо були слабі, щоб перейти потока Бесор.
1SAM|30|11|І знайшли вони в полі єгиптянина, і привели його до Давида, і дали йому хліба, а він їв, і напоїли його водою.
1SAM|30|12|І дали йому половину грудки сушених фіґ та дві в'язки родзинок. І він з'їв, і вернувся дух його до нього, бо він не їв хліба та не пив води три дні та три ночі.
1SAM|30|13|І запитав його Давид: Чий ти та звідкіля ти? А той відказав: Я єгипетський юнак, раб амаликитянина. Та покинув мене пан мій, бо я захворів три дні тому.
1SAM|30|14|Ми були вдерлися на південь керетеїв, і на той, що Юдин, та на південь Калева. А Ціклаґ ми спалили огнем.
1SAM|30|15|І сказав йому Давид: Чи не заведеш мене до тієї орди? А той відповів: Присягни мені Богом, що не вб'єш мене, і що не видаси мене в руку мого пана, то спроваджу тебе до тієї орди.
1SAM|30|16|І він спровадив його, аж ось вони розпорошені по поверхні всієї тієї землі, їдять та п'ють та святкують з приводу всієї тієї великої здобичі, що вони набрали з филистимського краю та з Краю Юдиного.
1SAM|30|17|І бив їх Давид від ранку аж до вечора наступного дня, і не втік із них ніхто, крім чотирьохсот чоловіка хлопців, що повсідали на верблюдів, і повтікали.
1SAM|30|18|І врятував Давид усе, що позабирав був Амалик. І обидві свої жінки Давид урятував.
1SAM|30|19|І не пропало їм нічого: усе, від малого й аж до великого, і аж до синів та дочок, і від здобичі, і аж до всього, що ті взяли були собі, усе вернув Давид!
1SAM|30|20|І взяв Давид усю худобу дрібну та худобу велику, а ті, що йшли перед тією чередою, говорили: Це Давидова здобич!
1SAM|30|21|Потому прийшов Давид до тих двохсот людей, що були слабі, щоб іти за Давидом, і що їх він лишив був при потоці Бесор, а вони повиходили назустріч Давидові та назустріч народові, що з ним. І підійшов Давид до народу, і запитався їх про мир.
1SAM|30|22|І стали говорити всі люди злі та негідні з тих людей, що ходили з Давидом, та й сказали: Вони не ходили з нами, тому не дамо їм зо здобичі, що ми відняли, бо кожному дамо тільки жінок його та синів його, нехай відведуть, і нехай ідуть!
1SAM|30|23|А Давид сказав: Не робіть так, браття мої, з тим, що дав нам Господь, і пильнував нас, і дав орду, що йшла на нас, у нашу руку.
1SAM|30|24|А хто послухає вас у такій речі? Бо яка частина того, хто ходив до бою, то така частина й того, хто сидів при речах, рівно поділять.
1SAM|30|25|І сталося від цього дня й далі, і зробив він це за постанову та за звичай для Ізраїля, і він існує аж до цього дня.
1SAM|30|26|І прийшов Давид до Ціклаґу, і послав зо здобичі Юдиним старшим, приятелям своїм, говорячи: Оце вам подарок зо здобичі Господніх ворогів,
1SAM|30|27|тим, що в Бет-Елі, і тим, що в Рамоті південнім, і тим, що в Яттері,
1SAM|30|28|і тим, що в Ароері, і тим, що в Сіфмоті, і тим, що в Ештемоа,
1SAM|30|29|і тим, що в Рахалі, і тим, що в містах Єрахмелеянина, і тим, що в містах Кенеянина,
1SAM|30|30|і тим, що в Хормі, і тим, що в Бор-Ашані, і тим, що в Атаху,
1SAM|30|31|і тим, що в Хевроні, і до всіх тих місць, куди ходив Давид, він та люди його.
1SAM|31|1|А филистимляни воювали з Ізраїлем. І побігли Ізраїлеві мужі перед филистимлянами, і падали трупами на горі Ґілбоа.
1SAM|31|2|І догнали филистимляни Саула та його синів. І повбивали филистимляни Йонатана й Авінадава та Малкі-Шуя, Саулових синів.
1SAM|31|3|І став бій тяжкий для Саула, і його знайшли лучники, він був дуже поранений тими лучниками.
1SAM|31|4|І сказав Саул до свого зброєноші: Витягни меча свого, і пробий мене ним, щоб не прийшли ці необрізані, і не пробили мене, і не знущалися надо мною! Та не хотів зброєноша, бо дуже боявся. Тоді взяв Саул меча, та й упав на нього!
1SAM|31|5|І побачив зброєноша, що помер Саул, і впав і він на свого меча, та й помер із ним.
1SAM|31|6|І помер того дня Саул і троє синів його та зброєноша, також усі люди разом.
1SAM|31|7|А ізраїльтяни, що мешкали на тім боці долини й на тім боці Йордану, коли побачили, що повтікали ізраїльтяни, і що померли Саул та сини його, покидали ті міста й повтікали, а филистимляни поприходили й осілися в них.
1SAM|31|8|І сталося другого дня, і прийшли филистимляни, щоб пообдирати трупи, та й знайшли Саула та трьох синів його, що лежали на горі Ґілбоа.
1SAM|31|9|І вони стяли йому голову, і поздирали зброю його, і послали в филистимські краї навколо, щоб сповістити в домах їхніх божків та народові.
1SAM|31|10|І вони поклали зброю його в домі Астарти, а тіло його прибили на мурі Бет-Шану.
1SAM|31|11|І почули мешканці ґілеадського Явешу про те, що филистимляни зробили Саулові,
1SAM|31|12|і встали всі хоробрі, і йшли всю ніч, і взяли Саулове тіло та тіла синів його з муру Бет-Шану, і прийшли до Явешу, та й спалили їх там.
1SAM|31|13|І взяли вони їхні кості, і поховали під тамариском в Явешу, та й постили сім день.
