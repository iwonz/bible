1PET|1|1|Petrus apostolus Iesu Christi electis advenis dispersionis Ponti Galatiae Cappadociae Asiae et Bithyniae
1PET|1|2|secundum praescientiam Dei Patris in sanctificatione Spiritus in oboedientiam et aspersionem sanguinis Iesu Christi gratia vobis et pax multiplicetur
1PET|1|3|benedictus Deus et Pater Domini nostri Iesu Christi qui secundum magnam misericordiam suam regeneravit nos in spem vivam per resurrectionem Iesu Christi ex mortuis
1PET|1|4|in hereditatem incorruptibilem et incontaminatam et inmarcescibilem conservatam in caelis in vobis
1PET|1|5|qui in virtute Dei custodimini per fidem in salutem paratam revelari in tempore novissimo
1PET|1|6|in quo exultatis modicum nunc si oportet contristati in variis temptationibus
1PET|1|7|ut probatum vestrae fidei multo pretiosius sit auro quod perit per ignem probato inveniatur in laudem et gloriam et honorem in revelatione Iesu Christi
1PET|1|8|quem cum non videritis diligitis in quem nunc quoque non videntes credentes autem exultatis laetitia inenarrabili et glorificata
1PET|1|9|reportantes finem fidei vestrae salutem animarum
1PET|1|10|de qua salute exquisierunt atque scrutati sunt prophetae qui de futura in vobis gratia prophetaverunt
1PET|1|11|scrutantes in quod vel quale tempus significaret in eis Spiritus Christi praenuntians eas quae in Christo sunt passiones et posteriores glorias
1PET|1|12|quibus revelatum est quia non sibi ipsis vobis autem ministrabant ea quae nunc nuntiata sunt vobis per eos qui evangelizaverunt vos Spiritu Sancto misso de caelo in quae desiderant angeli prospicere
1PET|1|13|propter quod succincti lumbos mentis vestrae sobrii perfecte sperate in eam quae offertur vobis gratiam in revelatione Iesu Christi
1PET|1|14|quasi filii oboedientiae non configurati prioribus ignorantiae vestrae desideriis
1PET|1|15|sed secundum eum qui vocavit vos sanctum et ipsi sancti in omni conversatione sitis
1PET|1|16|quoniam scriptum est sancti eritis quia ego sanctus sum
1PET|1|17|et si Patrem invocatis eum qui sine acceptione personarum iudicat secundum uniuscuiusque opus in timore incolatus vestri tempore conversamini
1PET|1|18|scientes quod non corruptibilibus argento vel auro redempti estis de vana vestra conversatione paternae traditionis
1PET|1|19|sed pretioso sanguine quasi agni incontaminati et inmaculati Christi
1PET|1|20|praecogniti quidem ante constitutionem mundi manifestati autem novissimis temporibus propter vos
1PET|1|21|qui per ipsum fideles estis in Deo qui suscitavit eum a mortuis et dedit ei gloriam ut fides vestra et spes esset in Deo
1PET|1|22|animas vestras castificantes in oboedientia caritatis in fraternitatis amore simplici ex corde invicem diligite adtentius
1PET|1|23|renati non ex semine corruptibili sed incorruptibili per verbum Dei vivi et permanentis
1PET|1|24|quia omnis caro ut faenum et omnis gloria eius tamquam flos faeni exaruit faenum et flos decidit
1PET|1|25|verbum autem Domini manet in aeternum hoc est autem verbum quod evangelizatum est in vos
1PET|2|1|deponentes igitur omnem malitiam et omnem dolum et simulationes et invidias et omnes detractiones
1PET|2|2|sicut modo geniti infantes rationale sine dolo lac concupiscite ut in eo crescatis in salutem
1PET|2|3|si gustastis quoniam dulcis Dominus
1PET|2|4|ad quem accedentes lapidem vivum ab hominibus quidem reprobatum a Deo autem electum honorificatum
1PET|2|5|et ipsi tamquam lapides vivi superaedificamini domus spiritalis sacerdotium sanctum offerre spiritales hostias acceptabiles Deo per Iesum Christum
1PET|2|6|propter quod continet in scriptura ecce pono in Sion lapidem summum angularem electum pretiosum et qui crediderit in eo non confundetur
1PET|2|7|vobis igitur honor credentibus non credentibus autem lapis quem reprobaverunt aedificantes hic factus est in caput anguli
1PET|2|8|et lapis offensionis et petra scandali qui offendunt verbo nec credunt in quod et positi sunt
1PET|2|9|vos autem genus electum regale sacerdotium gens sancta populus adquisitionis ut virtutes adnuntietis eius qui de tenebris vos vocavit in admirabile lumen suum
1PET|2|10|qui aliquando non populus nunc autem populus Dei qui non consecuti misericordiam nunc autem misericordiam consecuti
1PET|2|11|carissimi obsecro tamquam advenas et peregrinos abstinere vos a carnalibus desideriis quae militant adversus animam
1PET|2|12|conversationem vestram inter gentes habentes bonam ut in eo quod detractant de vobis tamquam de malefactoribus ex bonis operibus considerantes glorificent Deum in die visitationis
1PET|2|13|subiecti estote omni humanae creaturae propter Dominum sive regi quasi praecellenti
1PET|2|14|sive ducibus tamquam ab eo missis ad vindictam malefactorum laudem vero bonorum
1PET|2|15|quia sic est voluntas Dei ut benefacientes obmutescere faciatis inprudentium hominum ignorantiam
1PET|2|16|quasi liberi et non quasi velamen habentes malitiae libertatem sed sicut servi Dei
1PET|2|17|omnes honorate fraternitatem diligite Deum timete regem honorificate
1PET|2|18|servi subditi in omni timore dominis non tantum bonis et modestis sed etiam discolis
1PET|2|19|haec est enim gratia si propter conscientiam Dei sustinet quis tristitias patiens iniuste
1PET|2|20|quae enim gloria est si peccantes et colaphizati suffertis sed si benefacientes et patientes sustinetis haec est gratia apud Deum
1PET|2|21|in hoc enim vocati estis quia et Christus passus est pro vobis vobis relinquens exemplum ut sequamini vestigia eius
1PET|2|22|qui peccatum non fecit nec inventus est dolus in ore ipsius
1PET|2|23|qui cum malediceretur non maledicebat cum pateretur non comminabatur tradebat autem iudicanti se iniuste
1PET|2|24|qui peccata nostra ipse pertulit in corpore suo super lignum ut peccatis mortui iustitiae viveremus cuius livore sanati estis
1PET|2|25|eratis enim sicut oves errantes sed conversi estis nunc ad pastorem et episcopum animarum vestrarum
1PET|3|1|similiter mulieres subditae suis viris ut et si qui non credunt verbo per mulierum conversationem sine verbo lucri fiant
1PET|3|2|considerantes in timore castam conversationem vestram
1PET|3|3|quarum sit non extrinsecus capillaturae aut circumdatio auri aut indumenti vestimentorum cultus
1PET|3|4|sed qui absconditus cordis est homo in incorruptibilitate quieti et modesti spiritus quod est in conspectu Dei locuples
1PET|3|5|sic enim aliquando et sanctae mulieres sperantes in Deo ornabant se subiectae propriis viris
1PET|3|6|sicut Sarra oboediebat Abrahae dominum eum vocans cuius estis filiae benefacientes et non timentes ullam perturbationem
1PET|3|7|viri similiter cohabitantes secundum scientiam quasi infirmiori vaso muliebri inpertientes honorem tamquam et coheredibus gratiae vitae uti ne inpediantur orationes vestrae
1PET|3|8|in fine autem omnes unianimes conpatientes fraternitatis amatores misericordes humiles
1PET|3|9|non reddentes malum pro malo vel maledictum pro maledicto sed e contrario benedicentes quia in hoc vocati estis ut benedictionem hereditate possideatis
1PET|3|10|qui enim vult vitam diligere et videre dies bonos coerceat linguam suam a malo et labia eius ne loquantur dolum
1PET|3|11|declinet autem a malo et faciat bonum inquirat pacem et persequatur eam
1PET|3|12|quia oculi Domini super iustos et aures eius in preces eorum vultus autem Domini super facientes mala
1PET|3|13|et quis est qui vobis noceat si boni aemulatores fueritis
1PET|3|14|sed et si quid patimini propter iustitiam beati timorem autem eorum ne timueritis et non conturbemini
1PET|3|15|Dominum autem Christum sanctificate in cordibus vestris parati semper ad satisfactionem omni poscenti vos rationem de ea quae in vobis est spe
1PET|3|16|sed cum modestia et timore conscientiam habentes bonam ut in eo quod detrahunt vobis confundantur qui calumniantur vestram bonam in Christo conversationem
1PET|3|17|melius est enim benefacientes si velit voluntas Dei pati quam malefacientes
1PET|3|18|quia et Christus semel pro peccatis mortuus est iustus pro iniustis ut nos offerret Deo mortificatus carne vivificatus autem spiritu
1PET|3|19|in quo et his qui in carcere erant spiritibus veniens praedicavit
1PET|3|20|qui increduli fuerant aliquando quando expectabat Dei patientia in diebus Noe cum fabricaretur arca in qua pauci id est octo animae salvae factae sunt per aquam
1PET|3|21|quod et vos nunc similis formae salvos facit baptisma non carnis depositio sordium sed conscientiae bonae interrogatio in Deum per resurrectionem Iesu Christi
1PET|3|22|qui est in dextera Dei profectus in caelum subiectis sibi angelis et potestatibus et virtutibus
1PET|4|1|Christo igitur passo in carne et vos eadem cogitatione armamini quia qui passus est carne desiit a peccatis
1PET|4|2|ut iam non hominum desideriis sed voluntate Dei quod reliquum est in carne vivat temporis
1PET|4|3|sufficit enim praeteritum tempus ad voluntatem gentium consummandam qui ambulaverunt in luxuriis desideriis vinolentiis comesationibus potationibus et inlicitis idolorum cultibus
1PET|4|4|in quo peregrinantur non concurrentibus vobis in eandem luxuriae confusionem blasphemantes
1PET|4|5|qui reddent rationem ei qui paratus est iudicare vivos et mortuos
1PET|4|6|propter hoc enim et mortuis evangelizatum est ut iudicentur quidem secundum homines in carne vivant autem secundum Deum spiritu
1PET|4|7|omnium autem finis adpropinquavit estote itaque prudentes et vigilate in orationibus
1PET|4|8|ante omnia mutuam in vosmet ipsos caritatem continuam habentes quia caritas operit multitudinem peccatorum
1PET|4|9|hospitales invicem sine murmuratione
1PET|4|10|unusquisque sicut accepit gratiam in alterutrum illam administrantes sicut boni dispensatores multiformis gratiae Dei
1PET|4|11|si quis loquitur quasi sermones Dei si quis ministrat tamquam ex virtute quam administrat Deus ut in omnibus honorificetur Deus per Iesum Christum cui est gloria et imperium in saecula saeculorum amen
1PET|4|12|carissimi nolite peregrinari in fervore qui ad temptationem vobis fit quasi novi aliquid vobis contingat
1PET|4|13|sed communicantes Christi passionibus gaudete ut et in revelatione gloriae eius gaudeatis exultantes
1PET|4|14|si exprobramini in nomine Christi beati quoniam gloriae Dei Spiritus in vobis requiescit
1PET|4|15|nemo enim vestrum patiatur quasi homicida aut fur aut maledicus aut alienorum appetitor
1PET|4|16|si autem ut Christianus non erubescat glorificet autem Deum in isto nomine
1PET|4|17|quoniam tempus ut incipiat iudicium de domo Dei si autem primum a nobis qui finis eorum qui non credunt Dei evangelio
1PET|4|18|et si iustus vix salvatur impius et peccator ubi parebit
1PET|4|19|itaque et hii qui patiuntur secundum voluntatem Dei fideli creatori commendant animas suas in benefactis
1PET|5|1|seniores ergo qui in vobis sunt obsecro consenior et testis Christi passionum qui et eius quae in futuro revelanda est gloriae communicator
1PET|5|2|pascite qui est in vobis gregem Dei providentes non coacto sed spontanee secundum Deum neque turpis lucri gratia sed voluntarie
1PET|5|3|neque ut dominantes in cleris sed formae facti gregi et ex animo
1PET|5|4|et cum apparuerit princeps pastorum percipietis inmarcescibilem gloriae coronam
1PET|5|5|similiter adulescentes subditi estote senioribus omnes autem invicem humilitatem insinuate quia Deus superbis resistit humilibus autem dat gratiam
1PET|5|6|humiliamini igitur sub potenti manu Dei ut vos exaltet in tempore visitationis
1PET|5|7|omnem sollicitudinem vestram proicientes in eum quoniam ipsi cura est de vobis
1PET|5|8|sobrii estote vigilate quia adversarius vester diabolus tamquam leo rugiens circuit quaerens quem devoret
1PET|5|9|cui resistite fortes fide scientes eadem passionum ei quae in mundo est vestrae fraternitati fieri
1PET|5|10|Deus autem omnis gratiae qui vocavit nos in aeternam suam gloriam in Christo Iesu modicum passos ipse perficiet confirmabit solidabit
1PET|5|11|ipsi imperium in saecula saeculorum amen
1PET|5|12|per Silvanum vobis fidelem fratrem ut arbitror breviter scripsi obsecrans et contestans hanc esse veram gratiam Dei in qua state
1PET|5|13|salutat vos quae est in Babylone cumelecta et Marcus filius meus
1PET|5|14|salutate invicem in osculo sancto gratia vobis omnibus qui estis in Christo
