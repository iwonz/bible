DAN|1|1|猶大 王 約雅敬 在位第三年， 巴比倫 王 尼布甲尼撒 來到 耶路撒冷 ，將城圍困。
DAN|1|2|主將 猶大 王 約雅敬 和上帝殿中的一些器皿交在他的手中。他就把他們帶到 示拿 地他神明的廟裏，將器皿收入他神明的庫房中。
DAN|1|3|王吩咐太監長 亞施毗拿 ，從 以色列 人的王室後裔和貴族中帶進幾個人來，
DAN|1|4|就是沒有殘疾、相貌俊美、通達各樣學問 、知識聰明俱備、足能在王宮侍立的少年，要教他們 迦勒底 的文字和語言。
DAN|1|5|王從自己所用的膳和所飲的酒中，派給他們每日的分量，養育他們三年，好叫他們期滿以後侍立在王面前。
DAN|1|6|他們中間有 猶大 人 但以理 、 哈拿尼雅 、 米沙利 和 亞撒利雅 。
DAN|1|7|太監長給他們另外起名，稱 但以理 為 伯提沙撒 ，稱 哈拿尼雅 為 沙得拉 ，稱 米沙利 為 米煞 ，稱 亞撒利雅 為 亞伯尼歌 。
DAN|1|8|但以理 卻立志，不以王的膳和王所飲的酒玷污自己，於是懇求太監長容他不使自己玷污。
DAN|1|9|上帝使 但以理 在太監長眼前蒙恩，得憐憫。
DAN|1|10|太監長對 但以理 說：「我懼怕我主我王，他已經派給你們飲食，何必讓他見你們的面貌比你們同年齡的少年憔悴呢？這樣，你們就使我的頭在王那裏不保了。」
DAN|1|11|但以理 對太監長所派監管 但以理 、 哈拿尼雅 、 米沙利 、 亞撒利雅 的管理者說：
DAN|1|12|「請你考驗僕人們十天，給我們素菜吃，清水喝，
DAN|1|13|然後你親自觀察我們的面貌和那用王膳的少年的面貌；就照你所觀察的待你的僕人吧！」
DAN|1|14|管理者准許他們這件事，考驗他們十天。
DAN|1|15|過了十天，他們的身材看來比所有享用王膳的少年更加俊美健壯，
DAN|1|16|於是管理者撤去王派給他們用的膳和所飲的酒，只給他們素菜。
DAN|1|17|這四個少年，上帝在各樣文字學問上賜給他們知識和聰明； 但以理 又明白各樣異象和夢兆。
DAN|1|18|王吩咐帶他們進宮的日子到了，太監長就把他們帶到 尼布甲尼撒 面前。
DAN|1|19|王與他們談論，在所有少年中找不到人能與 但以理 、 哈拿尼雅 、 米沙利 、 亞撒利雅 相比，於是他們就在王面前侍立。
DAN|1|20|王考問他們一切智慧和聰明的事，發現他們比全國所有的術士和巫師勝過十倍。
DAN|1|21|到 居魯士 王元年， 但以理 還健在。
DAN|2|1|尼布甲尼撒 在位第二年，他做了很多夢，心裏煩亂，不能睡覺。
DAN|2|2|王吩咐人將術士、巫師、行邪術的和 迦勒底 人召來，要他們把王的夢告訴王；他們就來，站在王面前。
DAN|2|3|王對他們說：「我做了一個夢，心裏煩亂，想要知道這是甚麼夢。」
DAN|2|4|迦勒底 人用 亞蘭 話對王說：「願王萬歲！請將夢告訴僕人，我們就可以講解。」
DAN|2|5|王回答 迦勒底 人說：「這事我已決定，你們若不把夢和夢的解釋告訴我，就必被凌遲，你們的房屋必成糞堆；
DAN|2|6|但你們若能說出這個夢和夢的解釋，就必從我得到禮物、賞賜和殊榮。現在，你們要把夢和夢的解釋告訴我。」
DAN|2|7|他們再一次回答說：「請王將夢告訴僕人，我們就可以講解。」
DAN|2|8|王回答說：「我確實知道你們是故意拖延，因為你們知道這事我已決定。
DAN|2|9|你們若不將夢告訴我，只有一個辦法對待你們；因為你們彼此串通，向我胡言亂語，要等候情勢改變。現在，你們要將夢告訴我，讓我知道你們真能為我解夢。」
DAN|2|10|迦勒底 人回答王說：「世上沒有人能解釋王的事情；從來沒有君王、大臣、掌權者向術士、巫師，或 迦勒底 人問過這樣的事。
DAN|2|11|王所問的事很難，除了不與血肉之軀同住的上帝，沒有人能在王面前解釋。」
DAN|2|12|王因這事生氣，大大震怒，吩咐滅絕 巴比倫 所有的智慧人。
DAN|2|13|命令發出，智慧人將要被殺，人就尋找 但以理 和他的同伴，要殺他們。
DAN|2|14|王的護衛長 亞略 奉命去殺 巴比倫 的智慧人， 但以理 用婉言和智慧回應，
DAN|2|15|向王的大臣 亞略 說：「王的命令為何這樣緊急呢？」 亞略 就把事情告訴 但以理 。
DAN|2|16|於是 但以理 進去求王寬限，好為王解夢。
DAN|2|17|但以理 回到他的居所，把這事告訴他的同伴 哈拿尼雅 、 米沙利 、 亞撒利雅 ，
DAN|2|18|要他們祈求天上的上帝施憐憫，將這奧祕指明，免得 但以理 和他的同伴與 巴比倫 其餘的智慧人一同滅亡。
DAN|2|19|這奧祕就在夜間異象中顯明給 但以理 ， 但以理 就稱頌天上的上帝。
DAN|2|20|但以理 說： 「上帝的名是應當稱頌的，從亙古直到永遠！ 因為智慧和能力都屬乎他。
DAN|2|21|他改變時間、季節， 他廢王，立王； 將智慧賜給智慧人， 將知識賜給聰明人。
DAN|2|22|他顯明深奧隱祕的事， 洞悉幽暗中的一切， 光明也與他同住。
DAN|2|23|我列祖的上帝啊，我感謝你，讚美你， 因你將智慧才能賜給我， 我們所求問的現在你已指明給我， 把王的事給我們指明。」
DAN|2|24|於是， 但以理 進到王所派滅絕 巴比倫 智慧人的 亞略 那裏去，對他這樣說：「不要滅絕 巴比倫 的智慧人，求你領我到王面前，我可以為王解夢。」
DAN|2|25|亞略 就急忙領 但以理 到王面前，對王這樣說：「我在被擄的 猶大 人中找到一人，能將夢的解釋告訴王。」
DAN|2|26|王對那稱為 伯提沙撒 的 但以理 說：「你能將我所做的夢和夢的解釋告訴我嗎？」
DAN|2|27|但以理 回答王說：「王所問的那奧祕，智慧人、巫師、術士、觀兆的都不能告訴王，
DAN|2|28|只有那在天上的上帝能顯明奧祕。他已把日後將要發生的事指示 尼布甲尼撒 王。你在床上做的夢和你腦中的異象是這樣：
DAN|2|29|你，王啊，你在床上所思想的是關乎日後的事，那顯明奧祕的主已把將來要發生的事指示你。
DAN|2|30|至於我，那奧祕顯明給我，並非因我智慧勝過一切活著的人，而是為了讓王知道夢的解釋，知道你心裏的意念。
DAN|2|31|「你，王啊，你正觀看，看哪，有一個很大的像，這像甚高，極其光耀，立在你面前，形狀非常可怕。
DAN|2|32|這像的頭是純金的，胸膛和膀臂是銀的，腹部和腰是銅的，
DAN|2|33|腿是鐵的，腳是半鐵半泥的。
DAN|2|34|你正觀看，見有一塊非人手鑿出來的石頭打在它半鐵半泥的腳上，把腳砸碎；
DAN|2|35|於是鐵、泥、銅、銀、金都一同砸得粉碎，如夏天禾場上的糠秕，被風吹散，無處可尋。打碎這像的石頭成了一座大山，覆蓋全地。
DAN|2|36|「這就是那夢；我們要在王面前講解那夢。
DAN|2|37|你，王啊，你是諸王之王。天上的上帝已將國度、權勢、能力、尊榮都賜給你。
DAN|2|38|世人和走獸，並天空的飛鳥，不論居住何處，他都交在你的手中，令你掌管這一切。你就是那金的頭。
DAN|2|39|在你以後必興起另一國，不及於你；又有第三國如銅，必掌管全地。
DAN|2|40|第四國必堅壯如鐵，就像鐵能打碎砸碎一切；鐵怎樣壓碎一切，那國也必照樣打碎壓碎。
DAN|2|41|你既看見像的腳和腳趾頭，一半是陶匠的泥，一半是鐵，那國將來也必分裂。你既看見鐵和泥攙雜，那國也必有鐵的力量。
DAN|2|42|那腳趾頭既是半鐵半泥，那國也必半強半弱。
DAN|2|43|你既看見鐵和泥攙雜，他們必有混雜的後裔，卻不能彼此相合，正如鐵和泥不能相合。
DAN|2|44|當諸王在位的時候，天上的上帝必另立一個永不敗壞的國度，這國度必不歸給其他百姓，卻要打碎滅絕所有的國度，存立到永遠。
DAN|2|45|你既看見非人手鑿出來的一塊石頭從山而出，打碎鐵、銅、泥、銀、金，那就是至大的上帝把將來要發生的事給王指明。這夢是確實的，這解釋也是準確的。」
DAN|2|46|當時， 尼布甲尼撒 王臉伏於地，向 但以理 下拜，並且吩咐人給他奉上供物和香。
DAN|2|47|王對 但以理 說：「你既能講明這奧祕，你們的上帝誠然是萬神之神、萬王之主，是奧祕的啟示者。」
DAN|2|48|於是王使 但以理 高升，賞賜他極多的禮物，派他管理 巴比倫 全省，又立他為總理，掌管 巴比倫 所有的智慧人。
DAN|2|49|但以理 求王，王就派 沙得拉 、 米煞 、 亞伯尼歌 管理 巴比倫 省的事務，只是 但以理 仍在朝中侍立。
DAN|3|1|尼布甲尼撒 王造了一個金像，高六十肘，寬六肘，立在 巴比倫 省的 杜拉 平原。
DAN|3|2|尼布甲尼撒 王差人將總督、欽差、省長、參謀、財務、法官、地方官和各省的官員都召了來，為 尼布甲尼撒 王所立的像行開光禮。
DAN|3|3|於是總督、欽差、省長、參謀、財務、法官、地方官和各省的官員都聚集，站在 尼布甲尼撒 所立的像前，要為 尼布甲尼撒 王所立的像行開光禮。
DAN|3|4|那時傳令的大聲呼叫說：「各方、各國、各族 的人哪，有命令傳給你們：
DAN|3|5|你們一聽見角、號、琴、瑟、三角琴、鼓和各樣樂器的聲音，就當俯伏，拜 尼布甲尼撒 王所立的金像。
DAN|3|6|凡不俯伏下拜的，必立刻扔在烈火的窯中。」
DAN|3|7|因此百姓一聽見角、號、琴、瑟、三角琴 和各樣樂器的聲音，各方、各國、各族的人就都俯伏，拜 尼布甲尼撒 王所立的金像。
DAN|3|8|在那時，有幾個 迦勒底 人進前來控告 猶大 人。
DAN|3|9|他們對 尼布甲尼撒 王說：「願王萬歲！
DAN|3|10|你，王啊，你曾降旨，凡聽見角、號、琴、瑟、三角琴、鼓和各樣樂器聲音的，都當俯伏拜這金像。
DAN|3|11|凡不俯伏下拜的，必扔在烈火的窯中。
DAN|3|12|現在有幾個 猶大 人，就是王所派管理 巴比倫 省事務的 沙得拉 、 米煞 、 亞伯尼歌 ；王啊，這些人不理你的諭旨，不事奉你的神明，也不拜你所立的金像。」
DAN|3|13|當時， 尼布甲尼撒 大發烈怒，命令把 沙得拉 、 米煞 、 亞伯尼歌 帶過來；他們就把這幾個人帶到王面前。
DAN|3|14|尼布甲尼撒 對他們說：「 沙得拉 、 米煞 、 亞伯尼歌 ，你們不事奉我的神明，不拜我所立的金像，是真的嗎？
DAN|3|15|現在，你們若準備好，一聽見角、號、琴、瑟、三角琴、鼓和各樣樂器的聲音，就俯伏拜我所造的像；若不下拜，必立刻扔在烈火的窯中，有哪一個神明能救你們脫離我的手呢？」
DAN|3|16|沙得拉 、 米煞 、 亞伯尼歌 對王說：「 尼布甲尼撒 啊，這件事我們不必回答你，
DAN|3|17|即便如此，我們所事奉的上帝能將我們從烈火的窯中救出來。王啊，他必救我們脫離你的手；
DAN|3|18|即或不然，王啊，你當知道，我們絕不事奉你的神明，也不拜你所立的金像。」
DAN|3|19|當時， 尼布甲尼撒 怒氣填胸，向 沙得拉 、 米煞 、 亞伯尼歌 變了臉色，命令把窯燒熱，比平常熱七倍；
DAN|3|20|又命令他軍中的幾個壯士，把 沙得拉 、 米煞 、 亞伯尼歌 捆起來，扔在烈火的窯中。
DAN|3|21|這三人穿著內袍、外衣、頭巾和其他的衣服，被捆起來扔在烈火的窯中。
DAN|3|22|因為王的命令緊急，窯又非常熱，那抬 沙得拉 、 米煞 、 亞伯尼歌 的人都被火焰燒死。
DAN|3|23|但是這三個人， 沙得拉 、 米煞 、 亞伯尼歌 被捆綁著，掉進烈火的窯中。
DAN|3|24|那時， 尼布甲尼撒 王驚奇，急忙站起來，對謀士說：「我們捆起來扔在火裏的不是三個人嗎？」他們回答王說：「王啊，是的。」
DAN|3|25|王說：「看哪，我看見有四個人，並沒有捆綁，在火中行走，也沒有受傷；那第四個的相貌好像神明的兒子。」
DAN|3|26|於是 尼布甲尼撒 靠近烈火窯門，說：「至高上帝的僕人 沙得拉 、 米煞 、 亞伯尼歌 ，出來，來吧！」 沙得拉 、 米煞 、 亞伯尼歌 就從火中出來。
DAN|3|27|那些總督、欽差、省長和王的謀士一同聚集來看這三個人，見火不能傷他們的身體，頭髮沒有燒焦，衣裳也沒有變色，都沒有火燒過的氣味。
DAN|3|28|尼布甲尼撒 說：「 沙得拉 、 米煞 、 亞伯尼歌 的上帝是應當稱頌的！他差遣使者救護倚靠他的僕人，他們不遵王的命令，甚至捨身，在他們上帝以外不肯事奉敬拜別神。
DAN|3|29|現在我降旨，無論何方、何國、何族，凡有人毀謗 沙得拉 、 米煞 、 亞伯尼歌 的上帝，他必被凌遲，他的房屋必成糞堆，因為沒有別神能像這樣施行拯救。」
DAN|3|30|那時王在 巴比倫 省使 沙得拉 、 米煞 、 亞伯尼歌 高升。
DAN|4|1|尼布甲尼撒 王對住在全地各方、各國、各族的人說：「願你們大享平安！
DAN|4|2|我樂意宣揚至高上帝向我所行的神蹟奇事。
DAN|4|3|他的神蹟何其大！ 他的奇事何其盛！ 他的國度存到永遠； 他的權柄存到萬代！
DAN|4|4|「我－ 尼布甲尼撒 安居在家中，在宮裏享受榮華。
DAN|4|5|我做了一個夢，使我懼怕。我在床上的意念和腦中的異象，使我驚惶。
DAN|4|6|因此我降旨召 巴比倫 的智慧人全都到我面前，要他們將夢的解釋告訴我。
DAN|4|7|於是那些術士、巫師、 迦勒底 人、觀兆的都進來，我將那夢告訴他們，他們卻不能把夢的解釋告訴我。
DAN|4|8|最後， 但以理 ，就是按照我神明的名字稱為 伯提沙撒 的，來到我面前，他裏頭有神聖神明的靈，我將夢告訴他：
DAN|4|9|『術士的領袖 伯提沙撒 啊，我知道你裏頭有神聖神明的靈，甚麼奧祕都不能為難你。現在你要把我夢中所見的異象和夢的解釋告訴我 。』
DAN|4|10|「我在床上腦中的異象是這樣：我觀看，看哪，大地中間有一棵樹，極其高大。
DAN|4|11|那樹漸長，而且茁壯，高得頂天，從地極都能看見，
DAN|4|12|葉子華美，果子甚多，可作所有動物的食物；野地的走獸臥在蔭下，天空的飛鳥宿在枝上，凡有血肉的都從這樹得食物。
DAN|4|13|「我觀看，我在床上腦中的異象是這樣，看哪，有守望者，就是神聖的一位，從天而降，
DAN|4|14|大聲呼叫說：『砍倒這樹！砍下枝子！拔掉葉子！拋散果子！使走獸逃離樹下，飛鳥躲開樹枝。
DAN|4|15|樹的殘幹卻要留在地裏，在田野的青草中用鐵圈和銅圈套住。任他讓天上的露水滴濕，和地上的走獸一同吃草，
DAN|4|16|使他的心改變，不再是人的心，而給他一個獸心，使他經過七個時期 。
DAN|4|17|這是眾守望者所發的命令，是眾聖者所作的決定，好叫世人知道至高者在人的國中掌權，要將國賜給誰就賜給誰，並且立極卑微的人執掌國權。』
DAN|4|18|「這是我－ 尼布甲尼撒 王所做的夢。 伯提沙撒 啊，你要說明這夢的解釋；我國中所有的智慧人都不能把夢的解釋告訴我，惟獨你能，因你裏頭有神聖神明的靈。」
DAN|4|19|於是稱為 伯提沙撒 的 但以理 驚駭片時，心意驚惶。王說：「 伯提沙撒 啊，不要因夢和夢的解釋驚惶。」 伯提沙撒 回答說：「我主啊，願這夢歸給恨惡你的人，這夢的解釋歸給你的敵人。
DAN|4|20|你所見的樹漸長，而且茁壯，高得頂天，全地都能看見，
DAN|4|21|葉子華美，果子甚多，可作所有動物的食物；野地的走獸住在其下，天空的飛鳥宿在枝上。
DAN|4|22|「王啊，這成長又茁壯的樹就是你。你的威勢成長及於天，你的權柄達到地極。
DAN|4|23|王既看見一位神聖的守望者從天而降，說：『將這樹砍倒毀壞，樹的殘幹卻要留在地裏，在田野的青草中用鐵圈和銅圈套住。任他讓天上的露水滴濕，與野地的走獸一同吃草，直到經過七個時期。』
DAN|4|24|「王啊，夢的解釋就是這樣：臨到我主我王的事是出於至高者的命令。
DAN|4|25|你必被趕出離開世人，與野地的走獸同住，吃草如牛，讓天上的露水滴濕，且要經過七個時期，直等到你知道至高者在人的國中掌權，要將國賜給誰就賜給誰。
DAN|4|26|這使樹的殘幹存留的命令，是要等你知道天在掌權，你的國必定歸你。
DAN|4|27|王啊，求你悅納我的諫言，以施行公義除去罪過，以憐憫窮人除掉罪惡，或者你的平安可以延長。」
DAN|4|28|這些事都臨到 尼布甲尼撒 王。
DAN|4|29|過了十二個月，他在 巴比倫 王宮頂上散步。
DAN|4|30|王說：「這大 巴比倫 豈不是我用大能大力建為首都，要顯示我威嚴的榮耀嗎？」
DAN|4|31|這話還在王口中的時候，有聲音從天降下，說：「 尼布甲尼撒 王啊，有話對你說，你的國離開你了。
DAN|4|32|你必被趕出離開世人，與野地的走獸同住，吃草如牛，且要經過七個時期；等你知道至高者在人的國中掌權，要將國賜給誰就賜給誰。」
DAN|4|33|當時這話就應驗在 尼布甲尼撒 身上，他被趕出離開世人，吃草如牛，身體被天上的露水滴濕，頭髮長得像鷹的羽毛，指甲長得像鳥爪。
DAN|4|34|「時候到了，我－ 尼布甲尼撒 舉目望天，我的知識復歸於我，我就稱頌至高者，讚美尊敬活到永遠的上帝。 他的權柄存到永遠， 他的國度存到萬代。
DAN|4|35|地上所有的居民都算為虛無； 在天上萬軍和地上居民中， 他都憑自己的旨意行事。 無人能攔住他的手， 或問他說，你在做甚麼呢？
DAN|4|36|「那時，我的知識復歸於我，威嚴和光榮也復歸於我，使我的國度得榮耀，我的謀士和大臣也來朝見我。我又重建我的國度，更大的權勢加添在我身上。
DAN|4|37|現在我－ 尼布甲尼撒 讚美、尊崇、恭敬天上的王，因為他所行的全都信實，他所做的盡都公平。那行事驕傲的，他能降為卑。」
DAN|5|1|伯沙撒 王為他的一千大臣擺設盛筵，與這一千人飲酒。
DAN|5|2|伯沙撒 在歡飲之間，吩咐人將他父 尼布甲尼撒 從 耶路撒冷 聖殿所擄掠的金銀器皿拿來，好使王與大臣、王后、妃嬪用這器皿飲酒。
DAN|5|3|於是他們把聖殿，就是 耶路撒冷 上帝殿中所擄掠的金器皿拿來，王和大臣、王后、妃嬪就用這器皿飲酒。
DAN|5|4|他們飲酒，讚美金、銀、銅、鐵、木、石造的神明。
DAN|5|5|當時，忽然有人的指頭出現，在燈臺對面王宮粉刷的牆上寫字。王看見寫字的指頭，
DAN|5|6|就變了臉色，心意驚惶，腰骨好像脫節，雙膝彼此相碰，
DAN|5|7|大聲吩咐將巫師、 迦勒底 人和觀兆的領進來。王對 巴比倫 的智慧人說：「誰能讀這文字，並且向我講解它的意思，他必身穿紫袍，項帶金鏈，在我國中位列第三。」
DAN|5|8|於是王所有的智慧人都進前來，他們卻不能讀那文字，也不能為王講解它的意思。
DAN|5|9|伯沙撒 王就甚驚惶，臉色改變，他的大臣也都困惑。
DAN|5|10|太后 因王和他大臣所說的話，就進入宴會廳，說：「願王萬歲！你的心不要驚惶，臉不要變色。
DAN|5|11|在你國中有一人，他裏頭有神聖神明的靈，你父在世的日子，這人心中光明，又有聰明智慧，好像神明的智慧。你父 尼布甲尼撒 王，就是王的父，曾立他為術士、巫師、 迦勒底 人和觀兆者的領袖，
DAN|5|12|都因他有美好的靈性，又有知識聰明，能解夢，釋謎語，解疑惑。這人名叫 但以理 ， 尼布甲尼撒 王又稱他為 伯提沙撒 ，現在可以召他來，他必解明這意思。」
DAN|5|13|於是 但以理 被領到王面前。王問 但以理 說：「你就是我父王從 猶大 帶來、被擄的 猶大 人 但以理 嗎？
DAN|5|14|我聽說你裏頭有神明的靈，心中有光，又有聰明和高超的智慧。
DAN|5|15|現在智慧人和巫師都被帶到我面前，要叫他們讀這文字，為我講解它的意思；無奈他們都不能講解它的意思。
DAN|5|16|我聽說你能講解，能解疑惑；現在你若能讀這文字，為我講解它的意思，就必身穿紫袍，項戴金鏈，在我國中位列第三。」
DAN|5|17|但以理 回答王說：「你的禮物可以歸你自己，你的賞賜可以歸給別人；我卻要為王讀這文字，講解它的意思。
DAN|5|18|你，王啊，至高的上帝曾將國度、大權、榮耀、威嚴賜給你父 尼布甲尼撒 ；
DAN|5|19|因上帝所賜給他的大權，各方、各國、各族的人都在他面前恐懼戰兢，因他要殺就殺，要人活就活，要升就升，要降就降。
DAN|5|20|但他的心高傲，靈也剛愎，以致行事狂傲，就被革去國度的王位，奪走榮耀。
DAN|5|21|他被趕出離開世人，他的心變為獸心，與野驢同住，吃草如牛，身體被天上的露水滴濕，直到他知道，至高的上帝在人的國中掌權，憑自己的旨意立人治國。
DAN|5|22|伯沙撒 啊，你是他的兒子 ，你雖知道這一切，卻不謙卑自己，
DAN|5|23|竟向天上的主自高，差人將他殿中的器皿拿到你面前，你和大臣、王后、妃嬪用這器皿飲酒。你又讚美那不能看、不能聽、無知無識，用金、銀、銅、鐵、木、石造的神明，沒有將榮耀歸與那手中掌管你氣息，管理你一切行動的上帝。
DAN|5|24|於是從他那裏顯出指頭寫這文字。
DAN|5|25|「所寫的文字是：『彌尼，彌尼，提客勒，烏法珥新 。』
DAN|5|26|解釋是這樣：彌尼就是上帝數算你國的年日到此完畢。
DAN|5|27|提客勒就是你被秤在天平上，秤出你的虧欠來。
DAN|5|28|毗勒斯 就是你的國要分裂，歸給 瑪代 人和 波斯 人。」
DAN|5|29|於是 伯沙撒 下令，人就把紫袍給 但以理 穿上，把金鏈給他戴在頸項上，又傳令使他在國中位列第三。
DAN|5|30|當夜， 迦勒底 王 伯沙撒 被殺。
DAN|5|31|瑪代 人 大流士 年六十二歲，取了 迦勒底 國。
DAN|6|1|大流士 隨心所願，立了一百二十個總督，治理全國，
DAN|6|2|又在他們以上立總長三人， 但以理 也在其中；使總督在他們三人面前呈報，免得王受虧損。
DAN|6|3|這 但以理 因有卓越的靈性，超乎其餘的總長和總督，王想立他治理全國。
DAN|6|4|那時，總長和總督在治國的事務上尋找 但以理 的把柄，為要控告他；只是找不到任何的把柄和過失，因他忠心辦事，毫無錯誤過失。
DAN|6|5|那些人就說：「我們要找 但以理 的把柄，若不從他上帝的律法中下手，就尋不著。」
DAN|6|6|於是，總長和總督紛紛聚集來見王，說：「 大流士 王萬歲！
DAN|6|7|國中的總長、欽差、總督、謀士和省長彼此商議，求王下旨，立一條禁令，三十天之內，不拘何人，若在王以外，或向神明或向人求甚麼，就必扔在獅子坑中。
DAN|6|8|王啊，現在求你立這禁令，在這文件上簽署，使它不能更改；照 瑪代 人和 波斯 人的例，絕不更動。」
DAN|6|9|於是 大流士 王在這禁令的文件上簽署。
DAN|6|10|但以理 知道這文件已經簽署，就進自己的家，他家樓上的窗戶開向 耶路撒冷 。他一天三次，雙膝跪著，在他的上帝面前禱告感謝，像平常一樣。
DAN|6|11|於是，那些人紛紛聚集，發現 但以理 在他上帝面前祈禱懇求。
DAN|6|12|他們就進到王面前，向王提及禁令，說：「三十天之內不拘何人，若在王以外，或向神明或向人求甚麼，必被扔在獅子坑中，王不是在這禁令上簽署了嗎？」王回答說：「確有這事，照 瑪代 人和 波斯 人的例是不可更改的。」
DAN|6|13|他們對王說：「王啊，那被擄的 猶大 人 但以理 不理會你，也不遵守你簽署的禁令，竟一天三次祈禱。」
DAN|6|14|王聽見這話，就甚愁煩，一心要救 但以理 ，直到日落的時候，他還在籌劃解救他。
DAN|6|15|那些人就紛紛聚集到王那裏，對王說：「王啊，當知道 瑪代 人和 波斯 人有例，凡王所立的禁令和律例都不可更改。」
DAN|6|16|於是王下令，人就把 但以理 帶來，扔在獅子坑中。王對 但以理 說：「你經常事奉的上帝，他必拯救你。」
DAN|6|17|有人搬來一塊石頭放在坑口，王用自己的璽和大臣的印，封閉那坑，使懲辦 但以理 的事絕不更改。
DAN|6|18|王回到宮裏，終夜禁食，不讓人帶樂器 到他面前，他也失眠了。
DAN|6|19|次日黎明，王起來，急忙往獅子坑那裏去，
DAN|6|20|臨近坑邊，哀聲呼叫 但以理 。王對 但以理 說：「永生上帝的僕人 但以理 啊，你經常事奉的上帝能救你脫離獅子嗎？」
DAN|6|21|但以理 對王說：「願王萬歲！
DAN|6|22|我的上帝差遣使者封住獅子的口，叫獅子不傷我，因我在上帝面前無辜。王啊，在你面前我也沒有做過任何虧損的事。」
DAN|6|23|王因此就甚喜樂，吩咐把 但以理 從坑裏拉上來。於是 但以理 從坑裏被拉上來，身上毫無損傷，因為他信靠他的上帝。
DAN|6|24|王下令，把那些控告 但以理 的人和他們的妻子兒女都帶來，扔在獅子坑中。他們還沒有到坑底，獅子就制伏他們，咬碎他們的骨頭。
DAN|6|25|於是， 大流士 王傳旨給住在全地各方、各國、各族的人說：「願你們大享平安！
DAN|6|26|現在我降旨，我所統轄全國的人民，都要在 但以理 的上帝面前戰兢畏懼。 因為他是活的上帝， 永遠長存， 他的國度永不敗壞， 他的權柄永存無極！
DAN|6|27|他庇護，搭救， 在天上地下施行神蹟奇事， 救了 但以理 脫離獅子的口。」
DAN|6|28|如此，這 但以理 ，當 大流士 在位的時候和 波斯 的 居魯士 在位的時候，大享亨通。
DAN|7|1|巴比倫 王 伯沙撒 元年， 但以理 在床上做夢，腦中看見異象，就記錄這夢，述說其中的大意。
DAN|7|2|但以理 說： 我在夜間的異象中觀看，看哪，天上有四風，突然颳在大海之上。
DAN|7|3|有四隻巨獸從海裏上來，牠們各不相同：
DAN|7|4|頭一個像獅子，有鷹的翅膀；我正觀看的時候，牠的翅膀被拔去，牠從地上被扶起來，用兩腳站立，像人一樣，還給了牠人的心。
DAN|7|5|看哪，另有一獸如熊，就是第二獸，半身側立，口裏的牙齒中有三根獠牙 。有人吩咐這獸說：「起來，吞吃許多的肉。」
DAN|7|6|其後，我觀看，看哪，另有一獸如豹，背上有四個鳥的翅膀；這獸有四個頭，還給了牠權柄。
DAN|7|7|其後，我在夜間的異象中觀看，看哪，第四獸可怕可懼，極其強壯，有大鐵牙，吞吃嚼碎，剩下的用腳踐踏。這獸與前面所有的獸不同，牠有十隻角。
DAN|7|8|我正思考這些角的時候，看哪，其中又長出另一隻小角；先前的角中有三隻角在它面前連根被拔出。看哪，這角有眼，像人的眼，有口說誇大的話。
DAN|7|9|我正觀看的時候， 有寶座設立， 上面坐著亙古常在者。 他的衣服潔白如雪， 頭髮如純淨的羊毛。 寶座是火焰， 其輪為烈火。
DAN|7|10|有火如河湧出， 從他面前流出來； 事奉他的有千千， 在他面前侍立的有萬萬； 他坐著要行審判 ， 案卷都展開了。
DAN|7|11|於是我觀看，因這角說誇大的話，我正觀看的時候，那獸被殺，身體被毀，扔在火中焚燒。
DAN|7|12|其餘的獸，權柄都被奪去，生命卻得以延續，直到所定的時候和日期。
DAN|7|13|我在夜間的異象中觀看， 看哪，有一位像人子的， 駕著天上的雲而來， 被領到亙古常在者面前。
DAN|7|14|他得了權柄、榮耀、國度， 使各方、各國、各族的人都事奉他。 他的權柄是永遠的，不能廢去， 他的國度必不敗壞。
DAN|7|15|至於我－ 但以理 ，我的靈在我裏面憂傷，我腦中的異象使我驚惶。
DAN|7|16|我走近其中一位侍立者，問他這一切的實情。他就告訴我，使我知道這事的解釋：
DAN|7|17|這四隻巨獸就是將要在世上興起的四個王 。
DAN|7|18|然而，至高者的眾聖者必要得到這國度，並且擁有它，直到永遠，永永遠遠。
DAN|7|19|於是我想要更清楚知道第四獸的實情，牠與一切的獸不同，甚是可怕，有鐵牙銅爪，吞吃嚼碎，剩下的用腳踐踏；
DAN|7|20|頭上有十隻角和那另長出的一角，三隻角在這角面前掉落；這角有眼，有口說誇大的話，形狀比牠的同類更強。
DAN|7|21|我觀看，這角與眾聖者爭戰，勝了他們，
DAN|7|22|直到亙古常在者來到，為至高者的眾聖者伸冤，眾聖者得到國度的時候就到了。
DAN|7|23|那侍立者這樣說： 第四獸就是世上要興起的第四國， 與其他各國不同， 它要併吞全地， 並且踐踏嚼碎。
DAN|7|24|至於那十隻角，就是從這國中興起的十個王； 後來又興起另一王， 與先前的不相同， 他要制伏三個王。
DAN|7|25|他說話抵擋至高者， 折磨至高者的眾聖者， 又改變節期和律法。 眾聖者要交在他手中一年 、兩年、又半年。
DAN|7|26|然而，他坐著要行審判； 他的權柄要被奪去， 毀壞，滅絕，一直到底。
DAN|7|27|國度、權柄和天下諸國的大權 必賜給至高者的眾聖民。 他的國是永遠的國， 所有掌權的都必事奉他，順從他。
DAN|7|28|這事到此結束。我－ 但以理 因這些念頭甚是驚惶，臉色也變了，卻將這事記在心裏。
DAN|8|1|伯沙撒 王在位第三年，有異象向我－ 但以理 顯現，是在先前所見的異象之後。
DAN|8|2|我在異象中觀看，見自己在 以攔 省 書珊 的城堡中；我在異象中又見自己在 烏萊河 邊。
DAN|8|3|我舉目觀看，看哪，有一隻公綿羊站在河邊，牠有兩隻角，這兩角都高，一角高過另一角，後長出來的比較高。
DAN|8|4|我見那公綿羊向西、向北、向南牴撞，沒有任何獸在牠面前站立得住，沒有能逃脫牠手的；牠任意而行，自高自大。
DAN|8|5|我正思想的時候，看哪，有一隻公山羊從西而來，遍行全地，腳不著地。這山羊兩眼當中有一隻顯眼的角。
DAN|8|6|牠往我先前所見、站在河邊、有雙角的公綿羊那裏，以猛烈的怒氣向牠直闖。
DAN|8|7|我見公山羊靠近公綿羊，向牠發怒，攻擊牠，折斷牠的兩角。公綿羊在公山羊面前站立不住；牠把公綿羊撞倒在地，用腳踐踏，沒有能救公綿羊脫離牠手的。
DAN|8|8|這公山羊長得極其高大，正強壯的時候，那大角折斷了，從角的下面向天的四方 長出四隻顯眼的角來。
DAN|8|9|從四角中的一角又長出另一隻小角，向南、向東、向佳美之地，日漸壯大。
DAN|8|10|牠漸壯大，高及諸天萬象，把一些天象和星辰摔落在地，用腳踐踏。
DAN|8|11|牠自高自大 ，自以為高及萬象之君，牠除掉經常獻給君的祭，毀壞君的聖所。
DAN|8|12|因罪過的緣故，有軍隊和經常獻的祭交給牠。牠把真理拋在地上，任意而行 ，無往不利。
DAN|8|13|我聽見有一位聖者說話，又有一位聖者向那說話的聖者說：「這經常獻的祭、帶來荒涼的罪過、聖所與軍隊被踐踏的異象，要持續到幾時呢？」
DAN|8|14|他對我 說：「要到二千三百日，聖所就必潔淨 。」
DAN|8|15|我－ 但以理 見了這異象，想要明白其中的意思。看哪，有一位形狀像人的站在我面前。
DAN|8|16|我聽見 烏萊河 中有人聲呼叫說：「 加百列 啊，要使這人明白這異象。」
DAN|8|17|他就來到我所站的地方。他一來，我就驚慌，臉伏於地。他對我說：「人子啊，你要明白，因為這是關乎末後時期的異象。」
DAN|8|18|他對我說話的時候，我正沉睡，臉伏於地。他就摸我，扶我站起來。
DAN|8|19|他說：「看哪，我要指示你惱怒結束的時候必成的事，因為這是關乎末後指定的時期。
DAN|8|20|你所看見那有雙角的公綿羊就是 瑪代 王和 波斯 王。
DAN|8|21|那公山羊就是 希臘 王；兩眼當中的大角就是第一個王。
DAN|8|22|至於角折斷了，又從角的下面長出四隻角，意思就是有四個國要從這國興起，只是權勢都不及它。
DAN|8|23|這四國末期，惡貫滿盈的時候，必有一王興起，面貌兇惡，詭計多端。
DAN|8|24|他的權柄極大，卻不是因自己的能力；他要施行驚人的毀滅，無往不利，任意而行，又要毀滅強有力的人和眾聖民。
DAN|8|25|他用權術使手中的詭計成功；他的心自高自大，趁人無備的時候毀滅多人。他又起來攻擊萬君之君，至終卻非因人的手而遭毀滅。
DAN|8|26|所說二千三百日 的異象是真的，但你要將這異象封住，因為它關乎未來許多的日子。」
DAN|8|27|於是我－ 但以理 昏倒，病了數日，然後起來辦理王的事務。我因這異象驚駭不已，但還是不能了解。
DAN|9|1|瑪代 族 亞哈隨魯 的兒子 大流士 被立為王，統治 迦勒底 國元年，
DAN|9|2|就是他在位第一年，我－ 但以理 從書上得知，耶和華的話臨到 耶利米 先知，論 耶路撒冷 荒涼期滿的年數為七十年。
DAN|9|3|我面向主上帝，禁食，披麻蒙灰，懇切禱告祈求。
DAN|9|4|我向耶和華－我的上帝祈禱、認罪，說：「主啊，你是大而可畏的上帝，向愛主、守主誡命的人守約施慈愛。
DAN|9|5|我們犯罪作惡，行惡叛逆，偏離你的誡命典章，
DAN|9|6|沒有聽從你僕人眾先知奉你的名向我們君王、官長、祖先和這地所有百姓所說的話。
DAN|9|7|主啊，你是公義的，但我們 猶大 人和 耶路撒冷 的居民，並你所趕到各國的 以色列 眾人，不論遠近，因為背叛了你，臉上蒙羞，正如今日一樣。
DAN|9|8|耶和華啊，我們和我們的君王、官長、祖先因得罪了你，臉上就都蒙羞。
DAN|9|9|主－我們的上帝是憐憫饒恕人的，我們卻違背了他，
DAN|9|10|沒有聽從耶和華－我們上帝的話，沒有遵行他藉僕人眾先知向我們頒佈的律法。
DAN|9|11|以色列 眾人都犯了你的律法，偏離、不聽從你的話；因此，你僕人 摩西 律法上所寫的詛咒和誓言傾倒在我們身上，因我們得罪了上帝。
DAN|9|12|上帝使大災禍臨到我們，實現了警戒我們和審判我們官長的話；原來 耶路撒冷 所遭遇的災禍是普天之下未曾有過的。
DAN|9|13|這一切災禍臨到我們，是照 摩西 律法上所寫的，我們卻沒有求耶和華－我們上帝的恩惠，使我們回轉離開罪孽，明白你的真理。
DAN|9|14|所以耶和華特意使這災禍臨到我們，耶和華－我們的上帝在他所行的事上都是公義的；我們並沒有聽從他的話。
DAN|9|15|主－我們的上帝啊，你曾用大能的手領你的子民出 埃及 地，使自己得了名聲，正如今日一樣，現在，我們犯了罪，作了惡。
DAN|9|16|主啊，求你按你豐盛的公義，使你的怒氣和憤怒轉離你的城 耶路撒冷 ，就是你的聖山。因我們的罪惡和我們祖先的罪孽， 耶路撒冷 和你的子民被四圍的人羞辱。
DAN|9|17|我們的上帝啊，現在求你垂聽你僕人的祈禱懇求，為你自己的緣故使你的臉向荒涼的聖所發光。
DAN|9|18|我的上帝啊，求你側耳而聽，睜眼而看，眷顧我們那荒涼之地和稱為你名下的城。我們在你面前懇求，不是因自己的義，而是因你豐富的憐憫。
DAN|9|19|主啊，求你垂聽！主啊，求你赦免！主啊，求你側耳，求你實行！為你自己的緣故不要遲延。我的上帝啊，因這城和這民都是稱為你名下的。」
DAN|9|20|我正說話、禱告，承認我的罪和我百姓 以色列 的罪，為我上帝的聖山，在耶和華－我的上帝面前懇求；
DAN|9|21|我正在禱告中說話，先前在異象中所見的那位 加百列 ，約在獻晚祭的時候迅速飛到我這裏來。
DAN|9|22|他指教我說 ：「 但以理 啊，現在我來要使你有智慧，有聰明。
DAN|9|23|你剛開始懇求的時候，就有命令發出。現在我來告訴你，因你是蒙愛的；所以你要思想這事，明白這異象。
DAN|9|24|「為你百姓和你聖城，已經定了七十個七，要止住罪過，除淨罪惡，贖盡罪孽，引進永恆的公義，封住異象和預言，並膏至聖所 。
DAN|9|25|你當知道，當明白，從發出命令恢復並重建 耶路撒冷 ，直到受膏的君出現，必有七個七和六十二個七。 耶路撒冷城 連街帶濠都必在艱難中恢復並重建。
DAN|9|26|過了六十二個七，那受膏者 被剪除，一無所有；必有一王的百姓來毀滅這城和聖所，它的結局 必如洪水沖沒。必有戰爭，一直到末了，荒涼的事已經定了。
DAN|9|27|在一七之期，他必與許多人堅立盟約；一七之半，他必使獻祭與供獻止息。那施行毀滅的可憎之物必立在聖殿裏 ，直到所定的結局傾倒在那行毀滅者的身上。」
DAN|10|1|波斯 王 居魯士 第三年，有話指示那稱為 伯提沙撒 的 但以理 。這話是確實的，指著大戰爭； 但以理 明白這話，明白這異象。
DAN|10|2|那時，我－ 但以理 悲傷了三個七日；
DAN|10|3|美味我沒有吃，酒和肉沒有入我的口，也沒有用油抹我的身，直到滿了三個七日。
DAN|10|4|正月二十四日，我在 大河 ，就是 底格里斯河 邊，
DAN|10|5|舉目觀看，看哪，有一人身穿細麻衣，腰束 烏法 的純金腰帶。
DAN|10|6|他的身體如水蒼玉，面貌如閃電，眼目如火把，手臂和腳如明亮的銅，說話的聲音像眾人的聲音。
DAN|10|7|我－ 但以理 一人看見這異象，跟我一起的人沒有看見，卻有極大的戰兢落在他們身上，他們就逃跑躲避，
DAN|10|8|只剩下我一人。我看見這大異象就渾身無力，面容變色，毫無氣力。
DAN|10|9|我聽見他說話的聲音；一聽見他說話的聲音，我就沉睡，臉伏於地。
DAN|10|10|看哪，有一隻手摸我，使我膝蓋和手掌戰抖。
DAN|10|11|他對我說：「蒙愛的 但以理 啊，要思想我對你所說的話，只管站起來，因為我現在奉差遣來到你這裏。」他對我說這話，我就戰戰兢兢地站起來。
DAN|10|12|他說：「 但以理 啊，不要懼怕！因為自從第一日你立志要明白，又在你上帝面前刻苦自己，你的話已蒙應允；我就是因你的話而來。
DAN|10|13|但 波斯 國的領袖攔阻了我二十一天。看哪，天使長 中的一位 米迦勒 來幫助我，因為我被留在 波斯 諸王那裏。
DAN|10|14|現在我來，要使你明白你百姓日後必遭遇的事，因為這異象關乎未來的日子。」
DAN|10|15|他向我這樣說，我就臉面朝地，啞口無聲。
DAN|10|16|看哪，有一位形狀像人的，摸我的嘴唇，我就開口說話，向那站在我面前的說：「我主啊，因這異象使我感到劇痛，毫無氣力。
DAN|10|17|我主的僕人怎能跟我主說話呢？我現在渾身無力，毫無氣息。」
DAN|10|18|有一位形狀像人的再一次摸我，使我有力量。
DAN|10|19|他說：「蒙愛的人哪，不要懼怕，願你平安！你要剛強！要剛強！ 」他一對我說話，我就覺得有力量，說：「我主請說，因你使我有力量。」
DAN|10|20|他說：「你知道我為甚麼到你這裏來嗎？現在我要回去與 波斯 的領袖爭戰，我去了之後，看哪， 希臘 的領袖必來。
DAN|10|21|但我要將那記錄在真理之書上的話告訴你。除了你們的天使 米迦勒 之外，沒有人幫助我抵擋他們。」
DAN|11|1|「至於我，當 瑪代 的 大流士 元年，我曾起來扶助 米迦勒 ，使他堅強。
DAN|11|2|現在我要指示你確實的事。」 「看哪， 波斯 還有三個王要興起，第四王必富足遠勝諸王。他因富足成為強盛，就煽動各國攻擊 希臘 國。
DAN|11|3|必有一個勇敢的王興起，執掌大權，隨意而行。
DAN|11|4|他正興起的時候，他的國必瓦解，向天的四方 裂開，卻不歸他的後裔，也不如他當年統治的權威；他的國必被拔出，歸給他後裔之外的人。
DAN|11|5|「南方的王必強盛，他的將帥中必有一個比他更強，執掌權柄，權柄甚大。
DAN|11|6|過了幾年，他們必結盟，南方王的女兒必來到北方王那裏，使約生效；但這女子不能保留實力，王的力量 也未能存留。這女子、帶她來的、生她的 和當時扶助她的必被殺害 。
DAN|11|7|但從這女子的本家必另有一子 接續王位，他要率領軍隊進入北方王的堡壘，攻擊他們，而且得勝，
DAN|11|8|把他們的神像和鑄成的偶像，與金銀寶器都擄掠到 埃及 去。數年之內，他不去攻擊北方的王。
DAN|11|9|北方的王必侵入南方王的國土，但卻要撤回本地。
DAN|11|10|「北方王的兒子們必動干戈，招聚許多軍兵。他要前進，如洪水氾濫；要再度爭戰，直搗南方王的堡壘。
DAN|11|11|南方王必發烈怒，出來與北方王爭戰，擺列大軍；北方王的軍兵必敗在南方王的手下。
DAN|11|12|這大軍既被掃蕩，南方王的心就自高；他雖使萬人仆倒，卻不能保持勝利。
DAN|11|13|「北方王要再度擺列大軍，比先前更多。過了幾年，他必率領大軍，帶極多的裝備而來。
DAN|11|14|那時，必有許多人起來攻擊南方王，並且你百姓中的殘暴人要興起，應驗異象，他們卻要敗亡。
DAN|11|15|北方王必來建土堆攻取堅固城，南方的軍兵抵擋不住，就是精選的部隊也無力抵擋；
DAN|11|16|前來攻擊南方王的必任意而行，無人在北方王面前站立得住。他要站在那佳美之地，用手施行毀滅。
DAN|11|17|「他必定意傾全國之力而來，與南方王訂約，把自己的女兒 給南方王為妻，企圖敗壞他的國度。這計謀卻未得逞，自己也得不到好處。
DAN|11|18|其後北方王必轉頭，奪取許多海島。但有一將帥除掉北方王對人的羞辱，並且使羞辱歸到他自己身上。
DAN|11|19|他必轉頭回到本地的堡壘，卻要絆跌仆倒，歸於無有。
DAN|11|20|「那時，有一人興起接續他的王位，他為了王國的榮華，差官員橫征暴斂。這王過不多時就死了，不是因怒氣 ，也不是因戰役。」
DAN|11|21|「後來，有一個卑鄙的人興起接續他的王位，人未曾將國的尊榮給他，他卻趁人無備的時候前來，用詭詐奪取政權。
DAN|11|22|勢如洪水般的軍兵在他面前被沖沒，遭擊潰；立約的領袖也是如此。
DAN|11|23|他與人結盟之後，卻行詭詐。跟隨他的人雖不多，他卻日漸強盛。
DAN|11|24|他趁人無備的時候，來到國中極肥沃之地，做他祖宗和祖宗的祖宗未曾做過的事，瓜分擄物、掠物和財寶，又策劃進攻堡壘；然而這都是暫時的。
DAN|11|25|「他必奮勇向前，率領大軍攻擊南方王；南方王以極強的大軍迎戰，卻抵擋不住，因為有人設計謀害南方王。
DAN|11|26|吃王餉的使王敗壞，王的軍隊必被沖沒，仆倒被殺的甚多。
DAN|11|27|至於這二王，他們心懷惡計，同席吃飯卻彼此說謊，但計謀不成，因為結局要在指定的時期來到。
DAN|11|28|北方王必帶許多財寶回本地，但他的心反對聖約；他恣意橫行，回到本地。
DAN|11|29|「到了指定的時期，他必返回，侵入南方。這一次卻不像前一次，
DAN|11|30|因為 基提 的戰船要來攻擊他，他就喪膽而退。他惱恨聖約，恣意橫行，要回來善待那些背棄聖約的人。
DAN|11|31|他要興兵，這兵必褻瀆聖所，就是堡壘，除掉經常獻的祭，設立那施行毀滅的可憎之物。
DAN|11|32|他必用巧言奉承違背聖約的惡人；惟獨認識上帝的子民必剛強行事。
DAN|11|33|民間的智慧人必訓誨許多人，然而在一段日子裏，他們必因刀劍、火燒、擄掠、搶奪而仆倒。
DAN|11|34|他們仆倒的時候，會得到少許援助，卻有許多人用詭詐加入他們。
DAN|11|35|智慧人中有些人仆倒，為要使他們受熬煉，成為潔淨、潔白，直到末了；因為還有一段日子才到所定的時期。
DAN|11|36|「王必任意而行，自高自大，超過所有的神明，又用荒謬的話攻擊萬神之神。他必行事亨通，直到主的憤怒結束，因為所定的事必然實現。
DAN|11|37|他不顧他祖宗的神明，也不顧婦女所仰慕的神明，任何神明他都不顧；因為他自大，高過一切，
DAN|11|38|以敬奉堡壘的神明取而代之，用金、銀、寶石和珍寶敬奉他祖宗所不認識的神明。
DAN|11|39|他靠外邦神明的幫助，攻破最堅固的堡壘。凡承認他的，他要給他們許多尊榮，使他們管轄許多人，又分封土地作為報償。
DAN|11|40|「到末了，南方王要與北方王交戰。北方王要用戰車、騎兵和許多戰船，勢如暴風來攻擊他，又要侵入列國，如洪水氾濫。
DAN|11|41|他要侵入那佳美之地，許多國就被傾覆 ，但 以東 人、 摩押 人和大半的 亞捫 人必逃離他的手。
DAN|11|42|他要伸手攻擊列國，連 埃及 地也不得逃脫。
DAN|11|43|他要掌管 埃及 的金銀財寶和各樣珍寶， 路比 人和 古實 人都跟從他的腳步。
DAN|11|44|但從東方和北方必有消息傳來擾亂他，他就大發烈怒出去，要將許多人殺滅淨盡。
DAN|11|45|他要在海和榮美的聖山之間搭起王宮的帳幕；然而他的結局到了，無人能幫助他。」
DAN|12|1|「那時，保佑你百姓的天使長 米迦勒 必站起來，並且有大艱難，自從有國以來直到此時，未曾有過這樣的事。那時，你的百姓凡記錄在冊上的，必得拯救。
DAN|12|2|睡在地裏塵埃中的必有多人醒過來；其中有得永生的，有受羞辱永遠被憎惡的。
DAN|12|3|智慧人要發光，如同天上的光；那領許多人歸於義的必發光如星，直到永永遠遠。
DAN|12|4|但以理 啊，你要隱藏這話，封閉這書，直到末時。必有許多人往來奔跑 ，知識 就必增長。」
DAN|12|5|我－ 但以理 觀看，看哪，另有兩個人站立：一個在河這邊，一個在河那邊。
DAN|12|6|其中一個對那在河水之上、穿細麻衣的說：「這奇異的事要到幾時才應驗呢？」
DAN|12|7|我聽見那在河水之上、穿細麻衣的，向天舉起左右手，指著那活到永遠的起誓說：「要到一年 、兩年，又半年，粉碎聖民力量結束的時候，這一切的事就要應驗。」
DAN|12|8|我聽了卻不明白，就說：「我主啊，這些事的結局是怎樣呢？」
DAN|12|9|他說：「 但以理 ，去吧！因為這話已經隱藏封閉，直到末時。
DAN|12|10|必有許多人使自己潔淨、潔白，且受熬煉；但惡人仍必行惡，沒有一個惡人明白，惟獨智慧人能明白。
DAN|12|11|從除掉經常獻的祭，設立那施行毀滅的可憎之物的時候起，必有一千二百九十日。
DAN|12|12|那等候，直到一千三百三十五日的有福了。
DAN|12|13|「至於你，你要去等候結局。你必安息，到了末期，你必起來，享受你的福分。」
