MIC|1|1|The word of the LORD that came to Micah of Moresheth during the reigns of Jotham, Ahaz and Hezekiah, kings of Judah-the vision he saw concerning Samaria and Jerusalem.
MIC|1|2|Hear, O peoples, all of you, listen, O earth and all who are in it, that the Sovereign LORD may witness against you, the Lord from his holy temple.
MIC|1|3|Look! The LORD is coming from his dwelling place; he comes down and treads the high places of the earth.
MIC|1|4|The mountains melt beneath him and the valleys split apart, like wax before the fire, like water rushing down a slope.
MIC|1|5|All this is because of Jacob's transgression, because of the sins of the house of Israel. What is Jacob's transgression? Is it not Samaria? What is Judah's high place? Is it not Jerusalem?
MIC|1|6|"Therefore I will make Samaria a heap of rubble, a place for planting vineyards. I will pour her stones into the valley and lay bare her foundations.
MIC|1|7|All her idols will be broken to pieces; all her temple gifts will be burned with fire; I will destroy all her images. Since she gathered her gifts from the wages of prostitutes, as the wages of prostitutes they will again be used."
MIC|1|8|Because of this I will weep and wail; I will go about barefoot and naked. I will howl like a jackal and moan like an owl.
MIC|1|9|For her wound is incurable; it has come to Judah. It has reached the very gate of my people, even to Jerusalem itself.
MIC|1|10|Tell it not in Gath; weep not at all. In Beth Ophrah roll in the dust.
MIC|1|11|Pass on in nakedness and shame, you who live in Shaphir. Those who live in Zaanan will not come out. Beth Ezel is in mourning; its protection is taken from you.
MIC|1|12|Those who live in Maroth writhe in pain, waiting for relief, because disaster has come from the LORD, even to the gate of Jerusalem.
MIC|1|13|You who live in Lachish, harness the team to the chariot. You were the beginning of sin to the Daughter of Zion, for the transgressions of Israel were found in you.
MIC|1|14|Therefore you will give parting gifts to Moresheth Gath. The town of Aczib will prove deceptive to the kings of Israel.
MIC|1|15|I will bring a conqueror against you who live in Mareshah. He who is the glory of Israel will come to Adullam.
MIC|1|16|Shave your heads in mourning for the children in whom you delight; make yourselves as bald as the vulture, for they will go from you into exile.
MIC|2|1|Woe to those who plan iniquity, to those who plot evil on their beds! At morning's light they carry it out because it is in their power to do it.
MIC|2|2|They covet fields and seize them, and houses, and take them. They defraud a man of his home, a fellowman of his inheritance.
MIC|2|3|Therefore, the LORD says: "I am planning disaster against this people, from which you cannot save yourselves. You will no longer walk proudly, for it will be a time of calamity.
MIC|2|4|In that day men will ridicule you; they will taunt you with this mournful song: 'We are utterly ruined; my people's possession is divided up. He takes it from me! He assigns our fields to traitors.'"
MIC|2|5|Therefore you will have no one in the assembly of the LORD to divide the land by lot.
MIC|2|6|"Do not prophesy," their prophets say. "Do not prophesy about these things; disgrace will not overtake us."
MIC|2|7|Should it be said, O house of Jacob: "Is the Spirit of the LORD angry? Does he do such things?Do not my words do good to him whose ways are upright?
MIC|2|8|Lately my people have risen up like an enemy. You strip off the rich robe from those who pass by without a care, like men returning from battle.
MIC|2|9|You drive the women of my people from their pleasant homes. You take away my blessing from their children forever.
MIC|2|10|Get up, go away! For this is not your resting place, because it is defiled, it is ruined, beyond all remedy.
MIC|2|11|If a liar and deceiver comes and says, 'I will prophesy for you plenty of wine and beer,' he would be just the prophet for this people!
MIC|2|12|"I will surely gather all of you, O Jacob; I will surely bring together the remnant of Israel. I will bring them together like sheep in a pen, like a flock in its pasture; the place will throng with people.
MIC|2|13|One who breaks open the way will go up before them; they will break through the gate and go out. Their king will pass through before them, the LORD at their head."
MIC|3|1|Then I said, "Listen, you leaders of Jacob, you rulers of the house of Israel. Should you not know justice,
MIC|3|2|you who hate good and love evil; who tear the skin from my people and the flesh from their bones;
MIC|3|3|who eat my people's flesh, strip off their skin and break their bones in pieces; who chop them up like meat for the pan, like flesh for the pot?"
MIC|3|4|Then they will cry out to the LORD, but he will not answer them. At that time he will hide his face from them because of the evil they have done.
MIC|3|5|This is what the LORD says: "As for the prophets who lead my people astray, if one feeds them, they proclaim 'peace'; if he does not, they prepare to wage war against him.
MIC|3|6|Therefore night will come over you, without visions, and darkness, without divination. The sun will set for the prophets, and the day will go dark for them.
MIC|3|7|The seers will be ashamed and the diviners disgraced. They will all cover their faces because there is no answer from God."
MIC|3|8|But as for me, I am filled with power, with the Spirit of the LORD, and with justice and might, to declare to Jacob his transgression, to Israel his sin.
MIC|3|9|Hear this, you leaders of the house of Jacob, you rulers of the house of Israel, who despise justice and distort all that is right;
MIC|3|10|who build Zion with bloodshed, and Jerusalem with wickedness.
MIC|3|11|Her leaders judge for a bribe, her priests teach for a price, and her prophets tell fortunes for money. Yet they lean upon the LORD and say, "Is not the LORD among us? No disaster will come upon us."
MIC|3|12|Therefore because of you, Zion will be plowed like a field, Jerusalem will become a heap of rubble, the temple hill a mound overgrown with thickets.
MIC|4|1|In the last days the mountain of the LORD's temple will be established as chief among the mountains; it will be raised above the hills, and peoples will stream to it.
MIC|4|2|Many nations will come and say, "Come, let us go up to the mountain of the LORD, to the house of the God of Jacob. He will teach us his ways, so that we may walk in his paths." The law will go out from Zion, the word of the LORD from Jerusalem.
MIC|4|3|He will judge between many peoples and will settle disputes for strong nations far and wide. They will beat their swords into plowshares and their spears into pruning hooks. Nation will not take up sword against nation, nor will they train for war anymore.
MIC|4|4|Every man will sit under his own vine and under his own fig tree, and no one will make them afraid, for the LORD Almighty has spoken.
MIC|4|5|All the nations may walk in the name of their gods; we will walk in the name of the LORD our God for ever and ever. The LORD 's Plan
MIC|4|6|"In that day," declares the LORD, "I will gather the lame; I will assemble the exiles and those I have brought to grief.
MIC|4|7|I will make the lame a remnant, those driven away a strong nation. The LORD will rule over them in Mount Zion from that day and forever.
MIC|4|8|As for you, O watchtower of the flock, O stronghold of the Daughter of Zion, the former dominion will be restored to you; kingship will come to the Daughter of Jerusalem."
MIC|4|9|Why do you now cry aloud- have you no king? Has your counselor perished, that pain seizes you like that of a woman in labor?
MIC|4|10|Writhe in agony, O Daughter of Zion, like a woman in labor, for now you must leave the city to camp in the open field. You will go to Babylon; there you will be rescued. There the LORD will redeem you out of the hand of your enemies.
MIC|4|11|But now many nations are gathered against you. They say, "Let her be defiled, let our eyes gloat over Zion!"
MIC|4|12|But they do not know the thoughts of the LORD; they do not understand his plan, he who gathers them like sheaves to the threshing floor.
MIC|4|13|"Rise and thresh, O Daughter of Zion, for I will give you horns of iron; I will give you hoofs of bronze and you will break to pieces many nations." You will devote their ill-gotten gains to the LORD, their wealth to the Lord of all the earth.
MIC|5|1|Marshal your troops, O city of troops, for a siege is laid against us. They will strike Israel's ruler on the cheek with a rod.
MIC|5|2|"But you, Bethlehem Ephrathah, though you are small among the clans of Judah, out of you will come for me one who will be ruler over Israel, whose origins are from of old, from ancient times. "
MIC|5|3|Therefore Israel will be abandoned until the time when she who is in labor gives birth and the rest of his brothers return to join the Israelites.
MIC|5|4|He will stand and shepherd his flock in the strength of the LORD, in the majesty of the name of the LORD his God. And they will live securely, for then his greatness will reach to the ends of the earth.
MIC|5|5|And he will be their peace. When the Assyrian invades our land and marches through our fortresses, we will raise against him seven shepherds, even eight leaders of men.
MIC|5|6|They will rule the land of Assyria with the sword, the land of Nimrod with drawn sword. He will deliver us from the Assyrian when he invades our land and marches into our borders.
MIC|5|7|The remnant of Jacob will be in the midst of many peoples like dew from the LORD, like showers on the grass, which do not wait for man or linger for mankind.
MIC|5|8|The remnant of Jacob will be among the nations, in the midst of many peoples, like a lion among the beasts of the forest, like a young lion among flocks of sheep, which mauls and mangles as it goes, and no one can rescue.
MIC|5|9|Your hand will be lifted up in triumph over your enemies, and all your foes will be destroyed.
MIC|5|10|"In that day," declares the LORD, "I will destroy your horses from among you and demolish your chariots.
MIC|5|11|I will destroy the cities of your land and tear down all your strongholds.
MIC|5|12|I will destroy your witchcraft and you will no longer cast spells.
MIC|5|13|I will destroy your carved images and your sacred stones from among you; you will no longer bow down to the work of your hands.
MIC|5|14|I will uproot from among you your Asherah poles and demolish your cities.
MIC|5|15|I will take vengeance in anger and wrath upon the nations that have not obeyed me."
MIC|6|1|Listen to what the LORD says: "Stand up, plead your case before the mountains; let the hills hear what you have to say.
MIC|6|2|Hear, O mountains, the LORD's accusation; listen, you everlasting foundations of the earth. For the LORD has a case against his people; he is lodging a charge against Israel.
MIC|6|3|"My people, what have I done to you? How have I burdened you? Answer me.
MIC|6|4|I brought you up out of Egypt and redeemed you from the land of slavery. I sent Moses to lead you, also Aaron and Miriam.
MIC|6|5|My people, remember what Balak king of Moab counseled and what Balaam son of Beor answered. Remember your journey from Shittim to Gilgal, that you may know the righteous acts of the LORD."
MIC|6|6|With what shall I come before the LORD and bow down before the exalted God? Shall I come before him with burnt offerings, with calves a year old?
MIC|6|7|Will the LORD be pleased with thousands of rams, with ten thousand rivers of oil? Shall I offer my firstborn for my transgression, the fruit of my body for the sin of my soul?
MIC|6|8|He has showed you, O man, what is good. And what does the LORD require of you? To act justly and to love mercy and to walk humbly with your God.
MIC|6|9|Listen! The LORD is calling to the city- and to fear your name is wisdom- "Heed the rod and the One who appointed it.
MIC|6|10|Am I still to forget, O wicked house, your ill-gotten treasures and the short ephah, which is accursed?
MIC|6|11|Shall I acquit a man with dishonest scales, with a bag of false weights?
MIC|6|12|Her rich men are violent; her people are liars and their tongues speak deceitfully.
MIC|6|13|Therefore, I have begun to destroy you, to ruin you because of your sins.
MIC|6|14|You will eat but not be satisfied; your stomach will still be empty. You will store up but save nothing, because what you save I will give to the sword.
MIC|6|15|You will plant but not harvest; you will press olives but not use the oil on yourselves, you will crush grapes but not drink the wine.
MIC|6|16|You have observed the statutes of Omri and all the practices of Ahab's house, and you have followed their traditions. Therefore I will give you over to ruin and your people to derision; you will bear the scorn of the nations. "
MIC|7|1|What misery is mine! I am like one who gathers summer fruit at the gleaning of the vineyard; there is no cluster of grapes to eat, none of the early figs that I crave.
MIC|7|2|The godly have been swept from the land; not one upright man remains. All men lie in wait to shed blood; each hunts his brother with a net.
MIC|7|3|Both hands are skilled in doing evil; the ruler demands gifts, the judge accepts bribes, the powerful dictate what they desire- they all conspire together.
MIC|7|4|The best of them is like a brier, the most upright worse than a thorn hedge. The day of your watchmen has come, the day God visits you. Now is the time of their confusion.
MIC|7|5|Do not trust a neighbor; put no confidence in a friend. Even with her who lies in your embrace be careful of your words.
MIC|7|6|For a son dishonors his father, a daughter rises up against her mother, a daughter-in-law against her mother-in-law- a man's enemies are the members of his own household.
MIC|7|7|But as for me, I watch in hope for the LORD, I wait for God my Savior; my God will hear me.
MIC|7|8|Do not gloat over me, my enemy! Though I have fallen, I will rise. Though I sit in darkness, the LORD will be my light.
MIC|7|9|Because I have sinned against him, I will bear the LORD's wrath, until he pleads my case and establishes my right. He will bring me out into the light; I will see his righteousness.
MIC|7|10|Then my enemy will see it and will be covered with shame, she who said to me, "Where is the LORD your God?" My eyes will see her downfall; even now she will be trampled underfoot like mire in the streets.
MIC|7|11|The day for building your walls will come, the day for extending your boundaries.
MIC|7|12|In that day people will come to you from Assyria and the cities of Egypt, even from Egypt to the Euphrates and from sea to sea and from mountain to mountain.
MIC|7|13|The earth will become desolate because of its inhabitants, as the result of their deeds.
MIC|7|14|Shepherd your people with your staff, the flock of your inheritance, which lives by itself in a forest, in fertile pasturelands. Let them feed in Bashan and Gilead as in days long ago.
MIC|7|15|"As in the days when you came out of Egypt, I will show them my wonders."
MIC|7|16|Nations will see and be ashamed, deprived of all their power. They will lay their hands on their mouths and their ears will become deaf.
MIC|7|17|They will lick dust like a snake, like creatures that crawl on the ground. They will come trembling out of their dens; they will turn in fear to the LORD our God and will be afraid of you.
MIC|7|18|Who is a God like you, who pardons sin and forgives the transgression of the remnant of his inheritance? You do not stay angry forever but delight to show mercy.
MIC|7|19|You will again have compassion on us; you will tread our sins underfoot and hurl all our iniquities into the depths of the sea.
MIC|7|20|You will be true to Jacob, and show mercy to Abraham, as you pledged on oath to our fathers in days long ago.
