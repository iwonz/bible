TITUS|1|1|上帝的仆人、耶稣基督的使徒 保罗 ，为了使上帝的选民信从与认识合乎敬虔的真理—
TITUS|1|2|这真理是在盼望那无谎言的上帝在万古之先所应许的永生，
TITUS|1|3|到了适当的时机，藉着传扬福音，把他的道显明了；这传扬的责任是按着我们的救主上帝的命令交托给我的—
TITUS|1|4|我写信给在共同的信仰上作我真儿子的 提多 。愿恩惠、平安 从父上帝和我们的救主基督耶稣归给你！
TITUS|1|5|我从前把你留在 克里特 ，是要你将那没有办完的事都办妥，又照我所吩咐你的，在各城设立长老。
TITUS|1|6|若有无可指责的人，只作一个妇人的丈夫，儿女也是信主的，没有人告他们放荡，不受约束，就可以设立。
TITUS|1|7|监督既然是上帝的管家，必须无可指责、不自负、不暴躁、不酗酒、不好斗、不贪财；
TITUS|1|8|却要乐意接待外人、好善、克己、正直、圣洁、节制，
TITUS|1|9|坚守合乎教义的可靠之道，就能将健全的教导劝勉人，又能驳倒争辩的人。
TITUS|1|10|因为也有许多人不受约束，说空话欺哄人，尤其是那些奉割礼的人。
TITUS|1|11|这些人的口必须堵住，因为他们贪不义之财，将不该教导的事教导人，败坏人的全家。
TITUS|1|12|克里特 人中有一个本地的先知说：“ 克里特 人常说谎话，是恶兽，贪吃懒做。”
TITUS|1|13|这个见证是真的。为这缘故，你要严厉地责备他们，使他们在信仰上健全。
TITUS|1|14|不要听 犹太 人无稽的传说和背弃真理之人的命令。
TITUS|1|15|在洁净的人，凡物都洁净；在污秽不信的人，什么都不洁净，连心地和天良也都污秽了。
TITUS|1|16|他们宣称认识上帝，却在行为上否认他；他们是可憎恶的，是悖逆的，不配做任何好事。
TITUS|2|1|至于你，你所讲的总要合乎那健全的教导。
TITUS|2|2|劝老年人要有节制、端正、克己，在信心、爱心、耐心上都要健全。
TITUS|2|3|又要劝年长的妇女在操守上恭正，不说谗言，不作酒的奴隶，用善道教导人，
TITUS|2|4|好指教年轻的妇女爱丈夫，爱儿女，
TITUS|2|5|克己，贞洁，理家，善良，顺服自己的丈夫，免得上帝的道被毁谤。
TITUS|2|6|同样，要劝年轻人凡事克己。
TITUS|2|7|你要显出自己是好行为的榜样，在教导上要正直、庄重，
TITUS|2|8|言语健全，无可指责，使那反对的人，因说不出我们有什么不好而自觉羞愧。
TITUS|2|9|要劝仆人顺服自己的主人，凡事讨他的喜悦，不可顶撞他，
TITUS|2|10|不可私窃财物；要凡事显出完美的忠诚，好事事都能荣耀我们救主上帝的教导。
TITUS|2|11|因为，上帝救众人的恩典已经显明出来，
TITUS|2|12|训练我们除去不敬虔的心和世俗的情欲，在今世过克己、正直、敬虔的生活，
TITUS|2|13|等候福乐的盼望，并等候至大的上帝和我们的救主 耶稣基督的荣耀显现。
TITUS|2|14|他为我们的缘故舍己，为了要赎我们脱离一切罪恶，又洁净我们作他自己的子民，热心为善。
TITUS|2|15|这些事你要讲明，要充分运用你的职权劝勉人，责备人。不要让任何人轻看你。
TITUS|3|1|你要提醒众人，叫他们顺服执政的、掌权的，要服从，预备行各样善事。
TITUS|3|2|不要毁谤，不要争吵，要和气，对众人总要显出温柔。
TITUS|3|3|我们从前也是无知、悖逆、受迷惑，作各样私欲和宴乐的奴隶，在恶毒、嫉妒中度日，是可恨的，而且彼此相恨。
TITUS|3|4|但到了我们救主上帝的恩慈和慈爱显明的时候，
TITUS|3|5|他救了我们，并不是因我们自己所行的义，而是照他的怜悯，藉着重生的洗和圣灵的更新。
TITUS|3|6|圣灵就是上帝藉着我们的救主耶稣基督厚厚地浇灌在我们身上的，
TITUS|3|7|好让我们因他的恩得称为义，可以凭着永生的盼望成为后嗣 。
TITUS|3|8|这话是可信的。 我愿你坚持这些事，使那些已信上帝的人留心行善 。这都是美好且对人有益的。
TITUS|3|9|要远避愚拙的辩论、家谱、纷争和因律法而起的争辩，因为这都是虚妄无益的。
TITUS|3|10|分门结党的人，警戒过一两次后就要拒绝跟他来往；
TITUS|3|11|因为你知道这样的人已经背道，常常犯罪，自己定自己的罪了。
TITUS|3|12|我打发 亚提马 或 推基古 到你那里去的时候，你要赶紧往 尼哥坡里 来见我，因为我已经决定在那里过冬。
TITUS|3|13|你要赶紧给 西纳 律师和 亚波罗 送行，让他们没有缺乏。
TITUS|3|14|我们的人也该学习行善，帮助有迫切需要的人，这样才不会不结果子。
TITUS|3|15|跟我同在一起的人都向你问安。请代向在信仰上爱我们的人问安。愿恩惠与你们众人同在！
