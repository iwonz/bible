JER|1|1|Слова Иеремии, сына Хелкиина, из священников в Анафофе, в земле Вениаминовой,
JER|1|2|к которому было слово Господне во дни Иосии, сына Амонова, царя Иудейского, в тринадцатый год царствования его,
JER|1|3|и также во дни Иоакима, сына Иосиина, царя Иудейского, до конца одиннадцатого года Седекии, сына Иосиина, царя Иудейского, до переселения Иерусалима в пятом месяце.
JER|1|4|И было ко мне слово Господне:
JER|1|5|прежде нежели Я образовал тебя во чреве, Я познал тебя, и прежде нежели ты вышел из утробы, Я освятил тебя: пророком для народов поставил тебя.
JER|1|6|А я сказал: о, Господи Боже! я не умею говорить, ибо я еще молод.
JER|1|7|Но Господь сказал мне: не говори: "я молод"; ибо ко всем, к кому пошлю тебя, пойдешь, и все, что повелю тебе, скажешь.
JER|1|8|Не бойся их; ибо Я с тобою, чтобы избавлять тебя, сказал Господь.
JER|1|9|И простер Господь руку Свою, и коснулся уст моих, и сказал мне Господь: вот, Я вложил слова Мои в уста твои.
JER|1|10|Смотри, Я поставил тебя в сей день над народами и царствами, чтобы искоренять и разорять, губить и разрушать, созидать и насаждать.
JER|1|11|И было слово Господне ко мне: что видишь ты, Иеремия? Я сказал: вижу жезл миндального дерева.
JER|1|12|Господь сказал мне: ты верно видишь; ибо Я бодрствую над словом Моим, чтоб оно скоро исполнилось.
JER|1|13|И было слово Господне ко мне в другой раз: что видишь ты? Я сказал: вижу поддуваемый ветром кипящий котел, и лицо его со стороны севера.
JER|1|14|И сказал мне Господь: от севера откроется бедствие на всех обитателей сей земли.
JER|1|15|Ибо вот, Я призову все племена царств северных, говорит Господь, и придут они, и поставят каждый престол свой при входе в ворота Иерусалима, и вокруг всех стен его, и во всех городах Иудейских.
JER|1|16|И произнесу над ними суды Мои за все беззакония их, за то, что они оставили Меня, и воскуряли фимиам чужеземным богам и поклонялись делам рук своих.
JER|1|17|А ты препояшь чресла твои, и встань, и скажи им все, что Я повелю тебе; не малодушествуй пред ними, чтобы Я не поразил тебя в глазах их.
JER|1|18|И вот, Я поставил тебя ныне укрепленным городом и железным столбом и медною стеною на всей этой земле, против царей Иуды, против князей его, против священников его и против народа земли сей.
JER|1|19|Они будут ратовать против тебя, но не превозмогут тебя; ибо Я с тобою, говорит Господь, чтобы избавлять тебя.
JER|2|1|И было слово Господне ко мне:
JER|2|2|иди и возгласи в уши [дщери] Иерусалима: так говорит Господь: Я вспоминаю о дружестве юности твоей, о любви твоей, когда ты была невестою, когда последовала за Мною в пустыню, в землю незасеянную.
JER|2|3|Израиль [был] святынею Господа, начатком плодов Его; все поедавшие его были осуждаемы, бедствие постигало их, говорит Господь.
JER|2|4|Выслушайте слово Господне, дом Иаковлев и все роды дома Израилева!
JER|2|5|Так говорит Господь: какую неправду нашли во Мне отцы ваши, что удалились от Меня и пошли за суетою, и осуетились,
JER|2|6|и не сказали: "где Господь, Который вывел нас из земли Египетской, вел нас по пустыне, по земле пустой и необитаемой, по земле сухой, по земле тени смертной, по которой никто не ходил и где не обитал человек?"
JER|2|7|И Я ввел вас в землю плодоносную, чтобы вы питались плодами ее и добром ее; а вы вошли и осквернили землю Мою, и достояние Мое сделали мерзостью.
JER|2|8|Священники не говорили: "где Господь?", и учители закона не знали Меня, и пастыри отпали от Меня, и пророки пророчествовали во имя Ваала и ходили во след тех, которые не помогают.
JER|2|9|Поэтому Я еще буду судиться с вами, говорит Господь, и с сыновьями сыновей ваших буду судиться.
JER|2|10|Ибо пойдите на острова Хиттимские и посмотрите, и пошлите в Кидар и разведайте прилежно, и рассмотрите: было ли [там] что–нибудь подобное сему?
JER|2|11|переменил ли какой народ богов [своих], хотя они и не боги? а Мой народ променял славу свою на то, что не помогает.
JER|2|12|Подивитесь сему, небеса, и содрогнитесь, и ужаснитесь, говорит Господь.
JER|2|13|Ибо два зла сделал народ Мой: Меня, источник воды живой, оставили, и высекли себе водоемы разбитые, которые не могут держать воды.
JER|2|14|Разве Израиль раб? или он домочадец? почему он сделался добычею?
JER|2|15|Зарыкали на него молодые львы, подали голос свой и сделали землю его пустынею; города его сожжены, без жителей.
JER|2|16|И сыновья Мемфиса и Тафны объели темя твое.
JER|2|17|Не причинил ли ты себе это тем, что оставил Господа Бога твоего в то время, когда Он путеводил тебя?
JER|2|18|И ныне для чего тебе путь в Египет, чтобы пить воду из Нила? и для чего тебе путь в Ассирию, чтобы пить воду из реки ее?
JER|2|19|Накажет тебя нечестие твое, и отступничество твое обличит тебя; итак познай и размысли, как худо и горько то, что ты оставил Господа Бога твоего и страха Моего нет в тебе, говорит Господь Бог Саваоф.
JER|2|20|Ибо издавна Я сокрушил ярмо твое, разорвал узы твои, и ты говорил: "не буду служить [идолам]", а между тем на всяком высоком холме и под всяким ветвистым деревом ты блудодействовал.
JER|2|21|Я насадил тебя [как] благородную лозу, – самое чистое семя; как же ты превратилась у Меня в дикую отрасль чужой лозы?
JER|2|22|Посему, хотя бы ты умылся мылом и много употребил на себя щелоку, нечестие твое отмечено предо Мною, говорит Господь Бог.
JER|2|23|Как можешь ты сказать: "я не осквернил себя, я не ходил во след Ваала?" Посмотри на поведение твое в долине, познай, что делала ты, резвая верблюдица, рыщущая по путям твоим?
JER|2|24|Привыкшую к пустыне дикую ослицу, в страсти души своей глотающую воздух, кто может удержать? Все, ищущие ее, не утомятся: в ее месяце они найдут ее.
JER|2|25|Не давай ногам твоим истаптывать обувь, и гортани твоей – томиться жаждою. Но ты сказал: "не надейся, нет! ибо люблю чужих и буду ходить во след их".
JER|2|26|Как вор, когда поймают его, бывает осрамлен, так осрамил себя дом Израилев: они, цари их, князья их, и священники их, и пророки их, –
JER|2|27|говоря дереву: "ты мой отец", и камню: "ты родил меня"; ибо они оборотили ко Мне спину, а не лице; а во время бедствия своего будут говорить: "встань и спаси нас!"
JER|2|28|Где же боги твои, которых ты сделал себе? – пусть они встанут, если могут спасти тебя во время бедствия твоего; ибо сколько у тебя городов, столько и богов у тебя, Иуда.
JER|2|29|Для чего вам состязаться со Мною? – все вы согрешали против Меня, говорит Господь.
JER|2|30|Вотще поражал Я детей ваших: они не приняли вразумления; пророков ваших поядал меч ваш, как истребляющий лев.
JER|2|31|О, род! внемлите вы слову Господню: был ли Я пустынею для Израиля? был ли Я страною мрака? Зачем же народ Мой говорит: "мы сами себе господа; мы уже не придем к Тебе"?
JER|2|32|Забывает ли девица украшение свое и невеста – наряд свой? а народ Мой забыл Меня, – нет числа дням.
JER|2|33|Как искусно направляешь ты пути твои, чтобы снискать любовь! и для того даже к преступлениям приспособляла ты пути твои.
JER|2|34|Даже на полах одежды твоей находится кровь людей бедных, невинных, которых ты не застала при взломе, и, несмотря на все это,
JER|2|35|говоришь: "так как я невинна, то верно гнев Его отвратится от меня". Вот, Я буду судиться с тобою за то, что говоришь: "я не согрешила".
JER|2|36|Зачем ты так много бродишь, меняя путь твой? Ты так же будешь посрамлена и Египтом, как была посрамлена Ассириею;
JER|2|37|и от него ты выйдешь, положив руки на голову, потому что отверг Господь надежды твои, и не будешь иметь с ними успеха.
JER|3|1|Говорят: "если муж отпустит жену свою, и она отойдет от него и сделается женою другого мужа, то может ли она возвратиться к нему? Не осквернилась ли бы этим страна та?" А ты со многими любовниками блудодействовала, – и однако же возвратись ко Мне, говорит Господь.
JER|3|2|Подними глаза твои на высоты и посмотри, где не блудодействовали с тобою? У дороги сидела ты для них, как Аравитянин в пустыне, и осквернила землю блудом твоим и лукавством твоим.
JER|3|3|За то были удержаны дожди, и не было дождя позднего; но у тебя был лоб блудницы, ты отбросила стыд.
JER|3|4|Не будешь ли ты отныне взывать ко Мне: "Отец мой! Ты был путеводителем юности моей!
JER|3|5|Неужели всегда будет Он во гневе? и неужели вечно будет удерживать его в Себе?" Вот, что говоришь ты, а делаешь зло и преуспеваешь в нем.
JER|3|6|Господь сказал мне во дни Иосии царя: видел ли ты, что делала отступница, дочь Израиля? Она ходила на всякую высокую гору и под всякое ветвистое дерево и там блудодействовала.
JER|3|7|И после того, как она все это делала, Я говорил: "возвратись ко Мне"; но она не возвратилась; и видела [это] вероломная сестра ее Иудея.
JER|3|8|И Я видел, что, когда за все прелюбодейные действия отступницы, дочери Израиля, Я отпустил ее и дал ей разводное письмо, вероломная сестра ее Иудея не убоялась, а пошла и сама блудодействовала.
JER|3|9|И явным блудодейством она осквернила землю, и прелюбодействовала с камнем и деревом.
JER|3|10|Но при всем этом вероломная сестра ее Иудея не обратилась ко Мне всем сердцем своим, а только притворно, говорит Господь.
JER|3|11|И сказал мне Господь: отступница, [дочь] Израилева, оказалась правее, нежели вероломная Иудея.
JER|3|12|Иди и провозгласи слова сии к северу, и скажи: возвратись, отступница, [дочь] Израилева, говорит Господь. Я не изолью на вас гнева Моего; ибо Я милостив, говорит Господь, – не вечно буду негодовать.
JER|3|13|Признай только вину твою: ибо ты отступила от Господа Бога твоего и распутствовала с чужими под всяким ветвистым деревом, а гласа Моего вы не слушали, говорит Господь.
JER|3|14|Возвратитесь, дети–отступники, говорит Господь, потому что Я сочетался с вами, и возьму вас по одному из города, по два из племени, и приведу вас на Сион.
JER|3|15|И дам вам пастырей по сердцу Моему, которые будут пасти вас с знанием и благоразумием
JER|3|16|И будет, когда вы размножитесь и сделаетесь многоплодными на земле, в те дни, говорит Господь, не будут говорить более: "ковчег завета Господня"; он и на ум не придет, и не вспомнят о нем, и не будут приходить к нему, и его уже не будет.
JER|3|17|В то время назовут Иерусалим престолом Господа; и все народы ради имени Господа соберутся в Иерусалим и не будут более поступать по упорству злого сердца своего.
JER|3|18|В те дни придет дом Иудин к дому Израилеву, и пойдут вместе из земли северной в землю, которую Я дал в наследие отцам вашим.
JER|3|19|И говорил Я: как поставлю тебя в число детей и дам тебе вожделенную землю, прекраснейшее наследие множества народов? И сказал: ты будешь называть Меня отцом твоим и не отступишь от Меня.
JER|3|20|Но поистине, как жена вероломно изменяет другу своему, так вероломно поступили со Мною вы, дом Израилев, говорит Господь.
JER|3|21|Голос слышен на высотах, жалобный плач сынов Израиля о том, что они извратили путь свой, забыли Господа Бога своего.
JER|3|22|Возвратитесь, мятежные дети: Я исцелю вашу непокорность. – Вот, мы идем к Тебе, ибо Ты – Господь Бог наш.
JER|3|23|Поистине, напрасно надеялись мы на холмы и на множество гор; поистине, в Господе Боге нашем спасение Израилево!
JER|3|24|От юности нашей эта мерзость пожирала труды отцов наших, овец их и волов их, сыновей их и дочерей их.
JER|3|25|Мы лежим в стыде своем, и срам наш покрывает нас, потому что мы грешили пред Господом Богом нашим, – мы и отцы наши, от юности нашей и до сего дня, и не слушались голоса Господа Бога нашего.
JER|4|1|Если хочешь обратиться, Израиль, говорит Господь, ко Мне обратись; и если удалишь мерзости твои от лица Моего, то не будешь скитаться.
JER|4|2|И будешь клясться: "жив Господь!" в истине, суде и правде; и народы Им будут благословляться и Им хвалиться.
JER|4|3|Ибо так говорит Господь к мужам Иуды и Иерусалима: распашите себе новые нивы и не сейте между тернами.
JER|4|4|Обрежьте себя для Господа, и снимите крайнюю плоть с сердца вашего, мужи Иуды и жители Иерусалима, чтобы гнев Мой не открылся, как огонь, и не воспылал неугасимо по причине злых наклонностей ваших.
JER|4|5|Объявите в Иудее и разгласите в Иерусалиме, и говорите, и трубите трубою по земле; взывайте громко и говорите: "соберитесь, и пойдем в укрепленные города".
JER|4|6|Выставьте знамя к Сиону, бегите, не останавливайтесь, ибо Я приведу от севера бедствие и великую гибель.
JER|4|7|Выходит лев из своей чащи, и выступает истребитель народов: он выходит из своего места, чтобы землю твою сделать пустынею; города твои будут разорены, [останутся] без жителей.
JER|4|8|Посему препояшьтесь вретищем, плачьте и рыдайте, ибо ярость гнева Господня не отвратится от нас.
JER|4|9|И будет в тот день, говорит Господь, замрет сердце у царя и сердце у князей; и ужаснутся священники, и изумятся пророки.
JER|4|10|И сказал я: о, Господи Боже! Неужели Ты обольщал только народ сей и Иерусалим, говоря: "мир будет у вас"; а между тем меч доходит до души?
JER|4|11|В то время сказано будет народу сему и Иерусалиму: жгучий ветер несется с высот пустынных на путь дочери народа Моего, не для веяния и не для очищения;
JER|4|12|и придет ко Мне оттуда ветер сильнее сего, и Я произнесу суд над ними.
JER|4|13|Вот, поднимается он подобно облакам, и колесницы его – как вихрь, кони его быстрее орлов; горе нам! ибо мы будем разорены.
JER|4|14|Смой злое с сердца твоего, Иерусалим, чтобы спастись тебе: доколе будут гнездиться в тебе злочестивые мысли?
JER|4|15|Ибо уже несется голос от Дана и гибельная весть с горы Ефремовой:
JER|4|16|объявите народам, известите Иерусалим, что идут из дальней страны осаждающие и криками своими оглашают города Иудеи.
JER|4|17|Как сторожа полей, они обступают его кругом, ибо он возмутился против Меня, говорит Господь.
JER|4|18|Пути твои и деяния твои причинили тебе это; от твоего нечестия тебе так горько, что доходит до сердца твоего.
JER|4|19|Утроба моя! утроба моя! скорблю во глубине сердца моего, волнуется во мне сердце мое, не могу молчать; ибо ты слышишь, душа моя, звук трубы, тревогу брани.
JER|4|20|Беда за бедою: вся земля опустошается, внезапно разорены шатры мои, мгновенно – палатки мои.
JER|4|21|Долго ли мне видеть знамя, слушать звук трубы?
JER|4|22|Это от того, что народ Мой глуп, не знает Меня: неразумные они дети, и нет у них смысла; они умны на зло, но добра делать не умеют.
JER|4|23|Смотрю на землю, и вот, она разорена и пуста, – на небеса, и нет на них света.
JER|4|24|Смотрю на горы, и вот, они дрожат, и все холмы колеблются.
JER|4|25|Смотрю, и вот, нет человека, и все птицы небесные разлетелись.
JER|4|26|Смотрю, и вот, Кармил – пустыня, и все города его разрушены от лица Господа, от ярости гнева Его.
JER|4|27|Ибо так сказал Господь: вся земля будет опустошена, но совершенного истребления не сделаю.
JER|4|28|Восплачет о сем земля, и небеса помрачатся вверху, потому что Я сказал, Я определил, и не раскаюсь в том, и не отступлю от того.
JER|4|29|От шума всадников и стрелков разбегутся все города: они уйдут в густые леса и влезут на скалы; все города будут оставлены, и не будет в них ни одного жителя.
JER|4|30|А ты, опустошенная, что станешь делать? Хотя ты одеваешься в пурпур, хотя украшаешь себя золотыми нарядами, обрисовываешь глаза твои красками, но напрасно украшаешь себя: презрели тебя любовники, они ищут души твоей.
JER|4|31|Ибо Я слышу голос как бы женщины в родах, стон как бы рождающей в первый раз, голос дочери Сиона; она стонет, простирая руки свои: "о, горе мне! душа моя изнывает пред убийцами".
JER|5|1|Походите по улицам Иерусалима, и посмотрите, и разведайте, и поищите на площадях его, не найдете ли человека, нет ли соблюдающего правду, ищущего истины? Я пощадил бы [Иерусалим].
JER|5|2|Хотя и говорят они: "жив Господь!", но клянутся ложно.
JER|5|3|О, Господи! очи Твои не к истине ли [обращены]? Ты поражаешь их, а они не чувствуют боли; Ты истребляешь их, а они не хотят принять вразумления; лица свои сделали они крепче камня, не хотят обратиться.
JER|5|4|И сказал я [сам в себе]: это, может быть, бедняки; они глупы, потому что не знают пути Господня, закона Бога своего;
JER|5|5|пойду я к знатным и поговорю с ними, ибо они знают путь Господень, закон Бога своего. Но и они все сокрушили ярмо, расторгли узы.
JER|5|6|За то поразит их лев из леса, волк пустынный опустошит их, барс будет подстерегать у городов их: кто выйдет из них, будет растерзан; ибо умножились преступления их, усилились отступничества их.
JER|5|7|Как же Мне простить тебя за это? Сыновья твои оставили Меня и клянутся теми, которые не боги. Я насыщал их, а они прелюбодействовали и толпами ходили в домы блудниц.
JER|5|8|Это откормленные кони: каждый из них ржет на жену другого.
JER|5|9|Неужели Я не накажу за это? говорит Господь; и не отмстит ли душа Моя такому народу, как этот?
JER|5|10|Восходите на стены его и разрушайте, но не до конца; уничтожьте зубцы их, потому что они не Господни;
JER|5|11|ибо дом Израилев и дом Иудин поступили со Мною очень вероломно, говорит Господь:
JER|5|12|они солгали на Господа и сказали: "нет Его, и беда не придет на нас, и мы не увидим ни меча, ни голода.
JER|5|13|И пророки станут ветром, и слова [Господня] нет в них; над ними самими пусть это будет".
JER|5|14|Посему так говорит Господь Бог Саваоф: за то, что вы говорите такие слова, вот, Я сделаю слова Мои в устах твоих огнем, а этот народ – дровами, и этот [огонь] пожрет их.
JER|5|15|Вот, Я приведу на вас, дом Израилев, народ издалека, говорит Господь, народ сильный, народ древний, народ, которого языка ты не знаешь, и не будешь понимать, что он говорит.
JER|5|16|Колчан его – как открытый гроб; все они люди храбрые.
JER|5|17|И съедят они жатву твою и хлеб твой, съедят сыновей твоих и дочерей твоих, съедят овец твоих и волов твоих, съедят виноград твой и смоквы твои; разрушат мечом укрепленные города твои, на которые ты надеешься.
JER|5|18|Но и в те дни, говорит Господь, не истреблю вас до конца.
JER|5|19|И если вы скажете: "за что Господь, Бог наш, делает нам все это?", то отвечай: так как вы оставили Меня и служили чужим богам в земле своей, то будете служить чужим в земле не вашей.
JER|5|20|Объявите это в доме Иакова и возвестите в Иудее, говоря:
JER|5|21|выслушай это, народ глупый и неразумный, у которого есть глаза, а не видит, у которого есть уши, а не слышит:
JER|5|22|Меня ли вы не боитесь, говорит Господь, предо Мною ли не трепещете? Я положил песок границею морю, вечным пределом, которого не перейдет; и хотя волны его устремляются, но превозмочь не могут; хотя они бушуют, но переступить его не могут.
JER|5|23|А у народа сего сердце буйное и мятежное; они отступили и пошли;
JER|5|24|и не сказали в сердце своем: "убоимся Господа Бога нашего, Который дает нам дождь ранний и поздний в свое время, хранит для нас седмицы, назначенные для жатвы".
JER|5|25|Беззакония ваши отвратили это, и грехи ваши удалили от вас это доброе.
JER|5|26|Ибо между народом Моим находятся нечестивые: сторожат, как птицеловы, припадают к земле, ставят ловушки и уловляют людей.
JER|5|27|Как клетка, наполненная птицами, домы их полны обмана; чрез это они и возвысились и разбогатели,
JER|5|28|сделались тучны, жирны, переступили даже всякую меру во зле, не разбирают судебных дел, дел сирот; благоденствуют, и справедливому делу нищих не дают суда.
JER|5|29|Неужели Я не накажу за это? говорит Господь; и не отмстит ли душа Моя такому народу, как этот?
JER|5|30|Изумительное и ужасное совершается в сей земле:
JER|5|31|пророки пророчествуют ложь, и священники господствуют при посредстве их, и народ Мой любит это. Что же вы будете делать после всего этого?
JER|6|1|Бегите, дети Вениаминовы, из среды Иерусалима, и в Фекое трубите трубою и дайте знать огнем в Бефкареме, ибо от севера появляется беда и великая гибель.
JER|6|2|Разорю Я дочь Сиона, красивую и изнеженную.
JER|6|3|Пастухи со своими стадами придут к ней, раскинут палатки вокруг нее; каждый будет пасти свой участок.
JER|6|4|Приготовляйте против нее войну; вставайте и пойдем в полдень. Горе нам! день уже склоняется, распростираются вечерние тени.
JER|6|5|Вставайте, пойдем и ночью, и разорим чертоги ее!
JER|6|6|Ибо так говорит Господь Саваоф: рубите дерева и делайте насыпь против Иерусалима: этот город должен быть наказан; в нем всякое угнетение.
JER|6|7|Как источник извергает из себя воду, так он источает из себя зло: в нем слышно насилие и грабительство, пред лицем Моим всегда обиды и раны.
JER|6|8|Вразумись, Иерусалим, чтобы душа Моя не удалилась от тебя, чтоб Я не сделал тебя пустынею, землею необитаемою.
JER|6|9|Так говорит Господь Саваоф: до конца доберут остаток Израиля, как виноград; работай рукою твоею, как обиратель винограда, наполняя корзины.
JER|6|10|К кому мне говорить и кого увещевать, чтобы слушали? Вот, ухо у них необрезанное, и они не могут слушать; вот, слово Господне у них в посмеянии; оно неприятно им.
JER|6|11|Поэтому я преисполнен яростью Господнею, не могу держать ее в себе; изолью ее на детей на улице и на собрание юношей; взяты будут муж с женою, пожилой с отжившим лета.
JER|6|12|И домы их перейдут к другим, равно поля и жены; потому что Я простру руку Мою на обитателей сей земли, говорит Господь.
JER|6|13|Ибо от малого до большого, каждый из них предан корысти, и от пророка до священника – все действуют лживо;
JER|6|14|врачуют раны народа Моего легкомысленно, говоря: "мир! мир!", а мира нет.
JER|6|15|Стыдятся ли они, делая мерзости? нет, нисколько не стыдятся и не краснеют. За то падут между падшими, и во время посещения Моего будут повержены, говорит Господь.
JER|6|16|Так говорит Господь: остановитесь на путях ваших и рассмотрите, и расспросите о путях древних, где путь добрый, и идите по нему, и найдете покой душам вашим. Но они сказали: "не пойдем".
JER|6|17|И поставил Я стражей над вами, [сказав]: "слушайте звука трубы". Но они сказали: "не будем слушать".
JER|6|18|Итак слушайте, народы, и знай, собрание, что с ними будет.
JER|6|19|Слушай, земля: вот, Я приведу на народ сей пагубу, плод помыслов их; ибо они слов Моих не слушали и закон Мой отвергли.
JER|6|20|Для чего Мне ладан, который идет из Савы, и благовонный тростник из дальней страны? Всесожжения ваши неугодны, и жертвы ваши неприятны Мне.
JER|6|21|Посему так говорит Господь: вот, Я полагаю пред народом сим преткновения, и преткнутся о них отцы и дети вместе, сосед и друг его, и погибнут.
JER|6|22|Так говорит Господь: вот, идет народ от страны северной, и народ великий поднимается от краев земли;
JER|6|23|держат в руках лук и копье; они жестоки и немилосерды, голос их шумит, как море, и несутся на конях, выстроены, как один человек, чтобы сразиться с тобою, дочь Сиона.
JER|6|24|Мы услышали весть о них, и руки у нас опустились, скорбь объяла нас, муки, как женщину в родах.
JER|6|25|Не выходите в поле и не ходите по дороге, ибо меч неприятелей, ужас со всех сторон.
JER|6|26|Дочь народа моего! опояшь себя вретищем и посыпь себя пеплом; сокрушайся, как бы о смерти единственного сына, горько плачь; ибо внезапно придет на нас губитель.
JER|6|27|Башнею поставил Я тебя среди народа Моего, столпом, чтобы ты знал и следил путь их.
JER|6|28|Все они – упорные отступники, живут клеветою; это медь и железо, – все они развратители.
JER|6|29|Раздувальный мех обгорел, свинец истлел от огня: плавильщик плавил напрасно, ибо злые не отделились;
JER|6|30|отверженным серебром назовут их, ибо Господь отверг их.
JER|7|1|Слово, которое было к Иеремии от Господа:
JER|7|2|стань во вратах дома Господня и провозгласи там слово сие и скажи: слушайте слово Господне, все Иудеи, входящие сими вратами на поклонение Господу.
JER|7|3|Так говорит Господь Саваоф, Бог Израилев: исправьте пути ваши и деяния ваши, и Я оставлю вас жить на сем месте.
JER|7|4|Не надейтесь на обманчивые слова: "здесь храм Господень, храм Господень, храм Господень".
JER|7|5|Но если совсем исправите пути ваши и деяния ваши, если будете верно производить суд между человеком и соперником его,
JER|7|6|не будете притеснять иноземца, сироты и вдовы, и проливать невинной крови на месте сем, и не пойдете во след иных богов на беду себе, –
JER|7|7|то Я оставлю вас жить на месте сем, на этой земле, которую дал отцам вашим в роды родов.
JER|7|8|Вот, вы надеетесь на обманчивые слова, которые не принесут вам пользы.
JER|7|9|Как! вы крадете, убиваете и прелюбодействуете, и клянетесь во лжи и кадите Ваалу, и ходите во след иных богов, которых вы не знаете,
JER|7|10|и потом приходите и становитесь пред лицем Моим в доме сем, над которым наречено имя Мое, и говорите: "мы спасены", чтобы впредь делать все эти мерзости.
JER|7|11|Не соделался ли вертепом разбойников в глазах ваших дом сей, над которым наречено имя Мое? Вот, Я видел это, говорит Господь.
JER|7|12|Пойдите же на место Мое в Силом, где Я прежде назначил пребывать имени Моему, и посмотрите, что сделал Я с ним за нечестие народа Моего Израиля.
JER|7|13|И ныне, так как вы делаете все эти дела, говорит Господь, и Я говорил вам с раннего утра, а вы не слушали, и звал вас, а вы не отвечали, –
JER|7|14|то Я так же поступлю с домом [сим], над которым наречено имя Мое, на который вы надеетесь, и с местом, которое Я дал вам и отцам вашим, как поступил с Силомом.
JER|7|15|И отвергну вас от лица Моего, как отверг всех братьев ваших, все семя Ефремово.
JER|7|16|Ты же не проси за этот народ и не возноси за них молитвы и прошения, и не ходатайствуй предо Мною, ибо Я не услышу тебя.
JER|7|17|Не видишь ли, что они делают в городах Иудеи и на улицах Иерусалима?
JER|7|18|Дети собирают дрова, а отцы разводят огонь, и женщины месят тесто, чтобы делать пирожки для богини неба и совершать возлияния иным богам, чтобы огорчать Меня.
JER|7|19|Но Меня ли огорчают они? говорит Господь; не себя ли самих к стыду своему?
JER|7|20|Посему так говорит Господь Бог: вот, изливается гнев Мой и ярость Моя на место сие, на людей и на скот, и на дерева полевые и на плоды земли, и возгорится и не погаснет.
JER|7|21|Так говорит Господь Саваоф, Бог Израилев: всесожжения ваши прилагайте к жертвам вашим и ешьте мясо;
JER|7|22|ибо отцам вашим Я не говорил и не давал им заповеди в тот день, в который Я вывел их из земли Египетской, о всесожжении и жертве;
JER|7|23|но такую заповедь дал им: "слушайтесь гласа Моего, и Я буду вашим Богом, а вы будете Моим народом, и ходите по всякому пути, который Я заповедаю вам, чтобы вам было хорошо".
JER|7|24|Но они не послушали и не приклонили уха своего, и жили по внушению и упорству злого сердца своего, и стали ко Мне спиною, а не лицом.
JER|7|25|С того дня, как отцы ваши вышли из земли Египетской, до сего дня Я посылал к вам всех рабов Моих – пророков, посылал всякий день с раннего утра;
JER|7|26|но они не слушались Меня и не приклонили уха своего, а ожесточили выю свою, поступали хуже отцов своих.
JER|7|27|И когда ты будешь говорить им все эти слова, они тебя не послушают; и когда будешь звать их, они тебе не ответят.
JER|7|28|Тогда скажи им: вот народ, который не слушает гласа Господа Бога своего и не принимает наставления! Не стало у них истины, она отнята от уст их.
JER|7|29|Остриги волоса твои и брось, и подними плач на горах, ибо отверг Господь и оставил род, [навлекший] гнев Его.
JER|7|30|Ибо сыновья Иуды делают злое пред очами Моими, говорит Господь; поставили мерзости свои в доме, над которым наречено имя Мое, чтобы осквернить его;
JER|7|31|и устроили высоты Тофета в долине сыновей Енномовых, чтобы сожигать сыновей своих и дочерей своих в огне, чего Я не повелевал и что Мне на сердце не приходило.
JER|7|32|За то вот, приходят дни, говорит Господь, когда не будут более называть [место сие] Тофетом и долиною сыновей Енномовых, но долиною убийства, и в Тофете будут хоронить по недостатку места.
JER|7|33|И будут трупы народа сего пищею птицам небесным и зверям земным, и некому будет отгонять их.
JER|7|34|И прекращу в городах Иудеи и на улицах Иерусалима голос торжества и голос веселия, голос жениха и голос невесты; потому что земля эта будет пустынею.
JER|8|1|В то время, говорит Господь, выбросят кости царей Иуды, и кости князей его, и кости священников, и кости пророков, и кости жителей Иерусалима из гробов их;
JER|8|2|и раскидают их пред солнцем и луною и пред всем воинством небесным, которых они любили и которым служили и в след которых ходили, которых искали и которым поклонялись; не уберут их и не похоронят: они будут навозом на земле.
JER|8|3|И будут смерть предпочитать жизни все остальные, которые останутся от этого злого племени во всех местах, куда Я изгоню их, говорит Господь Саваоф.
JER|8|4|И скажи им: так говорит Господь: разве, упав, не встают и, совратившись с дороги, не возвращаются?
JER|8|5|Для чего этот народ, Иерусалим, находится в упорном отступничестве? они крепко держатся обмана и не хотят обратиться.
JER|8|6|Я наблюдал и слушал: не говорят они правды, никто не раскаивается в своем нечестии, никто не говорит: "что я сделал?"; каждый обращается на свой путь, как конь, бросающийся в сражение.
JER|8|7|И аист под небом знает свои определенные времена, и горлица, и ласточка, и журавль наблюдают время, когда им прилететь; а народ Мой не знает определения Господня.
JER|8|8|Как вы говорите: "мы мудры, и закон Господень у нас"? А вот, лживая трость книжников [и его] превращает в ложь.
JER|8|9|Посрамились мудрецы, смутились и запутались в сеть: вот, они отвергли слово Господне; в чем же мудрость их?
JER|8|10|За то жен их отдам другим, поля их – иным владетелям; потому что все они, от малого до большого, предались корыстолюбию; от пророка до священника – все действуют лживо.
JER|8|11|И врачуют рану дочери народа Моего легкомысленно, говоря: "мир, мир!", а мира нет.
JER|8|12|Стыдятся ли они, делая мерзости? нет, они нисколько не стыдятся и не краснеют. За то падут они между падшими; во время посещения их будут повержены, говорит Господь.
JER|8|13|До конца оберу их, говорит Господь, не останется ни одной виноградины на лозе, ни смоквы на смоковнице, и лист опадет, и что Я дал им, отойдет от них.
JER|8|14|"Что мы сидим? собирайтесь, пойдем в укрепленные города, и там погибнем; ибо Господь Бог наш определил нас на погибель и дает нам пить воду с желчью за то, что мы грешили пред Господом".
JER|8|15|Ждем мира, а ничего доброго нет, – времени исцеления, и вот ужасы.
JER|8|16|От Дана слышен храп коней его, от громкого ржания жеребцов его дрожит вся земля; и придут и истребят землю и все, что на ней, город и живущих в нем.
JER|8|17|Ибо вот, Я пошлю на вас змеев, василисков, против которых нет заговариванья, и они будут уязвлять вас, говорит Господь.
JER|8|18|Когда утешусь я в горести моей! сердце мое изныло во мне.
JER|8|19|Вот, слышу вопль дщери народа Моего из дальней страны: разве нет Господа на Сионе? разве нет Царя его на нем? – Зачем они подвигли Меня на гнев своими идолами, чужеземными, ничтожными?
JER|8|20|Прошла жатва, кончилось лето, а мы не спасены.
JER|8|21|О сокрушении дщери народа моего я сокрушаюсь, хожу мрачен, ужас объял меня.
JER|8|22|Разве нет бальзама в Галааде? разве нет там врача? Отчего же нет исцеления дщери народа моего?
JER|8|23|О, кто даст голове моей воду и глазам моим – источник слез! я плакал бы день и ночь о пораженных дщери народа моего.
JER|9|1|О, кто даст голове моей воду и глазам моим--источник слез! я плакал бы день и ночь о пораженных дщери народа моего.
JER|9|2|О, кто дал бы мне в пустыне пристанище путников! оставил бы я народ мой и ушел бы от них: ибо все они прелюбодеи, скопище вероломных.
JER|9|3|Как лук, напрягают язык свой для лжи, усиливаются на земле неправдою; ибо переходят от одного зла к другому, и Меня не знают, говорит Господь.
JER|9|4|Берегитесь каждый своего друга, и не доверяйте ни одному из своих братьев; ибо всякий брат ставит преткновение другому, и всякий друг разносит клеветы.
JER|9|5|Каждый обманывает своего друга, и правды не говорят: приучили язык свой говорить ложь, лукавствуют до усталости.
JER|9|6|Ты живешь среди коварства; по коварству они отрекаются знать Меня, говорит Господь.
JER|9|7|Посему так говорит Господь Саваоф: вот, Я расплавлю и испытаю их; ибо как иначе Мне поступать со дщерью народа Моего?
JER|9|8|Язык их – убийственная стрела, говорит коварно; устами своими говорят с ближним своим дружелюбно, а в сердце своем строят ему ковы.
JER|9|9|Неужели Я не накажу их за это? говорит Господь; не отмстит ли душа Моя такому народу, как этот?
JER|9|10|О горах подниму плач и вопль, и о степных пастбищах – рыдание, потому что они выжжены, так что никто там не проходит, и не слышно блеяния стад: от птиц небесных до скота – [все] рассеялись, ушли.
JER|9|11|И сделаю Иерусалим грудою камней, жилищем шакалов, и города Иудеи сделаю пустынею, без жителей.
JER|9|12|Есть ли такой мудрец, который понял бы это? И к кому говорят уста Господни – объяснил бы, за что погибла страна и выжжена, как пустыня, так что никто не проходит [по ней]?
JER|9|13|И сказал Господь: за то, что они оставили закон Мой, который Я постановил для них, и не слушали гласа Моего и не поступали по нему;
JER|9|14|а ходили по упорству сердца своего и во след Ваалов, как научили их отцы их.
JER|9|15|Посему так говорит Господь Саваоф, Бог Израилев: вот, Я накормлю их, этот народ, полынью, и напою их водою с желчью;
JER|9|16|и рассею их между народами, которых не знали ни они, ни отцы их, и пошлю вслед их меч, доколе не истреблю их.
JER|9|17|Так говорит Господь Саваоф: подумайте, и позовите плакальщиц, чтобы они пришли; пошлите за искусницами [в этом деле], чтобы они пришли.
JER|9|18|Пусть они поспешат и поднимут плач о нас, чтобы из глаз наших лились слезы, и с ресниц наших текла вода.
JER|9|19|Ибо голос плача слышен с Сиона: "как мы ограблены! мы жестоко посрамлены, ибо оставляем землю, потому что разрушили жилища наши".
JER|9|20|Итак слушайте, женщины, слово Господа, и да внимает ухо ваше слову уст Его; и учите дочерей ваших плачу, и одна другую – плачевным песням.
JER|9|21|Ибо смерть входит в наши окна, вторгается в чертоги наши, чтобы истребить детей с улицы, юношей с площадей.
JER|9|22|Скажи: так говорит Господь: и будут повержены трупы людей, как навоз на поле и как снопы позади жнеца, и некому будет собрать их.
JER|9|23|Так говорит Господь: да не хвалится мудрый мудростью своею, да не хвалится сильный силою своею, да не хвалится богатый богатством своим.
JER|9|24|Но хвалящийся хвались тем, что разумеет и знает Меня, что Я – Господь, творящий милость, суд и правду на земле; ибо только это благоугодно Мне, говорит Господь.
JER|9|25|Вот, приходят дни, говорит Господь, когда Я посещу всех обрезанных и необрезанных:
JER|9|26|Египет и Иудею, и Едома и сыновей Аммоновых, и Моава и всех стригущих волосы на висках, обитающих в пустыне; ибо все эти народы необрезаны, а весь дом Израилев с необрезанным сердцем.
JER|10|1|Слушайте слово, которое Господь говорит вам, дом Израилев.
JER|10|2|Так говорит Господь: не учитесь путям язычников и не страшитесь знамений небесных, которых язычники страшатся.
JER|10|3|Ибо уставы народов – пустота: вырубают дерево в лесу, обделывают его руками плотника при помощи топора,
JER|10|4|покрывают серебром и золотом, прикрепляют гвоздями и молотом, чтобы не шаталось.
JER|10|5|Они – как обточенный столп, и не говорят; их носят, потому что ходить не могут. Не бойтесь их, ибо они не могут причинить зла, но и добра делать не в силах.
JER|10|6|Нет подобного Тебе, Господи! Ты велик, и имя Твое велико могуществом.
JER|10|7|Кто не убоится Тебя, Царь народов? ибо Тебе [единому] принадлежит это; потому что между всеми мудрецами народов и во всех царствах их нет подобного Тебе.
JER|10|8|Все до одного они бессмысленны и глупы; пустое учение – это дерево.
JER|10|9|Разбитое в листы серебро привезено из Фарсиса, золото – из Уфаза, дело художника и рук плавильщика; одежда на них – гиацинт и пурпур: все это – дело людей искусных.
JER|10|10|А Господь Бог есть истина; Он есть Бог живый и Царь вечный. От гнева Его дрожит земля, и народы не могут выдержать негодования Его.
JER|10|11|Так говорите им: боги, которые не сотворили неба и земли, исчезнут с земли и из–под небес.
JER|10|12|Он сотворил землю силою Своею, утвердил вселенную мудростью Своею и разумом Своим распростер небеса.
JER|10|13|По гласу Его шумят воды на небесах, и Он возводит облака от краев земли, творит молнии среди дождя и изводит ветер из хранилищ Своих.
JER|10|14|Безумствует всякий человек в своем знании, срамит себя всякий плавильщик истуканом [своим], ибо выплавленное им есть ложь, и нет в нем духа.
JER|10|15|Это совершенная пустота, дело заблуждения; во время посещения их они исчезнут.
JER|10|16|Не такова, как их, доля Иакова; ибо [Бог его] есть Творец всего, и Израиль есть жезл наследия Его; имя Его – Господь Саваоф.
JER|10|17|Убирай с земли имущество твое, имеющая сидеть в осаде;
JER|10|18|ибо так говорит Господь: вот, Я выброшу жителей сей земли на сей раз и загоню их в тесное место, чтобы схватили их.
JER|10|19|Горе мне в моем сокрушении; мучительна рана моя, но я говорю [сам] [в себе]: "подлинно, это моя скорбь, и я буду нести ее;
JER|10|20|шатер мой опустошен, и все веревки мои порваны; дети мои ушли от меня, и нет их: некому уже раскинуть шатра моего и развесить ковров моих,
JER|10|21|ибо пастыри сделались бессмысленными и не искали Господа, а потому они и поступали безрассудно, и все стадо их рассеяно".
JER|10|22|Несется слух: вот он идет, и большой шум от страны северной, чтобы города Иудеи сделать пустынею, жилищем шакалов.
JER|10|23|Знаю, Господи, что не в воле человека путь его, что не во власти идущего давать направление стопам своим.
JER|10|24|Наказывай меня, Господи, но по правде, не во гневе Твоем, чтобы не умалить меня.
JER|10|25|Излей ярость Твою на народы, которые не знают Тебя, и на племена, которые не призывают имени Твоего; ибо они съели Иакова, пожрали его и истребили его, и жилище его опустошили.
JER|11|1|Слово, которое было к Иеремии от Господа:
JER|11|2|слушайте слова завета сего и скажите мужам Иуды и жителям Иерусалима;
JER|11|3|и скажи им: так говорит Господь, Бог Израилев: проклят человек, который не послушает слов завета сего,
JER|11|4|который Я заповедал отцам вашим, когда вывел их из земли Египетской, из железной печи, сказав: "слушайтесь гласа Моего и делайте все, что Я заповедаю вам, – и будете Моим народом, и Я буду вашим Богом,
JER|11|5|чтобы исполнить клятву, которою Я клялся отцам вашим – дать им землю, текущую молоком и медом, как это ныне". И отвечал я, сказав: аминь, Господи!
JER|11|6|И сказал мне Господь: провозгласи все сии слова в городах Иуды и на улицах Иерусалима и скажи: слушайте слова завета сего и исполняйте их.
JER|11|7|Ибо отцов ваших Я увещевал постоянно с того дня, как вывел их из земли Египетской, до сего дня; увещевал их с раннего утра, говоря: "слушайтесь гласа Моего".
JER|11|8|Но они не слушались и не приклоняли уха своего, а ходили каждый по упорству злого сердца своего: поэтому Я навел на них все сказанное в завете сем, который Я заповедал им исполнять, а они не исполняли.
JER|11|9|И сказал мне Господь: есть заговор между мужами Иуды и жителями Иерусалима:
JER|11|10|они опять обратились к беззакониям праотцев своих, которые отреклись слушаться слов Моих и пошли вослед чужих богов, служа им. Дом Израиля и дом Иуды нарушили завет Мой, который Я заключил с отцами их.
JER|11|11|Посему так говорит Господь: вот, Я наведу на них бедствие, от которого они не могут избавиться, и когда воззовут ко Мне, не услышу их.
JER|11|12|Тогда города Иуды и жители Иерусалима пойдут и воззовут к богам, которым они кадят; но они нисколько не помогут им во время бедствия их.
JER|11|13|Ибо сколько у тебя городов, столько и богов у тебя, Иуда, и сколько улиц в Иерусалиме, столько вы наставили жертвенников постыдному, жертвенников для каждения Ваалу.
JER|11|14|Ты же не проси за этот народ и не возноси за них молитвы и прошений; ибо Я не услышу, когда они будут взывать ко Мне в бедствии своем.
JER|11|15|Что возлюбленному Моему в доме Моем, когда в нем совершаются многие непотребства? и священные мяса не помогут тебе, когда, делая зло, ты радуешься.
JER|11|16|Зеленеющею маслиною, красующеюся приятными плодами, именовал тебя Господь. А ныне, при шуме сильного смятения, Он воспламенил огонь вокруг нее, и сокрушились ветви ее.
JER|11|17|Господь Саваоф, Который насадил тебя, изрек на тебя злое за зло дома Израилева и дома Иудина, которое они причинили себе тем, что подвигли Меня на гнев каждением Ваалу.
JER|11|18|Господь открыл мне, и я знаю; Ты показал мне деяния их.
JER|11|19|А я, как кроткий агнец, ведомый на заклание, и не знал, что они составляют замыслы против меня, [говоря]: "положим [ядовитое] дерево в пищу его и отторгнем его от земли живых, чтобы и имя его более не упоминалось".
JER|11|20|Но, Господи Саваоф, Судия праведный, испытующий сердца и утробы! дай увидеть мне мщение Твое над ними, ибо Тебе вверил я дело мое.
JER|11|21|Посему так говорит Господь о мужах Анафофа, ищущих души твоей и говорящих: "не пророчествуй во имя Господа, чтобы не умереть тебе от рук наших";
JER|11|22|посему так говорит Господь Саваоф: вот, Я посещу их: юноши [их] умрут от меча; сыновья их и дочери их умрут от голода.
JER|11|23|И остатка не будет от них; ибо Я наведу бедствие на мужей Анафофа в год посещения их.
JER|12|1|Праведен будешь Ты, Господи, если я стану судиться с Тобою; и однако же буду говорить с Тобою о правосудии: почему путь нечестивых благоуспешен, и все вероломные благоденствуют?
JER|12|2|Ты насадил их, и они укоренились, выросли и приносят плод. В устах их Ты близок, но далек от сердца их.
JER|12|3|А меня, Господи, Ты знаешь, видишь меня и испытываешь сердце мое, каково оно к Тебе. Отдели их, как овец на заклание, и приготовь их на день убиения.
JER|12|4|Долго ли будет сетовать земля, и трава на всех полях – сохнуть? скот и птицы гибнут за нечестие жителей ее, ибо они говорят: "Он не увидит, что с нами будет".
JER|12|5|Если ты с пешими бежал, и они утомили тебя, как же тебе состязаться с конями? и если в стране мирной ты был безопасен, то что будешь делать в наводнение Иордана?
JER|12|6|Ибо и братья твои и дом отца твоего, и они вероломно поступают с тобою, и они кричат вслед тебя громким голосом. Не верь им, когда они говорят тебе и доброе.
JER|12|7|Я оставил дом Мой; покинул удел Мой; самое любезное для души Моей отдал в руки врагов его.
JER|12|8|Удел Мой сделался для Меня как лев в лесу; возвысил на Меня голос свой: за то Я возненавидел его.
JER|12|9|Удел Мой стал у Меня, как разноцветная птица, на которую со всех сторон напали другие хищные птицы. Идите, собирайтесь, все полевые звери: идите пожирать его.
JER|12|10|Множество пастухов испортили Мой виноградник, истоптали ногами участок Мой; любимый участок Мой сделали пустою степью;
JER|12|11|сделали его пустынею, и в запустении он плачет предо Мною; вся земля опустошена, потому что ни один человек не прилагает этого к сердцу.
JER|12|12|На все горы в пустыне пришли опустошители; ибо меч Господа пожирает [все] от одного края земли до другого: нет мира ни для какой плоти.
JER|12|13|Они сеяли пшеницу, а пожали терны; измучились, и не получили никакой пользы; постыдитесь же таких прибытков ваших по причине пламенного гнева Господа.
JER|12|14|Так говорит Господь обо всех злых Моих соседях, нападающих на удел, который Я дал в наследие народу Моему, Израилю: вот, Я исторгну их из земли их, и дом Иудин исторгну из среды их.
JER|12|15|Но после того, как Я исторгну их, снова возвращу и помилую их, и приведу каждого в удел его и каждого в землю его.
JER|12|16|И если они научатся путям народа Моего, чтобы клясться именем Моим: "жив Господь!", как они научили народ Мой клясться Ваалом, то водворятся среди народа Моего.
JER|12|17|Если же не послушаются, то Я искореню и совершенно истреблю такой народ, говорит Господь.
JER|13|1|Так сказал мне Господь: пойди, купи себе льняной пояс и положи его на чресла твои, но в воду не клади его.
JER|13|2|И я купил пояс, по слову Господню, и положил его на чресла мои.
JER|13|3|И было ко мне слово Господне в другой раз, и сказано:
JER|13|4|возьми пояс, который ты купил, который на чреслах твоих, и встань, пойди к Евфрату и спрячь его там в расселине скалы.
JER|13|5|Я пошел и спрятал его у Евфрата, как повелел мне Господь.
JER|13|6|По прошествии же многих дней сказал мне Господь: встань, пойди к Евфрату и возьми оттуда пояс, который Я велел тебе спрятать там.
JER|13|7|И я пришел к Евфрату, выкопал и взял пояс из того места, где спрятал его, и вот, пояс был испорчен, ни к чему стал не годен.
JER|13|8|И было ко мне слово Господне:
JER|13|9|так говорит Господь: так сокрушу Я гордость Иуды и великую гордость Иерусалима.
JER|13|10|Этот негодный народ, который не хочет слушать слов Моих, живет по упорству сердца своего и ходит во след иных богов, чтобы служить им и поклоняться им, будет как этот пояс, который ни к чему не годен.
JER|13|11|Ибо, как пояс близко лежит к чреслам человека, так Я приблизил к Себе весь дом Израилев и весь дом Иудин, говорит Господь, чтобы они были Моим народом и Моею славою, хвалою и украшением; но они не послушались.
JER|13|12|Посему скажи им слово сие: так говорит Господь, Бог Израилев: всякий винный мех наполняется вином. Они скажут тебе: "разве мы не знаем, что всякий винный мех наполняется вином?"
JER|13|13|А ты скажи им: так говорит Господь: вот, Я наполню вином до опьянения всех жителей сей земли и царей, сидящих на престоле Давида, и священников, и пророков и всех жителей Иерусалима,
JER|13|14|и сокрушу их друг о друга, и отцов и сыновей вместе, говорит Господь; не пощажу и не помилую, и не пожалею истребить их.
JER|13|15|Слушайте и внимайте; не будьте горды, ибо Господь говорит.
JER|13|16|Воздайте славу Господу Богу вашему, доколе Он еще не навел темноты, и доколе еще ноги ваши не спотыкаются на горах мрака: тогда вы будете ожидать света, а Он обратит его в тень смерти и сделает тьмою.
JER|13|17|Если же вы не послушаете сего, то душа моя в сокровенных местах будет оплакивать гордость вашу, будет плакать горько, и глаза мои будут изливаться в слезах; потому что стадо Господне отведено будет в плен.
JER|13|18|Скажи царю и царице: смиритесь, сядьте пониже, ибо упал с головы вашей венец славы вашей.
JER|13|19|Южные города заперты, и некому отворять их; Иуда весь отводится в плен, отводится в плен весь совершенно.
JER|13|20|Поднимите глаза ваши и посмотрите на идущих от севера: где стадо, которое дано было тебе, прекрасное стадо твое?
JER|13|21|Что скажешь, [дочь Сиона], когда Он посетит тебя? Ты сама приучила их начальствовать над тобою; не схватят ли тебя боли, как рождающую женщину?
JER|13|22|И если скажешь в сердце твоем: "за что постигло меня это?" – За множество беззаконий твоих открыт подол у тебя, обнажены пяты твои.
JER|13|23|Может ли Ефиоплянин переменить кожу свою и барс – пятна свои? так и вы можете ли делать доброе, привыкнув делать злое?
JER|13|24|Поэтому развею их, как прах, разносимый ветром пустынным.
JER|13|25|Вот жребий твой, отмеренная тебе от Меня часть, говорит Господь, потому что ты забыла Меня и надеялась на ложь.
JER|13|26|За то будет поднят подол твой на лице твое, чтобы открылся срам твой.
JER|13|27|Видел Я прелюбодейство твое и неистовые похотения твои, твои непотребства и твои мерзости на холмах в поле. Горе тебе, Иерусалим! ты и после сего не очистишься. Доколе же?
JER|14|1|Слово Господа, которое было к Иеремии по случаю бездождия.
JER|14|2|Плачет Иуда, ворота его распались, почернели на земле, и вопль поднимается в Иерусалиме.
JER|14|3|Вельможи посылают слуг своих за водою; они приходят к колодезям и не находят воды; возвращаются с пустыми сосудами; пристыженные и смущенные, они покрывают свои головы.
JER|14|4|Так как почва растрескалась от того, что не было дождя на землю, то и земледельцы в смущении и покрывают свои головы.
JER|14|5|Даже и лань рождает на поле и оставляет [детей], потому что нет травы.
JER|14|6|И дикие ослы стоят на возвышенных местах и глотают, подобно шакалам, воздух; глаза их потускли, потому что нет травы.
JER|14|7|Хотя беззакония наши свидетельствуют против нас, но Ты, Господи, твори с нами ради имени Твоего; отступничество наше велико, согрешили мы пред Тобою.
JER|14|8|Надежда Израиля, Спаситель его во время скорби! Для чего Ты – как чужой в этой земле, как прохожий, который зашел переночевать?
JER|14|9|Для чего Ты – как человек изумленный, как сильный, не имеющий силы спасти? И однако же Ты, Господи, посреди нас, и Твое имя наречено над нами; не оставляй нас.
JER|14|10|Так говорит Господь народу сему: за то, что они любят бродить, не удерживают ног своих, за то Господь не благоволит к ним, припоминает ныне беззакония их и наказывает грехи их.
JER|14|11|И сказал мне Господь: ты не молись о народе сем во благо ему.
JER|14|12|Если они будут поститься, Я не услышу вопля их; и если вознесут всесожжение и дар, не приму их; но мечом и голодом, и моровою язвою истреблю их.
JER|14|13|Тогда сказал я: Господи Боже! вот, пророки говорят им: "не увидите меча, и голода не будет у вас, но постоянный мир дам вам на сем месте".
JER|14|14|И сказал мне Господь: пророки пророчествуют ложное именем Моим; Я не посылал их и не давал им повеления, и не говорил им; они возвещают вам видения ложные и гадания, и пустое и мечты сердца своего.
JER|14|15|Поэтому так говорит Господь о пророках: они пророчествуют именем Моим, а Я не посылал их; они говорят: "меча и голода не будет на сей земле": мечом и голодом будут истреблены эти пророки,
JER|14|16|и народ, которому они пророчествуют, разбросан будет по улицам Иерусалима от голода и меча, и некому будет хоронить их, – они и жены их, и сыновья их, и дочери их; и Я изолью на них зло их.
JER|14|17|И скажи им слово сие: да льются из глаз моих слезы ночь и день, и да не перестают; ибо великим поражением поражена дева, дочь народа моего, тяжким ударом.
JER|14|18|Выхожу я на поле, – и вот, убитые мечом; вхожу в город, – и вот истаевающие от голода; даже и пророк и священник бродят по земле бессознательно.
JER|14|19|Разве Ты совсем отверг Иуду? Разве душе Твоей опротивел Сион? Для чего поразил нас так, что нет нам исцеления? Ждем мира, и ничего доброго нет; ждем времени исцеления, и вот ужасы.
JER|14|20|Сознаем, Господи, нечестие наше, беззаконие отцов наших; ибо согрешили мы пред Тобою.
JER|14|21|Не отрини [нас] ради имени Твоего; не унижай престола славы Твоей: вспомни, не разрушай завета Твоего с нами.
JER|14|22|Есть ли между суетными [богами] языческими производящие дождь? или может ли небо [само собою] подавать ливень? не Ты ли это, Господи, Боже наш? На Тебя надеемся мы; ибо Ты творишь все это.
JER|15|1|И сказал мне Господь: хотя бы предстали пред лице Мое Моисей и Самуил, душа Моя не [приклонится] к народу сему; отгони [их] от лица Моего, пусть они отойдут.
JER|15|2|Если же скажут тебе: "куда нам идти?", то скажи им: так говорит Господь: кто [обречен] на смерть, иди на смерть; и кто под меч, – под меч; и кто на голод, – на голод; и кто в плен, – в плен.
JER|15|3|И пошлю на них четыре рода [казней], говорит Господь: меч, чтобы убивать, и псов, чтобы терзать, и птиц небесных и зверей полевых, чтобы пожирать и истреблять;
JER|15|4|и отдам их на озлобление всем царствам земли за Манассию, сына Езекии, царя Иудейского, за то, что он сделал в Иерусалиме.
JER|15|5|Ибо кто пожалеет о тебе, Иерусалим? и кто окажет сострадание к тебе? и кто зайдет к тебе спросить о твоем благосостоянии?
JER|15|6|Ты оставил Меня, говорит Господь, отступил назад; поэтому Я простру на тебя руку Мою и погублю тебя: Я устал миловать.
JER|15|7|Я развеваю их веялом за ворота земли; лишаю их детей, гублю народ Мой; но они не возвращаются с путей своих.
JER|15|8|Вдов их у Меня более, нежели песку в море; наведу на них, на мать юношей, опустошителя в полдень; нападет на них внезапно страх и ужас.
JER|15|9|Лежит в изнеможении родившая семерых, испускает дыхание свое; еще днем закатилось солнце ее, она постыжена и посрамлена. И остаток их предам мечу пред глазами врагов их, говорит Господь.
JER|15|10|"Горе мне, мать моя, что ты родила меня человеком, который спорит и ссорится со всею землею! никому не давал я в рост, и мне никто не давал в рост, [а] все проклинают меня".
JER|15|11|Господь сказал: конец твой будет хорош, и Я заставлю врага поступать с тобою хорошо во время бедствия и во время скорби.
JER|15|12|Может ли железо сокрушить железо северное и медь?
JER|15|13|Имущество твое и сокровища твои отдам на расхищение, без платы, за все грехи твои, во всех пределах твоих;
JER|15|14|и отправлю с врагами твоими в землю, которой ты не знаешь; ибо огонь возгорелся в гневе Моем, – будет пылать на вас.
JER|15|15|О, Господи! Ты знаешь [все]; вспомни обо мне и посети меня, и отмсти за меня гонителям моим; не погуби меня по долготерпению Твоему; Ты знаешь, что ради Тебя несу я поругание.
JER|15|16|Обретены слова Твои, и я съел их; и было слово Твое мне в радость и в веселие сердца моего; ибо имя Твое наречено на мне, Господи, Боже Саваоф.
JER|15|17|Не сидел я в собрании смеющихся и не веселился: под тяготеющею на мне рукою Твоею я сидел одиноко, ибо Ты исполнил меня негодования.
JER|15|18|За что так упорна болезнь моя, и рана моя так неисцельна, что отвергает врачевание? Неужели Ты будешь для меня как бы обманчивым источником, неверною водою?
JER|15|19|На сие так сказал Господь: если ты обратишься, то Я восставлю тебя, и будешь предстоять пред лицем Моим; и если извлечешь драгоценное из ничтожного, то будешь как Мои уста. Они сами будут обращаться к тебе, а не ты будешь обращаться к ним.
JER|15|20|И сделаю тебя для этого народа крепкою медною стеною; они будут ратовать против тебя, но не одолеют тебя, ибо Я с тобою, чтобы спасать и избавлять тебя, говорит Господь.
JER|15|21|И спасу тебя от руки злых и избавлю тебя от руки притеснителей.
JER|16|1|И было ко мне слово Господне:
JER|16|2|не бери себе жены, и пусть не будет у тебя ни сыновей, ни дочерей на месте сем.
JER|16|3|Ибо так говорит Господь о сыновьях и дочерях, которые родятся на месте сем, и о матерях их, которые родят их, и об отцах их, которые произведут их на сей земле:
JER|16|4|тяжкими смертями умрут они и не будут ни оплаканы, ни похоронены; будут навозом на поверхности земли; мечом и голодом будут истреблены, и трупы их будут пищею птицам небесным и зверям земным.
JER|16|5|Ибо так говорит Господь: не входи в дом сетующих и не ходи плакать и жалеть с ними; ибо Я отнял от этого народа, говорит Господь, мир Мой и милость и сожаление.
JER|16|6|И умрут великие и малые на земле сей; и не будут погребены, и не будут оплакивать их, ни терзать себя, ни стричься ради них.
JER|16|7|И не будут преломлять для них хлеб в печали, в утешение об умершем; и не подадут им чаши утешения, чтобы пить по отце их и матери их.
JER|16|8|Не ходи также и в дом пиршества, чтобы сидеть с ними, есть и пить;
JER|16|9|ибо так говорит Господь Саваоф, Бог Израилев: вот, Я прекращу на месте сем в глазах ваших и во дни ваши голос радости и голос веселья, голос жениха и голос невесты.
JER|16|10|Когда ты перескажешь народу сему все эти слова, и они скажут тебе: "за что изрек на нас Господь все это великое бедствие, и какая наша неправда, и какой наш грех, которым согрешили мы пред Господом Богом нашим?" –
JER|16|11|тогда скажи им: за то, что отцы ваши оставили Меня, говорит Господь, и пошли вослед иных богов, и служили им, и поклонялись им, а Меня оставили, и закона Моего не хранили.
JER|16|12|А вы поступаете еще хуже отцов ваших и живете каждый по упорству злого сердца своего, чтобы не слушать Меня.
JER|16|13|За это выброшу вас из земли сей в землю, которой не знали ни вы, ни отцы ваши, и там будете служить иным богам день и ночь; ибо Я не окажу вам милосердия.
JER|16|14|Посему вот, приходят дни, говорит Господь, когда не будут уже говорить: "жив Господь, Который вывел сынов Израилевых из земли Египетской";
JER|16|15|но: "жив Господь, Который вывел сынов Израилевых из земли северной и из всех земель, в которые изгнал их": ибо возвращу их в землю их, которую Я дал отцам их.
JER|16|16|Вот, Я пошлю множество рыболовов, говорит Господь, и будут ловить их; а потом пошлю множество охотников, и они погонят их со всякой горы, и со всякого холма, и из ущелий скал.
JER|16|17|Ибо очи Мои на всех путях их; они не скрыты от лица Моего, и неправда их не сокрыта от очей Моих.
JER|16|18|И воздам им прежде всего за неправду их и за сугубый грех их, потому что осквернили землю Мою, трупами гнусных своих и мерзостями своими наполнили наследие Мое.
JER|16|19|Господи, сила моя и крепость моя и прибежище мое в день скорби! к Тебе придут народы от краев земли и скажут: "только ложь наследовали наши отцы, пустоту и то, в чем никакой нет пользы".
JER|16|20|Может ли человек сделать себе богов, которые впрочем не боги?
JER|16|21|Посему, вот Я покажу им ныне, покажу им руку Мою и могущество Мое, и узнают, что имя Мое – Господь.
JER|17|1|Грех Иуды написан железным резцом, алмазным острием начертан на скрижали сердца их и на рогах жертвенников их.
JER|17|2|Как о сыновьях своих, воспоминают они о жертвенниках своих и дубравах своих у зеленых дерев, на высоких холмах.
JER|17|3|Гору Мою в поле, имущество твое и все сокровища твои отдам на расхищение, и все высоты твои – за грехи во всех пределах твоих.
JER|17|4|И ты чрез себя лишишься наследия твоего, которое Я дал тебе, и отдам тебя в рабство врагам твоим, в землю, которой ты не знаешь, потому что вы воспламенили огонь гнева Моего; он будет гореть вовеки.
JER|17|5|Так говорит Господь: проклят человек, который надеется на человека и плоть делает своею опорою, и которого сердце удаляется от Господа.
JER|17|6|Он будет как вереск в пустыне и не увидит, когда придет доброе, и поселится в местах знойных в степи, на земле бесплодной, необитаемой.
JER|17|7|Благословен человек, который надеется на Господа, и которого упование – Господь.
JER|17|8|Ибо он будет как дерево, посаженное при водах и пускающее корни свои у потока; не знает оно, когда приходит зной; лист его зелен, и во время засухи оно не боится и не перестает приносить плод.
JER|17|9|Лукаво сердце [человеческое] более всего и крайне испорчено; кто узнает его?
JER|17|10|Я, Господь, проникаю сердце и испытываю внутренности, чтобы воздать каждому по пути его и по плодам дел его.
JER|17|11|Куропатка садится на яйца, которых не несла; таков приобретающий богатство неправдою: он оставит его на половине дней своих, и глупцом останется при конце своем.
JER|17|12|Престол славы, возвышенный от начала, есть место освящения нашего.
JER|17|13|Ты, Господи, надежда Израилева; все, оставляющие Тебя, посрамятся. "Отступающие от Меня будут написаны на прахе, потому что оставили Господа, источник воды живой".
JER|17|14|Исцели меня, Господи, и исцелен буду; спаси меня, и спасен буду; ибо Ты хвала моя.
JER|17|15|Вот, они говорят мне: "где слово Господне? пусть оно придет!"
JER|17|16|Я не спешил быть пастырем у Тебя и не желал бедственного дня, Ты это знаешь; что вышло из уст моих, открыто пред лицем Твоим.
JER|17|17|Не будь страшен для меня, Ты – надежда моя в день бедствия.
JER|17|18|Пусть постыдятся гонители мои, а я не буду постыжен; пусть они вострепещут, а я буду бестрепетен; наведи на них день бедствия и сокруши их сугубым сокрушением.
JER|17|19|Так сказал мне Господь: пойди и стань в воротах сынов народа, которыми входят цари Иудейские и которыми они выходят, и во всех воротах Иерусалимских,
JER|17|20|и говори им: слушайте слово Господне, цари Иудейские, и вся Иудея, и все жители Иерусалима, входящие сими воротами.
JER|17|21|Так говорит Господь: берегите души свои и не носите нош в день субботний и не вносите их воротами Иерусалимскими,
JER|17|22|и не выносите нош из домов ваших в день субботний, и не занимайтесь никакою работою, но святите день субботний так, как Я заповедал отцам вашим,
JER|17|23|которые впрочем не послушались и не приклонили уха своего, но сделались жестоковыйными, чтобы не слушать и не принимать наставления.
JER|17|24|И если вы послушаете Меня в том, говорит Господь, чтобы не носить нош воротами сего города в день субботний и чтобы святить субботу, не занимаясь в этот день никакою работою,
JER|17|25|то воротами сего города будут входить цари и князья, сидящие на престоле Давида, ездящие на колесницах и на конях, они и князья их, Иудеи и жители Иерусалима, и город сей будет обитаем вечно.
JER|17|26|И будут приходить из городов Иудейских, и из окрестностей Иерусалима, и из земли Вениаминовой, и с равнины и с гор и с юга, и приносить всесожжение и жертву, и хлебное приношение, и ливан, и благодарственные жертвы в дом Господень.
JER|17|27|А если не послушаете Меня в том, чтобы святить день субботний и не носить нош, входя в ворота Иерусалима в день субботний, то возжгу огонь в воротах его, и он пожрет чертоги Иерусалима и не погаснет.
JER|18|1|Слово, которое было к Иеремии от Господа:
JER|18|2|встань и сойди в дом горшечника, и там Я возвещу тебе слова Мои.
JER|18|3|И сошел я в дом горшечника, и вот, он работал свою работу на кружале.
JER|18|4|И сосуд, который горшечник делал из глины, развалился в руке его; и он снова сделал из него другой сосуд, какой горшечнику вздумалось сделать.
JER|18|5|И было слово Господне ко мне:
JER|18|6|не могу ли Я поступить с вами, дом Израилев, подобно горшечнику сему? говорит Господь. Вот, что глина в руке горшечника, то вы в Моей руке, дом Израилев.
JER|18|7|Иногда Я скажу о каком–либо народе и царстве, что искореню, сокрушу и погублю его;
JER|18|8|но если народ этот, на который Я это изрек, обратится от своих злых дел, Я отлагаю то зло, которое помыслил сделать ему.
JER|18|9|А иногда скажу о каком–либо народе и царстве, что устрою и утвержу его;
JER|18|10|но если он будет делать злое пред очами Моими и не слушаться гласа Моего, Я отменю то добро, которым хотел облагодетельствовать его.
JER|18|11|Итак скажи мужам Иуды и жителям Иерусалима: так говорит Господь: вот, Я готовлю вам зло и замышляю против вас; итак обратитесь каждый от злого пути своего и исправьте пути ваши и поступки ваши.
JER|18|12|Но они говорят: "не надейся; мы будем жить по своим помыслам и будем поступать каждый по упорству злого своего сердца".
JER|18|13|Посему так говорит Господь: спросите между народами, слыхал ли кто подобное сему? крайне гнусные дела совершила дева Израилева.
JER|18|14|Оставляет ли снег Ливанский скалу горы? и иссякают ли из других мест текущие холодные воды?
JER|18|15|А народ Мой оставил Меня; они кадят суетным, споткнулись на путях своих, оставили пути древние, чтобы ходить по стезям пути непроложенного,
JER|18|16|чтобы сделать землю свою ужасом, всегдашним посмеянием, так что каждый, проходящий по ней, изумится и покачает головою своею.
JER|18|17|Как восточным ветром развею их пред лицем врага; спиною, а не лицем обращусь к ним в день бедствия их.
JER|18|18|А они сказали: "придите, составим замысел против Иеремии; ибо не исчез же закон у священника и совет у мудрого, и слово у пророка; придите, сразим его языком и не будем внимать словам его".
JER|18|19|Внемли мне, Господи, и услышь голос моих противников.
JER|18|20|Должно ли воздавать злом за добро? а они роют яму душе моей. Вспомни, что я стою пред лицем Твоим, чтобы говорить за них доброе, чтобы отвратить от них гнев Твой.
JER|18|21|Итак предай сыновей их голоду и подвергни их мечу; да будут жены их бездетными и вдовами, и мужья их да будут поражены смертью, и юноши их умерщвлены мечом на войне.
JER|18|22|Да будет слышен вопль из домов их, когда приведешь на них полки внезапно; ибо они роют яму, чтобы поймать меня, и тайно расставили сети для ног моих.
JER|18|23|Но Ты, Господи, знаешь все замыслы их против меня, чтобы умертвить меня; не прости неправды их и греха их не изгладь пред лицем Твоим; да будут они низвержены пред Тобою; поступи с ними во время гнева Твоего.
JER|19|1|Так сказал Господь: пойди и купи глиняный кувшин у горшечника; и возьми с собою старейших из народа и из старейшин священнических,
JER|19|2|и выйди в долину сыновей Енномовых, которая у ворот Харшиф, и провозгласи там слова, которые скажу тебе,
JER|19|3|и скажи: слушайте слово Господне, цари Иудейские и жители Иерусалима! так говорит Господь Саваоф, Бог Израилев: вот, Я наведу бедствие на место сие, – о котором кто услышит, у того зазвенит в ушах,
JER|19|4|за то, что они оставили Меня и чужим сделали место сие и кадят на нем иным богам, которых не знали ни они, ни отцы их, ни цари Иудейские; наполнили место сие кровью невинных
JER|19|5|и устроили высоты Ваалу, чтобы сожигать сыновей своих огнем во всесожжение Ваалу, чего Я не повелевал и не говорил, и что на мысль не приходило Мне;
JER|19|6|за то вот, приходят дни, говорит Господь, когда место сие не будет более называться Тофетом или долиною сыновей Енномовых, но долиною убиения.
JER|19|7|И уничтожу совет Иуды и Иерусалима на месте сем и сражу их мечом пред лицем врагов их и рукою ищущих души их, и отдам трупы их в пищу птицам небесным и зверям земным.
JER|19|8|И сделаю город сей ужасом и посмеянием; каждый, проходящий через него, изумится и посвищет, смотря на все язвы его.
JER|19|9|И накормлю их плотью сыновей их и плотью дочерей их; и будет каждый есть плоть своего ближнего, находясь в осаде и тесноте, когда стеснят их враги их и ищущие души их.
JER|19|10|И разбей кувшин пред глазами тех мужей, которые придут с тобою,
JER|19|11|и скажи им: так говорит Господь Саваоф: так сокрушу Я народ сей и город сей, как сокрушен горшечников сосуд, который уже не может быть восстановлен, и будут хоронить их в Тофете, по недостатку места для погребения.
JER|19|12|Так поступлю с местом сим, говорит Господь, и с жителями его; и город сей сделаю подобным Тофету.
JER|19|13|И домы Иерусалима и домы царей Иудейских будут, как место Тофет, нечистыми, потому что на кровлях всех домов кадят всему воинству небесному и совершают возлияния богам чужим.
JER|19|14|И пришел Иеремия с Тофета, куда Господь посылал его пророчествовать, и стал на дворе дома Господня и сказал всему народу:
JER|19|15|так говорит Господь Саваоф, Бог Израилев: вот, Я наведу на город сей и на все города его все то бедствие, которое изрек на него, потому что они жестоковыйны и не слушают слов Моих.
JER|20|1|Когда Пасхор, сын Еммеров, священник, он же и надзиратель в доме Господнем, услышал, что Иеремия пророчески произнес слова сии,
JER|20|2|то ударил Пасхор Иеремию пророка и посадил его в колоду, которая была у верхних ворот Вениаминовых при доме Господнем.
JER|20|3|Но на другой день Пасхор выпустил Иеремию из колоды, и Иеремия сказал ему: не "Пасхор" нарек Господь имя тебе, но "Магор Миссавив".
JER|20|4|Ибо так говорит Господь: вот, Я сделаю тебя ужасом для тебя самого и для всех друзей твоих, и падут они от меча врагов своих, и твои глаза увидят это. И всего Иуду предам в руки царя Вавилонского, и отведет их в Вавилон и поразит их мечом.
JER|20|5|И предам все богатство этого города и все стяжание его, и все драгоценности его; и все сокровища царей Иудейских отдам в руки врагов их, и разграбят их и возьмут, и отправят их в Вавилон.
JER|20|6|И ты, Пасхор, и все живущие в доме твоем, пойдете в плен; и придешь в Вавилон, и там умрешь, и там будешь похоронен, ты и все друзья твои, которым ты пророчествовал ложно.
JER|20|7|Ты влек меня, Господи, – и я увлечен; Ты сильнее меня – и превозмог, и я каждый день в посмеянии, всякий издевается надо мною.
JER|20|8|Ибо лишь только начну говорить я, – кричу о насилии, вопию о разорении, потому что слово Господне обратилось в поношение мне и в повседневное посмеяние.
JER|20|9|И подумал я: "не буду я напоминать о Нем и не буду более говорить во имя Его"; но было в сердце моем, как бы горящий огонь, заключенный в костях моих, и я истомился, удерживая его, и не мог.
JER|20|10|Ибо я слышал толки многих: угрозы вокруг; "заявите, [говорили] [они], и мы сделаем донос". Все, жившие со мною в мире, сторожат за мною, не споткнусь ли я: "может быть, [говорят], он попадется, и мы одолеем его и отмстим ему".
JER|20|11|Но со мною Господь, как сильный ратоборец; поэтому гонители мои споткнутся и не одолеют; сильно посрамятся, потому что поступали неразумно; посрамление будет вечное, никогда не забудется.
JER|20|12|Господи сил! Ты испытываешь праведного и видишь внутренность и сердце. Да увижу я мщение Твое над ними, ибо Тебе вверил я дело мое.
JER|20|13|Пойте Господу, хвалите Господа, ибо Он спасает душу бедного от руки злодеев. –
JER|20|14|Проклят день, в который я родился! день, в который родила меня мать моя, да не будет благословен!
JER|20|15|Проклят человек, который принес весть отцу моему и сказал: "у тебя родился сын", [и] тем очень обрадовал его.
JER|20|16|И да будет с тем человеком, что с городами, которые разрушил Господь и не пожалел; да слышит он утром вопль и в полдень рыдание
JER|20|17|за то, что он не убил меня в самой утробе – так, чтобы мать моя была мне гробом, и чрево ее оставалось вечно беременным.
JER|20|18|Для чего вышел я из утробы, чтобы видеть труды и скорби, и чтобы дни мои исчезали в бесславии?
JER|21|1|Слово, которое было к Иеремии от Господа, когда царь Седекия прислал к нему Пасхора, сына Молхиина, и Софонию, сына Маасеи священника, сказать [ему]:
JER|21|2|"вопроси о нас Господа, ибо Навуходоносор, царь Вавилонский, воюет против нас; может быть, Господь сотворит с нами что–либо такое, как все чудеса Его, чтобы тот отступил от нас".
JER|21|3|И сказал им Иеремия: так скажите Седекии:
JER|21|4|так говорит Господь, Бог Израилев: вот, Я обращу назад воинские орудия, которые в руках ваших, которыми вы сражаетесь с царем Вавилонским и с Халдеями, осаждающими вас вне стены, и соберу оные посреди города сего;
JER|21|5|и Сам буду воевать против вас рукою простертою и мышцею крепкою, во гневе и в ярости и в великом негодовании;
JER|21|6|и поражу живущих в сем городе – и людей и скот; от великой язвы умрут они.
JER|21|7|А после того, говорит Господь, Седекию, царя Иудейского, слуг его и народ, и оставшихся в городе сем от моровой язвы, меча и голода, предам в руки Навуходоносора, царя Вавилонского, и в руки врагов их и в руки ищущих души их; и он поразит их острием меча и не пощадит их, и не пожалеет и не помилует.
JER|21|8|И народу сему скажи: так говорит Господь: вот, Я предлагаю вам путь жизни и путь смерти:
JER|21|9|кто останется в этом городе, тот умрет от меча и голода и моровой язвы; а кто выйдет и предастся Халдеям, осаждающим вас, тот будет жив, и душа его будет ему вместо добычи;
JER|21|10|ибо Я обратил лице Мое против города сего, говорит Господь, на зло, а не на добро; он будет предан в руки царя Вавилонского, и тот сожжет его огнем.
JER|21|11|И дому царя Иудейского [скажи]: слушайте слово Господне:
JER|21|12|дом Давидов! так говорит Господь: с раннего утра производите суд и спасайте обижаемого от руки обидчика, чтобы ярость Моя не вышла, как огонь, и не разгорелась по причине злых дел ваших до того, что никто не погасит.
JER|21|13|Вот, Я – против тебя, жительница долины, скала равнины, говорит Господь, – против вас, которые говорите: "кто выступит против нас и кто войдет в жилища наши?"
JER|21|14|Но Я посещу вас по плодам дел ваших, говорит Господь, и зажгу огонь в лесу вашем, и пожрет все вокруг него.
JER|22|1|Так сказал Господь: сойди в дом царя Иудейского и произнеси слово сие
JER|22|2|и скажи: выслушай слово Господне, царь Иудейский, сидящий на престоле Давидовом, ты, и слуги твои, и народ твой, входящие сими воротами.
JER|22|3|Так говорит Господь: производите суд и правду и спасайте обижаемого от руки притеснителя, не обижайте и не тесните пришельца, сироты и вдовы, и невинной крови не проливайте на месте сем.
JER|22|4|Ибо если вы будете исполнять слово сие, то будут входить воротами дома сего цари, сидящие вместо Давида на престоле его, ездящие на колеснице и на конях, сами и слуги их и народ их.
JER|22|5|А если не послушаете слов сих, то Мною клянусь, говорит Господь, что дом сей сделается пустым.
JER|22|6|Ибо так говорит Господь дому царя Иудейского: Галаад ты у Меня, вершина Ливана; но Я сделаю тебя пустынею и города необитаемыми
JER|22|7|и приготовлю против тебя истребителей, каждого со своими орудиями, и срубят лучшие кедры твои и бросят в огонь.
JER|22|8|И многие народы будут проходить через город сей и говорить друг другу: "за что Господь так поступил с этим великим городом?"
JER|22|9|И скажут в ответ: "за то, что они оставили завет Господа Бога своего и поклонялись иным богам и служили им".
JER|22|10|Не плачьте об умершем и не жалейте о нем; но горько плачьте об отходящем в плен, ибо он уже не возвратится и не увидит родной страны своей.
JER|22|11|Ибо так говорит Господь о Саллуме, сыне Иосии, царе Иудейском, который царствовал после отца своего, Иосии, и который вышел из сего места: он уже не возвратится сюда,
JER|22|12|но умрет в том месте, куда отвели его пленным, и более не увидит земли сей.
JER|22|13|Горе тому, кто строит дом свой неправдою и горницы свои беззаконием, кто заставляет ближнего своего работать даром и не отдает ему платы его,
JER|22|14|кто говорит: "построю себе дом обширный и горницы просторные", – и прорубает себе окна, и обшивает кедром, и красит красною краскою.
JER|22|15|Думаешь ли ты быть царем, потому что заключил себя в кедр? отец твой ел и пил, но производил суд и правду, и потому ему было хорошо.
JER|22|16|Он разбирал дело бедного и нищего, и потому ему хорошо было. Не это ли значит знать Меня? говорит Господь.
JER|22|17|Но твои глаза и твое сердце обращены только к твоей корысти и к пролитию невинной крови, к тому, чтобы делать притеснение и насилие.
JER|22|18|Посему так говорит Господь о Иоакиме, сыне Иосии, царе Иудейском: не будут оплакивать его: "увы, брат мой!" и: "увы, сестра!" Не будут оплакивать его: "увы, государь!" и: "увы, его величие!"
JER|22|19|Ослиным погребением будет он погребен; вытащат его и бросят далеко за ворота Иерусалима.
JER|22|20|Взойди на Ливан и кричи, и на Васане возвысь голос твой и кричи с Аварима, ибо сокрушены все друзья твои.
JER|22|21|Я говорил тебе во время благоденствия твоего; но ты сказал: "не послушаю". Таково было поведение твое с самой юности твоей, что ты не слушал гласа Моего.
JER|22|22|Всех пастырей твоих унесет ветер, и друзья твои пойдут в плен; и тогда ты будешь постыжен и посрамлен за все злодеяния твои.
JER|22|23|Живущий на Ливане, гнездящийся на кедрах! как жалок будешь ты, когда постигнут тебя муки, как боли женщины в родах!
JER|22|24|Живу Я, сказал Господь: если бы Иехония, сын Иоакима, царь Иудейский, был перстнем на правой руке Моей, то и отсюда Я сорву тебя
JER|22|25|и отдам тебя в руки ищущих души твоей и в руки тех, которых ты боишься, в руки Навуходоносора, царя Вавилонского, и в руки Халдеев,
JER|22|26|и выброшу тебя и твою мать, которая родила тебя, в чужую страну, где вы не родились, и там умрете;
JER|22|27|а в землю, куда душа их будет желать возвратиться, туда не возвратятся.
JER|22|28|"Неужели этот человек, Иехония, есть создание презренное, отверженное? или он – сосуд непотребный? за что они выброшены – он и племя его, и брошены в страну, которой не знали?"
JER|22|29|О, земля, земля, земля! слушай слово Господне.
JER|22|30|Так говорит Господь: запишите человека сего лишенным детей, человеком злополучным во дни свои, потому что никто уже из племени его не будет сидеть на престоле Давидовом и владычествовать в Иудее.
JER|23|1|Горе пастырям, которые губят и разгоняют овец паствы Моей! говорит Господь.
JER|23|2|Посему так говорит Господь, Бог Израилев, к пастырям, пасущим народ Мой: вы рассеяли овец Моих, и разогнали их, и не смотрели за ними; вот, Я накажу вас за злые деяния ваши, говорит Господь.
JER|23|3|И соберу остаток стада Моего из всех стран, куда Я изгнал их, и возвращу их во дворы их; и будут плодиться и размножаться.
JER|23|4|И поставлю над ними пастырей, которые будут пасти их, и они уже не будут бояться и пугаться, и не будут теряться, говорит Господь.
JER|23|5|Вот, наступают дни, говорит Господь, и восставлю Давиду Отрасль праведную, и воцарится Царь, и будет поступать мудро, и будет производить суд и правду на земле.
JER|23|6|Во дни Его Иуда спасется и Израиль будет жить безопасно; и вот имя Его, которым будут называть Его: "Господь оправдание наше!"
JER|23|7|Посему, вот наступают дни, говорит Господь, когда уже не будут говорить: "жив Господь, Который вывел сынов Израилевых из земли Египетской",
JER|23|8|но: "жив Господь, Который вывел и Который привел племя дома Израилева из земли северной и из всех земель, куда Я изгнал их", и будут жить на земле своей.
JER|23|9|О пророках. Сердце мое во мне раздирается, все кости мои сотрясаются; я – как пьяный, как человек, которого одолело вино, ради Господа и ради святых слов Его,
JER|23|10|потому что земля наполнена прелюбодеями, потому что плачет земля от проклятия; засохли пастбища пустыни, и стремление их – зло, и сила их – неправда,
JER|23|11|ибо и пророк и священник – лицемеры; даже в доме Моем Я нашел нечестие их, говорит Господь.
JER|23|12|За то путь их будет для них, как скользкие места в темноте: их толкнут, и они упадут там; ибо Я наведу на них бедствие, год посещения их, говорит Господь.
JER|23|13|И в пророках Самарии Я видел безумие; они пророчествовали именем Ваала, и ввели в заблуждение народ Мой, Израиля.
JER|23|14|Но в пророках Иерусалима вижу ужасное: они прелюбодействуют и ходят во лжи, поддерживают руки злодеев, чтобы никто не обращался от своего нечестия; все они предо Мною – как Содом, и жители его – как Гоморра.
JER|23|15|Посему так говорит Господь Саваоф о пророках: вот, Я накормлю их полынью и напою их водою с желчью, ибо от пророков Иерусалимских нечестие распространилось на всю землю.
JER|23|16|Так говорит Господь Саваоф: не слушайте слов пророков, пророчествующих вам: они обманывают вас, рассказывают мечты сердца своего, [а] не от уст Господних.
JER|23|17|Они постоянно говорят пренебрегающим Меня: "Господь сказал: мир будет у вас". И всякому, поступающему по упорству своего сердца, говорят: "не придет на вас беда".
JER|23|18|Ибо кто стоял в совете Господа и видел и слышал слово Его? Кто внимал слову Его и услышал?
JER|23|19|Вот, идет буря Господня с яростью, буря грозная, и падет на главу нечестивых.
JER|23|20|Гнев Господа не отвратится, доколе Он не совершит и доколе не выполнит намерений сердца Своего; в последующие дни вы ясно уразумеете это.
JER|23|21|Я не посылал пророков сих, а они сами побежали; Я не говорил им, а они пророчествовали.
JER|23|22|Если бы они стояли в Моем совете, то объявили бы народу Моему слова Мои и отводили бы их от злого пути их и от злых дел их.
JER|23|23|Разве Я – Бог [только] вблизи, говорит Господь, а не Бог и вдали?
JER|23|24|Может ли человек скрыться в тайное место, где Я не видел бы его? говорит Господь. Не наполняю ли Я небо и землю? говорит Господь.
JER|23|25|Я слышал, что говорят пророки, Моим именем пророчествующие ложь. Они говорят: "мне снилось, мне снилось".
JER|23|26|Долго ли это будет в сердце пророков, пророчествующих ложь, пророчествующих обман своего сердца?
JER|23|27|Думают ли они довести народ Мой до забвения имени Моего посредством снов своих, которые они пересказывают друг другу, как отцы их забыли имя Мое из–за Ваала?
JER|23|28|Пророк, который видел сон, пусть и рассказывает его как сон; а у которого Мое слово, тот пусть говорит слово Мое верно. Что общего у мякины с чистым зерном? говорит Господь.
JER|23|29|Слово Мое не подобно ли огню, говорит Господь, и не подобно ли молоту, разбивающему скалу?
JER|23|30|Посему, вот Я – на пророков, говорит Господь, которые крадут слова Мои друг у друга.
JER|23|31|Вот, Я – на пророков, говорит Господь, которые действуют своим языком, а говорят: "Он сказал".
JER|23|32|Вот, Я – на пророков ложных снов, говорит Господь, которые рассказывают их и вводят народ Мой в заблуждение своими обманами и обольщением, тогда как Я не посылал их и не повелевал им, и они никакой пользы не приносят народу сему, говорит Господь.
JER|23|33|Если спросит у тебя народ сей, или пророк, или священник: "какое бремя от Господа?", то скажи им: "какое бремя? Я покину вас, говорит Господь".
JER|23|34|Если пророк, или священник, или народ скажет: "бремя от Господа", Я накажу того человека и дом его.
JER|23|35|Так говорите друг другу и брат брату: "что ответил Господь?" или: "что сказал Господь?"
JER|23|36|А этого слова: "бремя от Господа", впредь не употребляйте: ибо бременем будет [такому] человеку слово его, потому что вы извращаете слова живаго Бога, Господа Саваофа Бога нашего.
JER|23|37|Так говори пророку: "что ответил тебе Господь?" или: "что сказал Господь?"
JER|23|38|А если вы еще будете говорить: "бремя от Господа", то так говорит Господь: за то, что вы говорите слово сие: "бремя от Господа", тогда как Я послал сказать вам: "не говорите: бремя от Господа", –
JER|23|39|за то, вот, Я забуду вас вовсе и оставлю вас, и город сей, который Я дал вам и отцам вашим, отвергну от лица Моего
JER|23|40|и положу на вас поношение вечное и бесславие вечное, которое не забудется.
JER|24|1|Господь показал мне: и вот, две корзины со смоквами поставлены пред храмом Господним, после того, как Навуходоносор, царь Вавилонский, вывел из Иерусалима пленными Иехонию, сына Иоакимова, царя Иудейского, и князей Иудейских с плотниками и кузнецами и привел их в Вавилон:
JER|24|2|одна корзина была со смоквами весьма хорошими, каковы бывают смоквы ранние, а другая корзина – со смоквами весьма худыми, которых по негодности [их] нельзя есть.
JER|24|3|И сказал мне Господь: что видишь ты, Иеремия? Я сказал: смоквы, смоквы хорошие – весьма хороши, а худые – весьма худы, так что их нельзя есть, потому что они очень нехороши.
JER|24|4|И было ко мне слово Господне:
JER|24|5|так говорит Господь, Бог Израилев: подобно этим смоквам хорошим Я признаю хорошими переселенцев Иудейских, которых Я послал из сего места в землю Халдейскую;
JER|24|6|и обращу на них очи Мои во благо им и возвращу их в землю сию, и устрою их, а не разорю, и насажду их, а не искореню;
JER|24|7|и дам им сердце, чтобы знать Меня, что Я Господь, и они будут Моим народом, а Я буду их Богом; ибо они обратятся ко Мне всем сердцем своим.
JER|24|8|А о худых смоквах, которых и есть нельзя по негодности [их], так говорит Господь: таким Я сделаю Седекию, царя Иудейского, и князей его и прочих Иерусалимлян, остающихся в земле сей и живущих в земле Египетской;
JER|24|9|и отдам их на озлобление и на злострадание во всех царствах земных, в поругание, в притчу, в посмеяние и проклятие во всех местах, куда Я изгоню их.
JER|24|10|И пошлю на них меч, голод и моровую язву, доколе не истреблю их с земли, которую Я дал им и отцам их.
JER|25|1|Слово, которое было к Иеремии о всем народе Иудейском, в четвертый год Иоакима, сына Иосии, царя Иудейского, – это был первый год Навуходоносора, царя Вавилонского, –
JER|25|2|и которое пророк Иеремия произнес ко всему народу Иудейскому и ко всем жителям Иерусалима и сказал:
JER|25|3|от тринадцатого года Иосии, сына Амонова, царя Иудейского, до сего дня, вот уже двадцать три года, было ко мне слово Господне, и я с раннего утра говорил вам, – и вы не слушали.
JER|25|4|Господь посылал к вам всех рабов Своих, пророков, с раннего утра посылал, – и вы не слушали и не приклоняли уха своего, чтобы слушать.
JER|25|5|Вам говорили: "обратитесь каждый от злого пути своего и от злых дел своих и живите на земле, которую Господь дал вам и отцам вашим из века в век;
JER|25|6|и не ходите во след иных богов, чтобы служить им и поклоняться им, и не прогневляйте Меня делами рук своих, и не сделаю вам зла".
JER|25|7|Но вы не слушали Меня, говорит Господь, прогневляя Меня делами рук своих, на зло себе.
JER|25|8|Посему так говорит Господь Саваоф: за то, что вы не слушали слов Моих,
JER|25|9|вот, Я пошлю и возьму все племена северные, говорит Господь, и пошлю к Навуходоносору, царю Вавилонскому, рабу Моему, и приведу их на землю сию и на жителей ее и на все окрестные народы; и совершенно истреблю их и сделаю их ужасом и посмеянием и вечным запустением.
JER|25|10|И прекращу у них голос радости и голос веселия, голос жениха и голос невесты, звук жерновов и свет светильника.
JER|25|11|И вся земля эта будет пустынею и ужасом; и народы сии будут служить царю Вавилонскому семьдесят лет.
JER|25|12|И будет: когда исполнится семьдесят лет, накажу царя Вавилонского и тот народ, говорит Господь, за их нечестие, и землю Халдейскую, и сделаю ее вечною пустынею.
JER|25|13|И совершу над тою землею все слова Мои, которые Я произнес на нее, все написанное в сей книге, что Иеремия пророчески изрек на все народы.
JER|25|14|Ибо и их поработят многочисленные народы и цари великие; и Я воздам им по их поступкам и по делам рук их.
JER|25|15|Ибо так сказал мне Господь, Бог Израилев: возьми из руки Моей чашу сию с вином ярости и напой из нее все народы, к которым Я посылаю тебя.
JER|25|16|И они выпьют, и будут шататься и обезумеют при виде меча, который Я пошлю на них.
JER|25|17|И взял я чашу из руки Господней и напоил из нее все народы, к которым послал меня Господь:
JER|25|18|Иерусалим и города Иудейские, и царей его и князей его, чтоб опустошить их и сделать ужасом, посмеянием и проклятием, как и видно ныне,
JER|25|19|фараона, царя Египетского, и слуг его, и князей его и весь народ его,
JER|25|20|и весь смешанный народ, и всех царей земли Уца, и всех царей земли Филистимской, и Аскалон, и Газу, и Екрон, и остатки Азота,
JER|25|21|Едома, и Моава, и сыновей Аммоновых,
JER|25|22|и всех царей Тира, и всех царей Сидона, и царей островов, которые за морем,
JER|25|23|Дедана, и Фему, и Буза, и всех, стригущих волосы на висках,
JER|25|24|и всех царей Аравии, и всех царей народов разноплеменных, живущих в пустыне,
JER|25|25|всех царей Зимврии, и всех царей Елама, и всех царей Мидии,
JER|25|26|и всех царей севера, близких друг к другу и дальних, и все царства земные, которые на лице земли, а царь Сесаха выпьет после них.
JER|25|27|И скажи им: так говорит Господь Саваоф, Бог Израилев: пейте и опьянейте, и изрыгните и падите, и не вставайте при виде меча, который Я пошлю на вас.
JER|25|28|Если же они будут отказываться брать чашу из руки твоей, чтобы пить, то скажи им: так говорит Господь Саваоф: вы непременно будете пить.
JER|25|29|Ибо вот на город сей, на котором наречено имя Мое, Я начинаю наводить бедствие; и вы ли останетесь ненаказанными? Нет, не останетесь ненаказанными; ибо Я призываю меч на всех живущих на земле, говорит Господь Саваоф.
JER|25|30|Посему прореки на них все слова сии и скажи им: Господь возгремит с высоты и из жилища святыни Своей подаст глас Свой; страшно возгремит на селение Свое; как топчущие в точиле, воскликнет на всех живущих на земле.
JER|25|31|Шум дойдет до концов земли, ибо у Господа состязание с народами: Он будет судиться со всякою плотью, нечестивых Он предаст мечу, говорит Господь.
JER|25|32|Так говорит Господь Саваоф: вот, бедствие пойдет от народа к народу, и большой вихрь поднимется от краев земли.
JER|25|33|И будут пораженные Господом в тот день от конца земли до конца земли, не будут оплаканы и не будут прибраны и похоронены, навозом будут на лице земли.
JER|25|34|Рыдайте, пастыри, и стенайте, и посыпайте себя прахом, вожди стада; ибо исполнились дни ваши для заклания и рассеяния вашего, и падете, как дорогой сосуд.
JER|25|35|И не будет убежища пастырям и спасения вождям стада.
JER|25|36|Слышен вопль пастырей и рыдание вождей стада, ибо опустошил Господь пажить их.
JER|25|37|Истребляются мирные селения от ярости гнева Господня.
JER|25|38|Он оставил жилище Свое, как лев; и земля их сделалась пустынею от ярости опустошителя и от пламенного гнева Его.
JER|26|1|В начале царствования Иоакима, сына Иосии, царя Иудейского, было такое слово от Господа:
JER|26|2|так говорит Господь: стань на дворе дома Господня и скажи ко всем городам Иудеи, приходящим на поклонение в дом Господень, все те слова, какие повелю тебе сказать им; не убавь ни слова.
JER|26|3|Может быть, они послушают и обратятся каждый от злого пути своего, и тогда Я отменю то бедствие, которое думаю сделать им за злые деяния их.
JER|26|4|И скажи им: так говорит Господь: если вы не послушаетесь Меня в том, чтобы поступать по закону Моему, который Я дал вам,
JER|26|5|чтобы внимать словам рабов Моих, пророков, которых Я посылаю к вам, посылаю с раннего утра, и которых вы не слушаете, –
JER|26|6|то с домом сим Я сделаю то же, что с Силомом, и город сей предам на проклятие всем народам земли.
JER|26|7|Священники и пророки и весь народ слушали Иеремию, когда он говорил сии слова в доме Господнем.
JER|26|8|И когда Иеремия сказал все, что Господь повелел ему сказать всему народу, тогда схватили его священники и пророки и весь народ, и сказали: "ты должен умереть;
JER|26|9|зачем ты пророчествуешь именем Господа и говоришь: дом сей будет как Силом, и город сей опустеет, [останется] без жителей?" И собрался весь народ против Иеремии в доме Господнем.
JER|26|10|Когда услышали об этом князья Иудейские, то пришли из дома царя к дому Господню и сели у входа в новые ворота [дома] Господня.
JER|26|11|Тогда священники и пророки так сказали князьям и всему народу: "смертный приговор этому человеку! потому что он пророчествует против города сего, как вы слышали своими ушами".
JER|26|12|И сказал Иеремия всем князьям и всему народу: "Господь послал меня пророчествовать против дома сего и против города сего все те слова, которые вы слышали;
JER|26|13|итак исправьте пути ваши и деяния ваши и послушайтесь гласа Господа Бога вашего, и Господь отменит бедствие, которое изрек на вас;
JER|26|14|а что до меня, вот – я в ваших руках; делайте со мною, что в глазах ваших покажется хорошим и справедливым;
JER|26|15|только твердо знайте, что если вы умертвите меня, то невинную кровь возложите на себя и на город сей и на жителей его; ибо истинно Господь послал меня к вам сказать все те слова в уши ваши".
JER|26|16|Тогда князья и весь народ сказали священникам и пророкам: "этот человек не подлежит смертному приговору, потому что он говорил нам именем Господа Бога нашего".
JER|26|17|И из старейшин земли встали некоторые и сказали всему народному собранию:
JER|26|18|"Михей Морасфитянин пророчествовал во дни Езекии, царя Иудейского, и сказал всему народу Иудейскому: так говорит Господь Саваоф: Сион будет вспахан, как поле, и Иерусалим сделается грудою развалин, и гора дома сего – лесистым холмом.
JER|26|19|Умертвили ли его за это Езекия, царь Иудейский, и весь Иуда? Не убоялся ли он Господа и не умолял ли Господа? и Господь отменил бедствие, которое изрек на них; а мы хотим сделать большое зло душам нашим?
JER|26|20|Пророчествовал также именем Господа некто Урия, сын Шемаии, из Кариаф–Иарима, – и пророчествовал против города сего и против земли сей точно такими же словами, как Иеремия.
JER|26|21|Когда услышал слова его царь Иоаким и все вельможи его и все князья, то искал царь умертвить его. Услышав об этом, Урия убоялся и убежал, и удалился в Египет.
JER|26|22|Но царь Иоаким и в Египет послал людей: Елнафана, сына Ахборова, и других с ним.
JER|26|23|И вывели Урию из Египта и привели его к царю Иоакиму, и он умертвил его мечом и бросил труп его, где были простонародные гробницы.
JER|26|24|Но рука Ахикама, сына Сафанова, была за Иеремию, чтобы не отдавать его в руки народа на убиение".
JER|27|1|В начале царствования Иоакима, сына Иосии, царя Иудейского, было слово сие к Иеремии от Господа:
JER|27|2|так сказал мне Господь: сделай себе узы и ярмо и возложи их себе на выю;
JER|27|3|и пошли такие же к царю Идумейскому, и к царю Моавитскому, и к царю сыновей Аммоновых, и к царю Тира, и к царю Сидона, через послов, пришедших в Иерусалим к Седекии, царю Иудейскому;
JER|27|4|и накажи им сказать государям их: так говорит Господь Саваоф, Бог Израилев: так скажите государям вашим:
JER|27|5|Я сотворил землю, человека и животных, которые на лице земли, великим могуществом Моим и простертою мышцею Моею, и отдал ее, кому Мне благоугодно было.
JER|27|6|И ныне Я отдаю все земли сии в руку Навуходоносора, царя Вавилонского, раба Моего, и даже зверей полевых отдаю ему на служение.
JER|27|7|И все народы будут служить ему и сыну его и сыну сына его, доколе не придет время и его земле и ему самому; и будут служить ему народы многие и цари великие.
JER|27|8|И если какой народ и царство не захочет служить ему, Навуходоносору, царю Вавилонскому, и не подклонит выи своей под ярмо царя Вавилонского, – этот народ Я накажу мечом, голодом и моровою язвою, говорит Господь, доколе не истреблю их рукою его.
JER|27|9|И вы не слушайте своих пророков и своих гадателей, и своих сновидцев, и своих волшебников, и своих звездочетов, которые говорят вам: "не будете служить царю Вавилонскому".
JER|27|10|Ибо они пророчествуют вам ложь, чтобы удалить вас из земли вашей, и чтобы Я изгнал вас и вы погибли.
JER|27|11|Народ же, который подклонит выю свою под ярмо царя Вавилонского и станет служить ему, Я оставлю на земле своей, говорит Господь, и он будет возделывать ее и жить на ней.
JER|27|12|И Седекии, царю Иудейскому, я говорил всеми сими словами и сказал: подклоните выю свою под ярмо царя Вавилонского и служите ему и народу его, и будете живы.
JER|27|13|Зачем умирать тебе и народу твоему от меча, голода и моровой язвы, как изрек Господь о том народе, который не будет служить царю Вавилонскому?
JER|27|14|И не слушайте слов пророков, которые говорят вам: "не будете служить царю Вавилонскому"; ибо они пророчествуют вам ложь.
JER|27|15|Я не посылал их, говорит Господь; и они ложно пророчествуют именем Моим, чтоб Я изгнал вас и чтобы вы погибли, – вы и пророки ваши, пророчествующие вам.
JER|27|16|И священникам и всему народу сему я говорил: так говорит Господь: не слушайте слов пророков ваших, которые пророчествуют вам и говорят: "вот, скоро возвращены будут из Вавилона сосуды дома Господня"; ибо они пророчествуют вам ложь.
JER|27|17|Не слушайте их, служите царю Вавилонскому и живите; зачем доводить город сей до опустошения?
JER|27|18|А если они пророки, и если у них есть слово Господне, то пусть ходатайствуют пред Господом Саваофом, чтобы сосуды, остающиеся в доме Господнем и в доме царя Иудейского и в Иерусалиме, не перешли в Вавилон.
JER|27|19|Ибо так говорит Господь Саваоф о столбах и о [медном] море и о подножиях и о прочих вещах, оставшихся в этом городе,
JER|27|20|которых Навуходоносор, царь Вавилонский, не взял, когда Иехонию, сына Иоакима, царя Иудейского, и всех знатных Иудеев и Иерусалимлян вывел из Иерусалима в Вавилон,
JER|27|21|ибо так говорит Господь Саваоф, Бог Израилев, о сосудах, оставшихся в доме Господнем и в доме царя Иудейского и в Иерусалиме:
JER|27|22|они будут отнесены в Вавилон и там останутся до того дня, когда Я посещу их, говорит Господь, и выведу их и возвращу их на место сие.
JER|28|1|В тот же год, в начале царствования Седекии, царя Иудейского, в четвертый год, в пятый месяц, Анания, сын Азура, пророк из Гаваона, говорил мне в доме Господнем пред глазами священников и всего народа и сказал:
JER|28|2|так говорит Господь Саваоф, Бог Израилев: сокрушу ярмо царя Вавилонского;
JER|28|3|через два года Я возвращу на место сие все сосуды дома Господня, которые Навуходоносор, царь Вавилонский, взял из сего места и перенес их в Вавилон;
JER|28|4|и Иехонию, сына Иоакима, царя Иудейского, и всех пленных Иудеев, пришедших в Вавилон, Я возвращу на место сие, говорит Господь; ибо сокрушу ярмо царя Вавилонского.
JER|28|5|И сказал Иеремия пророк пророку Анании пред глазами священников и пред глазами всего народа, стоявших в доме Господнем, –
JER|28|6|и сказал Иеремия пророк: да будет так, да сотворит сие Господь! да исполнит Господь слова твои, какие ты произнес о возвращении из Вавилона сосудов дома Господня и всех пленников на место сие!
JER|28|7|Только выслушай слово сие, которое я скажу вслух тебе и вслух всего народа:
JER|28|8|пророки, которые издавна были прежде меня и прежде тебя, предсказывали многим землям и великим царствам войну и бедствие и мор.
JER|28|9|Если какой пророк предсказывал мир, то тогда только он признаваем был за пророка, которого истинно послал Господь, когда сбывалось слово того пророка.
JER|28|10|Тогда пророк Анания взял ярмо с выи Иеремии пророка и сокрушил его.
JER|28|11|И сказал Анания пред глазами всего народа сии слова: так говорит Господь: так сокрушу ярмо Навуходоносора, царя Вавилонского, через два года, [сняв его] с выи всех народов. И пошел Иеремия своею дорогою.
JER|28|12|И было слово Господне к Иеремии после того, как пророк Анания сокрушил ярмо с выи пророка Иеремии:
JER|28|13|иди и скажи Анании: так говорит Господь: ты сокрушил ярмо деревянное, и сделаешь вместо него ярмо железное.
JER|28|14|Ибо так говорит Господь Саваоф, Бог Израилев: железное ярмо возложу на выю всех этих народов, чтобы они работали Навуходоносору, царю Вавилонскому, и они будут служить ему, и даже зверей полевых Я отдал ему.
JER|28|15|И сказал пророк Иеремия пророку Анании: послушай, Анания: Господь тебя не посылал, и ты обнадеживаешь народ сей ложно.
JER|28|16|Посему так говорит Господь: вот, Я сброшу тебя с лица земли; в этом же году ты умрешь, потому что ты говорил вопреки Господу.
JER|28|17|И умер пророк Анания в том же году, в седьмом месяце.
JER|29|1|И вот слова письма, которое пророк Иеремия послал из Иерусалима к остатку старейшин между переселенцами и к священникам, и к пророкам, и ко всему народу, которых Навуходоносор вывел из Иерусалима в Вавилон, –
JER|29|2|после того, как вышли из Иерусалима царь Иехония и царица и евнухи, князья Иудеи и Иерусалима, и плотники и кузнецы, –
JER|29|3|через Елеасу, сына Сафанова, и Гемарию, сына Хелкиина, которых Седекия, царь Иудейский, посылал в Вавилон к Навуходоносору, царю Вавилонскому:
JER|29|4|так говорит Господь Саваоф, Бог Израилев, всем пленникам, которых Я переселил из Иерусалима в Вавилон:
JER|29|5|стройте домы и живите [в них], и разводите сады и ешьте плоды их;
JER|29|6|берите жен и рождайте сыновей и дочерей; и сыновьям своим берите жен и дочерей своих отдавайте в замужество, чтобы они рождали сыновей и дочерей, и размножайтесь там, а не умаляйтесь;
JER|29|7|и заботьтесь о благосостоянии города, в который Я переселил вас, и молитесь за него Господу; ибо при благосостоянии его и вам будет мир.
JER|29|8|Ибо так говорит Господь Саваоф, Бог Израилев: да не обольщают вас пророки ваши, которые среди вас, и гадатели ваши; и не слушайте снов ваших, которые вам снятся;
JER|29|9|ложно пророчествуют они вам именем Моим; Я не посылал их, говорит Господь.
JER|29|10|Ибо так говорит Господь: когда исполнится вам в Вавилоне семьдесят лет, тогда Я посещу вас и исполню доброе слово Мое о вас, чтобы возвратить вас на место сие.
JER|29|11|Ибо [только] Я знаю намерения, какие имею о вас, говорит Господь, намерения во благо, а не на зло, чтобы дать вам будущность и надежду.
JER|29|12|И воззовете ко Мне, и пойдете и помолитесь Мне, и Я услышу вас;
JER|29|13|и взыщете Меня и найдете, если взыщете Меня всем сердцем вашим.
JER|29|14|И буду Я найден вами, говорит Господь, и возвращу вас из плена и соберу вас из всех народов и из всех мест, куда Я изгнал вас, говорит Господь, и возвращу вас в то место, откуда переселил вас.
JER|29|15|Вы говорите: "Господь воздвиг нам пророков и в Вавилоне".
JER|29|16|Так говорит Господь о царе, сидящем на престоле Давидовом, и о всем народе, живущем в городе сем, о братьях ваших, которые не отведены с вами в плен, –
JER|29|17|так говорит [о них] Господь Саваоф: вот, Я пошлю на них меч, голод и моровую язву, и сделаю их такими, как негодные смоквы, которых нельзя есть по негодности [их];
JER|29|18|и буду преследовать их мечом, голодом и моровою язвою, и предам их на озлобление всем царствам земли, на проклятие и ужас, на посмеяние и поругание между всеми народами, куда Я изгоню их,
JER|29|19|за то, что они не слушали слов Моих, говорит Господь, с которыми Я посылал к ним рабов Моих, пророков, посылал с раннего утра, но они не слушали, говорит Господь.
JER|29|20|А вы, все переселенцы, которых Я послал из Иерусалима в Вавилон, слушайте слово Господне:
JER|29|21|так говорит Господь Саваоф, Бог Израилев, об Ахаве, сыне Колии, и о Седекии, сыне Маасеи, которые пророчествуют вам именем Моим ложь: вот, Я предам их в руки Навуходоносора, царя Вавилонского, и он умертвит их пред вашими глазами.
JER|29|22|И принято будет от них всеми переселенцами Иудейскими, которые в Вавилоне, проклинать так: "да соделает тебе Господь то же, что Седекии и Ахаву", которых царь Вавилонский изжарил на огне
JER|29|23|за то, что они делали гнусное в Израиле: прелюбодействовали с женами ближних своих и именем Моим говорили ложь, чего Я не повелевал им; Я знаю это, и Я свидетель, говорит Господь.
JER|29|24|И Шемаии Нехеламитянину скажи:
JER|29|25|так говорит Господь Саваоф, Бог Израилев: за то, что ты посылал письма от имени своего ко всему народу, который в Иерусалиме, и к священнику Софонии, сыну Маасеи, и ко всем священникам, и писал:
JER|29|26|"Господь поставил тебя священником вместо священника Иодая, чтобы ты был между блюстителями в доме Господнем за всяким человеком, неистовствующим и пророчествующим, и чтобы ты сажал такого в темницу и в колоду:
JER|29|27|почему же ты не запретишь Иеремии Анафофскому пророчествовать у вас?
JER|29|28|Ибо он и к нам в Вавилон прислал сказать: плен будет продолжителен: стройте домы и живите в них; разводите сады и ешьте плоды их".
JER|29|29|Когда Софония священник прочитал это письмо вслух пророка Иеремии,
JER|29|30|тогда было слово Господне к Иеремии:
JER|29|31|пошли ко всем переселенцам сказать: так говорит Господь о Шемаии Нехеламитянине: за то, что Шемаия у вас пророчествует, а Я не посылал его, и обнадеживает вас ложно, –
JER|29|32|за то, так говорит Господь: вот, Я накажу Шемаию Нехеламитянина и племя его; не будет от него человека, живущего среди народа сего, и не увидит он того добра, которое Я сделаю народу Моему, говорит Господь; ибо он говорил вопреки Господу.
JER|30|1|Слово, которое было к Иеремии от Господа:
JER|30|2|так говорит Господь, Бог Израилев: напиши себе все слова, которые Я говорил тебе, в книгу.
JER|30|3|Ибо вот, наступают дни, говорит Господь, когда Я возвращу из плена народ Мой, Израиля и Иуду, говорит Господь; и приведу их опять в ту землю, которую дал отцам их, и они будут владеть ею.
JER|30|4|И вот те слова, которые сказал Господь об Израиле и Иуде.
JER|30|5|Так сказал Господь: голос смятения и ужаса слышим мы, а не мира.
JER|30|6|Спросите и рассудите: рождает ли мужчина? Почему же Я вижу у каждого мужчины руки на чреслах его, как у женщины в родах, и лица у всех бледные?
JER|30|7|О, горе! велик тот день, не было подобного ему; это – бедственное время для Иакова, но он будет спасен от него.
JER|30|8|И будет в тот день, говорит Господь Саваоф: сокрушу ярмо его, которое на вые твоей, и узы твои разорву; и не будут уже служить чужеземцам,
JER|30|9|но будут служить Господу Богу своему и Давиду, царю своему, которого Я восстановлю им.
JER|30|10|И ты, раб Мой Иаков, не бойся, говорит Господь, и не страшись, Израиль; ибо вот, Я спасу тебя из далекой страны и племя твое из земли пленения их; и возвратится Иаков и будет жить спокойно и мирно, и никто не будет устрашать его,
JER|30|11|ибо Я с тобою, говорит Господь, чтобы спасать тебя: Я совершенно истреблю все народы, среди которых рассеял тебя, а тебя не истреблю; Я буду наказывать тебя в мере, но ненаказанным не оставлю тебя.
JER|30|12|Ибо так говорит Господь: рана твоя неисцельна, язва твоя жестока;
JER|30|13|никто не заботится о деле твоем, чтобы заживить рану твою; целебного врачевства нет для тебя;
JER|30|14|все друзья твои забыли тебя, не ищут тебя; ибо Я поразил тебя ударами неприятельскими, жестоким наказанием за множество беззаконий твоих, потому что грехи твои умножились.
JER|30|15|Что вопиешь ты о ранах твоих, о жестокости болезни твоей? по множеству беззаконий твоих Я сделал тебе это, потому что грехи твои умножились.
JER|30|16|Но все пожирающие тебя будут пожраны; и все враги твои, все сами пойдут в плен, и опустошители твои будут опустошены, и всех грабителей твоих предам грабежу.
JER|30|17|Я обложу тебя пластырем и исцелю тебя от ран твоих, говорит Господь. Тебя называли отверженным, говоря: "вот Сион, о котором никто не спрашивает";
JER|30|18|так говорит Господь: вот, возвращу плен шатров Иакова и селения его помилую; и город опять будет построен на холме своем, и храм устроится по–прежнему.
JER|30|19|И вознесутся из них благодарение и голос веселящихся; и Я умножу их, и не будут умаляться, и прославлю их, и не будут унижены.
JER|30|20|И сыновья его будут, как прежде, и сонм его будет предстоять предо Мною, и накажу всех притеснителей его.
JER|30|21|И будет вождь его из него самого, и владыка его произойдет из среды его; и Я приближу его, и он приступит ко Мне; ибо кто отважится сам собою приблизиться ко Мне? говорит Господь.
JER|30|22|И вы будете Моим народом, и Я буду вам Богом.
JER|30|23|Вот, яростный вихрь идет от Господа, вихрь грозный; он падет на голову нечестивых.
JER|30|24|Пламенный гнев Господа не отвратится, доколе Он не совершит и не выполнит намерений сердца Своего. В последние дни уразумеете это.
JER|31|1|В то время, говорит Господь, Я буду Богом всем племенам Израилевым, а они будут Моим народом.
JER|31|2|Так говорит Господь: народ, уцелевший от меча, нашел милость в пустыне; иду успокоить Израиля.
JER|31|3|Издали явился мне Господь и сказал: любовью вечною Я возлюбил тебя и потому простер к тебе благоволение.
JER|31|4|Я снова устрою тебя, и ты будешь устроена, дева Израилева, снова будешь украшаться тимпанами твоими и выходить в хороводе веселящихся;
JER|31|5|снова разведешь виноградники на горах Самарии; виноградари, которые будут разводить их, сами будут и пользоваться ими.
JER|31|6|Ибо будет день, когда стражи на горе Ефремовой провозгласят: "вставайте, и взойдем на Сион к Господу Богу нашему".
JER|31|7|Ибо так говорит Господь: радостно пойте об Иакове и восклицайте пред главою народов: провозглашайте, славьте и говорите: "спаси, Господи, народ твой, остаток Израиля!"
JER|31|8|Вот, Я приведу их из страны северной и соберу их с краев земли; слепой и хромой, беременная и родильница вместе с ними, – великий сонм возвратится сюда.
JER|31|9|Они пошли со слезами, а Я поведу их с утешением; поведу их близ потоков вод дорогою ровною, на которой не споткнутся; ибо Я – отец Израилю, и Ефрем – первенец Мой.
JER|31|10|Слушайте слово Господне, народы, и возвестите островам отдаленным и скажите: "Кто рассеял Израиля, Тот и соберет его, и будет охранять его, как пастырь стадо свое";
JER|31|11|ибо искупит Господь Иакова и избавит его от руки того, кто был сильнее его.
JER|31|12|И придут они, и будут торжествовать на высотах Сиона; и стекутся к благостыне Господа, к пшенице и вину и елею, к агнцам и волам; и душа их будет как напоенный водою сад, и они не будут уже более томиться.
JER|31|13|Тогда девица будет веселиться в хороводе, и юноши и старцы вместе; и изменю печаль их на радость и утешу их, и обрадую их после скорби их.
JER|31|14|И напитаю душу священников туком, и народ Мой насытится благами Моими, говорит Господь.
JER|31|15|Так говорит Господь: голос слышен в Раме, вопль и горькое рыдание; Рахиль плачет о детях своих и не хочет утешиться о детях своих, ибо их нет.
JER|31|16|Так говорит Господь: удержи голос твой от рыдания и глаза твои от слез, ибо есть награда за труд твой, говорит Господь, и возвратятся они из земли неприятельской.
JER|31|17|И есть надежда для будущности твоей, говорит Господь, и возвратятся сыновья твои в пределы свои.
JER|31|18|Слышу Ефрема плачущего: "Ты наказал меня, и я наказан, как телец неукротимый; обрати меня, и обращусь, ибо Ты Господь Бог мой.
JER|31|19|Когда я был обращен, я каялся, и когда был вразумлен, бил себя по бедрам; я был постыжен, я был смущен, потому что нес бесславие юности моей".
JER|31|20|Не дорогой ли у Меня сын Ефрем? не любимое ли дитя? ибо, как только заговорю о нем, всегда с любовью воспоминаю о нем; внутренность Моя возмущается за него; умилосержусь над ним, говорит Господь.
JER|31|21|Поставь себе путевые знаки, поставь себе столбы, обрати сердце твое на дорогу, на путь, по которому ты шла; возвращайся, дева Израилева, возвращайся в сии города твои.
JER|31|22|Долго ли тебе скитаться, отпадшая дочь? Ибо Господь сотворит на земле нечто новое: жена спасет мужа.
JER|31|23|Так говорит Господь Саваоф, Бог Израилев: впредь, когда Я возвращу плен их, будут говорить на земле Иуды и в городах его сие слово: "да благословит тебя Господь, жилище правды, гора святая!"
JER|31|24|И поселится на ней Иуда и все города его вместе, земледельцы и ходящие со стадами.
JER|31|25|Ибо Я напою душу утомленную и насыщу всякую душу скорбящую.
JER|31|26|При этом я пробудился и посмотрел, и сон мой был приятен мне.
JER|31|27|Вот, наступают дни, говорит Господь, когда Я засею дом Израилев и дом Иудин семенем человека и семенем скота.
JER|31|28|И как Я наблюдал за ними, искореняя и сокрушая, и разрушая и погубляя, и повреждая, так буду наблюдать за ними, созидая и насаждая, говорит Господь.
JER|31|29|В те дни уже не будут говорить: "отцы ели кислый виноград, а у детей на зубах оскомина",
JER|31|30|но каждый будет умирать за свое собственное беззаконие; кто будет есть кислый виноград, у того на зубах и оскомина будет.
JER|31|31|Вот наступают дни, говорит Господь, когда Я заключу с домом Израиля и с домом Иуды новый завет,
JER|31|32|не такой завет, какой Я заключил с отцами их в тот день, когда взял их за руку, чтобы вывести их из земли Египетской; тот завет Мой они нарушили, хотя Я оставался в союзе с ними, говорит Господь.
JER|31|33|Но вот завет, который Я заключу с домом Израилевым после тех дней, говорит Господь: вложу закон Мой во внутренность их и на сердцах их напишу его, и буду им Богом, а они будут Моим народом.
JER|31|34|И уже не будут учить друг друга, брат брата, и говорить: "познайте Господа", ибо все сами будут знать Меня, от малого до большого, говорит Господь, потому что Я прощу беззакония их и грехов их уже не воспомяну более.
JER|31|35|Так говорит Господь, Который дал солнце для освещения днем, уставы луне и звездам для освещения ночью, Который возмущает море, так что волны его ревут; Господь Саваоф – имя Ему.
JER|31|36|Если сии уставы перестанут действовать предо Мною, говорит Господь, то и племя Израилево перестанет быть народом предо Мною навсегда.
JER|31|37|Так говорит Господь: если небо может быть измерено вверху, и основания земли исследованы внизу, то и Я отвергну все племя Израилево за все то, что они делали, говорит Господь.
JER|31|38|Вот, наступают дни, говорит Господь, когда город устроен будет во славу Господа от башни Анамеила до ворот угольных,
JER|31|39|и землемерная вервь пойдет далее прямо до холма Гарива и обойдет Гоаф.
JER|31|40|И вся долина трупов и пепла, и все поле до потока Кедрона, до угла конских ворот к востоку, будет святынею Господа; не разрушится и не распадется вовеки.
JER|32|1|Слово, которое было от Господа к Иеремии в десятый год Седекии, царя Иудейского; этот год был восемнадцатым годом Навуходоносора.
JER|32|2|Тогда войско царя Вавилонского осаждало Иерусалим, и Иеремия пророк был заключен во дворе стражи, который был при доме царя Иудейского.
JER|32|3|Седекия, царь Иудейский, заключил его туда, сказав: "зачем ты пророчествуешь и говоришь: так говорит Господь: вот, Я отдаю город сей в руки царя Вавилонского, и он возьмет его;
JER|32|4|и Седекия, царь Иудейский, не избегнет от рук Халдеев, но непременно предан будет в руки царя Вавилонского, и будет говорить с ним устами к устам, и глаза его увидят глаза его;
JER|32|5|и он отведет Седекию в Вавилон, где он и будет, доколе не посещу его, говорит Господь. Если вы будете воевать с Халдеями, то не будете иметь успеха?"
JER|32|6|И сказал Иеремия: таково было ко мне слово Господне:
JER|32|7|вот Анамеил, сын Саллума, дяди твоего, идет к тебе сказать: "купи себе поле мое, которое в Анафофе, потому что по праву родства тебе надлежит купить его".
JER|32|8|И Анамеил, сын дяди моего, пришел ко мне, по слову Господню, во двор стражи и сказал мне: "купи поле мое, которое в Анафофе, в земле Вениаминовой, ибо право наследства твое и право выкупа твое; купи себе". Тогда я узнал, что это было слово Господне.
JER|32|9|И купил я поле у Анамеила, сына дяди моего, которое в Анафофе, и отвесил ему семь сиклей серебра и десять сребренников;
JER|32|10|и записал в книгу и запечатал ее, и пригласил к тому свидетелей и отвесил серебро на весах.
JER|32|11|И взял я купчую запись, как запечатанную по закону и уставу, так и открытую;
JER|32|12|и отдал эту купчую запись Варуху, сыну Нирии, сына Маасеи, в глазах Анамеила, сына дяди моего, и в глазах свидетелей, подписавших эту купчую запись, в глазах всех Иудеев, сидевших на дворе стражи;
JER|32|13|и заповедал Варуху в присутствии их:
JER|32|14|так говорит Господь Саваоф, Бог Израилев: возьми сии записи, эту купчую запись, которая запечатана, и эту запись открытую, и положи их в глиняный сосуд, чтобы они оставались там многие дни.
JER|32|15|Ибо так говорит Господь Саваоф, Бог Израилев: домы и поля и виноградники будут снова покупаемы в земле сей.
JER|32|16|И, передав купчую запись Варуху, сыну Нирии, я помолился Господу:
JER|32|17|"о, Господи Боже! Ты сотворил небо и землю великою силою Твоею и простертою мышцею; для Тебя ничего нет невозможного;
JER|32|18|Ты являешь милость тысячам и за беззаконие отцов воздаешь в недро детям их после них: Боже великий, сильный, Которому имя Господь Саваоф!
JER|32|19|Великий в совете и сильный в делах, Которого очи отверсты на все пути сынов человеческих, чтобы воздавать каждому по путям его и по плодам дел его,
JER|32|20|Который совершил чудеса и знамения в земле Египетской, [и] [совершаешь] до сего дня и в Израиле и между всеми людьми, и соделал Себе имя, как в сей день,
JER|32|21|и вывел народ Твой Израиля из земли Египетской знамениями и чудесами, и рукою сильною и мышцею простертою, при великом ужасе,
JER|32|22|и дал им землю сию, которую дать им клятвенно обещал отцам их, землю, текущую молоком и медом.
JER|32|23|Они вошли и завладели ею, но не стали слушать гласа Твоего и поступать по закону Твоему, не стали делать того, что Ты заповедал им делать, и за то Ты навел на них все это бедствие.
JER|32|24|Вот, насыпи достигают до города, чтобы взять его; и город от меча и голода и моровой язвы отдается в руки Халдеев, воюющих против него; что Ты говорил, то и исполняется, и вот, Ты видишь это.
JER|32|25|А Ты, Господи Боже, сказал мне: "купи себе поле за серебро и пригласи свидетелей, тогда как город отдается в руки Халдеев".
JER|32|26|И было слово Господне к Иеремии:
JER|32|27|вот, Я Господь, Бог всякой плоти; есть ли что невозможное для Меня?
JER|32|28|Посему так говорит Господь: вот, Я отдаю город сей в руки Халдеев и в руки Навуходоносора, царя Вавилонского, и он возьмет его,
JER|32|29|и войдут Халдеи, осаждающие сей город, зажгут город огнем и сожгут его и домы, на кровлях которых возносились курения Ваалу и возливаемы были возлияния чужим богам, чтобы прогневлять Меня.
JER|32|30|Ибо сыновья Израилевы и сыновья Иудины только зло делали пред очами Моими от юности своей; сыновья Израилевы только прогневляли Меня делами рук своих, говорит Господь.
JER|32|31|И как бы для гнева Моего и ярости Моей существовал город сей с самого дня построения его до сего дня, чтобы Я отверг его от лица Моего
JER|32|32|за все зло сыновей Израиля и сыновей Иуды, какое они к прогневлению Меня делали, они, цари их, князья их, священники их и пророки их, и мужи Иуды и жители Иерусалима.
JER|32|33|Они оборотились ко Мне спиною, а не лицем; и когда Я учил их, с раннего утра учил, они не хотели принять наставления,
JER|32|34|и в доме, над которым наречено имя Мое, поставили мерзости свои, оскверняя его.
JER|32|35|Устроили капища Ваалу в долине сыновей Енномовых, чтобы проводить через огонь сыновей своих и дочерей своих в честь Молоху, чего Я не повелевал им, и Мне на ум не приходило, чтобы они делали эту мерзость, вводя в грех Иуду.
JER|32|36|И однако же ныне так говорит Господь, Бог Израилев, об этом городе, о котором вы говорите: "он предается в руки царя Вавилонского мечом и голодом и моровою язвою", –
JER|32|37|вот, Я соберу их из всех стран, в которые изгнал их во гневе Моем и в ярости Моей и в великом негодовании, и возвращу их на место сие и дам им безопасное житие.
JER|32|38|Они будут Моим народом, а Я буду им Богом.
JER|32|39|И дам им одно сердце и один путь, чтобы боялись Меня во все дни [жизни], ко благу своему и благу детей своих после них.
JER|32|40|И заключу с ними вечный завет, по которому Я не отвращусь от них, чтобы благотворить им, и страх Мой вложу в сердца их, чтобы они не отступали от Меня.
JER|32|41|И буду радоваться о них, благотворя им, и насажду их на земле сей твердо, от всего сердца Моего и от всей души Моей.
JER|32|42|Ибо так говорит Господь: как Я навел на народ сей все это великое зло, так наведу на них все благо, какое Я изрек о них.
JER|32|43|И будут покупать поля в земле сей, о которой вы говорите: "это пустыня, без людей и без скота; она отдана в руки Халдеям";
JER|32|44|будут покупать поля за серебро и вносить в записи, и запечатывать и приглашать свидетелей – в земле Вениаминовой и в окрестностях Иерусалима, и в городах Иуды и в городах нагорных, и в городах низменных и в городах южных; ибо возвращу плен их, говорит Господь.
JER|33|1|И было слово Господне к Иеремии вторично, когда он еще содержался во дворе стражи:
JER|33|2|Так говорит Господь, Который сотворил [землю], Господь, Который устроил и утвердил ее, – Господь имя Ему:
JER|33|3|воззови ко Мне – и Я отвечу тебе, покажу тебе великое и недоступное, чего ты не знаешь.
JER|33|4|Ибо так говорит Господь, Бог Израилев, о домах города сего и о домах царей Иудейских, которые разрушаются для завалов и для сражения
JER|33|5|пришедшими воевать с Халдеями, чтобы наполнить домы трупами людей, которых Я поражу во гневе Моем и в ярости Моей, и за все беззакония которых Я сокрыл лице Мое от города сего.
JER|33|6|Вот, Я приложу ему пластырь и целебные средства, и уврачую их, и открою им обилие мира и истины,
JER|33|7|и возвращу плен Иуды и плен Израиля и устрою их, как вначале,
JER|33|8|и очищу их от всего нечестия их, которым они грешили предо Мною, и прощу все беззакония их, которыми они грешили предо Мною и отпали от Меня.
JER|33|9|И будет для меня [Иерусалим] радостным именем, похвалою и честью пред всеми народами земли, которые услышат о всех благах, какие Я сделаю ему, и изумятся и затрепещут от всех благодеяний и всего благоденствия, которое Я доставлю ему.
JER|33|10|Так говорит Господь: на этом месте, о котором вы говорите: "оно пусто, без людей и без скота", – в городах Иудейских и на улицах Иерусалима, которые пусты, без людей, без жителей, без скота,
JER|33|11|опять будет слышен голос радости и голос веселья, голос жениха и голос невесты, голос говорящих: "славьте Господа Саваофа, ибо благ Господь, ибо вовек милость Его", и голос приносящих жертву благодарения в доме Господнем; ибо Я возвращу плененных сей земли в прежнее состояние, говорит Господь.
JER|33|12|Так говорит Господь Саваоф: на этом месте, которое пусто, без людей, без скота, и во всех городах его опять будут жилища пастухов, которые будут покоить стада.
JER|33|13|В городах нагорных, в городах низменных и в городах южных, и в земле Вениаминовой, и в окрестностях Иерусалима, и в городах Иуды опять будут проходить стада под рукою считающего, говорит Господь.
JER|33|14|Вот, наступят дни, говорит Господь, когда Я выполню то доброе слово, которое изрек о доме Израилевом и о доме Иудином.
JER|33|15|В те дни и в то время возращу Давиду Отрасль праведную, и будет производить суд и правду на земле.
JER|33|16|В те дни Иуда будет спасен и Иерусалим будет жить безопасно, и нарекут имя Ему: "Господь оправдание наше!"
JER|33|17|Ибо так говорит Господь: не прекратится у Давида муж, сидящий на престоле дома Израилева,
JER|33|18|и у священников–левитов не будет недостатка в муже пред лицем Моим, во все дни возносящем всесожжение и сожигающем приношения и совершающем жертвы.
JER|33|19|И было слово Господне к Иеремии:
JER|33|20|так говорит Господь: если можете разрушить завет Мой о дне и завет Мой о ночи, чтобы день и ночь не приходили в свое время,
JER|33|21|то может быть разрушен и завет Мой с рабом Моим Давидом, так что не будет у него сына, царствующего на престоле его, и также с левитами–священниками, служителями Моими.
JER|33|22|Как неисчислимо небесное воинство и неизмерим песок морской, так размножу племя Давида, раба Моего, и левитов, служащих Мне.
JER|33|23|И было слово Господне к Иеремии:
JER|33|24|не видишь ли, что народ этот говорит: "те два племени, которые избрал Господь, Он отверг?" и чрез это они презирают народ Мой, как бы он уже не был народом в глазах их.
JER|33|25|Так говорит Господь: если завета Моего о дне и ночи и уставов неба и земли Я не утвердил,
JER|33|26|то и племя Иакова и Давида, раба Моего, отвергну, чтобы не брать более владык из его племени для племени Авраама, Исаака и Иакова; ибо возвращу плен их и помилую их.
JER|34|1|Слово, которое было к Иеремии от Господа, когда Навуходоносор, царь Вавилонский, и все войско его и все царства земли, подвластные руке его, и все народы воевали против Иерусалима и против всех городов его:
JER|34|2|так говорит Господь, Бог Израилев: иди и скажи Седекии, царю Иудейскому, и скажи ему: так говорит Господь: вот, Я отдаю город сей в руки царя Вавилонского, и он сожжет его огнем;
JER|34|3|и ты не избежишь от руки его, но непременно будешь взят и предан в руки его, и глаза твои увидят глаза царя Вавилонского, и уста его будут говорить твоим устам, и пойдешь в Вавилон.
JER|34|4|Впрочем слушай слово Господне, Седекия, царь Иудейский! так говорит Господь о тебе: ты не умрешь от меча;
JER|34|5|ты умрешь в мире, и как для отцов твоих, прежних царей, которые были прежде тебя, сожигали [при погребении благовония], так сожгут и для тебя и оплачут тебя: "увы, государь!", ибо Я изрек это слово, говорит Господь.
JER|34|6|Иеремия пророк все слова сии пересказал Седекии, царю Иудейскому, в Иерусалиме.
JER|34|7|Между тем войско царя Вавилонского воевало против Иерусалима и против всех городов Иудейских, которые еще оставались, против Лахиса и Азеки; ибо из городов Иудейских сии только оставались, как города укрепленные.
JER|34|8|Слово, которое было к Иеремии от Господа после того, как царь Седекия заключил завет со всем народом, бывшим в Иерусалиме, чтобы объявить свободу,
JER|34|9|чтобы каждый отпустил на волю раба своего и рабу свою, Еврея и Евреянку, чтобы никто из них не держал в рабстве Иудея, брата своего.
JER|34|10|И послушались все князья и весь народ, которые вступили в завет, чтобы отпустить каждому раба своего и каждому рабу свою на волю, чтобы не держать их впредь в рабах, – и послушались и отпустили;
JER|34|11|но после того, раздумавши, стали брать назад рабов и рабынь, которых отпустили на волю, и принудили их быть рабами и рабынями.
JER|34|12|И было слово Господне к Иеремии от Господа:
JER|34|13|так говорит Господь, Бог Израилев: Я заключил завет с отцами вашими, когда вывел их из земли Египетской, из дома рабства, и сказал:
JER|34|14|"в конце седьмого года отпускайте каждый брата своего, Еврея, который продал себя тебе; пусть он работает тебе шесть лет, а потом отпусти его от себя на волю"; но отцы ваши не послушали Меня и не приклонили уха своего.
JER|34|15|Вы ныне обратились и поступили справедливо пред очами Моими, объявив каждый свободу ближнему своему, и заключили предо Мною завет в доме, над которым наречено имя Мое;
JER|34|16|но потом раздумали и обесславили имя Мое, и возвратили к себе каждый раба своего и каждый рабу свою, которых отпустили на волю, куда душе их угодно, и принуждаете их быть у вас рабами и рабынями.
JER|34|17|Посему так говорит Господь: вы не послушались Меня в том, чтобы каждый объявил свободу брату своему и ближнему своему; за то вот Я, говорит Господь, объявляю вам свободу подвергнуться мечу, моровой язве и голоду, и отдам вас на озлобление во все царства земли;
JER|34|18|и отдам преступивших завет Мой и не устоявших в словах завета, который они заключили пред лицем Моим, рассекши тельца надвое и пройдя между рассеченными частями его,
JER|34|19|князей Иудейских и князей Иерусалимских, евнухов и священников и весь народ земли, проходивший между рассеченными частями тельца, –
JER|34|20|отдам их в руки врагов их и в руки ищущих души их, и трупы их будут пищею птицам небесным и зверям земным.
JER|34|21|И Седекию, царя Иудейского, и князей его отдам в руки врагов их и в руки ищущих души их и в руки войска царя Вавилонского, которое отступило от вас.
JER|34|22|Вот, Я дам повеление, говорит Господь, и возвращу их к этому городу, и они нападут на него, и возьмут его, и сожгут его огнем, и города Иудеи сделаю пустынею необитаемою.
JER|35|1|Слово, которое было к Иеремии от Господа во дни Иоакима, сына Иосии, царя Иудейского:
JER|35|2|иди в дом Рехавитов и поговори с ними, и приведи их в дом Господень, в одну из комнат, и дай им пить вина.
JER|35|3|Я взял Иазанию, сына Иеремии, сына Авацинии, и братьев его, и всех сыновей его и весь дом Рехавитов,
JER|35|4|и привел их в дом Господень, в комнату сынов Анана, сына Годолии, человека Божия, которая подле комнаты князей, над комнатою Маасеи, сына Селлумова, стража у входа;
JER|35|5|и поставил перед сынами дома Рехавитов полные чаши вина и стаканы и сказал им: пейте вино.
JER|35|6|Но они сказали: мы вина не пьем; потому что Ионадав, сын Рехава, отец наш, дал нам заповедь, сказав: "не пейте вина ни вы, ни дети ваши, вовеки;
JER|35|7|и домов не стройте, и семян не сейте, и виноградников не разводите, и не имейте их, но живите в шатрах во все дни [жизни] вашей, чтобы вам долгое время прожить на той земле, где вы странниками".
JER|35|8|И мы послушались голоса Ионадава, сына Рехавова, отца нашего, во всем, что он завещал нам, чтобы не пить вина во все дни наши, – мы и жены наши, и сыновья наши и дочери наши, –
JER|35|9|и чтобы не строить домов для жительства нашего; и у нас нет ни виноградников, ни полей, ни посева;
JER|35|10|а живем в шатрах и во всем слушаемся и делаем все, что заповедал нам Ионадав, отец наш.
JER|35|11|Когда же Навуходоносор, царь Вавилонский, пришел в землю сию, мы сказали: "пойдем, уйдем в Иерусалим от войска Халдеев и от войска Арамеев", и вот, мы живем в Иерусалиме.
JER|35|12|И было слово Господне к Иеремии:
JER|35|13|так говорит Господь Саваоф, Бог Израилев: иди и скажи мужам Иуды и жителям Иерусалима: неужели вы не возьмете из этого наставление для себя, чтобы слушаться слов Моих? говорит Господь.
JER|35|14|Слова Ионадава, сына Рехавова, который завещал сыновьям своим не пить вина, выполняются, и они не пьют до сего дня, потому что слушаются завещания отца своего; а Я непрестанно говорил вам, говорил с раннего утра, и вы не послушались Меня.
JER|35|15|Я посылал к вам всех рабов Моих, пророков, посылал с раннего утра, и говорил: "обратитесь каждый от злого пути своего и исправьте поведение ваше, и не ходите во след иных богов, чтобы служить им; и будете жить на этой земле, которую Я дал вам и отцам вашим"; но вы не приклонили уха своего и не послушались Меня.
JER|35|16|Так как сыновья Ионадава, сына Рехавова, выполняют заповедь отца своего, которую он заповедал им, а народ сей не слушает Меня,
JER|35|17|посему так говорит Господь Бог Саваоф, Бог Израилев: вот, Я наведу на Иудею и на всех жителей Иерусалима все то зло, которое Я изрек на них, потому что Я говорил им, а они не слушались, звал их, а они не отвечали.
JER|35|18|А дому Рехавитов сказал Иеремия: так говорит Господь Саваоф, Бог Израилев: за то, что вы послушались завещания Ионадава, отца вашего, и храните все заповеди его и во всем поступаете, как он завещал вам, –
JER|35|19|за то, так говорит Господь Саваоф, Бог Израилев: не отнимется у Ионадава, сына Рехавова, муж, предстоящий пред лицем Моим во все дни.
JER|36|1|В четвертый год Иоакима, сына Иосии, царя Иудейского, было такое слово к Иеремии от Господа:
JER|36|2|возьми себе книжный свиток и напиши в нем все слова, которые Я говорил тебе об Израиле и об Иуде и о всех народах с того дня, как Я начал говорить тебе, от дней Иосии до сего дня;
JER|36|3|может быть, дом Иудин услышит о всех бедствиях, какие Я помышляю сделать им, чтобы они обратились каждый от злого пути своего, чтобы Я простил неправду их и грех их.
JER|36|4|И призвал Иеремия Варуха, сына Нирии, и написал Варух в книжный свиток из уст Иеремии все слова Господа, которые Он говорил ему.
JER|36|5|И приказал Иеремия Варуху и сказал: я заключен и не могу идти в дом Господень;
JER|36|6|итак иди ты и прочитай написанные тобою в свитке с уст моих слова Господни вслух народа в доме Господнем в день поста, также и вслух всех Иудеев, пришедших из городов своих, прочитай их;
JER|36|7|может быть, они вознесут смиренное моление пред лице Господа и обратятся каждый от злого пути своего; ибо велик гнев и негодование, которое объявил Господь на народ сей.
JER|36|8|Варух, сын Нирии, сделал все, что приказал ему пророк Иеремия, чтобы слова Господни, написанные в свитке, прочитать в доме Господнем.
JER|36|9|В пятый год Иоакима, сына Иосии, царя Иудейского, в девятом месяце объявили пост пред лицем Господа всему народу в Иерусалиме и всему народу, пришедшему в Иерусалим из городов Иудейских.
JER|36|10|И прочитал Варух написанные в свитке слова Иеремии в доме Господнем, в комнате Гемарии, сына Сафанова, писца, на верхнем дворе, у входа в новые ворота дома Господня, вслух всего народа.
JER|36|11|Михей, сын Гемарии, сына Сафанова, слышал все слова Господни, [написанные] в свитке,
JER|36|12|и сошел в дом царя, в комнату царского писца, и вот, там сидели все князья: Елисам, царский писец, и Делаия, сын Семаия, и Елнафан, сын Ахбора, и Гемария, сын Сафана, и Седекия, сын Анании, и все князья;
JER|36|13|и пересказал им Михей все слова, которые он слышал, когда Варух читал свиток вслух народа.
JER|36|14|Тогда все князья послали к Варуху Иегудия, сына Нафании, сына Селемии, сына Хусии, сказать ему: свиток, который ты читал вслух народа, возьми в руку твою и приди. И взял Варух, сын Нирии, свиток в руку свою и пришел к ним.
JER|36|15|Они сказали ему: сядь, и прочитай нам вслух. И прочитал Варух вслух им.
JER|36|16|Когда они выслушали все слова, то с ужасом посмотрели друг на друга и сказали Варуху: мы непременно перескажем все сии слова царю.
JER|36|17|И спросили Варуха: скажи же нам, как ты написал все слова сии из уст его?
JER|36|18|И сказал им Варух: он произносил мне устами своими все сии слова, а я чернилами писал их в этот свиток.
JER|36|19|Тогда сказали князья Варуху: пойди, скройся, ты и Иеремия, чтобы никто не знал, где вы.
JER|36|20|И пошли они к царю во дворец, а свиток оставили в комнате Елисама, царского писца, и пересказали вслух царя все слова сии.
JER|36|21|Царь послал Иегудия принести свиток, и он взял его из комнаты Елисама, царского писца; и читал его Иегудий вслух царя и вслух всех князей, стоявших подле царя.
JER|36|22|Царь в то время, в девятом месяце, сидел в зимнем доме, и перед ним горела жаровня.
JER|36|23|Когда Иегудий прочитывал три или четыре столбца, [царь] отрезывал их писцовым ножичком и бросал на огонь в жаровне, доколе не уничтожен был весь свиток на огне, который был в жаровне.
JER|36|24|И не убоялись, и не разодрали одежд своих ни царь, ни все слуги его, слышавшие все слова сии.
JER|36|25|Хотя Елнафан и Делаия и Гемария упрашивали царя не сожигать свитка, но он не послушал их.
JER|36|26|И приказал царь Иерамеилу, сыну царя, и Сераии, сыну Азриилову, и Селемии, сыну Авдиилову, взять Варуха писца и Иеремию пророка; но Господь сокрыл их.
JER|36|27|И было слово Господне к Иеремии, после того как царь сожег свиток и слова, которые Варух написал из уст Иеремии, и сказано ему:
JER|36|28|возьми себе опять другой свиток и напиши в нем все прежние слова, какие были в первом свитке, который сожег Иоаким, царь Иудейский;
JER|36|29|а царю Иудейскому Иоакиму скажи: так говорит Господь: ты сожег свиток сей, сказав: "зачем ты написал в нем: непременно придет царь Вавилонский и разорит землю сию, и истребит на ней людей и скот?"
JER|36|30|за это, так говорит Господь об Иоакиме, царе Иудейском: не будет от него сидящего на престоле Давидовом, и труп его будет брошен на зной дневной и на холод ночной;
JER|36|31|и посещу его и племя его и слуг его за неправду их, и наведу на них и на жителей Иерусалима и на мужей Иуды все зло, которое Я изрек на них, а они не слушали.
JER|36|32|И взял Иеремия другой свиток и отдал его Варуху писцу, сыну Нирии, и он написал в нем из уст Иеремии все слова того свитка, который сожег Иоаким, царь Иудейский, на огне; и еще прибавлено к ним много подобных тем слов.
JER|37|1|Вместо Иехонии, сына Иоакима, царствовал Седекия, сын Иосии, которого Навуходоносор, царь Вавилонский, поставил царем в земле Иудейской.
JER|37|2|Ни он, ни слуги его, ни народ страны не слушали слов Господа, которые говорил Он чрез Иеремию пророка.
JER|37|3|Царь Седекия послал Иегухала, сына Селемии, и Софонию, сына Маасеи, священника, к Иеремии пророку сказать: помолись о нас Господу Богу нашему.
JER|37|4|Иеремия тогда еще свободно входил и выходил среди народа, потому что не заключили его в дом темничный.
JER|37|5|Между тем войско фараоново выступило из Египта, и Халдеи, осаждавшие Иерусалим, услышав весть о том, отступили от Иерусалима.
JER|37|6|И было слово Господне к Иеремии пророку:
JER|37|7|так говорит Господь, Бог Израилев: так скажите царю Иудейскому, пославшему вас ко Мне вопросить Меня: вот, войско фараоново, которое шло к вам на помощь, возвратится в землю свою, в Египет;
JER|37|8|а Халдеи снова придут и будут воевать против города сего, и возьмут его и сожгут его огнем.
JER|37|9|Так говорит Господь: не обманывайте себя, говоря: "непременно отойдут от нас Халдеи", ибо они не отойдут;
JER|37|10|если бы вы даже разбили все войско Халдеев, воюющих против вас, и остались бы у них только раненые, то и те встали бы, каждый из палатки своей, и сожгли бы город сей огнем.
JER|37|11|В то время, как войско Халдейское отступило от Иерусалима, по причине войска фараонова,
JER|37|12|Иеремия пошел из Иерусалима, чтобы уйти в землю Вениаминову, скрываясь оттуда среди народа.
JER|37|13|Но когда он был в воротах Вениаминовых, бывший там начальник стражи, по имени Иреия, сын Селемии, сына Анании, задержал Иеремию пророка, сказав: ты хочешь перебежать к Халдеям?
JER|37|14|Иеремия сказал: это ложь; я не хочу перебежать к Халдеям. Но он не послушал его, и взял Иреия Иеремию и привел его к князьям.
JER|37|15|Князья озлобились на Иеремию и били его, и заключили его в темницу, в дом Ионафана писца, потому что сделали его темницею.
JER|37|16|Когда Иеремия вошел в темницу и подвал, и пробыл там Иеремия много дней, –
JER|37|17|царь Седекия послал и взял его. И спрашивал его царь в доме своем тайно и сказал: нет ли слова от Господа? Иеремия сказал: есть; и сказал: ты будешь предан в руки царя Вавилонского.
JER|37|18|И сказал Иеремия царю Седекии: чем я согрешил перед тобою и перед слугами твоими, и перед народом сим, что вы посадили меня в темницу?
JER|37|19|и где ваши пророки, которые пророчествовали вам, говоря: "царь Вавилонский не пойдет против вас и против земли сей"?
JER|37|20|И ныне послушай, государь мой царь, да падет прошение мое пред лице твое; не возвращай меня в дом Ионафана писца, чтобы мне не умереть там.
JER|37|21|И дал повеление царь Седекия, чтобы заключили Иеремию во дворе стражи и давали ему по куску хлеба на день из улицы хлебопеков, доколе не истощился весь хлеб в городе; и так оставался Иеремия во дворе стражи.
JER|38|1|И услышали Сафатия, сын Матфана, и Годолия, сын Пасхора, и Юхал, сын Селемии, и Пасхор, сын Малхии, слова, которые Иеремия произнес ко всему народу, говоря:
JER|38|2|так говорит Господь: кто останется в этом городе, умрет от меча, голода и моровой язвы; а кто выйдет к Халдеям, будет жив, и душа его будет ему вместо добычи, и он останется жив.
JER|38|3|Так говорит Господь: непременно предан будет город сей в руки войска царя Вавилонского, и он возьмет его.
JER|38|4|Тогда князья сказали царю: да будет этот человек предан смерти, потому что он ослабляет руки воинов, которые остаются в этом городе, и руки всего народа, говоря к ним такие слова; ибо этот человек не благоденствия желает народу сему, а бедствия.
JER|38|5|И сказал царь Седекия: вот, он в ваших руках, потому что царь ничего не может делать вопреки вам.
JER|38|6|Тогда взяли Иеремию и бросили его в яму Малхии, сына царя, которая была во дворе стражи, и опустили Иеремию на веревках; в яме той не было воды, а только грязь, и погрузился Иеремия в грязь.
JER|38|7|И услышал Авдемелех Ефиоплянин, один из евнухов, находившихся в царском доме, что Иеремию посадили в яму; а царь сидел тогда у ворот Вениаминовых.
JER|38|8|И вышел Авдемелех из дома царского и сказал царю:
JER|38|9|государь мой царь! худо сделали эти люди, так поступив с Иеремиею пророком, которого бросили в яму; он умрет там от голода, потому что нет более хлеба в городе.
JER|38|10|Царь дал приказание Авдемелеху Ефиоплянину, сказав: возьми с собою отсюда тридцать человек и вытащи Иеремию пророка из ямы, доколе он не умер.
JER|38|11|Авдемелех взял людей с собою и вошел в дом царский под кладовую, и взял оттуда старых негодных тряпок и старых негодных лоскутьев и опустил их на веревках в яму к Иеремии.
JER|38|12|И сказал Авдемелех Ефиоплянин Иеремии: подложи эти старые брошенные тряпки и лоскутья под мышки рук твоих, под веревки. И сделал так Иеремия.
JER|38|13|И потащили Иеремию на веревках и вытащили его из ямы; и оставался Иеремия во дворе стражи.
JER|38|14|Тогда царь Седекия послал и призвал Иеремию пророка к себе, при третьем входе в дом Господень, и сказал царь Иеремии: я у тебя спрошу нечто; не скрой от меня ничего.
JER|38|15|И сказал Иеремия Седекии: если я открою тебе, не предашь ли ты меня смерти? и если дам тебе совет, ты не послушаешь меня.
JER|38|16|И клялся царь Седекия Иеремии тайно, говоря: жив Господь, Который сотворил нам душу сию, не предам тебя смерти и не отдам в руки этих людей, которые ищут души твоей.
JER|38|17|Тогда Иеремия сказал Седекии: так говорит Господь Бог Саваоф, Бог Израилев: если ты выйдешь к князьям царя Вавилонского, то жива будет душа твоя, и этот город не будет сожжен огнем, и ты будешь жив, и дом твой;
JER|38|18|а если не выйдешь к князьям царя Вавилонского, то этот город будет предан в руки Халдеев, и они сожгут его огнем, и ты не избежишь от рук их.
JER|38|19|И сказал царь Седекия Иеремии: я боюсь Иудеев, которые перешли к Халдеям, чтобы [Халдеи] не предали меня в руки их, и чтобы те не надругались надо мною.
JER|38|20|И сказал Иеремия: не предадут; послушай гласа Господа в том, что я говорю тебе, и хорошо тебе будет, и жива будет душа твоя.
JER|38|21|А если ты не захочешь выйти, то вот слово, которое открыл мне Господь:
JER|38|22|вот, все жены, которые остались в доме царя Иудейского, отведены будут к князьям царя Вавилонского, и скажут они: "тебя обольстили и превозмогли друзья твои; ноги твои погрузились в грязь, и они удалились от тебя".
JER|38|23|И всех жен твоих и детей твоих отведут к Халдеям, и ты не избежишь от рук их; но будешь взят рукою царя Вавилонского, и сделаешь то, что город сей будет сожжен огнем.
JER|38|24|И сказал Седекия Иеремии: никто не должен знать этих слов, и тогда ты не умрешь;
JER|38|25|и если услышат князья, что я разговаривал с тобою, и придут к тебе, и скажут тебе: "скажи нам, что говорил ты царю, не скрой от нас, и мы не предадим тебя смерти, – и также что говорил тебе царь",
JER|38|26|то скажи им: "я повергнул пред лице царя прошение мое, чтобы не возвращать меня в дом Ионафана, чтобы не умереть там".
JER|38|27|И пришли все князья к Иеремии и спрашивали его, и он сказал им согласно со всеми словами, какие царь велел [сказать], и они молча оставили его, потому что не узнали сказанного царю.
JER|38|28|И оставался Иеремия во дворе стражи до того дня, в который был взят Иерусалим. И Иерусалим был взят.
JER|39|1|В девятый год Седекии, царя Иудейского, в десятый месяц, пришел Навуходоносор, царь Вавилонский, со всем войском своим к Иерусалиму, и обложили его.
JER|39|2|А в одиннадцатый год Седекии, в четвертый месяц, в девятый день месяца город был взят.
JER|39|3|И вошли [в него] все князья царя Вавилонского, и расположились в средних воротах, Нергал–Шарецер, Самгар–Нево, Сарсехим, начальник евнухов, Нергал–Шарецер, начальник магов, и все остальные князья царя Вавилонского.
JER|39|4|Когда Седекия, царь Иудейский, и все военные люди увидели их, – побежали, и ночью вышли из города через царский сад в ворота между двумя стенами и пошли по дороге равнины.
JER|39|5|Но войско Халдейское погналось за ними; и настигли Седекию на равнинах Иерихонских; и взяли его и отвели к Навуходоносору, царю Вавилонскому, в Ривлу, в землю Емаф, где он произнес суд над ним.
JER|39|6|И заколол царь Вавилонский сыновей Седекии в Ривле перед его глазами, и всех вельмож Иудейских заколол царь Вавилонский;
JER|39|7|а Седекии выколол глаза и заковал его в оковы, чтобы отвести его в Вавилон.
JER|39|8|Дом царя и домы народа сожгли Халдеи огнем, и стены Иерусалима разрушили.
JER|39|9|А остаток народа, остававшийся в городе, и перебежчиков, которые перешли к нему, и прочий оставшийся народ Навузардан, начальник телохранителей, переселил в Вавилон.
JER|39|10|Бедных же из народа, которые ничего не имели, Навузардан, начальник телохранителей, оставил в Иудейской земле и дал им тогда же виноградники и поля.
JER|39|11|А о Иеремии Навуходоносор, царь Вавилонский, дал такое повеление Навузардану, начальнику телохранителей:
JER|39|12|возьми его и имей его во внимании, и не делай ему ничего худого, но поступай с ним так, как он скажет тебе.
JER|39|13|И послал Навузардан, начальник телохранителей, и Навузазван, начальник евнухов, и Нергал–Шарецер, начальник магов, и все князья царя Вавилонского
JER|39|14|послали и взяли Иеремию со двора стражи, и поручили его Годолии, сыну Ахикама, сына Сафанова, отвести его домой. И он остался жить среди народа.
JER|39|15|К Иеремии, когда он еще содержался во дворе темничном, было слово Господне:
JER|39|16|иди, скажи Авдемелеху Ефиоплянину: так говорит Господь Саваоф, Бог Израилев: вот, Я исполню слова Мои о городе сем во зло, а не в добро ему, и они сбудутся в тот день перед глазами твоими;
JER|39|17|но тебя Я избавлю в тот день, говорит Господь, и не будешь предан в руки людей, которых ты боишься.
JER|39|18|Я избавлю тебя, и ты не падешь от меча, и душа твоя останется у тебя вместо добычи, потому что ты на Меня возложил упование, сказал Господь.
JER|40|1|Слово, которое было к Иеремии от Господа, после того как Навузардан, начальник телохранителей, отпустил его из Рамы, где он взял его скованного цепями среди прочих пленных Иерусалимлян и Иудеев, переселяемых в Вавилон.
JER|40|2|Начальник телохранителей взял Иеремию и сказал ему: Господь Бог твой изрек это бедствие на место сие,
JER|40|3|и навел его Господь и сделал то, что сказал; потому что вы согрешили пред Господом и не слушались гласа Его, за то и постигло вас это.
JER|40|4|Итак вот, я освобождаю тебя сегодня от цепей, которые на руках твоих: если тебе угодно идти со мною в Вавилон, иди, и я буду иметь попечение о тебе; а если не угодно тебе идти со мною в Вавилон, оставайся. Вот, вся земля перед тобою; куда тебе угодно, и куда нравится идти, туда и иди.
JER|40|5|Когда он еще не отошел, сказал [Навузардан]: пойди к Годолии, сыну Ахикама, сына Сафанова, которого царь Вавилонский поставил начальником над городами Иудейскими, и оставайся с ним среди народа; или иди, куда нравится тебе идти. И дал ему начальник телохранителей продовольствие и подарок и отпустил его.
JER|40|6|И пришел Иеремия к Годолии, сыну Ахикама, в Массифу, и жил с ним среди народа, остававшегося в стране.
JER|40|7|Когда все военачальники, бывшие в поле, они и люди их, услышали, что царь Вавилонский поставил Годолию, сына Ахикама, начальником над страною и поручил ему мужчин и женщин, и детей, и тех из бедных страны, которые не были переселены в Вавилон;
JER|40|8|тогда пришли к Годолии в Массифу и Исмаил, сын Нафании, и Иоанан и Ионафан, сыновья Карея, и Сераия, сын Фанасмефа, и сыновья Офи из Нетофафы, и Иезония, сын Махафы, они и дружина их.
JER|40|9|Годолия, сын Ахикама, сына Сафанова, клялся им и людям их, говоря: не бойтесь служить Халдеям, оставайтесь на земле и служите царю Вавилонскому, и будет вам хорошо;
JER|40|10|а я останусь в Массифе, чтобы предстательствовать пред лицем Халдеев, которые будут приходить к нам; вы же собирайте вино и летние плоды, и масло и убирайте в сосуды ваши, и живите в городах ваших, которые заняли.
JER|40|11|Также все Иудеи, которые находились в земле Моавитской и между сыновьями Аммона и в Идумее, и во всех странах, услышали, что царь Вавилонский оставил часть Иудеев и поставил над ними Годолию, сына Ахикама, сына Сафана:
JER|40|12|и возвратились все сии Иудеи из всех мест, куда были изгнаны, и пришли в землю Иудейскую к Годолии в Массифу, и собрали вина и летних плодов очень много.
JER|40|13|Между тем Иоанан, сын Карея, и все военные начальники, бывшие в поле, пришли к Годолии в Массифу
JER|40|14|и сказали ему: знаешь ли ты, что Ваалис, царь сыновей Аммоновых, прислал Исмаила, сына Нафании, чтобы убить тебя? Но Годолия, сын Ахикама, не поверил им.
JER|40|15|Тогда Иоанан, сын Карея, сказал Годолии тайно в Массифе: позволь мне, я пойду и убью Исмаила, сына Нафании, и никто не узнает; зачем допускать, чтобы он убил тебя, и чтобы все Иудеи, собравшиеся к тебе, рассеялись, и чтобы погиб остаток Иуды?
JER|40|16|Но Годолия, сын Ахикама, сказал Иоанану, сыну Карея: не делай этого, ибо ты неправду говоришь об Исмаиле.
JER|41|1|И было в седьмой месяц, Исмаил, сын Нафании, сына Елисама из племени царского, и вельможи царя и десять человек с ним пришли к Годолии, сыну Ахикама, в Массифу, и там они ели вместе хлеб в Массифе.
JER|41|2|И встал Исмаил, сын Нафании, и десять человек, которые были с ним, и поразили Годолию, сына Ахикама, сына Сафанова, мечом и умертвили того, которого царь Вавилонский поставил начальником над страною.
JER|41|3|Также убил Исмаил и всех Иудеев, которые были с ним, с Годолиею, в Массифе, и находившихся там Халдеев, людей военных.
JER|41|4|На другой день по убиении Годолии, когда никто не знал об этом,
JER|41|5|пришли из Сихема, Силома и Самарии восемьдесят человек с обритыми бородами и в разодранных одеждах, и изранив себя, с дарами и ливаном в руках для принесения их в дом Господень.
JER|41|6|Исмаил, сын Нафании, вышел из Массифы навстречу им, идя и плача, и, встретившись с ними, сказал им: идите к Годолии, сыну Ахикама.
JER|41|7|И как только они вошли в средину города, Исмаил, сын Нафании, убил их и [бросил] в ров, он и бывшие с ним люди.
JER|41|8|Но нашлись между ними десять человек, которые сказали Исмаилу: не умерщвляй нас, ибо у нас есть в поле скрытые кладовые с пшеницею и ячменем, и маслом и медом. И он удержался и не умертвил их с другими братьями их.
JER|41|9|Ров же, куда бросил Исмаил все трупы людей, которых он убил из–за Годолии, был тот самый, который сделал царь Аса, боясь Ваасы, царя Израильского; его наполнил Исмаил, сын Нафании, убитыми.
JER|41|10|И захватил Исмаил весь остаток народа, бывшего в Массифе, дочерей царя и весь остававшийся в Массифе народ, который Навузардан, начальник телохранителей, поручил Годолии, сыну Ахикама, и захватил их Исмаил, сын Нафании, и отправился к сыновьям Аммоновым.
JER|41|11|Но когда Иоанан, сын Карея, и все бывшие с ним военные начальники услышали о всех злодеяниях, какие совершил Исмаил, сын Нафании,
JER|41|12|взяли всех людей и пошли сразиться с Исмаилом, сыном Нафании, и настигли его у больших вод, в Гаваоне.
JER|41|13|И когда весь народ, бывший у Исмаила, увидел Иоанана, сына Карея, и всех бывших с ним военных начальников, обрадовался;
JER|41|14|и отворотился весь народ, который Исмаил увел в плен из Массифы, и обратился и пошел к Иоанану, сыну Карея;
JER|41|15|а Исмаил, сын Нафании, убежал от Иоанана с восемью человеками и ушел к сыновьям Аммоновым.
JER|41|16|Тогда Иоанан, сын Карея, и все бывшие с ним военные начальники взяли из Массифы весь оставшийся народ, который он освободил от Исмаила, сына Нафании, после того как тот убил Годолию, сына Ахикама, мужчин, военных людей, и жен, и детей, и евнухов, которых он вывел из Гаваона;
JER|41|17|и пошли, и остановились в селении Химам, близ Вифлеема, чтобы уйти в Египет
JER|41|18|от Халдеев, ибо они боялись их, потому что Исмаил, сын Нафании, убил Годолию, сына Ахикама, которого царь Вавилонский поставил начальником над страною.
JER|42|1|И приступили все военные начальники, и Иоанан, сын Карея, и Иезания, сын Гошаии, и весь народ от малого до большого,
JER|42|2|и сказали Иеремии пророку: да падет пред лице твое прошение наше, помолись о нас Господу Богу твоему обо всем этом остатке, ибо из многого осталось нас мало, как глаза твои видят нас,
JER|42|3|чтобы Господь, Бог твой, указал нам путь, по которому нам идти, и то, что нам делать.
JER|42|4|И сказал им Иеремия пророк: слышу, помолюсь Господу Богу вашему по словам вашим, и все, что ответит вам Господь, объявлю вам, не скрою от вас ни слова.
JER|42|5|Они сказали Иеремии: Господь да будет между нами свидетелем верным и истинным в том, что мы точно выполним все то, с чем пришлет тебя к нам Господь Бог Твой:
JER|42|6|хорошо ли, худо ли то будет, но гласа Господа Бога нашего, к Которому посылаем тебя, послушаемся, чтобы нам было хорошо, когда будем послушны гласу Господа Бога нашего.
JER|42|7|По прошествии десяти дней было слово Господне к Иеремии.
JER|42|8|Он позвал к себе Иоанана, сына Карея, и всех бывших с ним военных начальников и весь народ, от малого и до большого,
JER|42|9|и сказал им: так говорит Господь, Бог Израилев, к Которому вы посылали меня, чтобы повергнуть пред Ним моление ваше:
JER|42|10|если останетесь на земле сей, то Я устрою вас и не разорю, насажду вас и не искореню, ибо Я сожалею о том бедствии, какое сделал вам.
JER|42|11|Не бойтесь царя Вавилонского, которого вы боитесь; не бойтесь его, говорит Господь, ибо Я с вами, чтобы спасать вас и избавлять вас от руки его.
JER|42|12|И явлю к вам милость, и он умилостивится к вам и возвратит вас в землю вашу.
JER|42|13|Если же вы скажете: "не хотим жить в этой земле", и не послушаетесь гласа Господа Бога вашего, говоря:
JER|42|14|"нет, мы пойдем в землю Египетскую, где войны не увидим и трубного голоса не услышим, и голодать не будем, и там будем жить";
JER|42|15|то выслушайте ныне слово Господне, вы, остаток Иуды: так говорит Господь Саваоф, Бог Израилев: если вы решительно обратите лица ваши, чтобы идти в Египет, и пойдете, чтобы жить там,
JER|42|16|то меч, которого вы боитесь, настигнет вас там, в земле Египетской, и голод, которого вы страшитесь, будет всегда следовать за вами там, в Египте, и там умрете.
JER|42|17|И все, которые обратят лице свое, чтобы идти в Египет и там жить, умрут от меча, голода и моровой язвы, и ни один из них не останется и не избежит того бедствия, которое Я наведу на них.
JER|42|18|Ибо так говорит Господь Саваоф, Бог Израилев: как излился гнев Мой и ярость Моя на жителей Иерусалима, так изольется ярость Моя на вас, когда войдете в Египет, и вы будете проклятием и ужасом, и поруганием и поношением, и не увидите более места сего.
JER|42|19|К вам, остаток Иуды, изрек Господь: "не ходите в Египет"; твердо знайте, что я ныне предостерегал вас,
JER|42|20|ибо вы погрешили против себя самих: вы послали меня к Господу Богу нашему сказав: "помолись о нас Господу Богу нашему и все, что скажет Господь Бог наш, объяви нам, и мы сделаем".
JER|42|21|Я объявил вам ныне; но вы не послушали гласа Господа Бога нашего и всего того, с чем Он послал меня к вам.
JER|42|22|Итак знайте, что вы умрете от меча, голода и моровой язвы в том месте, куда хотите идти, чтобы жить там.
JER|43|1|Когда Иеремия передал всему народу все слова Господа Бога их, все те слова, с которыми Господь, Бог их, послал его к ним,
JER|43|2|тогда сказал Азария, сын Осаии, и Иоанан, сын Карея, и все дерзкие люди сказали Иеремии: неправду ты говоришь, не посылал тебя Господь Бог наш сказать: "не ходите в Египет, чтобы жить там";
JER|43|3|а Варух, сын Нирии, возбуждает тебя против нас, чтобы предать нас в руки Халдеев, чтобы они умертвили нас или отвели нас пленными в Вавилон.
JER|43|4|И не послушал Иоанан, сын Карея, и все военные начальники и весь народ гласа Господа, чтобы остаться в земле Иудейской.
JER|43|5|И взял Иоанан, сын Карея, и все военные начальники весь остаток Иудеев, которые возвратились из всех народов, куда они были изгнаны, чтобы жить в земле Иудейской,
JER|43|6|мужей и жен, и детей, и дочерей царя, и всех тех, которых Навузардан, начальник телохранителей, оставил с Годолиею, сыном Ахикама, сына Сафанова, и Иеремию пророка, и Варуха, сына Нирии;
JER|43|7|и пошли в землю Египетскую, ибо не послушали гласа Господня, и дошли до Тафниса.
JER|43|8|И было слово Господне к Иеремии в Тафнисе:
JER|43|9|возьми в руки свои большие камни и скрой их в смятой глине при входе в дом фараона в Тафнисе, пред глазами Иудеев,
JER|43|10|и скажи им: так говорит Господь Саваоф, Бог Израилев: вот, Я пошлю и возьму Навуходоносора, царя Вавилонского, раба Моего, и поставлю престол его на этих камнях, скрытых Мною, и раскинет он над ним великолепный шатер свой
JER|43|11|и придет, и поразит землю Египетскую: кто [обречен] на смерть, тот [предан будет] смерти; и кто в плен, [пойдет] в плен; и кто под меч, под меч.
JER|43|12|И зажгу огонь в капищах богов Египтян; и он сожжет оные, а их пленит, и оденется в землю Египетскую, как пастух надевает на себя одежду свою, и выйдет оттуда спокойно,
JER|43|13|и сокрушит статуи в Бефсамисе, что в земле Египетской, и капища богов Египетских сожжет огнем.
JER|44|1|Слово, которое было к Иеремии о всех Иудеях, живущих в земле Египетской, поселившихся в Магдоле и Тафнисе, и в Нофе, и в земле Пафрос:
JER|44|2|так говорит Господь Саваоф, Бог Израилев: вы видели все бедствие, какое Я навел на Иерусалим и на все города Иудейские; вот, они теперь пусты, и никто не живет в них,
JER|44|3|за нечестие их, которое они делали, прогневляя Меня, ходя кадить и служить иным богам, которых не знали ни они, ни вы, ни отцы ваши.
JER|44|4|Я посылал к вам всех рабов Моих, пророков, посылал с раннего утра, чтобы сказать: "не делайте этого мерзкого дела, которое Я ненавижу".
JER|44|5|Но они не слушали и не приклонили уха своего, чтобы обратиться от своего нечестия, не кадить иным богам.
JER|44|6|И излилась ярость Моя и гнев Мой и разгорелась в городах Иудеи и на улицах Иерусалима; и они сделались развалинами и пустынею, как видите ныне.
JER|44|7|И ныне так говорит Господь Бог Саваоф, Бог Израилев: зачем вы делаете это великое зло душам вашим, истребляя у себя мужей и жен, взрослых детей и младенцев из среды Иудеи, чтобы не оставить у себя остатка,
JER|44|8|прогневляя Меня изделием рук своих, каждением иным богам в земле Египетской, куда вы пришли жить, чтобы погубить себя и сделаться проклятием и поношением у всех народов земли?
JER|44|9|Разве вы забыли нечестие отцов ваших и нечестие царей Иудейских, ваше собственное нечестие и нечестие жен ваших, какое они делали в земле Иудейской и на улицах Иерусалима?
JER|44|10|Не смирились они и до сего дня, и не боятся и не поступают по закону Моему и по уставам Моим, которые Я дал вам и отцам вашим.
JER|44|11|Посему так говорит Господь Саваоф, Бог Израилев: вот, Я обращу против вас лице Мое на погибель и на истребление всей Иудеи
JER|44|12|и возьму оставшихся Иудеев, которые обратили лице свое, чтобы идти в землю Египетскую и жить там, и все они будут истреблены, падут в земле Египетской; мечом и голодом будут истреблены; от малого и до большого умрут от меча и голода, и будут проклятием и ужасом, поруганием и поношением.
JER|44|13|Посещу живущих в земле Египетской, как Я посетил Иерусалим, мечом, голодом и моровою язвою,
JER|44|14|и никто не избежит и не уцелеет из остатка Иудеев, пришедших в землю Египетскую, чтобы пожить там и потом возвратиться в землю Иудейскую, куда они всею душею желают возвратиться, чтобы жить там; никто не возвратится, кроме тех, которые убегут оттуда.
JER|44|15|И отвечали Иеремии все мужья, знавшие, что жены их кадят иным богам, и все жены, стоявшие [там] в большом множестве, и весь народ, живший в земле Египетской, в Пафросе, и сказали:
JER|44|16|слова, которое ты говорил нам именем Господа, мы не слушаем от тебя;
JER|44|17|но непременно будем делать все то, что вышло из уст наших, чтобы кадить богине неба и возливать ей возлияния, как мы делали, мы и отцы наши, цари наши и князья наши, в городах Иудеи и на улицах Иерусалима, потому что тогда мы были сыты и счастливы и беды не видели.
JER|44|18|А с того времени, как перестали мы кадить богине неба и возливать ей возлияния, терпим во всем недостаток и гибнем от меча и голода.
JER|44|19|И когда мы кадили богине неба и возливали ей возлияния, то разве без ведома мужей наших делали мы ей пирожки с изображением ее и возливали ей возлияния?
JER|44|20|Тогда сказал Иеремия всему народу, мужьям и женам, и всему народу, который так отвечал ему:
JER|44|21|не это ли каждение, которое совершали вы в городах Иудейских и на улицах Иерусалима, вы и отцы ваши, цари ваши и князья ваши, и народ страны, воспомянул Господь? И не оно ли взошло Ему на сердце?
JER|44|22|Господь не мог более терпеть злых дел ваших и мерзостей, какие вы делали; поэтому и сделалась земля ваша пустынею и ужасом, и проклятием, без жителей, как видите ныне.
JER|44|23|Так как вы, совершая то курение, грешили пред Господом и не слушали гласа Господа, и не поступали по закону Его и по установлениям Его, и по повелениям Его, то и постигло вас это бедствие, как видите ныне.
JER|44|24|И сказал Иеремия всему народу и всем женам: слушайте слово Господне, все Иудеи, которые в земле Египетской:
JER|44|25|так говорит Господь Саваоф, Бог Израилев: вы и жены ваши, что устами своими говорили, то и руками своими делали; вы говорите: "станем выполнять обеты наши, какие мы обещали, чтобы кадить богине неба и возливать ей возлияние", – твердо держитесь обетов ваших и в точности исполняйте обеты ваши.
JER|44|26|За то выслушайте слово Господне, все Иудеи, живущие в земле Египетской: вот, Я поклялся великим именем Моим, говорит Господь, что не будет уже на всей земле Египетской произносимо имя Мое устами какого–либо Иудея, говорящего: "жив Господь Бог!"
JER|44|27|Вот, Я буду наблюдать над вами к погибели, а не к добру; и все Иудеи, которые в земле Египетской, будут погибать от меча и голода, доколе совсем не истребятся.
JER|44|28|Только малое число избежавших от меча возвратится из земли Египетской в землю Иудейскую, и узнают все оставшиеся Иудеи, которые пришли в землю Египетскую, чтобы пожить там, чье слово сбудется: Мое или их.
JER|44|29|И вот вам знамение, говорит Господь, что Я посещу вас на сем месте, чтобы вы знали, что сбудутся слова Мои о вас на погибель вам.
JER|44|30|Так говорит Господь: вот, Я отдам фараона Вафрия, царя Египетского, в руки врагов его и в руки ищущих души его, как отдал Седекию, царя Иудейского, в руки Навуходоносора, царя Вавилонского, врага его и искавшего души его.
JER|45|1|Слово, которое пророк Иеремия сказал Варуху, сыну Нирии, когда он написал слова сии из уст Иеремии в книгу, в четвертый год Иоакима, сына Иосии, царя Иудейского:
JER|45|2|так говорит Господь, Бог Израилев, к тебе, Варух:
JER|45|3|ты говоришь: "горе мне! ибо Господь приложил скорбь к болезни моей; я изнемог от вздохов моих, и не нахожу покоя".
JER|45|4|Так скажи ему: так говорит Господь: вот, что Я построил, разрушу, и что насадил, искореню, – всю эту землю.
JER|45|5|А ты просишь себе великого: не проси; ибо вот, Я наведу бедствие на всякую плоть, говорит Господь, а тебе вместо добычи оставлю душу твою во всех местах, куда ни пойдешь.
JER|46|1|Слово Господне, которое было к Иеремии пророку о народах [языческих]:
JER|46|2|о Египте, о войске фараона Нехао, царя Египетского, которое было при реке Евфрате в Кархемисе, и которое поразил Навуходоносор, царь Вавилонский, в четвертый год Иоакима, сына Иосии, царя Иудейского.
JER|46|3|Готовьте щиты и копья, и вступайте в сражение:
JER|46|4|седлайте коней и садитесь, всадники, и становитесь в шлемах; точите копья, облекайтесь в брони.
JER|46|5|Почему же, вижу Я, они оробели и обратились назад? и сильные их поражены, и бегут не оглядываясь; отвсюду ужас, говорит Господь.
JER|46|6|Не убежит быстроногий, и не спасется сильный; на севере, у реки Евфрата, они споткнутся и падут.
JER|46|7|Кто это поднимается, как река, и, как потоки, волнуются воды его?
JER|46|8|Египет поднимается, как река, и, как потоки, взволновались воды его, и говорит: "поднимусь и покрою землю, погублю город и жителей его".
JER|46|9|Садитесь на коней, и мчитесь, колесницы, и выступайте, сильные Ефиопляне и Ливияне, вооруженные щитом, и Лидяне, держащие луки и натягивающие их;
JER|46|10|ибо день сей у Господа Бога Саваофа есть день отмщения, чтобы отмстить врагам Его; и меч будет пожирать, и насытится и упьется кровью их; ибо это Господу Богу Саваофу будет жертвоприношение в земле северной, при реке Евфрате.
JER|46|11|Пойди в Галаад и возьми бальзама, дева, дочь Египта; напрасно ты будешь умножать врачевства, нет для тебя исцеления.
JER|46|12|Услышали народы о посрамлении твоем, и вопль твой наполнил землю; ибо сильный столкнулся с сильным, и оба вместе пали.
JER|46|13|Слово, которое сказал Господь пророку Иеремии о нашествии Навуходоносора, царя Вавилонского, чтобы поразить землю Египетскую:
JER|46|14|возвестите в Египте и дайте знать в Магдоле, и дайте знать в Нофе и Тафнисе; скажите: "становись и готовься, ибо меч пожирает окрестности твои".
JER|46|15|Отчего сильный твой опрокинут? – Не устоял, потому что Господь погнал его.
JER|46|16|Он умножил падающих, даже падали один на другого и говорили: "вставай и возвратимся к народу нашему в родную нашу землю от губительного меча".
JER|46|17|А там кричат: "фараон, царь Египта, смутился; он пропустил условленное время".
JER|46|18|Живу Я, говорит Царь, Которого имя Господь Саваоф: как Фавор среди гор и как Кармил при море, [так верно] придет он.
JER|46|19|Готовь себе нужное для переселения, дочь – жительница Египта, ибо Ноф будет опустошен, разорен, останется без жителя.
JER|46|20|Египет – прекрасная телица; но погибель от севера идет, идет.
JER|46|21|И наемники его среди него, как откормленные тельцы, – и сами обратились назад, побежали все, не устояли, потому что пришел на них день погибели их, время посещения их.
JER|46|22|Голос его несется, как змеиный; они идут с войском, придут на него с топорами, как дровосеки;
JER|46|23|вырубят лес его, говорит Господь, ибо они несметны; их более, нежели саранчи, и нет числа им.
JER|46|24|Посрамлена дочь Египта, предана в руки народа северного.
JER|46|25|Господь Саваоф, Бог Израилев, говорит: вот, Я посещу Аммона, который в Но, и фараона и Египет, и богов его и царей его, фараона и надеющихся на него;
JER|46|26|и предам их в руки ищущих души их и в руки Навуходоносора, царя Вавилонского, и в руки рабов его; но после того будет он населен, как в прежние дни, говорит Господь.
JER|46|27|Ты же не бойся, раб мой Иаков, и не страшись, Израиль: ибо вот, Я спасу тебя из далекой страны и семя твое из земли плена их; и возвратится Иаков, и будет жить спокойно и мирно, и никто не будет устрашать его.
JER|46|28|Не бойся, раб Мой Иаков, говорит Господь: ибо Я с тобою; Я истреблю все народы, к которым Я изгнал тебя, а тебя не истреблю, а только накажу тебя в мере; ненаказанным же не оставлю тебя.
JER|47|1|Слово Господа, которое было к пророку Иеремии о Филистимлянах, прежде нежели фараон поразил Газу.
JER|47|2|Так говорит Господь: вот, поднимаются воды с севера и сделаются наводняющим потоком, и потопят землю и все, что наполняет ее, город и живущих в нем; тогда возопиют люди, и зарыдают все обитатели страны.
JER|47|3|От шумного топота копыт сильных коней его, от стука колесниц его, от звука колес его, отцы не оглянутся на детей своих, потому что руки у них опустятся
JER|47|4|от того дня, который придет истребить всех Филистимлян, отнять у Тира и Сидона всех остальных помощников, ибо Господь разорит Филистимлян, остаток острова Кафтора.
JER|47|5|Оплешивела Газа, гибнет Аскалон, остаток долины их.
JER|47|6|Доколе будешь посекать, о, меч Господень! доколе ты не успокоишься? возвратись в ножны твои, перестань и успокойся.
JER|47|7|Но как тебе успокоиться, когда Господь дал повеление против Аскалона и против берега морского? туда Он направил его.
JER|48|1|О Моаве так говорит Господь Саваоф, Бог Израилев: горе Нево! он опустошен; Кариафаим посрамлен и взят; Мизгав посрамлен и сокрушен.
JER|48|2|Нет более славы Моава; в Есевоне замышляют против него зло: "пойдем, истребим его из числа народов". И ты, Мадмена, погибнешь; меч следует за тобою.
JER|48|3|Слышен вопль от Оронаима, опустошение и разрушение великое.
JER|48|4|Сокрушен Моав; вопль подняли дети его.
JER|48|5|На восхождении в Лухит плач за плачем поднимается; и на спуске с Оронаима неприятель слышит вопль о разорении.
JER|48|6|Бегите, спасайте жизнь свою, и будьте подобны обнаженному дереву в пустыне.
JER|48|7|Так как ты надеялся на дела твои и на сокровища твои, то и ты будешь взят, и Хамос пойдет в плен вместе со своими священниками и своими князьями.
JER|48|8|И придет опустошитель на всякий город, и город не уцелеет; и погибнет долина, и опустеет равнина, как сказал Господь.
JER|48|9|Дайте крылья Моаву, чтобы он мог улететь; города его будут пустынею, потому что некому будет жить в них.
JER|48|10|Проклят, кто дело Господне делает небрежно, и проклят, кто удерживает меч Его от крови!
JER|48|11|Моав от юности своей был в покое, сидел на дрожжах своих и не был переливаем из сосуда с сосуд, и в плен не ходил; от того оставался в нем вкус его, и запах его не изменялся.
JER|48|12|Посему вот, приходят дни, говорит Господь, когда Я пришлю к нему переливателей, которые перельют его и опорожнят сосуды его, и разобьют кувшины его.
JER|48|13|И постыжен будет Моав ради Хамоса, как дом Израилев постыжен был ради Вефиля, надежды своей.
JER|48|14|Как вы говорите: "мы люди храбрые и крепкие для войны"?
JER|48|15|Опустошен Моав, и города его горят, и отборные юноши его пошли на заклание, говорит Царь, – Господь Саваоф имя Его.
JER|48|16|Близка погибель Моава, и сильно спешит бедствие его.
JER|48|17|Пожалейте о нем все соседи его и все, знающие имя его, скажите: "как сокрушен жезл силы, посох славы!"
JER|48|18|Сойди с высоты величия и сиди в жажде, дочь – обитательница Дивона, ибо опустошитель Моава придет к тебе и разорит укрепления твои.
JER|48|19|Стань у дороги и смотри, обитательница Ароера, спрашивай бегущего и спасающегося: "что сделалось?"
JER|48|20|Посрамлен Моав, ибо сокрушен; рыдайте и вопите, объявите в Арноне, что опустошен Моав.
JER|48|21|И суд пришел на равнины, на Халон и на Иаацу, и на Мофаф,
JER|48|22|и на Дивон и на Нево, и на Бет–Дивлафаим,
JER|48|23|и на Кариафаим и на Бет–Гамул, и на Бет–Маон,
JER|48|24|и на Кериоф, и на Восор, и на все города земли Моавитской, дальние и ближние.
JER|48|25|Отсечен рог Моава, и мышца его сокрушена, говорит Господь.
JER|48|26|Напойте его пьяным, ибо он вознесся против Господа; и пусть Моав валяется в блевотине своей, и сам будет посмеянием.
JER|48|27|Не был ли в посмеянии у тебя Израиль? разве он между ворами был пойман, что ты, бывало, лишь только заговоришь о нем, качаешь головою?
JER|48|28|Оставьте города и живите на скалах, жители Моава, и будьте как голуби, которые делают гнезда во входе в пещеру.
JER|48|29|Слыхали мы о гордости Моава, гордости чрезмерной, о его высокомерии и его надменности, и кичливости его и превозношении сердца его.
JER|48|30|Знаю Я дерзость его, говорит Господь, но это ненадежно; пустые слова его: не так сделают.
JER|48|31|Поэтому буду рыдать о Моаве и вопить о всем Моаве; будут воздыхать о мужах Кирхареса.
JER|48|32|Буду плакать о тебе, виноградник Севамский, плачем Иазера; отрасли твои простирались за море, достигали до озера Иазера; опустошитель напал на летние плоды твои и на зрелый виноград.
JER|48|33|Радость и веселье отнято от Кармила и от земли Моава. Я положу конец вину в точилах; не будут более топтать в них с песнями; крик брани будет, а не крик радости.
JER|48|34|От вопля Есевона до Елеалы и до Иаацы они поднимут голос свой от Сигора до Оронаима, до третьей Эглы, ибо и воды Нимрима иссякнут.
JER|48|35|Истреблю у Моава, говорит Господь, приносящих жертвы на высотах и кадящих богам его.
JER|48|36|От того сердце мое стонет о Моаве, как свирель; о жителях Кирхареса стонет сердце мое, как свирель, ибо богатства, ими приобретенные, погибли:
JER|48|37|у каждого голова гола и у каждого борода умалена; у всех на руках царапины и на чреслах вретище.
JER|48|38|На всех кровлях Моава и на улицах его общий плач, ибо Я сокрушил Моава, как непотребный сосуд, говорит Господь.
JER|48|39|"Как сокрушен он!" будут говорить рыдая; "как Моав покрылся стыдом, обратив тыл!". И будет Моав посмеянием и ужасом для всех окружающих его,
JER|48|40|ибо так говорит Господь: вот, как орел, налетит он и распрострет крылья свои над Моавом.
JER|48|41|Города будут взяты, и крепости завоеваны, и сердце храбрых Моавитян будет в тот день, как сердце женщины, мучимой родами.
JER|48|42|И истреблен будет Моав из числа народов, потому что он восстал против Господа.
JER|48|43|Ужас и яма и петля – для тебя, житель Моава, сказал Господь.
JER|48|44|Кто убежит от ужаса, упадет в яму; а кто выйдет из ямы, попадет в петлю, ибо Я наведу на него, на Моава, годину посещения их, говорит Господь.
JER|48|45|Под тенью Есевона остановились бегущие, обессилев; но огонь вышел из Есевона и пламя из среды Сигона, и пожрет бок Моава и темя сыновей мятежных.
JER|48|46|Горе тебе, Моав! погиб народ Хамоса, ибо сыновья твои взяты в плен, и дочери твои – в пленение.
JER|48|47|Но в последние дни возвращу плен Моава, говорит Господь. Доселе суд на Моава.
JER|49|1|О сыновьях Аммоновых так говорит Господь: разве нет сыновей у Израиля? разве нет у него наследника? Почему же Малхом завладел Гадом, и народ его живет в городах его?
JER|49|2|Посему вот, наступают дни, говорит Господь, когда в Равве сыновей Аммоновых слышен будет крик брани, и сделается она грудою развалин, и города ее будут сожжены огнем, и овладеет Израиль теми, которые владели им, говорит Господь.
JER|49|3|Рыдай, Есевон, ибо опустошен Гай; кричите, дочери Раввы, опояшьтесь вретищем, плачьте и скитайтесь по огородам, ибо Малхом пойдет в плен вместе со священниками и князьями своими.
JER|49|4|Что хвалишься долинами? Потечет долина твоя кровью, вероломная дочь, надеющаяся на сокровища свои, [говорящая]: "кто придет ко мне?"
JER|49|5|Вот, Я наведу на тебя ужас со всех окрестностей твоих, говорит Господь Бог Саваоф; разбежитесь, кто куда, и никто не соберет разбежавшихся.
JER|49|6|Но после того Я возвращу плен сыновей Аммоновых, говорит Господь.
JER|49|7|О Едоме так говорит Господь Саваоф: разве нет более мудрости в Фемане? [разве] не стало совета у разумных? разве оскудела мудрость их?
JER|49|8|Бегите, обратив тыл, скрывайтесь в пещерах, жители Дедана, ибо погибель Исава Я наведу на него, – время посещения Моего.
JER|49|9|Если бы обиратели винограда пришли к тебе, то верно оставили бы несколько недобранных ягод. И если бы воры [пришли] ночью, то они похитили бы, сколько им нужно.
JER|49|10|А Я донага оберу Исава, открою потаенные места его, и скрыться он не может. Истреблено будет племя его, и братья его и соседи его; и не будет его.
JER|49|11|Оставь сирот твоих, Я поддержу жизнь их, и вдовы твои пусть надеются на Меня.
JER|49|12|Ибо так говорит Господь: вот и те, которым не суждено было пить чашу, непременно будут пить ее, и ты ли останешься ненаказанным? Нет, не останешься ненаказанным, но непременно будешь пить [чашу].
JER|49|13|Ибо Мною клянусь, говорит Господь, что ужасом, посмеянием, пустынею и проклятием будет Восор, и все города его сделаются вечными пустынями.
JER|49|14|Я слышал слух от Господа, и посол послан к народам сказать: соберитесь и идите против него, и поднимайтесь на войну.
JER|49|15|Ибо вот, Я сделаю тебя малым между народами, презренным между людьми.
JER|49|16|Грозное положение твое и надменность сердца твоего обольстили тебя, живущего в расселинах скал и занимающего вершины холмов. Но, хотя бы ты, как орел, высоко свил гнездо твое, и оттуда низрину тебя, говорит Господь.
JER|49|17|И будет Едом ужасом; всякий, проходящий мимо, изумится и посвищет, [смотря] на все язвы его.
JER|49|18|Как ниспровергнуты Содом и Гоморра и соседние города их, говорит Господь, так [и] там ни один человек не будет жить, и сын человеческий не остановится в нем.
JER|49|19|Вот, восходит он, как лев, от возвышения Иордана на укрепленные жилища; но Я заставлю их поспешно уйти из [Идумеи], и кто избран, того поставлю над нею. Ибо кто подобен Мне? и кто потребует ответа от Меня? и какой пастырь противостанет Мне?
JER|49|20|Итак выслушайте определение Господа, какое Он поставил об Едоме, и намерения Его, какие Он имеет о жителях Фемана: истинно, самые малые из стад повлекут их и опустошат жилища их.
JER|49|21|От шума падения их потрясется земля, и отголосок крика их слышен будет у Чермного моря.
JER|49|22|Вот, как орел поднимется он, и полетит, и распустит крылья свои над Восором; и сердце храбрых Идумеян будет в тот день, как сердце женщины в родах.
JER|49|23|О Дамаске. – Посрамлены Емаф и Арпад, ибо, услышав скорбную весть, они уныли; тревога на море, успокоиться не могут.
JER|49|24|Оробел Дамаск и обратился в бегство; страх овладел им; боль и муки схватили его, как женщину в родах.
JER|49|25|Как не уцелел город славы, город радости моей?
JER|49|26|Итак падут юноши его на улицах его, и все воины погибнут в тот день, говорит Господь Саваоф.
JER|49|27|И зажгу огонь в стенах Дамаска, и истребит чертоги Венадада.
JER|49|28|О Кидаре и о царствах Асорских, которые поразил Навуходоносор, царь Вавилонский, так говорит Господь: вставайте, выступайте против Кидара, и опустошайте сыновей востока!
JER|49|29|Шатры их и овец их возьмут себе, и покровы их и всю утварь их, и верблюдов их возьмут, и будут кричать им: "ужас отовсюду!"
JER|49|30|Бегите, уходите скорее, сокройтесь в пропасти, жители Асора, говорит Господь, ибо Навуходоносор, царь Вавилонский, сделал решение о вас и составил против вас замысел.
JER|49|31|Вставайте, выступайте против народа мирного, живущего беспечно, говорит Господь; ни дверей, ни запоров нет у него, живут поодиночке.
JER|49|32|Верблюды их [отданы] будут в добычу, и множество стад их – на расхищение; и рассею их по всем ветрам, этих стригущих волосы на висках, и со всех сторон их наведу на них гибель, говорит Господь.
JER|49|33|И будет Асор жилищем шакалов, вечною пустынею; человек не будет жить там, и сын человеческий не будет останавливаться в нем.
JER|49|34|Слово Господа, которое было к Иеремии пророку против Елама, в начале царствования Седекии, царя Иудейского:
JER|49|35|так говорит Господь Саваоф: вот, Я сокрушу лук Елама, главную силу их.
JER|49|36|И наведу на Елам четыре ветра от четырех краев неба и развею их по всем этим ветрам, и не будет народа, к которому не пришли бы изгнанные Еламиты.
JER|49|37|И поражу Еламитян страхом пред врагами их и пред ищущими души их; и наведу на них бедствие, гнев Мой, говорит Господь, и пошлю вслед их меч, доколе не истреблю их.
JER|49|38|И поставлю престол Мой в Еламе, и истреблю там царя и князей, говорит Господь.
JER|49|39|Но в последние дни возвращу плен Елама, говорит Господь.
JER|50|1|Слово, которое изрек Господь о Вавилоне и о земле Халдеев чрез Иеремию пророка:
JER|50|2|возвестите и разгласите между народами, и поднимите знамя, объявите, не скрывайте, говорите: "Вавилон взят, Вил посрамлен, Меродах сокрушен, истуканы его посрамлены, идолы его сокрушены".
JER|50|3|Ибо от севера поднялся против него народ, который сделает землю его пустынею, и никто не будет жить там, от человека до скота, все двинутся и уйдут.
JER|50|4|В те дни и в то время, говорит Господь, придут сыновья Израилевы, они и сыновья Иудины вместе, будут ходить и плакать, и взыщут Господа Бога своего.
JER|50|5|Будут спрашивать о пути к Сиону, и, обращая к нему лица, [будут] [говорить]: "идите и присоединитесь к Господу союзом вечным, который не забудется".
JER|50|6|Народ Мой был как погибшие овцы; пастыри их совратили их с пути, разогнали их по горам; скитались они с горы на холм, забыли ложе свое.
JER|50|7|Все, которые находили их, пожирали их, и притеснители их говорили: "мы не виноваты, потому что они согрешили пред Господом, пред жилищем правды и пред Господом, надеждою отцов их".
JER|50|8|Бегите из среды Вавилона, и уходите из Халдейской земли, и будьте как козлы впереди стада овец.
JER|50|9|Ибо вот, Я подниму и приведу на Вавилон сборище великих народов от земли северной, и расположатся против него, и он будет взят; стрелы у них, как у искусного воина, не возвращаются даром.
JER|50|10|И Халдея сделается добычею их; и опустошители ее насытятся, говорит Господь.
JER|50|11|Ибо вы веселились, вы торжествовали, расхитители наследия Моего; прыгали от радости, как телица на траве, и ржали, как боевые кони.
JER|50|12|В большом стыде будет мать ваша, покраснеет родившая вас; вот будущность тех народов – пустыня, сухая земля и степь.
JER|50|13|От гнева Господа она сделается необитаемою, и вся она будет пуста; всякий проходящий чрез Вавилон изумится и посвищет, смотря на все язвы его.
JER|50|14|Выстройтесь в боевой порядок вокруг Вавилона; все, натягивающие лук, стреляйте в него, не жалейте стрел, ибо он согрешил против Господа.
JER|50|15|Поднимите крик против него со всех сторон; он подал руку свою; пали твердыни его, рушились стены его, ибо это – возмездие Господа; отмщайте ему; как он поступал, так и вы поступайте с ним.
JER|50|16|Истребите в Вавилоне [и] сеющего и действующего серпом во время жатвы; от страха губительного меча пусть каждый возвратится к народу своему, и каждый пусть бежит в землю свою.
JER|50|17|Израиль – рассеянное стадо; львы разогнали [его]; прежде объедал его царь Ассирийский, а сей последний, Навуходоносор, царь Вавилонский, и кости его сокрушил.
JER|50|18|Посему так говорит Господь Саваоф, Бог Израилев: вот, Я посещу царя Вавилонского и землю его, как посетил царя Ассирийского.
JER|50|19|И возвращу Израиля на пажить его, и будет он пастись на Кармиле и Васане, и душа его насытится на горе Ефремовой и в Галааде.
JER|50|20|В те дни и в то время, говорит Господь, будут искать неправды Израилевой, и не будет ее, и грехов Иуды, и не найдется их; ибо прощу тех, которых оставлю [в живых].
JER|50|21|Иди на нее, на землю возмутительную, и накажи жителей ее; опустошай и истребляй все за ними, говорит Господь, и сделай все, что Я повелел тебе.
JER|50|22|Шум брани на земле и великое разрушение!
JER|50|23|Как разбит и сокрушен молот всей земли! Как Вавилон сделался ужасом между народами!
JER|50|24|Я расставил сети для тебя, и ты пойман, Вавилон, не предвидя того; ты найден и схвачен, потому что восстал против Господа.
JER|50|25|Господь открыл хранилище Свое и взял [из него] сосуды гнева Своего, потому что у Господа Бога Саваофа есть дело в земле Халдейской.
JER|50|26|Идите на нее со всех краев, растворяйте житницы ее, топчите ее как снопы, совсем истребите ее, чтобы ничего от нее не осталось.
JER|50|27|Убивайте всех волов ее, пусть идут на заклание; горе им! ибо пришел день их, время посещения их.
JER|50|28|[Слышен] голос бегущих и спасающихся из земли Вавилонской, чтобы возвестить на Сионе о мщении Господа Бога нашего, о мщении за храм Его.
JER|50|29|Созовите против Вавилона стрельцов; все, напрягающие лук, расположитесь станом вокруг него, чтобы никто не спасся из него; воздайте ему по делам его; как он поступал, так поступите и с ним, ибо он вознесся против Господа, против Святаго Израилева.
JER|50|30|За то падут юноши его на улицах его, и все воины его истреблены будут в тот день, говорит Господь.
JER|50|31|Вот, Я – на тебя, гордыня, говорит Господь Бог Саваоф; ибо пришел день твой, время посещения твоего.
JER|50|32|И споткнется гордыня, и упадет, и никто не поднимет его; и зажгу огонь в городах его, и пожрет все вокруг него.
JER|50|33|Так говорит Господь Саваоф: угнетены сыновья Израиля, как и сыновья Иуды, и все, пленившие их, крепко держат их и не хотят отпустить их.
JER|50|34|Но Искупитель их силен, Господь Саваоф имя Его; Он разберет дело их, чтобы успокоить землю и привести в трепет жителей Вавилона.
JER|50|35|Меч на Халдеев, говорит Господь, и на жителей Вавилона, и на князей его, и на мудрых его;
JER|50|36|меч на обаятелей, и они обезумеют; меч на воинов его, и они оробеют;
JER|50|37|меч на коней его и на колесницы его и на все разноплеменные народы среди него, и они будут как женщины; меч на сокровища его, и они будут расхищены;
JER|50|38|засуха на воды его, и они иссякнут; ибо это земля истуканов, и они обезумеют от идольских страшилищ.
JER|50|39|И поселятся там степные звери с шакалами, и будут жить на ней страусы, и не будет обитаема во веки и населяема в роды родов.
JER|50|40|Как ниспровержены Богом Содом и Гоморра и соседние города их, говорит Господь, так [и] тут ни один человек не будет жить, и сын человеческий не будет останавливаться.
JER|50|41|Вот, идет народ от севера, и народ великий, и многие цари поднимаются от краев земли;
JER|50|42|держат в руках лук и копье; они жестоки и немилосерды; голос их шумен, как море; несутся на конях, выстроились как один человек, чтобы сразиться с тобою, дочь Вавилона.
JER|50|43|Услышал царь Вавилонский весть о них, и руки у него опустились; скорбь объяла его, муки, как женщину в родах.
JER|50|44|Вот, восходит он, как лев, от возвышения Иордана на укрепленные жилища; но Я заставлю их поспешно уйти из него, и, кто избран, тому вверю его. Ибо кто подобен Мне? и кто потребует от Меня ответа? И какой пастырь противостанет Мне?
JER|50|45|Итак выслушайте определение Господа, какое Он постановил о Вавилоне, и намерения Его, какие Он имеет о земле Халдейской: истинно, самые малые из стад повлекут их; истинно, он опустошит жилища их с ними.
JER|50|46|От шума взятия Вавилона потрясется земля, и вопль будет слышен между народами.
JER|51|1|Так говорит Господь: вот, Я подниму на Вавилон и на живущих среди него противников Моих.
JER|51|2|И пошлю на Вавилон веятелей, и развеют его, и опустошат землю его; ибо в день бедствия нападут на него со всех сторон.
JER|51|3|Пусть стрелец напрягает лук против напрягающего [лук] и на величающегося бронею своею; и не щадите юношей его, истребите все войско его.
JER|51|4|Пораженные пусть падут на земле Халдейской, и пронзенные – на дорогах ее.
JER|51|5|Ибо не овдовел Израиль и Иуда от Бога Своего, Господа Саваофа; хотя земля их полна грехами пред Святым Израилевым.
JER|51|6|Бегите из среды Вавилона и спасайте каждый душу свою, чтобы не погибнуть от беззакония его, ибо это время отмщения у Господа, Он воздает ему воздаяние.
JER|51|7|Вавилон был золотою чашею в руке Господа, опьянявшею всю землю; народы пили из нее вино и безумствовали.
JER|51|8|Внезапно пал Вавилон и разбился; рыдайте о нем, возьмите бальзама для раны его: может быть, он исцелеет.
JER|51|9|Врачевали мы Вавилон, но не исцелился; оставьте его, и пойдем каждый в свою землю, потому что приговор о нем достиг до небес и поднялся до облаков.
JER|51|10|Господь вывел на свет правду нашу; пойдем и возвестим на Сионе дело Господа Бога нашего.
JER|51|11|Острите стрелы, наполняйте колчаны; Господь возбудил дух царей Мидийских, потому что у Него есть намерение против Вавилона, чтобы истребить его, ибо это есть отмщение Господа, отмщение за храм Его.
JER|51|12|Против стен Вавилона поднимите знамя, усильте надзор, расставьте сторожей, приготовьте засады, ибо, как Господь помыслил, так и сделает, что изрек на жителей Вавилона.
JER|51|13|О, ты, живущий при водах великих, изобилующий сокровищами! пришел конец твой, мера жадности твоей.
JER|51|14|Господь Саваоф поклялся Самим Собою: истинно говорю, что наполню тебя людьми, как саранчою, и поднимут крик против тебя.
JER|51|15|Он сотворил землю силою Своею, утвердил вселенную мудростью Своею и разумом Своим распростер небеса.
JER|51|16|По гласу Его шумят воды на небесах, и Он возводит облака от краев земли, творит молнии среди дождя и изводит ветер из хранилищ Своих.
JER|51|17|Безумствует всякий человек в своем знании, срамит себя всякий плавильщик истуканом своим, ибо истукан его есть ложь, и нет в нем духа.
JER|51|18|Это совершенная пустота, дело заблуждения; во время посещения их они исчезнут.
JER|51|19|Не такова, как их, доля Иакова, ибо [Бог его] есть Творец всего, и [Израиль] есть жезл наследия Его, имя Его – Господь Саваоф.
JER|51|20|Ты у Меня – молот, оружие воинское; тобою Я поражал народы и тобою разорял царства;
JER|51|21|тобою поражал коня и всадника его и тобою поражал колесницу и возницу ее;
JER|51|22|тобою поражал мужа и жену, тобою поражал и старого и молодого, тобою поражал и юношу и девицу;
JER|51|23|и тобою поражал пастуха и стадо его, тобою поражал и земледельца и рабочий скот его, тобою поражал и областеначальников и градоправителей.
JER|51|24|И воздам Вавилону и всем жителям Халдеи за все то зло, какое они делали на Сионе в глазах ваших, говорит Господь.
JER|51|25|Вот, Я – на тебя, гора губительная, говорит Господь, разоряющая всю землю, и простру на тебя руку Мою, и низрину тебя со скал, и сделаю тебя горою обгорелою.
JER|51|26|И не возьмут из тебя камня для углов и камня для основания, но вечно будешь запустением, говорит Господь.
JER|51|27|Поднимите знамя на земле, трубите трубою среди народов, вооружите против него народы, созовите на него царства Араратские, Минийские и Аскеназские, поставьте вождя против него, наведите коней, как страшную саранчу.
JER|51|28|Вооружите против него народы, царей Мидии, областеначальников ее и всех градоправителей ее, и всю землю, подвластную ей.
JER|51|29|Трясется земля и трепещет, ибо исполняются над Вавилоном намерения Господа сделать землю Вавилонскую пустынею, без жителей.
JER|51|30|Перестали сражаться сильные Вавилонские, сидят в укреплениях своих; истощилась сила их, сделались как женщины, жилища их сожжены, затворы их сокрушены.
JER|51|31|Гонец бежит навстречу гонцу, и вестник навстречу вестнику, чтобы возвестить царю Вавилонскому, что город его взят со всех концов,
JER|51|32|и броды захвачены, и ограды сожжены огнем, и воины поражены страхом.
JER|51|33|Ибо так говорит Господь Саваоф, Бог Израилев: дочь Вавилона подобна гумну во время молотьбы на нем; еще немного, и наступит время жатвы ее.
JER|51|34|Пожирал меня и грыз меня Навуходоносор, царь Вавилонский; сделал меня пустым сосудом; поглощал меня, как дракон; наполнял чрево свое сластями моими, извергал меня.
JER|51|35|Обида моя и плоть моя – на Вавилоне, скажет обитательница Сиона, и кровь моя – на жителях Халдеи, скажет Иерусалим.
JER|51|36|Посему так говорит Господь: вот, Я вступлюсь в твое дело и отмщу за тебя, и осушу море его, и иссушу каналы его.
JER|51|37|И Вавилон будет грудою развалин, жилищем шакалов, ужасом и посмеянием, без жителей.
JER|51|38|Как львы зарыкают все они, и заревут как щенки львиные.
JER|51|39|Во время разгорячения их сделаю им пир и упою их, чтобы они повеселились и заснули вечным сном, и не пробуждались, говорит Господь.
JER|51|40|Сведу их как ягнят на заклание, как овнов с козлами.
JER|51|41|Как взят Сесах, и завоевана слава всей земли! Как сделался Вавилон ужасом между народами!
JER|51|42|Устремилось на Вавилон море; он покрыт множеством волн его.
JER|51|43|Города его сделались пустыми, землею сухою, степью, землею, где не живет ни один человек и где не проходит сын человеческий.
JER|51|44|И посещу Вила в Вавилоне, и исторгну из уст его проглоченное им, и народы не будут более стекаться к нему, даже и стены Вавилонские падут.
JER|51|45|Выходи из среды его, народ Мой, и спасайте каждый душу свою от пламенного гнева Господа.
JER|51|46|Да не ослабевает сердце ваше, и не бойтесь слуха, который будет слышен на земле; слух придет в [один] год, и потом в [другой] год, и на земле [будет] насилие, властелин [восстанет] на властелина.
JER|51|47|Посему вот, приходят дни, когда Я посещу идолов Вавилона, и вся земля его будет посрамлена, и все пораженные его падут среди него.
JER|51|48|И восторжествуют над Вавилоном небо и земля и все, что на них; ибо от севера придут к нему опустошители, говорит Господь.
JER|51|49|Как Вавилон повергал пораженных Израильтян, так в Вавилоне будут повержены пораженные всей страны.
JER|51|50|Спасшиеся от меча, уходите, не останавливайтесь, вспомните издали о Господе, и да взойдет Иерусалим на сердце ваше.
JER|51|51|Стыдно нам было, когда мы слышали ругательство: бесчестие покрывало лица наши, когда чужеземцы пришли во святилище дома Господня.
JER|51|52|За то вот, приходят дни, говорит Господь, когда Я посещу истуканов его, и по всей земле его будут стонать раненые.
JER|51|53|Хотя бы Вавилон возвысился до небес, и хотя бы он на высоте укрепил твердыню свою; [но] от Меня придут к нему опустошители, говорит Господь.
JER|51|54|[Пронесется] гул вопля от Вавилона и великое разрушение – от земли Халдейской,
JER|51|55|ибо Господь опустошит Вавилон и положит конец горделивому голосу в нем. Зашумят волны их как большие воды, раздастся шумный голос их.
JER|51|56|Ибо придет на него, на Вавилон, опустошитель, и взяты будут ратоборцы его, сокрушены будут луки их; ибо Господь, Бог воздаяний, воздаст воздаяние.
JER|51|57|И напою допьяна князей его и мудрецов его, областеначальников его, и градоправителей его, и воинов его, и заснут сном вечным, и не пробудятся, говорит Царь – Господь Саваоф имя Его.
JER|51|58|Так говорит Господь Саваоф: толстые стены Вавилона до основания будут разрушены, и высокие ворота его будут сожжены огнем; итак напрасно трудились народы, и племена мучили себя для огня.
JER|51|59|Слово, которое пророк Иеремия заповедал Сераии, сыну Нирии, сыну Маасеи, когда он отправлялся в Вавилон с Седекиею, царем Иудейским, в четвертый год его царствования; Сераия был главный постельничий.
JER|51|60|Иеремия вписал в одну книгу все бедствия, какие должны были придти на Вавилон, все сии речи, написанные на Вавилон.
JER|51|61|И сказал Иеремия Сераии: когда ты придешь в Вавилон, то смотри, прочитай все сии речи,
JER|51|62|и скажи: "Господи! Ты изрек о месте сем, что истребишь его так, что не останется в нем ни человека, ни скота, но оно будет вечною пустынею".
JER|51|63|И когда окончишь чтение сей книги, привяжи к ней камень и брось ее в средину Евфрата,
JER|51|64|и скажи: "так погрузится Вавилон и не восстанет от того бедствия, которое Я наведу на него, и они совершенно изнемогут". Доселе речи Иеремии.
JER|52|1|Седекия был двадцати одного года, когда начал царствовать, и царствовал в Иерусалиме одиннадцать лет; имя матери его – Хамуталь, дочь Иеремии из Ливны.
JER|52|2|И он делал злое в очах Господа, все то, что делал Иоаким;
JER|52|3|посему гнев Господа был над Иерусалимом и Иудою до того, что Он отверг их от лица Своего; и Седекия отложился от царя Вавилонского.
JER|52|4|И было, в девятый год его царствования, в десятый месяц, в десятый день месяца, пришел Навуходоносор, царь Вавилонский, сам и все войско его, к Иерусалиму, и обложили его, и устроили вокруг него насыпи.
JER|52|5|И находился город в осаде до одиннадцатого года царя Седекии.
JER|52|6|В четвертом месяце, в девятый день месяца, голод в городе усилился, и не было хлеба у народа земли.
JER|52|7|Сделан был пролом в город, и побежали все военные, и вышли из города ночью воротами, находящимися между двумя стенами, подле царского сада, и пошли дорогою степи; Халдеи же были вокруг города.
JER|52|8|Войско Халдейское погналось за царем, и настигли Седекию на равнинах Иерихонских, и все войско его разбежалось от него.
JER|52|9|И взяли царя, и привели его к царю Вавилонскому, в Ривлу, в землю Емаф, где он произнес над ним суд.
JER|52|10|И заколол царь Вавилонский сыновей Седекии пред глазами его, и всех князей Иудейских заколол в Ривле.
JER|52|11|А Седекии выколол глаза и велел оковать его медными оковами; и отвел его царь Вавилонский в Вавилон и посадил его в дом стражи до дня смерти его.
JER|52|12|В пятый месяц, в десятый день месяца, – это был девятнадцатый год царя Навуходоносора, царя Вавилонского, – пришел Навузардан, начальник телохранителей, предстоявший пред царем Вавилонским, в Иерусалим
JER|52|13|и сожег дом Господень, и дом царя, и все домы в Иерусалиме, и все домы большие сожег огнем.
JER|52|14|И все войско Халдейское, бывшее с начальником телохранителей, разрушило все стены вокруг Иерусалима.
JER|52|15|Бедных из народа и прочий народ, остававшийся в городе, и переметчиков, которые передались царю Вавилонскому, и вообще остаток простого народа Навузардан, начальник телохранителей, выселил.
JER|52|16|Только несколько из бедного народа земли Навузардан, начальник телохранителей, оставил для виноградников и земледелия.
JER|52|17|И столбы медные, которые были в доме Господнем, и подставы, и медное море, которое в доме Господнем, изломали Халдеи и отнесли всю медь их в Вавилон.
JER|52|18|И тазы, и лопатки, и ножи, и чаши, и ложки, и все медные сосуды, которые употребляемы были при Богослужении, взяли;
JER|52|19|и блюда, и щипцы, и чаши, и котлы, и лампады, и фимиамники, и кружки, что было золотое – золотое, и что было серебряное – серебряное, взял начальник телохранителей;
JER|52|20|также два столба, одно море и двенадцать медных волов, которые служили подставами, которые царь Соломон сделал в доме Господнем, – меди во всех этих вещах невозможно было взвесить.
JER|52|21|Столбы сии были каждый столб в восемнадцать локтей вышины, и шнурок в двенадцать локтей обнимал его, а толщина стенок его внутри пустого, в четыре перста.
JER|52|22|И венец на нем медный, а высота венца пять локтей; и сетка и гранатовые яблоки вокруг были все медные; то же и на другом столбе с гранатовыми яблоками.
JER|52|23|Гранатовых яблоков было по всем сторонам девяносто шесть; всех яблоков вокруг сетки сто.
JER|52|24|Начальник телохранителей взял также Сераию первосвященника и Цефанию, второго священника, и трех сторожей порога.
JER|52|25|И из города взял одного евнуха, который был начальником над военными людьми, и семь человек предстоявших лицу царя, которые находились в городе, и главного писца в войске, записывавшего в войско народ земли, и шестьдесят человек из народа страны, найденных в городе.
JER|52|26|И взял их Навузардан, начальник телохранителей, и отвел их к царю Вавилонскому в Ривлу.
JER|52|27|И поразил их царь Вавилонский и умертвил их в Ривле, в земле Емаф; и выселен был Иуда из земли своей.
JER|52|28|Вот народ, который выселил Навуходоносор: в седьмой год три тысячи двадцать три Иудея;
JER|52|29|в восемнадцатый год Навуходоносора из Иерусалима [выселено] восемьсот тридцать две души;
JER|52|30|в двадцать третий год Навуходоносора Навузардан, начальник телохранителей, выселил Иудеев семьсот сорок пять душ: всего четыре тысячи шестьсот душ.
JER|52|31|В тридцать седьмой год после переселения Иоакима, царя Иудейского, в двенадцатый месяц, в двадцать пятый день месяца, Евильмеродах, царь Вавилонский, в первый год царствования своего, возвысил Иоакима, царя Иудейского, и вывел его из темничного дома.
JER|52|32|И беседовал с ним дружелюбно, и поставил престол его выше престола царей, которые были у него в Вавилоне;
JER|52|33|и переменил темничные одежды его, и он всегда у него обедал во все дни жизни своей.
JER|52|34|И содержание его, содержание постоянное, выдаваемо было ему от царя изо дня в день до дня смерти его, во все дни жизни его.
