NEH|1|1|The words of Nehemiah the son of Hacaliah. Now it happened in the month of Chislev, in the twentieth year, as I was in Susa the capital,
NEH|1|2|that Hanani, one of my brothers, came with certain men from Judah. And I asked them concerning the Jews who escaped, who had survived the exile, and concerning Jerusalem.
NEH|1|3|And they said to me, "The remnant there in the province who had survived the exile is in great trouble and shame. The wall of Jerusalem is broken down, and its gates are destroyed by fire."
NEH|1|4|As soon as I heard these words I sat down and wept and mourned for days, and I continued fasting and praying before the God of heaven.
NEH|1|5|And I said, "O LORD God of heaven, the great and awesome God who keeps covenant and steadfast love with those who love him and keep his commandments,
NEH|1|6|let your ear be attentive and your eyes open, to hear the prayer of your servant that I now pray before you day and night for the people of Israel your servants, confessing the sins of the people of Israel, which we have sinned against you. Even I and my father's house have sinned.
NEH|1|7|We have acted very corruptly against you and have not kept the commandments, the statutes, and the rules that you commanded your servant Moses.
NEH|1|8|Remember the word that you commanded your servant Moses, saying, 'If you are unfaithful, I will scatter you among the peoples,
NEH|1|9|but if you return to me and keep my commandments and do them, though your dispersed be under the farthest skies, I will gather them from there and bring them to the place that I have chosen, to make my name dwell there.'
NEH|1|10|They are your servants and your people, whom you have redeemed by your great power and by your strong hand.
NEH|1|11|O Lord, let your ear be attentive to the prayer of your servant, and to the prayer of your servants who delight to fear your name, and give success to your servant today, and grant him mercy in the sight of this man." Now I was cupbearer to the king.
NEH|2|1|In the month of Nisan, in the twentieth year of King Artaxerxes, when wine was before him, I took up the wine and gave it to the king. Now I had not been sad in his presence.
NEH|2|2|And the king said to me, "Why is your face sad, seeing you are not sick? This is nothing but sadness of the heart." Then I was very much afraid.
NEH|2|3|I said to the king, "Let the king live forever! Why should not my face be sad, when the city, the place of my fathers' graves, lies in ruins, and its gates have been destroyed by fire?"
NEH|2|4|Then the king said to me, "What are you requesting?" So I prayed to the God of heaven.
NEH|2|5|And I said to the king, "If it pleases the king, and if your servant has found favor in your sight, that you send me to Judah, to the city of my fathers' graves, that I may rebuild it."
NEH|2|6|And the king said to me (the queen sitting beside him), "How long will you be gone, and when will you return?" So it pleased the king to send me when I had given him a time.
NEH|2|7|And I said to the king, "If it pleases the king, let letters be given me to the governors of the province Beyond the River, that they may let me pass through until I come to Judah,
NEH|2|8|and a letter to Asaph, the keeper of the king's forest, that he may give me timber to make beams for the gates of the fortress of the temple, and for the wall of the city, and for the house that I shall occupy." And the king granted me what I asked, for the good hand of my God was upon me.
NEH|2|9|Then I came to the governors of the province Beyond the River and gave them the king's letters. Now the king had sent with me officers of the army and horsemen.
NEH|2|10|But when Sanballat the Horonite and Tobiah, the Ammonite servant, heard this, it displeased them greatly that someone had come to seek the welfare of the people of Israel.
NEH|2|11|So I went to Jerusalem and was there three days.
NEH|2|12|Then I arose in the night, I and a few men with me. And I told no one what my God had put into my heart to do for Jerusalem. There was no animal with me but the one on which I rode.
NEH|2|13|I went out by night by the Valley Gate to the Dragon Spring and to the Dung Gate, and I inspected the walls of Jerusalem that were broken down and its gates that had been destroyed by fire.
NEH|2|14|Then I went on to the Fountain Gate and to the King's Pool, but there was no room for the animal that was under me to pass.
NEH|2|15|Then I went up in the night by the valley and inspected the wall, and I turned back and entered by the Valley Gate, and so returned.
NEH|2|16|And the officials did not know where I had gone or what I was doing, and I had not yet told the Jews, the priests, the nobles, the officials, and the rest who were to do the work.
NEH|2|17|Then I said to them, "You see the trouble we are in, how Jerusalem lies in ruins with its gates burned. Come, let us build the wall of Jerusalem, that we may no longer suffer derision."
NEH|2|18|And I told them of the hand of my God that had been upon me for good, and also of the words that the king had spoken to me. And they said, "Let us rise up and build." So they strengthened their hands for the good work.
NEH|2|19|But when Sanballat the Horonite and Tobiah the Ammonite servant and Geshem the Arab heard of it, they jeered at us and despised us and said, "What is this thing that you are doing? Are you rebelling against the king?"
NEH|2|20|Then I replied to them, "The God of heaven will make us prosper, and we his servants will arise and build, but you have no portion or right or claim in Jerusalem."
NEH|3|1|Then Eliashib the high priest rose up with his brothers the priests, and they built the Sheep Gate. They consecrated it and set its doors. They consecrated it as far as the Tower of the Hundred, as far as the Tower of Hananel.
NEH|3|2|And next to him the men of Jericho built. And next to them Zaccur the son of Imri built.
NEH|3|3|The sons of Hassenaah built the Fish Gate. They laid its beams and set its doors, its bolts, and its bars.
NEH|3|4|And next to them Meremoth the son of Uriah, son of Hakkoz repaired. And next to them Meshullam the son of Berechiah, son of Meshezabel repaired. And next to them Zadok the son of Baana repaired.
NEH|3|5|And next to them the Tekoites repaired, but their nobles would not stoop to serve their Lord.
NEH|3|6|Joiada the son of Paseah and Meshullam the son of Besodeiah repaired the Gate of Yeshanah. They laid its beams and set its doors, its bolts, and its bars.
NEH|3|7|And next to them repaired Melatiah the Gibeonite and Jadon the Meronothite, the men of Gibeon and of Mizpah, the seat of the governor of the province Beyond the River.
NEH|3|8|Next to them Uzziel the son of Harhaiah, goldsmiths, repaired. Next to him Hananiah, one of the perfumers, repaired, and they restored Jerusalem as far as the Broad Wall.
NEH|3|9|Next to them Rephaiah the son of Hur, ruler of half the district of Jerusalem, repaired.
NEH|3|10|Next to them Jedaiah the son of Harumaph repaired opposite his house. And next to him Hattush the son of Hashabneiah repaired.
NEH|3|11|Malchijah the son of Harim and Hasshub the son of Pahath-moab repaired another section and the Tower of the Ovens.
NEH|3|12|Next to him Shallum the son of Hallohesh, ruler of half the district of Jerusalem, repaired, he and his daughters.
NEH|3|13|Hanun and the inhabitants of Zanoah repaired the Valley Gate. They rebuilt it and set its doors, its bolts, and its bars, and repaired a thousand cubits of the wall, as far as the Dung Gate.
NEH|3|14|Malchijah the son of Rechab, ruler of the district of Beth-haccherem, repaired the Dung Gate. He rebuilt it and set its doors, its bolts, and its bars.
NEH|3|15|And Shallum the son of Col-hozeh, ruler of the district of Mizpah, repaired the Fountain Gate. He rebuilt it and covered it and set its doors, its bolts, and its bars. And he built the wall of the Pool of Shelah of the king's garden, as far as the stairs that go down from the City of David.
NEH|3|16|After him Nehemiah the son of Azbuk, ruler of half the district of Beth-zur, repaired to a point opposite the tombs of David, as far as the artificial pool, and as far as the house of the mighty men.
NEH|3|17|After him the Levites repaired: Rehum the son of Bani. Next to him Hashabiah, ruler of half the district of Keilah, repaired for his district.
NEH|3|18|After him their brothers repaired: Bavvai the son of Henadad, ruler of half the district of Keilah.
NEH|3|19|Next to him Ezer the son of Jeshua, ruler of Mizpah, repaired another section opposite the ascent to the armory at the buttress.
NEH|3|20|After him Baruch the son of Zabbai repaired another section from the buttress to the door of the house of Eliashib the high priest.
NEH|3|21|After him Meremoth the son of Uriah, son of Hakkoz repaired another section from the door of the house of Eliashib to the end of the house of Eliashib.
NEH|3|22|After him the priests, the men of the surrounding area, repaired.
NEH|3|23|After them Benjamin and Hasshub repaired opposite their house. After them Azariah the son of Maaseiah, son of Ananiah repaired beside his own house.
NEH|3|24|After him Binnui the son of Henadad repaired another section, from the house of Azariah to the buttress
NEH|3|25|and to the corner. Palal the son of Uzai repaired opposite the buttress and the tower projecting from the upper house of the king at the court of the guard. After him Pedaiah the son of Parosh
NEH|3|26|and the temple servants living on Ophel repaired to a point opposite the Water Gate on the east and the projecting tower.
NEH|3|27|After him the Tekoites repaired another section opposite the great projecting tower as far as the wall of Ophel.
NEH|3|28|Above the Horse Gate the priests repaired, each one opposite his own house.
NEH|3|29|After them Zadok the son of Immer repaired opposite his own house. After him Shemaiah the son of Shecaniah, the keeper of the East Gate, repaired.
NEH|3|30|After him Hananiah the son of Shelemiah and Hanun the sixth son of Zalaph repaired another section. After him Meshullam the son of Berechiah repaired opposite his chamber.
NEH|3|31|After him Malchijah, one of the goldsmiths, repaired as far as the house of the temple servants and of the merchants, opposite the Muster Gate, and to the upper chamber of the corner.
NEH|3|32|And between the upper chamber of the corner and the Sheep Gate the goldsmiths and the merchants repaired.
NEH|4|1|Now when Sanballat heard that we were building the wall, he was angry and greatly enraged, and he jeered at the Jews.
NEH|4|2|And he said in the presence of his brothers and of the army of Samaria, "What are these feeble Jews doing? Will they restore it for themselves? Will they sacrifice? Will they finish up in a day? Will they revive the stones out of the heaps of rubbish, and burned ones at that?"
NEH|4|3|Tobiah the Ammonite was beside him, and he said, "Yes, what they are building- if a fox goes up on it he will break down their stone wall!"
NEH|4|4|Hear, O our God, for we are despised. Turn back their taunt on their own heads and give them up to be plundered in a land where they are captives.
NEH|4|5|Do not cover their guilt, and let not their sin be blotted out from your sight, for they have provoked you to anger in the presence of the builders.
NEH|4|6|So we built the wall. And all the wall was joined together to half its height, for the people had a mind to work.
NEH|4|7|But when Sanballat and Tobiah and the Arabs and the Ammonites and the Ashdodites heard that the repairing of the walls of Jerusalem was going forward and that the breaches were beginning to be closed, they were very angry.
NEH|4|8|And they all plotted together to come and fight against Jerusalem and to cause confusion in it.
NEH|4|9|And we prayed to our God and set a guard as a protection against them day and night.
NEH|4|10|In Judah it was said, "The strength of those who bear the burdens is failing. There is too much rubble. By ourselves we will not be able to rebuild the wall."
NEH|4|11|And our enemies said, "They will not know or see till we come among them and kill them and stop the work."
NEH|4|12|At that time the Jews who lived near them came from all directions and said to us ten times, "You must return to us."
NEH|4|13|So in the lowest parts of the space behind the wall, in open places, I stationed the people by their clans, with their swords, their spears, and their bows.
NEH|4|14|And I looked and arose and said to the nobles and to the officials and to the rest of the people, "Do not be afraid of them. Remember the Lord, who is great and awesome, and fight for your brothers, your sons, your daughters, your wives, and your homes."
NEH|4|15|When our enemies heard that it was known to us and that God had frustrated their plan, we all returned to the wall, each to his work.
NEH|4|16|From that day on, half of my servants worked on construction, and half held the spears, shields, bows, and coats of mail. And the leaders stood behind the whole house of Judah,
NEH|4|17|who were building on the wall. Those who carried burdens were loaded in such a way that each labored on the work with one hand and held his weapon with the other.
NEH|4|18|And each of the builders had his sword strapped at his side while he built. The man who sounded the trumpet was beside me.
NEH|4|19|And I said to the nobles and to the officials and to the rest of the people, "The work is great and widely spread, and we are separated on the wall, far from one another.
NEH|4|20|In the place where you hear the sound of the trumpet, rally to us there. Our God will fight for us."
NEH|4|21|So we labored at the work, and half of them held the spears from the break of dawn until the stars came out.
NEH|4|22|I also said to the people at that time, "Let every man and his servant pass the night within Jerusalem, that they may be a guard for us by night and may labor by day."
NEH|4|23|So neither I nor my brothers nor my servants nor the men of the guard who followed me, none of us took off our clothes; each kept his weapon at his right hand.
NEH|5|1|Now there arose a great outcry of the people and of their wives against their Jewish brothers.
NEH|5|2|For there were those who said, "With our sons and our daughters, we are many. So let us get grain, that we may eat and keep alive."
NEH|5|3|There were also those who said, "We are mortgaging our fields, our vineyards, and our houses to get grain because of the famine."
NEH|5|4|And there were those who said, "We have borrowed money for the king's tax on our fields and our vineyards.
NEH|5|5|Now our flesh is as the flesh of our brothers, our children are as their children. Yet we are forcing our sons and our daughters to be slaves, and some of our daughters have already been enslaved, but it is not in our power to help it, for other men have our fields and our vineyards."
NEH|5|6|I was very angry when I heard their outcry and these words.
NEH|5|7|I took counsel with myself, and I brought charges against the nobles and the officials. I said to them, "You are exacting interest, each from his brother." And I held a great assembly against them
NEH|5|8|and said to them, "We, as far as we are able, have bought back our Jewish brothers who have been sold to the nations, but you even sell your brothers that they may be sold to us!" They were silent and could not find a word to say.
NEH|5|9|So I said, "The thing that you are doing is not good. Ought you not to walk in the fear of our God to prevent the taunts of the nations our enemies?
NEH|5|10|Moreover, I and my brothers and my servants are lending them money and grain. Let us abandon this exacting of interest.
NEH|5|11|Return to them this very day their fields, their vineyards, their olive orchards, and their houses, and the percentage of money, grain, wine, and oil that you have been exacting from them."
NEH|5|12|Then they said, "We will restore these and require nothing from them. We will do as you say." And I called the priests and made them swear to do as they had promised.
NEH|5|13|I also shook out the fold of my garment and said, "So may God shake out every man from his house and from his labor who does not keep this promise. So may he be shaken out and emptied." And all the assembly said "Amen" and praised the LORD. And the people did as they had promised.
NEH|5|14|Moreover, from the time that I was appointed to be their governor in the land of Judah, from the twentieth year to the thirty-second year of Artaxerxes the king, twelve years, neither I nor my brothers ate the food allowance of the governor.
NEH|5|15|The former governors who were before me laid heavy burdens on the people and took from them for their daily ration forty shekels of silver. Even their servants lorded it over the people. But I did not do so, because of the fear of God.
NEH|5|16|I also persevered in the work on this wall, and we acquired no land, and all my servants were gathered there for the work.
NEH|5|17|Moreover, there were at my table 150 men, Jews and officials, besides those who came to us from the nations that were around us.
NEH|5|18|Now what was prepared at my expense for each day was one ox and six choice sheep and birds, and every ten days all kinds of wine in abundance. Yet for all this I did not demand the food allowance of the governor, because the service was too heavy on this people.
NEH|5|19|Remember for my good, O my God, all that I have done for this people.
NEH|6|1|Now when Sanballat and Tobiah and Geshem the Arab and the rest of our enemies heard that I had built the wall and that there was no breach left in it (although up to that time I had not set up the doors in the gates),
NEH|6|2|Sanballat and Geshem sent to me, saying, "Come and let us meet together at Hakkephirim in the plain of Ono." But they intended to do me harm.
NEH|6|3|And I sent messengers to them, saying, "I am doing a great work and I cannot come down. Why should the work stop while I leave it and come down to you?"
NEH|6|4|And they sent to me four times in this way, and I answered them in the same manner.
NEH|6|5|In the same way Sanballat for the fifth time sent his servant to me with an open letter in his hand.
NEH|6|6|In it was written, "It is reported among the nations, and Geshem also says it, that you and the Jews intend to rebel; that is why you are building the wall. And according to these reports you wish to become their king.
NEH|6|7|And you have also set up prophets to proclaim concerning you in Jerusalem, 'There is a king in Judah.' And now the king will hear of these reports. So now come and let us take counsel together."
NEH|6|8|Then I sent to him, saying, "No such things as you say have been done, for you are inventing them out of your own mind."
NEH|6|9|For they all wanted to frighten us, thinking, "Their hands will drop from the work, and it will not be done." But now, O God, strengthen my hands.
NEH|6|10|Now when I went into the house of Shemaiah the son of Delaiah, son of Mehetabel, who was confined to his home, he said, "Let us meet together in the house of God, within the temple. Let us close the doors of the temple, for they are coming to kill you. They are coming to kill you by night."
NEH|6|11|But I said, "Should such a man as I run away? And what man such as I could go into the temple and live? I will not go in."
NEH|6|12|And I understood and saw that God had not sent him, but he had pronounced the prophecy against me because Tobiah and Sanballat had hired him.
NEH|6|13|For this purpose he was hired, that I should be afraid and act in this way and sin, and so they could give me a bad name in order to taunt me.
NEH|6|14|Remember Tobiah and Sanballat, O my God, according to these things that they did, and also the prophetess Noadiah and the rest of the prophets who wanted to make me afraid.
NEH|6|15|So the wall was finished on the twenty-fifth day of the month Elul, in fifty-two days.
NEH|6|16|And when all our enemies heard of it, all the nations around us were afraid and fell greatly in their own esteem, for they perceived that this work had been accomplished with the help of our God.
NEH|6|17|Moreover, in those days the nobles of Judah sent many letters to Tobiah, and Tobiah's letters came to them.
NEH|6|18|For many in Judah were bound by oath to him, because he was the son-in-law of Shecaniah the son of Arah: and his son Jehohanan had taken the daughter of Meshullam the son of Berechiah as his wife.
NEH|6|19|Also they spoke of his good deeds in my presence and reported my words to him. And Tobiah sent letters to make me afraid.
NEH|7|1|Now when the wall had been built and I had set up the doors, and the gatekeepers, the singers, and the Levites had been appointed,
NEH|7|2|I gave my brother Hanani and Hananiah the governor of the castle charge over Jerusalem, for he was a more faithful and God-fearing man than many.
NEH|7|3|And I said to them, "Let not the gates of Jerusalem be opened until the sun is hot. And while they are still standing guard, let them shut and bar the doors. Appoint guards from among the inhabitants of Jerusalem, some at their guard posts and some in front of their own homes."
NEH|7|4|The city was wide and large, but the people within it were few, and no houses had been rebuilt.
NEH|7|5|Then my God put it into my heart to assemble the nobles and the officials and the people to be enrolled by genealogy. And I found the book of the genealogy of those who came up at the first, and I found written in it:
NEH|7|6|These were the people of the province who came up out of the captivity of those exiles whom Nebuchadnezzar the king of Babylon had carried into exile. They returned to Jerusalem and Judah, each to his town.
NEH|7|7|They came with Zerubbabel, Jeshua, Nehemiah, Azariah, Raamiah, Nahamani, Mordecai, Bilshan, Mispereth, Bigvai, Nehum, Baanah. The number of the men of the people of Israel:
NEH|7|8|the sons of Parosh, 2,172.
NEH|7|9|The sons of Shephatiah, 372.
NEH|7|10|The sons of Arah, 652.
NEH|7|11|The sons of Pahath-moab, namely the sons of Jeshua and Joab, 2,818.
NEH|7|12|The sons of Elam, 1,254.
NEH|7|13|The sons of Zattu, 845.
NEH|7|14|The sons of Zaccai, 760.
NEH|7|15|The sons of Binnui, 648.
NEH|7|16|The sons of Bebai, 628.
NEH|7|17|The sons of Azgad, 2,322.
NEH|7|18|The sons of Adonikam, 667.
NEH|7|19|The sons of Bigvai, 2,067.
NEH|7|20|The sons of Adin, 655.
NEH|7|21|The sons of Ater, namely of Hezekiah, 98.
NEH|7|22|The sons of Hashum, 328.
NEH|7|23|The sons of Bezai, 324.
NEH|7|24|The sons of Hariph, 112.
NEH|7|25|The sons of Gibeon, 95.
NEH|7|26|The men of Bethlehem and Netophah, 188.
NEH|7|27|The men of Anathoth, 128.
NEH|7|28|The men of Beth-azmaveth, 42.
NEH|7|29|The men of Kiriath-jearim, Chephirah, and Beeroth, 743.
NEH|7|30|The men of Ramah and Geba, 621.
NEH|7|31|The men of Michmas, 122.
NEH|7|32|The men of Bethel and Ai, 123.
NEH|7|33|The men of the other Nebo, 52.
NEH|7|34|The sons of the other Elam, 1,254.
NEH|7|35|The sons of Harim, 320.
NEH|7|36|The sons of Jericho, 345.
NEH|7|37|The sons of Lod, Hadid, and Ono, 721.
NEH|7|38|The sons of Senaah, 3,930.
NEH|7|39|The priests: the sons of Jedaiah, namely the house of Jeshua, 973.
NEH|7|40|The sons of Immer, 1,052.
NEH|7|41|The sons of Pashhur, 1,247.
NEH|7|42|The sons of Harim, 1,017.
NEH|7|43|The Levites: the sons of Jeshua, namely of Kadmiel of the sons of Hodevah, 74.
NEH|7|44|The singers: the sons of Asaph, 148.
NEH|7|45|The gatekeepers: the sons of Shallum, the sons of Ater, the sons of Talmon, the sons of Akkub, the sons of Hatita, the sons of Shobai, 138.
NEH|7|46|The temple servants: the sons of Ziha, the sons of Hasupha, the sons of Tabbaoth,
NEH|7|47|the sons of Keros, the sons of Sia, the sons of Padon,
NEH|7|48|the sons of Lebana, the sons of Hagaba, the sons of Shalmai,
NEH|7|49|the sons of Hanan, the sons of Giddel, the sons of Gahar,
NEH|7|50|the sons of Reaiah, the sons of Rezin, the sons of Nekoda,
NEH|7|51|the sons of Gazzam, the sons of Uzza, the sons of Paseah,
NEH|7|52|the sons of Besai, the sons of Meunim, the sons of Nephushesim,
NEH|7|53|the sons of Bakbuk, the sons of Hakupha, the sons of Harhur,
NEH|7|54|the sons of Bazlith, the sons of Mehida, the sons of Harsha,
NEH|7|55|the sons of Barkos, the sons of Sisera, the sons of Temah,
NEH|7|56|the sons of Neziah, the sons of Hatipha.
NEH|7|57|The sons of Solomon's servants: the sons of Sotai, the sons of Sophereth, the sons of Perida,
NEH|7|58|the sons of Jaala, the sons of Darkon, the sons of Giddel,
NEH|7|59|the sons of Shephatiah, the sons of Hattil, the sons of Pochereth-hazzebaim, the sons of Amon.
NEH|7|60|All the temple servants and the sons of Solomon's servants were 392.
NEH|7|61|The following were those who came up from Tel-melah, Tel-harsha, Cherub, Addon, and Immer, but they could not prove their fathers' houses nor their descent, whether they belonged to Israel:
NEH|7|62|the sons of Delaiah, the sons of Tobiah, the sons of Nekoda, 642.
NEH|7|63|Also, of the priests: the sons of Hobaiah, the sons of Hakkoz, the sons of Barzillai (who had taken a wife of the daughters of Barzillai the Gileadite and was called by their name).
NEH|7|64|These sought their registration among those enrolled in the genealogies, but it was not found there, so they were excluded from the priesthood as unclean.
NEH|7|65|The governor told them that they were not to partake of the most holy food until a priest with Urim and Thummim should arise.
NEH|7|66|The whole assembly together was 42,360,
NEH|7|67|besides their male and female servants, of whom there were 7,337. And they had 245 singers, male and female.
NEH|7|68|Their horses were 736, their mules 245,
NEH|7|69|their camels 435, and their donkeys 6,720.
NEH|7|70|Now some of the heads of fathers' houses gave to the work. The governor gave to the treasury 1,000 darics of gold, 50 basins, 30 priests' garments and 500 minas of silver.
NEH|7|71|And some of the heads of fathers' houses gave into the treasury of the work 20,000 darics of gold and 2,200 minas of silver.
NEH|7|72|And what the rest of the people gave was 20,000 darics of gold, 2,000 minas of silver, and 67 priests' garments.
NEH|7|73|So the priests, the Levites, the gatekeepers, the singers, some of the people, the temple servants, and all Israel, lived in their towns. And when the seventh month had come, the people of Israel were in their towns.
NEH|8|1|And all the people gathered as one man into the square before the Water Gate. And they told Ezra the scribe to bring the Book of the Law of Moses that the LORD had commanded Israel.
NEH|8|2|So Ezra the priest brought the Law before the assembly, both men and women and all who could understand what they heard, on the first day of the seventh month.
NEH|8|3|And he read from it facing the square before the Water Gate from early morning until midday, in the presence of the men and the women and those who could understand. And the ears of all the people were attentive to the Book of the Law.
NEH|8|4|And Ezra the scribe stood on a wooden platform that they had made for the purpose. And beside him stood Mattithiah, Shema, Anaiah, Uriah, Hilkiah, and Maaseiah on his right hand, and Pedaiah, Mishael, Malchijah, Hashum, Hashbaddanah, Zechariah, and Meshullam on his left hand.
NEH|8|5|And Ezra opened the book in the sight of all the people, for he was above all the people, and as he opened it all the people stood.
NEH|8|6|And Ezra blessed the LORD, the great God, and all the people answered, "Amen, Amen," lifting up their hands. And they bowed their heads and worshiped the LORD with their faces to the ground.
NEH|8|7|Also Jeshua, Bani, Sherebiah, Jamin, Akkub, Shabbethai, Hodiah, Maaseiah, Kelita, Azariah, Jozabad, Hanan, Pelaiah, the Levites, helped the people to understand the Law, while the people remained in their places.
NEH|8|8|They read from the book, from the Law of God, clearly, and they gave the sense, so that the people understood the reading.
NEH|8|9|And Nehemiah, who was the governor, and Ezra the priest and scribe, and the Levites who taught the people said to all the people, "This day is holy to the LORD your God; do not mourn or weep." For all the people wept as they heard the words of the Law.
NEH|8|10|Then he said to them, "Go your way. Eat the fat and drink sweet wine and send portions to anyone who has nothing ready, for this day is holy to our Lord. And do not be grieved, for the joy of the LORD is your strength."
NEH|8|11|So the Levites calmed all the people, saying, "Be quiet, for this day is holy; do not be grieved."
NEH|8|12|And all the people went their way to eat and drink and to send portions and to make great rejoicing, because they had understood the words that were declared to them.
NEH|8|13|On the second day the heads of fathers' houses of all the people, with the priests and the Levites, came together to Ezra the scribe in order to study the words of the Law.
NEH|8|14|And they found it written in the Law that the LORD had commanded by Moses that the people of Israel should dwell in booths during the feast of the seventh month,
NEH|8|15|and that they should proclaim it and publish it in all their towns and in Jerusalem, "Go out to the hills and bring branches of olive, wild olive, myrtle, palm, and other leafy trees to make booths, as it is written."
NEH|8|16|So the people went out and brought them and made booths for themselves, each on his roof, and in their courts and in the courts of the house of God, and in the square at the Water Gate and in the square at the Gate of Ephraim.
NEH|8|17|And all the assembly of those who had returned from the captivity made booths and lived in the booths, for from the days of Jeshua the son of Nun to that day the people of Israel had not done so. And there was very great rejoicing.
NEH|8|18|And day by day, from the first day to the last day, he read from the Book of the Law of God. They kept the feast seven days, and on the eighth day there was a solemn assembly, according to the rule.
NEH|9|1|Now on the twenty-fourth day of this month the people of Israel were assembled with fasting and in sackcloth, and with earth on their heads.
NEH|9|2|And the Israelites separated themselves from all foreigners and stood and confessed their sins and the iniquities of their fathers.
NEH|9|3|And they stood up in their place and read from the Book of the Law of the LORD their God for a quarter of the day; for another quarter of it they made confession and worshiped the LORD their God.
NEH|9|4|On the stairs of the Levites stood Jeshua, Bani, Kadmiel, Shebaniah, Bunni, Sherebiah, Bani, and Chenani; and they cried with a loud voice to the LORD their God.
NEH|9|5|Then the Levites, Jeshua, Kadmiel, Bani, Hashabneiah, Sherebiah, Hodiah, Shebaniah, and Pethahiah, said, "Stand up and bless the LORD your God from everlasting to everlasting. Blessed be your glorious name, which is exalted above all blessing and praise.
NEH|9|6|"You are the LORD, you alone. You have made heaven, the heaven of heavens, with all their host, the earth and all that is on it, the seas and all that is in them; and you preserve all of them; and the host of heaven worships you.
NEH|9|7|You are the LORD, the God who chose Abram and brought him out of Ur of the Chaldeans and gave him the name Abraham.
NEH|9|8|You found his heart faithful before you, and made with him the covenant to give to his offspring the land of the Canaanite, the Hittite, the Amorite, the Perizzite, the Jebusite, and the Girgashite. And you have kept your promise, for you are righteous.
NEH|9|9|"And you saw the affliction of our fathers in Egypt and heard their cry at the Red Sea,
NEH|9|10|and performed signs and wonders against Pharaoh and all his servants and all the people of his land, for you knew that they acted arrogantly against our fathers. And you made a name for yourself, as it is to this day.
NEH|9|11|And you divided the sea before them, so that they went through the midst of the sea on dry land, and you cast their pursuers into the depths, as a stone into mighty waters.
NEH|9|12|By a pillar of cloud you led them in the day, and by a pillar of fire in the night to light for them the way in which they should go.
NEH|9|13|You came down on Mount Sinai and spoke with them from heaven and gave them right rules and true laws, good statutes and commandments,
NEH|9|14|and you made known to them your holy Sabbath and commanded them commandments and statutes and a law by Moses your servant.
NEH|9|15|You gave them bread from heaven for their hunger and brought water for them out of the rock for their thirst, and you told them to go in to possess the land that you had sworn to give them.
NEH|9|16|"But they and our fathers acted presumptuously and stiffened their neck and did not obey your commandments.
NEH|9|17|They refused to obey and were not mindful of the wonders that you performed among them, but they stiffened their neck and appointed a leader to return to their slavery in Egypt. But you are a God ready to forgive, gracious and merciful, slow to anger and abounding in steadfast love, and did not forsake them.
NEH|9|18|Even when they had made for themselves a golden calf and said, 'This is your God who brought you up out of Egypt,' and had committed great blasphemies,
NEH|9|19|you in your great mercies did not forsake them in the wilderness. The pillar of cloud to lead them in the way did not depart from them by day, nor the pillar of fire by night to light for them the way by which they should go.
NEH|9|20|You gave your good Spirit to instruct them and did not withhold your manna from their mouth and gave them water for their thirst.
NEH|9|21|Forty years you sustained them in the wilderness, and they lacked nothing. Their clothes did not wear out and their feet did not swell.
NEH|9|22|"And you gave them kingdoms and peoples and allotted to them every corner. So they took possession of the land of Sihon king of Heshbon and the land of Og king of Bashan.
NEH|9|23|You multiplied their children as the stars of heaven, and you brought them into the land that you had told their fathers to enter and possess.
NEH|9|24|So the descendants went in and possessed the land, and you subdued before them the inhabitants of the land, the Canaanites, and gave them into their hand, with their kings and the peoples of the land, that they might do with them as they would.
NEH|9|25|And they captured fortified cities and a rich land, and took possession of houses full of all good things, cisterns already hewn, vineyards, olive orchards and fruit trees in abundance. So they ate and were filled and became fat and delighted themselves in your great goodness.
NEH|9|26|"Nevertheless, they were disobedient and rebelled against you and cast your law behind their back and killed your prophets, who had warned them in order to turn them back to you, and they committed great blasphemies.
NEH|9|27|Therefore you gave them into the hand of their enemies, who made them suffer. And in the time of their suffering they cried out to you and you heard them from heaven, and according to your great mercies you gave them saviors who saved them from the hand of their enemies.
NEH|9|28|But after they had rest they did evil again before you, and you abandoned them to the hand of their enemies, so that they had dominion over them. Yet when they turned and cried to you, you heard from heaven, and many times you delivered them according to your mercies.
NEH|9|29|And you warned them in order to turn them back to your law. Yet they acted presumptuously and did not obey your commandments, but sinned against your rules, which if a person does them, he shall live by them, and turned a stubborn shoulder and stiffened their neck and would not obey.
NEH|9|30|Many years you bore with them and warned them by your Spirit through your prophets. Yet they would not give ear. Therefore you gave them into the hand of the peoples of the lands.
NEH|9|31|Nevertheless, in your great mercies you did not make an end of them or forsake them, for you are a gracious and merciful God.
NEH|9|32|"Now, therefore, our God, the great, the mighty, and the awesome God, who keeps covenant and steadfast love, let not all the hardship seem little to you that has come upon us, upon our kings, our princes, our priests, our prophets, our fathers, and all your people, since the time of the kings of Assyria until this day.
NEH|9|33|Yet you have been righteous in all that has come upon us, for you have dealt faithfully and we have acted wickedly.
NEH|9|34|Our kings, our princes, our priests, and our fathers have not kept your law or paid attention to your commandments and your warnings that you gave them.
NEH|9|35|Even in their own kingdom, enjoying your great goodness that you gave them, and in the large and rich land that you set before them, they did not serve you or turn from their wicked works.
NEH|9|36|Behold, we are slaves this day; in the land that you gave to our fathers to enjoy its fruit and its good gifts, behold, we are slaves.
NEH|9|37|And its rich yield goes to the kings whom you have set over us because of our sins. They rule over our bodies and over our livestock as they please, and we are in great distress.
NEH|9|38|"Because of all this we make a firm covenant in writing; on the sealed document are the names of our princes, our Levites, and our priests."
NEH|10|1|On the seals are the names of Nehemiah the governor, the son of Hacaliah, Zedekiah,
NEH|10|2|Seraiah, Azariah, Jeremiah,
NEH|10|3|Pashhur, Amariah, Malchijah,
NEH|10|4|Hattush, Shebaniah, Malluch,
NEH|10|5|Harim, Meremoth, Obadiah,
NEH|10|6|Daniel, Ginnethon, Baruch,
NEH|10|7|Meshullam, Abijah, Mijamin,
NEH|10|8|Maaziah, Bilgai, Shemaiah; these are the priests.
NEH|10|9|And the Levites: Jeshua the son of Azaniah, Binnui of the sons of Henadad, Kadmiel;
NEH|10|10|and their brothers, Shebaniah, Hodiah, Kelita, Pelaiah, Hanan,
NEH|10|11|Mica, Rehob, Hashabiah,
NEH|10|12|Zaccur, Sherebiah, Shebaniah,
NEH|10|13|Hodiah, Bani, Beninu.
NEH|10|14|The chiefs of the people: Parosh, Pahath-moab, Elam, Zattu, Bani,
NEH|10|15|Bunni, Azgad, Bebai,
NEH|10|16|Adonijah, Bigvai, Adin,
NEH|10|17|Ater, Hezekiah, Azzur,
NEH|10|18|Hodiah, Hashum, Bezai,
NEH|10|19|Hariph, Anathoth, Nebai,
NEH|10|20|Magpiash, Meshullam, Hezir,
NEH|10|21|Meshezabel, Zadok, Jaddua,
NEH|10|22|Pelatiah, Hanan, Anaiah,
NEH|10|23|Hoshea, Hananiah, Hasshub,
NEH|10|24|Hallohesh, Pilha, Shobek,
NEH|10|25|Rehum, Hashabnah, Maaseiah,
NEH|10|26|Ahiah, Hanan, Anan,
NEH|10|27|Malluch, Harim, Baanah.
NEH|10|28|The rest of the people, the priests, the Levites, the gatekeepers, the singers, the temple servants, and all who have separated themselves from the peoples of the lands to the Law of God, their wives, their sons, their daughters, all who have knowledge and understanding,
NEH|10|29|join with their brothers, their nobles, and enter into a curse and an oath to walk in God's Law that was given by Moses the servant of God, and to observe and do all the commandments of the LORD our Lord and his rules and his statutes.
NEH|10|30|"We will not give our daughters to the peoples of the land or take their daughters for our sons.
NEH|10|31|And if the peoples of the land bring in goods or any grain on the Sabbath day to sell, we will not buy from them on the Sabbath or on a holy day. And we will forego the crops of the seventh year and the exaction of every debt.
NEH|10|32|"We also take on ourselves the obligation to give yearly a third part of a shekel for the service of the house of our God:
NEH|10|33|for the showbread, the regular grain offering, the regular burnt offering, the Sabbaths, the new moons, the appointed feasts, the holy things, and the sin offerings to make atonement for Israel, and for all the work of the house of our God.
NEH|10|34|We, the priests, the Levites, and the people, have likewise cast lots for the wood offering, to bring it into the house of our God, according to our fathers' houses, at times appointed, year by year, to burn on the altar of the LORD our God, as it is written in the Law.
NEH|10|35|We obligate ourselves to bring the firstfruits of our ground and the firstfruits of all fruit of every tree, year by year, to the house of the LORD;
NEH|10|36|also to bring to the house of our God, to the priests who minister in the house of our God, the firstborn of our sons and of our cattle, as it is written in the Law, and the firstborn of our herds and of our flocks;
NEH|10|37|and to bring the first of our dough, and our contributions, the fruit of every tree, the wine and the oil, to the priests, to the chambers of the house of our God; and to bring to the Levites the tithes from our ground, for it is the Levites who collect the tithes in all our towns where we labor.
NEH|10|38|And the priest, the son of Aaron, shall be with the Levites when the Levites receive the tithes. And the Levites shall bring up the tithe of the tithes to the house of our God, to the chambers of the storehouse.
NEH|10|39|For the people of Israel and the sons of Levi shall bring the contribution of grain, wine, and oil to the chambers, where the vessels of the sanctuary are, as well as the priests who minister, and the gatekeepers and the singers. We will not neglect the house of our God."
NEH|11|1|Now the leaders of the people lived in Jerusalem. And the rest of the people cast lots to bring one out of ten to live in Jerusalem the holy city, while nine out of ten remained in the other towns.
NEH|11|2|And the people blessed all the men who willingly offered to live in Jerusalem.
NEH|11|3|These are the chiefs of the province who lived in Jerusalem; but in the towns of Judah everyone lived on his property in their towns: Israel, the priests, the Levites, the temple servants, and the descendants of Sol-omon's servants.
NEH|11|4|And in Jerusalem lived certain of the sons of Judah and of the sons of Benjamin. Of the sons of Judah: Athaiah the son of Uzziah, son of Zechariah, son of Amariah, son of Shephatiah, son of Mahalalel, of the sons of Perez;
NEH|11|5|and Maaseiah the son of Baruch, son of Col-hozeh, son of Hazaiah, son of Adaiah, son of Joiarib, son of Zechariah, son of the Shilonite.
NEH|11|6|All the sons of Perez who lived in Jerusalem were 468 valiant men.
NEH|11|7|And these are the sons of Benjamin: Sallu the son of Meshullam, son of Joed, son of Pedaiah, son of Kolaiah, son of Maaseiah, son of Ithiel, son of Jeshaiah,
NEH|11|8|and his brothers, men of valor, 928.
NEH|11|9|Joel the son of Zichri was their overseer; and Judah the son of Hassenuah was second over the city.
NEH|11|10|Of the priests: Jedaiah the son of Joiarib, Jachin,
NEH|11|11|Seraiah the son of Hilkiah, son of Meshullam, son of Zadok, son of Meraioth, son of Ahitub, ruler of the house of God,
NEH|11|12|and their brothers who did the work of the house, 822; and Adaiah the son of Jeroham, son of Pelaliah, son of Amzi, son of Zechariah, son of Pashhur, son of Malchijah,
NEH|11|13|and his brothers, heads of fathers' houses, 242; and Amashsai, the son of Azarel, son of Ahzai, son of Meshillemoth, son of Immer,
NEH|11|14|and their brothers, mighty men of valor, 128; their overseer was Zabdiel the son of Haggedolim.
NEH|11|15|And of the Levites: Shemaiah the son of Hasshub, son of Azrikam, son of Hashabiah, son of Bunni;
NEH|11|16|and Shabbethai and Jozabad, of the chiefs of the Levites, who were over the outside work of the house of God;
NEH|11|17|and Mattaniah the son of Mica, son of Zabdi, son of Asaph, who was the leader of the praise, who gave thanks, and Bakbukiah, the second among his brothers; and Abda the son of Shammua, son of Galal, son of Jeduthun.
NEH|11|18|All the Levites in the holy city were 284.
NEH|11|19|The gatekeepers, Akkub, Talmon and their brothers, who kept watch at the gates, were 172.
NEH|11|20|And the rest of Israel, and of the priests and the Levites, were in all the towns of Judah, every one in his inheritance.
NEH|11|21|But the temple servants lived on Ophel; and Ziha and Gishpa were over the temple servants.
NEH|11|22|The overseer of the Levites in Jerusalem was Uzzi the son of Bani, son of Hashabiah, son of Mattaniah, son of Mica, of the sons of Asaph, the singers, over the work of the house of God.
NEH|11|23|For there was a command from the king concerning them, and a fixed provision for the singers, as every day required.
NEH|11|24|And Pethahiah the son of Meshezabel, of the sons of Zerah the son of Judah, was at the king's side in all matters concerning the people.
NEH|11|25|And as for the villages, with their fields, some of the people of Judah lived in Kiriath-arba and its villages, and in Dibon and its villages, and in Jekabzeel and its villages,
NEH|11|26|and in Jeshua and in Moladah and Beth-pelet,
NEH|11|27|in Hazar-shual, in Beersheba and its villages,
NEH|11|28|in Ziklag, in Meconah and its villages,
NEH|11|29|in En-rimmon, in Zorah, in Jarmuth,
NEH|11|30|Zanoah, Adullam, and their villages, Lachish and its fields, and Azekah and its villages. So they encamped from Beersheba to the valley of Hinnom.
NEH|11|31|The people of Benjamin also lived from Geba onward, at Michmash, Aija, Bethel and its villages,
NEH|11|32|Anathoth, Nob, Ananiah,
NEH|11|33|Hazor, Ramah, Gittaim,
NEH|11|34|Hadid, Zeboim, Neballat,
NEH|11|35|Lod, and Ono, the valley of craftsmen.
NEH|11|36|And certain divisions of the Levites in Judah were assigned to Benjamin.
NEH|12|1|These are the priests and the Levites who came up with Zerubbabel the son of Shealtiel, and Jeshua: Seraiah, Jeremiah, Ezra,
NEH|12|2|Amariah, Malluch, Hattush,
NEH|12|3|Shecaniah, Rehum, Meremoth,
NEH|12|4|Iddo, Gin-nethoi, Abijah,
NEH|12|5|Mijamin, Maadiah, Bilgah,
NEH|12|6|Shemaiah, Joiarib, Jedaiah,
NEH|12|7|Sallu, Amok, Hilkiah, Jedaiah. These were the chiefs of the priests and of their brothers in the days of Jeshua.
NEH|12|8|And the Levites: Jeshua, Binnui, Kadmiel, Sherebiah, Judah, and Mattaniah, who with his brothers was in charge of the songs of thanksgiving.
NEH|12|9|And Bakbukiah and Unni and their brothers stood opposite them in the service.
NEH|12|10|And Jeshua was the father of Joiakim, Joiakim the father of Eliashib, Eliashib the father of Joiada,
NEH|12|11|Joiada the father of Jonathan, and Jonathan the father of Jaddua.
NEH|12|12|And in the days of Joiakim were priests, heads of fathers' houses: of Seraiah, Meraiah; of Jeremiah, Hananiah;
NEH|12|13|of Ezra, Meshullam; of Amariah, Jehohanan;
NEH|12|14|of Malluchi, Jonathan; of Shebaniah, Joseph;
NEH|12|15|of Harim, Adna; of Meraioth, Helkai;
NEH|12|16|of Iddo, Zechariah; of Ginnethon, Meshullam;
NEH|12|17|of Abijah, Zichri; of Miniamin, of Moadiah, Piltai;
NEH|12|18|of Bilgah, Shammua; of Shemaiah, Jehonathan;
NEH|12|19|of Joiarib, Mattenai; of Jedaiah, Uzzi;
NEH|12|20|of Sallai, Kallai; of Amok, Eber;
NEH|12|21|of Hilkiah, Hashabiah; of Jedaiah, Nethanel.
NEH|12|22|In the days of Eliashib, Joiada, Johanan, and Jaddua, the Levites were recorded as heads of fathers' houses; so too were the priests in the reign of Darius the Persian.
NEH|12|23|As for the sons of Levi, their heads of fathers' houses were written in the Book of the Chronicles until the days of Johanan the son of Eliashib.
NEH|12|24|And the chiefs of the Levites: Hashabiah, Sherebiah, and Jeshua the son of Kadmiel, with their brothers who stood opposite them, to praise and to give thanks, according to the commandment of David the man of God, watch by watch.
NEH|12|25|Mattaniah, Bakbukiah, Obadiah, Meshullam, Talmon, and Akkub were gatekeepers standing guard at the storehouses of the gates.
NEH|12|26|These were in the days of Joiakim the son of Jeshua son of Jozadak, and in the days of Nehemiah the governor and of Ezra, the priest and scribe.
NEH|12|27|And at the dedication of the wall of Jerusalem they sought the Levites in all their places, to bring them to Jerusalem to celebrate the dedication with gladness, with thanksgivings and with singing, with cymbals, harps, and lyres.
NEH|12|28|And the sons of the singers gathered together from the district surrounding Jerusalem and from the villages of the Netophathites;
NEH|12|29|also from Beth-gilgal and from the region of Geba and Azmaveth, for the singers had built for themselves villages around Jerusalem.
NEH|12|30|And the priests and the Levites purified themselves, and they purified the people and the gates and the wall.
NEH|12|31|Then I brought the leaders of Judah up onto the wall and appointed two great choirs that gave thanks. One went to the south on the wall to the Dung Gate.
NEH|12|32|And after them went Hoshaiah and half of the leaders of Judah,
NEH|12|33|and Azariah, Ezra, Meshullam,
NEH|12|34|Judah, Benjamin, Shemaiah, and Jeremiah,
NEH|12|35|and certain of the priests' sons with trumpets: Zechariah the son of Jonathan, son of Shemaiah, son of Mattaniah, son of Micaiah, son of Zaccur, son of Asaph;
NEH|12|36|and his relatives, Shemaiah, Azarel, Milalai, Gilalai, Maai, Nethanel, Judah, and Hanani, with the musical instruments of David the man of God. And Ezra the scribe went before them.
NEH|12|37|At the Fountain Gate they went up straight before them by the stairs of the city of David, at the ascent of the wall, above the house of David, to the Water Gate on the east.
NEH|12|38|The other choir of those who gave thanks went to the north, and I followed them with half of the people, on the wall, above the Tower of the Ovens, to the Broad Wall,
NEH|12|39|and above the Gate of Ephraim, and by the Gate of Yeshanah, and by the Fish Gate and the Tower of Hananel and the Tower of the Hundred, to the Sheep Gate; and they came to a halt at the Gate of the Guard.
NEH|12|40|So both choirs of those who gave thanks stood in the house of God, and I and half of the officials with me;
NEH|12|41|and the priests Eliakim, Maaseiah, Miniamin, Micaiah, Elioenai, Zechariah, and Hananiah, with trumpets;
NEH|12|42|and Maaseiah, Shemaiah, Eleazar, Uzzi, Jehohanan, Malchijah, Elam, and Ezer. And the singers sang with Jezrahiah as their leader.
NEH|12|43|And they offered great sacrifices that day and rejoiced, for God had made them rejoice with great joy; the women and children also rejoiced. And the joy of Jerusalem was heard far away.
NEH|12|44|On that day men were appointed over the storerooms, the contributions, the firstfruits, and the tithes, to gather into them the portions required by the Law for the priests and for the Levites according to the fields of the towns, for Judah rejoiced over the priests and the Levites who ministered.
NEH|12|45|And they performed the service of their God and the service of purification, as did the singers and the gatekeepers, according to the command of David and his son Solomon.
NEH|12|46|For long ago in the days of David and Asaph there were directors of the singers, and there were songs of praise and thanksgiving to God.
NEH|12|47|And all Israel in the days of Zerubbabel and in the days of Nehemiah gave the daily portions for the singers and the gatekeepers; and they set apart that which was for the Levites; and the Levites set apart that which was for the sons of Aaron.
NEH|13|1|On that day they read from the Book of Moses in the hearing of the people. And in it was found written that no Ammonite or Moabite should ever enter the assembly of God,
NEH|13|2|for they did not meet the people of Israel with bread and water, but hired Balaam against them to curse them- yet our God turned the curse into a blessing.
NEH|13|3|As soon as the people heard the law, they separated from Israel all those of foreign descent.
NEH|13|4|Now before this, Eliashib the priest, who was appointed over the chambers of the house of our God, and who was related to Tobiah,
NEH|13|5|prepared for Tobiah a large chamber where they had previously put the grain offering, the frankincense, the vessels, and the tithes of grain, wine, and oil, which were given by commandment to the Levites, singers, and gatekeepers, and the contributions for the priests.
NEH|13|6|While this was taking place, I was not in Jerusalem, for in the thirty-second year of Artaxerxes king of Babylon I went to the king. And after some time I asked leave of the king
NEH|13|7|and came to Jerusalem, and I then discovered the evil that Eliashib had done for Tobiah, preparing for him a chamber in the courts of the house of God.
NEH|13|8|And I was very angry, and I threw all the household furniture of Tobiah out of the chamber.
NEH|13|9|Then I gave orders, and they cleansed the chambers, and I brought back there the vessels of the house of God, with the grain offering and the frankincense.
NEH|13|10|I also found out that the portions of the Levites had not been given to them, so that the Levites and the singers, who did the work, had fled each to his field.
NEH|13|11|So I confronted the officials and said, "Why is the house of God forsaken?" And I gathered them together and set them in their stations.
NEH|13|12|Then all Judah brought the tithe of the grain, wine, and oil into the storehouses.
NEH|13|13|And I appointed as treasurers over the storehouses Shelemiah the priest, Zadok the scribe, and Pedaiah of the Levites, and as their assistant Hanan the son of Zaccur, son of Mattaniah, for they were considered reliable, and their duty was to distribute to their brothers.
NEH|13|14|Remember me, O my God, concerning this, and do not wipe out my good deeds that I have done for the house of my God and for his service.
NEH|13|15|In those days I saw in Judah people treading winepresses on the Sabbath, and bringing in heaps of grain and loading them on donkeys, and also wine, grapes, figs, and all kinds of loads, which they brought into Jerusalem on the Sabbath day. And I warned them on the day when they sold food.
NEH|13|16|Tyrians also, who lived in the city, brought in fish and all kinds of goods and sold them on the Sabbath to the people of Judah, in Jerusalem itself!
NEH|13|17|Then I confronted the nobles of Judah and said to them, "What is this evil thing that you are doing, profaning the Sabbath day?
NEH|13|18|Did not your fathers act in this way, and did not our God bring all this disaster on us and on this city? Now you are bringing more wrath on Israel by profaning the Sabbath."
NEH|13|19|As soon as it began to grow dark at the gates of Jerusalem before the Sabbath, I commanded that the doors should be shut and gave orders that they should not be opened until after the Sabbath. And I stationed some of my servants at the gates, that no load might be brought in on the Sabbath day.
NEH|13|20|Then the merchants and sellers of all kinds of wares lodged outside Jerusalem once or twice.
NEH|13|21|But I warned them and said to them, "Why do you lodge outside the wall? If you do so again, I will lay hands on you." From that time on they did not come on the Sabbath.
NEH|13|22|Then I commanded the Levites that they should purify themselves and come and guard the gates, to keep the Sabbath day holy. Remember this also in my favor, O my God, and spare me according to the greatness of your steadfast love.
NEH|13|23|In those days also I saw the Jews who had married women of Ashdod, Ammon, and Moab.
NEH|13|24|And half of their children spoke the language of Ashdod, and they could not speak the language of Judah, but the language of each people.
NEH|13|25|And I confronted them and cursed them and beat some of them and pulled out their hair. And I made them take oath in the name of God, saying, "You shall not give your daughters to their sons, or take their daughters for your sons or for yourselves.
NEH|13|26|Did not Solomon king of Israel sin on account of such women? Among the many nations there was no king like him, and he was beloved by his God, and God made him king over all Israel. Nevertheless, foreign women made even him to sin.
NEH|13|27|Shall we then listen to you and do all this great evil and act treacherously against our God by marrying foreign women?"
NEH|13|28|And one of the sons of Jehoiada, the son of Eliashib the high priest, was the son-in-law of Sanballat the Horonite. Therefore I chased him from me.
NEH|13|29|Remember them, O my God, because they have desecrated the priesthood and the covenant of the priesthood and the Levites.
NEH|13|30|Thus I cleansed them from everything foreign, and I established the duties of the priests and Levites, each in his work;
NEH|13|31|and I provided for the wood offering at appointed times, and for the firstfruits. Remember me, O my God, for good.
