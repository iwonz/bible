JOSH|1|1|After the death of Moses the servant of the LORD, the LORD said to Joshua son of Nun, Moses' aide:
JOSH|1|2|"Moses my servant is dead. Now then, you and all these people, get ready to cross the Jordan River into the land I am about to give to them-to the Israelites.
JOSH|1|3|I will give you every place where you set your foot, as I promised Moses.
JOSH|1|4|Your territory will extend from the desert to Lebanon, and from the great river, the Euphrates-all the Hittite country-to the Great Sea on the west.
JOSH|1|5|No one will be able to stand up against you all the days of your life. As I was with Moses, so I will be with you; I will never leave you nor forsake you.
JOSH|1|6|"Be strong and courageous, because you will lead these people to inherit the land I swore to their forefathers to give them.
JOSH|1|7|Be strong and very courageous. Be careful to obey all the law my servant Moses gave you; do not turn from it to the right or to the left, that you may be successful wherever you go.
JOSH|1|8|Do not let this Book of the Law depart from your mouth; meditate on it day and night, so that you may be careful to do everything written in it. Then you will be prosperous and successful.
JOSH|1|9|Have I not commanded you? Be strong and courageous. Do not be terrified; do not be discouraged, for the LORD your God will be with you wherever you go."
JOSH|1|10|So Joshua ordered the officers of the people:
JOSH|1|11|"Go through the camp and tell the people, 'Get your supplies ready. Three days from now you will cross the Jordan here to go in and take possession of the land the LORD your God is giving you for your own.'"
JOSH|1|12|But to the Reubenites, the Gadites and the half-tribe of Manasseh, Joshua said,
JOSH|1|13|"Remember the command that Moses the servant of the LORD gave you: 'The LORD your God is giving you rest and has granted you this land.'
JOSH|1|14|Your wives, your children and your livestock may stay in the land that Moses gave you east of the Jordan, but all your fighting men, fully armed, must cross over ahead of your brothers. You are to help your brothers
JOSH|1|15|until the LORD gives them rest, as he has done for you, and until they too have taken possession of the land that the LORD your God is giving them. After that, you may go back and occupy your own land, which Moses the servant of the LORD gave you east of the Jordan toward the sunrise."
JOSH|1|16|Then they answered Joshua, "Whatever you have commanded us we will do, and wherever you send us we will go.
JOSH|1|17|Just as we fully obeyed Moses, so we will obey you. Only may the LORD your God be with you as he was with Moses.
JOSH|1|18|Whoever rebels against your word and does not obey your words, whatever you may command them, will be put to death. Only be strong and courageous!"
JOSH|2|1|Then Joshua son of Nun secretly sent two spies from Shittim. "Go, look over the land," he said, "especially Jericho." So they went and entered the house of a prostitute named Rahab and stayed there.
JOSH|2|2|The king of Jericho was told, "Look! Some of the Israelites have come here tonight to spy out the land."
JOSH|2|3|So the king of Jericho sent this message to Rahab: "Bring out the men who came to you and entered your house, because they have come to spy out the whole land."
JOSH|2|4|But the woman had taken the two men and hidden them. She said, "Yes, the men came to me, but I did not know where they had come from.
JOSH|2|5|At dusk, when it was time to close the city gate, the men left. I don't know which way they went. Go after them quickly. You may catch up with them."
JOSH|2|6|(But she had taken them up to the roof and hidden them under the stalks of flax she had laid out on the roof.)
JOSH|2|7|So the men set out in pursuit of the spies on the road that leads to the fords of the Jordan, and as soon as the pursuers had gone out, the gate was shut.
JOSH|2|8|Before the spies lay down for the night, she went up on the roof
JOSH|2|9|and said to them, "I know that the LORD has given this land to you and that a great fear of you has fallen on us, so that all who live in this country are melting in fear because of you.
JOSH|2|10|We have heard how the LORD dried up the water of the Red Sea for you when you came out of Egypt, and what you did to Sihon and Og, the two kings of the Amorites east of the Jordan, whom you completely destroyed.
JOSH|2|11|When we heard of it, our hearts melted and everyone's courage failed because of you, for the LORD your God is God in heaven above and on the earth below.
JOSH|2|12|Now then, please swear to me by the LORD that you will show kindness to my family, because I have shown kindness to you. Give me a sure sign
JOSH|2|13|that you will spare the lives of my father and mother, my brothers and sisters, and all who belong to them, and that you will save us from death."
JOSH|2|14|"Our lives for your lives!" the men assured her. "If you don't tell what we are doing, we will treat you kindly and faithfully when the LORD gives us the land."
JOSH|2|15|So she let them down by a rope through the window, for the house she lived in was part of the city wall.
JOSH|2|16|Now she had said to them, "Go to the hills so the pursuers will not find you. Hide yourselves there three days until they return, and then go on your way."
JOSH|2|17|The men said to her, "This oath you made us swear will not be binding on us
JOSH|2|18|unless, when we enter the land, you have tied this scarlet cord in the window through which you let us down, and unless you have brought your father and mother, your brothers and all your family into your house.
JOSH|2|19|If anyone goes outside your house into the street, his blood will be on his own head; we will not be responsible. As for anyone who is in the house with you, his blood will be on our head if a hand is laid on him.
JOSH|2|20|But if you tell what we are doing, we will be released from the oath you made us swear."
JOSH|2|21|"Agreed," she replied. "Let it be as you say." So she sent them away and they departed. And she tied the scarlet cord in the window.
JOSH|2|22|When they left, they went into the hills and stayed there three days, until the pursuers had searched all along the road and returned without finding them.
JOSH|2|23|Then the two men started back. They went down out of the hills, forded the river and came to Joshua son of Nun and told him everything that had happened to them.
JOSH|2|24|They said to Joshua, "The LORD has surely given the whole land into our hands; all the people are melting in fear because of us."
JOSH|3|1|Early in the morning Joshua and all the Israelites set out from Shittim and went to the Jordan, where they camped before crossing over.
JOSH|3|2|After three days the officers went throughout the camp,
JOSH|3|3|giving orders to the people: "When you see the ark of the covenant of the LORD your God, and the priests, who are Levites, carrying it, you are to move out from your positions and follow it.
JOSH|3|4|Then you will know which way to go, since you have never been this way before. But keep a distance of about a thousand yards between you and the ark; do not go near it."
JOSH|3|5|Joshua told the people, "Consecrate yourselves, for tomorrow the LORD will do amazing things among you."
JOSH|3|6|Joshua said to the priests, "Take up the ark of the covenant and pass on ahead of the people." So they took it up and went ahead of them.
JOSH|3|7|And the LORD said to Joshua, "Today I will begin to exalt you in the eyes of all Israel, so they may know that I am with you as I was with Moses.
JOSH|3|8|Tell the priests who carry the ark of the covenant: 'When you reach the edge of the Jordan's waters, go and stand in the river.'"
JOSH|3|9|Joshua said to the Israelites, "Come here and listen to the words of the LORD your God.
JOSH|3|10|This is how you will know that the living God is among you and that he will certainly drive out before you the Canaanites, Hittites, Hivites, Perizzites, Girgashites, Amorites and Jebusites.
JOSH|3|11|See, the ark of the covenant of the Lord of all the earth will go into the Jordan ahead of you.
JOSH|3|12|Now then, choose twelve men from the tribes of Israel, one from each tribe.
JOSH|3|13|And as soon as the priests who carry the ark of the LORD -the Lord of all the earth-set foot in the Jordan, its waters flowing downstream will be cut off and stand up in a heap."
JOSH|3|14|So when the people broke camp to cross the Jordan, the priests carrying the ark of the covenant went ahead of them.
JOSH|3|15|Now the Jordan is at flood stage all during harvest. Yet as soon as the priests who carried the ark reached the Jordan and their feet touched the water's edge,
JOSH|3|16|the water from upstream stopped flowing. It piled up in a heap a great distance away, at a town called Adam in the vicinity of Zarethan, while the water flowing down to the Sea of the Arabah (the Salt Sea ) was completely cut off. So the people crossed over opposite Jericho.
JOSH|3|17|The priests who carried the ark of the covenant of the LORD stood firm on dry ground in the middle of the Jordan, while all Israel passed by until the whole nation had completed the crossing on dry ground.
JOSH|4|1|When the whole nation had finished crossing the Jordan, the LORD said to Joshua,
JOSH|4|2|"Choose twelve men from among the people, one from each tribe,
JOSH|4|3|and tell them to take up twelve stones from the middle of the Jordan from right where the priests stood and to carry them over with you and put them down at the place where you stay tonight."
JOSH|4|4|So Joshua called together the twelve men he had appointed from the Israelites, one from each tribe,
JOSH|4|5|and said to them, "Go over before the ark of the LORD your God into the middle of the Jordan. Each of you is to take up a stone on his shoulder, according to the number of the tribes of the Israelites,
JOSH|4|6|to serve as a sign among you. In the future, when your children ask you, 'What do these stones mean?'
JOSH|4|7|tell them that the flow of the Jordan was cut off before the ark of the covenant of the LORD. When it crossed the Jordan, the waters of the Jordan were cut off. These stones are to be a memorial to the people of Israel forever."
JOSH|4|8|So the Israelites did as Joshua commanded them. They took twelve stones from the middle of the Jordan, according to the number of the tribes of the Israelites, as the LORD had told Joshua; and they carried them over with them to their camp, where they put them down.
JOSH|4|9|Joshua set up the twelve stones that had been in the middle of the Jordan at the spot where the priests who carried the ark of the covenant had stood. And they are there to this day.
JOSH|4|10|Now the priests who carried the ark remained standing in the middle of the Jordan until everything the LORD had commanded Joshua was done by the people, just as Moses had directed Joshua. The people hurried over,
JOSH|4|11|and as soon as all of them had crossed, the ark of the LORD and the priests came to the other side while the people watched.
JOSH|4|12|The men of Reuben, Gad and the half-tribe of Manasseh crossed over, armed, in front of the Israelites, as Moses had directed them.
JOSH|4|13|About forty thousand armed for battle crossed over before the LORD to the plains of Jericho for war.
JOSH|4|14|That day the LORD exalted Joshua in the sight of all Israel; and they revered him all the days of his life, just as they had revered Moses.
JOSH|4|15|Then the LORD said to Joshua,
JOSH|4|16|"Command the priests carrying the ark of the Testimony to come up out of the Jordan."
JOSH|4|17|So Joshua commanded the priests, "Come up out of the Jordan."
JOSH|4|18|And the priests came up out of the river carrying the ark of the covenant of the LORD. No sooner had they set their feet on the dry ground than the waters of the Jordan returned to their place and ran at flood stage as before.
JOSH|4|19|On the tenth day of the first month the people went up from the Jordan and camped at Gilgal on the eastern border of Jericho.
JOSH|4|20|And Joshua set up at Gilgal the twelve stones they had taken out of the Jordan.
JOSH|4|21|He said to the Israelites, "In the future when your descendants ask their fathers, 'What do these stones mean?'
JOSH|4|22|tell them, 'Israel crossed the Jordan on dry ground.'
JOSH|4|23|For the LORD your God dried up the Jordan before you until you had crossed over. The LORD your God did to the Jordan just what he had done to the Red Sea when he dried it up before us until we had crossed over.
JOSH|4|24|He did this so that all the peoples of the earth might know that the hand of the LORD is powerful and so that you might always fear the LORD your God."
JOSH|5|1|Now when all the Amorite kings west of the Jordan and all the Canaanite kings along the coast heard how the LORD had dried up the Jordan before the Israelites until we had crossed over, their hearts melted and they no longer had the courage to face the Israelites.
JOSH|5|2|At that time the LORD said to Joshua, "Make flint knives and circumcise the Israelites again."
JOSH|5|3|So Joshua made flint knives and circumcised the Israelites at Gibeath Haaraloth.
JOSH|5|4|Now this is why he did so: All those who came out of Egypt-all the men of military age-died in the desert on the way after leaving Egypt.
JOSH|5|5|All the people that came out had been circumcised, but all the people born in the desert during the journey from Egypt had not.
JOSH|5|6|The Israelites had moved about in the desert forty years until all the men who were of military age when they left Egypt had died, since they had not obeyed the LORD. For the LORD had sworn to them that they would not see the land that he had solemnly promised their fathers to give us, a land flowing with milk and honey.
JOSH|5|7|So he raised up their sons in their place, and these were the ones Joshua circumcised. They were still uncircumcised because they had not been circumcised on the way.
JOSH|5|8|And after the whole nation had been circumcised, they remained where they were in camp until they were healed.
JOSH|5|9|Then the LORD said to Joshua, "Today I have rolled away the reproach of Egypt from you." So the place has been called Gilgal to this day.
JOSH|5|10|On the evening of the fourteenth day of the month, while camped at Gilgal on the plains of Jericho, the Israelites celebrated the Passover.
JOSH|5|11|The day after the Passover, that very day, they ate some of the produce of the land: unleavened bread and roasted grain.
JOSH|5|12|The manna stopped the day after they ate this food from the land; there was no longer any manna for the Israelites, but that year they ate of the produce of Canaan.
JOSH|5|13|Now when Joshua was near Jericho, he looked up and saw a man standing in front of him with a drawn sword in his hand. Joshua went up to him and asked, "Are you for us or for our enemies?"
JOSH|5|14|"Neither," he replied, "but as commander of the army of the LORD I have now come." Then Joshua fell facedown to the ground in reverence, and asked him, "What message does my Lord have for his servant?"
JOSH|5|15|The commander of the LORD's army replied, "Take off your sandals, for the place where you are standing is holy." And Joshua did so.
JOSH|6|1|Now Jericho was tightly shut up because of the Israelites. No one went out and no one came in.
JOSH|6|2|Then the LORD said to Joshua, "See, I have delivered Jericho into your hands, along with its king and its fighting men.
JOSH|6|3|March around the city once with all the armed men. Do this for six days.
JOSH|6|4|Have seven priests carry trumpets of rams' horns in front of the ark. On the seventh day, march around the city seven times, with the priests blowing the trumpets.
JOSH|6|5|When you hear them sound a long blast on the trumpets, have all the people give a loud shout; then the wall of the city will collapse and the people will go up, every man straight in."
JOSH|6|6|So Joshua son of Nun called the priests and said to them, "Take up the ark of the covenant of the LORD and have seven priests carry trumpets in front of it."
JOSH|6|7|And he ordered the people, "Advance! March around the city, with the armed guard going ahead of the ark of the LORD."
JOSH|6|8|When Joshua had spoken to the people, the seven priests carrying the seven trumpets before the LORD went forward, blowing their trumpets, and the ark of the LORD's covenant followed them.
JOSH|6|9|The armed guard marched ahead of the priests who blew the trumpets, and the rear guard followed the ark. All this time the trumpets were sounding.
JOSH|6|10|But Joshua had commanded the people, "Do not give a war cry, do not raise your voices, do not say a word until the day I tell you to shout. Then shout!"
JOSH|6|11|So he had the ark of the LORD carried around the city, circling it once. Then the people returned to camp and spent the night there.
JOSH|6|12|Joshua got up early the next morning and the priests took up the ark of the LORD.
JOSH|6|13|The seven priests carrying the seven trumpets went forward, marching before the ark of the LORD and blowing the trumpets. The armed men went ahead of them and the rear guard followed the ark of the LORD, while the trumpets kept sounding.
JOSH|6|14|So on the second day they marched around the city once and returned to the camp. They did this for six days.
JOSH|6|15|On the seventh day, they got up at daybreak and marched around the city seven times in the same manner, except that on that day they circled the city seven times.
JOSH|6|16|The seventh time around, when the priests sounded the trumpet blast, Joshua commanded the people, "Shout! For the LORD has given you the city!
JOSH|6|17|The city and all that is in it are to be devoted to the LORD. Only Rahab the prostitute and all who are with her in her house shall be spared, because she hid the spies we sent.
JOSH|6|18|But keep away from the devoted things, so that you will not bring about your own destruction by taking any of them. Otherwise you will make the camp of Israel liable to destruction and bring trouble on it.
JOSH|6|19|All the silver and gold and the articles of bronze and iron are sacred to the LORD and must go into his treasury."
JOSH|6|20|When the trumpets sounded, the people shouted, and at the sound of the trumpet, when the people gave a loud shout, the wall collapsed; so every man charged straight in, and they took the city.
JOSH|6|21|They devoted the city to the LORD and destroyed with the sword every living thing in it-men and women, young and old, cattle, sheep and donkeys.
JOSH|6|22|Joshua said to the two men who had spied out the land, "Go into the prostitute's house and bring her out and all who belong to her, in accordance with your oath to her."
JOSH|6|23|So the young men who had done the spying went in and brought out Rahab, her father and mother and brothers and all who belonged to her. They brought out her entire family and put them in a place outside the camp of Israel.
JOSH|6|24|Then they burned the whole city and everything in it, but they put the silver and gold and the articles of bronze and iron into the treasury of the LORD's house.
JOSH|6|25|But Joshua spared Rahab the prostitute, with her family and all who belonged to her, because she hid the men Joshua had sent as spies to Jericho-and she lives among the Israelites to this day.
JOSH|6|26|At that time Joshua pronounced this solemn oath: "Cursed before the LORD is the man who undertakes to rebuild this city, Jericho: "At the cost of his firstborn son will he lay its foundations; at the cost of his youngest will he set up its gates."
JOSH|6|27|So the LORD was with Joshua, and his fame spread throughout the land.
JOSH|7|1|But the Israelites acted unfaithfully in regard to the devoted things; Achan son of Carmi, the son of Zimri, the son of Zerah, of the tribe of Judah, took some of them. So the LORD's anger burned against Israel.
JOSH|7|2|Now Joshua sent men from Jericho to Ai, which is near Beth Aven to the east of Bethel, and told them, "Go up and spy out the region." So the men went up and spied out Ai.
JOSH|7|3|When they returned to Joshua, they said, "Not all the people will have to go up against Ai. Send two or three thousand men to take it and do not weary all the people, for only a few men are there."
JOSH|7|4|So about three thousand men went up; but they were routed by the men of Ai,
JOSH|7|5|who killed about thirty-six of them. They chased the Israelites from the city gate as far as the stone quarries and struck them down on the slopes. At this the hearts of the people melted and became like water.
JOSH|7|6|Then Joshua tore his clothes and fell facedown to the ground before the ark of the LORD, remaining there till evening. The elders of Israel did the same, and sprinkled dust on their heads.
JOSH|7|7|And Joshua said, "Ah, Sovereign LORD, why did you ever bring this people across the Jordan to deliver us into the hands of the Amorites to destroy us? If only we had been content to stay on the other side of the Jordan!
JOSH|7|8|O Lord, what can I say, now that Israel has been routed by its enemies?
JOSH|7|9|The Canaanites and the other people of the country will hear about this and they will surround us and wipe out our name from the earth. What then will you do for your own great name?"
JOSH|7|10|The LORD said to Joshua, "Stand up! What are you doing down on your face?
JOSH|7|11|Israel has sinned; they have violated my covenant, which I commanded them to keep. They have taken some of the devoted things; they have stolen, they have lied, they have put them with their own possessions.
JOSH|7|12|That is why the Israelites cannot stand against their enemies; they turn their backs and run because they have been made liable to destruction. I will not be with you anymore unless you destroy whatever among you is devoted to destruction.
JOSH|7|13|"Go, consecrate the people. Tell them, 'Consecrate yourselves in preparation for tomorrow; for this is what the LORD, the God of Israel, says: That which is devoted is among you, O Israel. You cannot stand against your enemies until you remove it.
JOSH|7|14|"'In the morning, present yourselves tribe by tribe. The tribe that the LORD takes shall come forward clan by clan; the clan that the LORD takes shall come forward family by family; and the family that the LORD takes shall come forward man by man.
JOSH|7|15|He who is caught with the devoted things shall be destroyed by fire, along with all that belongs to him. He has violated the covenant of the LORD and has done a disgraceful thing in Israel!'"
JOSH|7|16|Early the next morning Joshua had Israel come forward by tribes, and Judah was taken.
JOSH|7|17|The clans of Judah came forward, and he took the Zerahites. He had the clan of the Zerahites come forward by families, and Zimri was taken.
JOSH|7|18|Joshua had his family come forward man by man, and Achan son of Carmi, the son of Zimri, the son of Zerah, of the tribe of Judah, was taken.
JOSH|7|19|Then Joshua said to Achan, "My son, give glory to the LORD, the God of Israel, and give him the praise. Tell me what you have done; do not hide it from me."
JOSH|7|20|Achan replied, "It is true! I have sinned against the LORD, the God of Israel. This is what I have done:
JOSH|7|21|When I saw in the plunder a beautiful robe from Babylonia, two hundred shekels of silver and a wedge of gold weighing fifty shekels, I coveted them and took them. They are hidden in the ground inside my tent, with the silver underneath."
JOSH|7|22|So Joshua sent messengers, and they ran to the tent, and there it was, hidden in his tent, with the silver underneath.
JOSH|7|23|They took the things from the tent, brought them to Joshua and all the Israelites and spread them out before the LORD.
JOSH|7|24|Then Joshua, together with all Israel, took Achan son of Zerah, the silver, the robe, the gold wedge, his sons and daughters, his cattle, donkeys and sheep, his tent and all that he had, to the Valley of Achor.
JOSH|7|25|Joshua said, "Why have you brought this trouble on us? The LORD will bring trouble on you today." Then all Israel stoned him, and after they had stoned the rest, they burned them.
JOSH|7|26|Over Achan they heaped up a large pile of rocks, which remains to this day. Then the LORD turned from his fierce anger. Therefore that place has been called the Valley of Achor ever since.
JOSH|8|1|Then the LORD said to Joshua, "Do not be afraid; do not be discouraged. Take the whole army with you, and go up and attack Ai. For I have delivered into your hands the king of Ai, his people, his city and his land.
JOSH|8|2|You shall do to Ai and its king as you did to Jericho and its king, except that you may carry off their plunder and livestock for yourselves. Set an ambush behind the city."
JOSH|8|3|So Joshua and the whole army moved out to attack Ai. He chose thirty thousand of his best fighting men and sent them out at night
JOSH|8|4|with these orders: "Listen carefully. You are to set an ambush behind the city. Don't go very far from it. All of you be on the alert.
JOSH|8|5|I and all those with me will advance on the city, and when the men come out against us, as they did before, we will flee from them.
JOSH|8|6|They will pursue us until we have lured them away from the city, for they will say, 'They are running away from us as they did before.' So when we flee from them,
JOSH|8|7|you are to rise up from ambush and take the city. The LORD your God will give it into your hand.
JOSH|8|8|When you have taken the city, set it on fire. Do what the LORD has commanded. See to it; you have my orders."
JOSH|8|9|Then Joshua sent them off, and they went to the place of ambush and lay in wait between Bethel and Ai, to the west of Ai-but Joshua spent that night with the people.
JOSH|8|10|Early the next morning Joshua mustered his men, and he and the leaders of Israel marched before them to Ai.
JOSH|8|11|The entire force that was with him marched up and approached the city and arrived in front of it. They set up camp north of Ai, with the valley between them and the city.
JOSH|8|12|Joshua had taken about five thousand men and set them in ambush between Bethel and Ai, to the west of the city.
JOSH|8|13|They had the soldiers take up their positions-all those in the camp to the north of the city and the ambush to the west of it. That night Joshua went into the valley.
JOSH|8|14|When the king of Ai saw this, he and all the men of the city hurried out early in the morning to meet Israel in battle at a certain place overlooking the Arabah. But he did not know that an ambush had been set against him behind the city.
JOSH|8|15|Joshua and all Israel let themselves be driven back before them, and they fled toward the desert.
JOSH|8|16|All the men of Ai were called to pursue them, and they pursued Joshua and were lured away from the city.
JOSH|8|17|Not a man remained in Ai or Bethel who did not go after Israel. They left the city open and went in pursuit of Israel.
JOSH|8|18|Then the LORD said to Joshua, "Hold out toward Ai the javelin that is in your hand, for into your hand I will deliver the city." So Joshua held out his javelin toward Ai.
JOSH|8|19|As soon as he did this, the men in the ambush rose quickly from their position and rushed forward. They entered the city and captured it and quickly set it on fire.
JOSH|8|20|The men of Ai looked back and saw the smoke of the city rising against the sky, but they had no chance to escape in any direction, for the Israelites who had been fleeing toward the desert had turned back against their pursuers.
JOSH|8|21|For when Joshua and all Israel saw that the ambush had taken the city and that smoke was going up from the city, they turned around and attacked the men of Ai.
JOSH|8|22|The men of the ambush also came out of the city against them, so that they were caught in the middle, with Israelites on both sides. Israel cut them down, leaving them neither survivors nor fugitives.
JOSH|8|23|But they took the king of Ai alive and brought him to Joshua.
JOSH|8|24|When Israel had finished killing all the men of Ai in the fields and in the desert where they had chased them, and when every one of them had been put to the sword, all the Israelites returned to Ai and killed those who were in it.
JOSH|8|25|Twelve thousand men and women fell that day-all the people of Ai.
JOSH|8|26|For Joshua did not draw back the hand that held out his javelin until he had destroyed all who lived in Ai.
JOSH|8|27|But Israel did carry off for themselves the livestock and plunder of this city, as the LORD had instructed Joshua.
JOSH|8|28|So Joshua burned Ai and made it a permanent heap of ruins, a desolate place to this day.
JOSH|8|29|He hung the king of Ai on a tree and left him there until evening. At sunset, Joshua ordered them to take his body from the tree and throw it down at the entrance of the city gate. And they raised a large pile of rocks over it, which remains to this day.
JOSH|8|30|Then Joshua built on Mount Ebal an altar to the LORD, the God of Israel,
JOSH|8|31|as Moses the servant of the LORD had commanded the Israelites. He built it according to what is written in the Book of the Law of Moses-an altar of uncut stones, on which no iron tool had been used. On it they offered to the LORD burnt offerings and sacrificed fellowship offerings.
JOSH|8|32|There, in the presence of the Israelites, Joshua copied on stones the law of Moses, which he had written.
JOSH|8|33|All Israel, aliens and citizens alike, with their elders, officials and judges, were standing on both sides of the ark of the covenant of the LORD, facing those who carried it-the priests, who were Levites. Half of the people stood in front of Mount Gerizim and half of them in front of Mount Ebal, as Moses the servant of the LORD had formerly commanded when he gave instructions to bless the people of Israel.
JOSH|8|34|Afterward, Joshua read all the words of the law-the blessings and the curses-just as it is written in the Book of the Law.
JOSH|8|35|There was not a word of all that Moses had commanded that Joshua did not read to the whole assembly of Israel, including the women and children, and the aliens who lived among them.
JOSH|9|1|Now when all the kings west of the Jordan heard about these things-those in the hill country, in the western foothills, and along the entire coast of the Great Sea as far as Lebanon (the kings of the Hittites, Amorites, Canaanites, Perizzites, Hivites and Jebusites)-
JOSH|9|2|they came together to make war against Joshua and Israel.
JOSH|9|3|However, when the people of Gibeon heard what Joshua had done to Jericho and Ai,
JOSH|9|4|they resorted to a ruse: They went as a delegation whose donkeys were loaded with worn-out sacks and old wineskins, cracked and mended.
JOSH|9|5|The men put worn and patched sandals on their feet and wore old clothes. All the bread of their food supply was dry and moldy.
JOSH|9|6|Then they went to Joshua in the camp at Gilgal and said to him and the men of Israel, "We have come from a distant country; make a treaty with us."
JOSH|9|7|The men of Israel said to the Hivites, "But perhaps you live near us. How then can we make a treaty with you?"
JOSH|9|8|"We are your servants," they said to Joshua. But Joshua asked, "Who are you and where do you come from?"
JOSH|9|9|They answered: "Your servants have come from a very distant country because of the fame of the LORD your God. For we have heard reports of him: all that he did in Egypt,
JOSH|9|10|and all that he did to the two kings of the Amorites east of the Jordan-Sihon king of Heshbon, and Og king of Bashan, who reigned in Ashtaroth.
JOSH|9|11|And our elders and all those living in our country said to us, 'Take provisions for your journey; go and meet them and say to them, "We are your servants; make a treaty with us."'
JOSH|9|12|This bread of ours was warm when we packed it at home on the day we left to come to you. But now see how dry and moldy it is.
JOSH|9|13|And these wineskins that we filled were new, but see how cracked they are. And our clothes and sandals are worn out by the very long journey."
JOSH|9|14|The men of Israel sampled their provisions but did not inquire of the LORD.
JOSH|9|15|Then Joshua made a treaty of peace with them to let them live, and the leaders of the assembly ratified it by oath.
JOSH|9|16|Three days after they made the treaty with the Gibeonites, the Israelites heard that they were neighbors, living near them.
JOSH|9|17|So the Israelites set out and on the third day came to their cities: Gibeon, Kephirah, Beeroth and Kiriath Jearim.
JOSH|9|18|But the Israelites did not attack them, because the leaders of the assembly had sworn an oath to them by the LORD, the God of Israel. The whole assembly grumbled against the leaders,
JOSH|9|19|but all the leaders answered, "We have given them our oath by the LORD, the God of Israel, and we cannot touch them now.
JOSH|9|20|This is what we will do to them: We will let them live, so that wrath will not fall on us for breaking the oath we swore to them."
JOSH|9|21|They continued, "Let them live, but let them be woodcutters and water carriers for the entire community." So the leaders' promise to them was kept.
JOSH|9|22|Then Joshua summoned the Gibeonites and said, "Why did you deceive us by saying, 'We live a long way from you,' while actually you live near us?
JOSH|9|23|You are now under a curse: You will never cease to serve as woodcutters and water carriers for the house of my God."
JOSH|9|24|They answered Joshua, "Your servants were clearly told how the LORD your God had commanded his servant Moses to give you the whole land and to wipe out all its inhabitants from before you. So we feared for our lives because of you, and that is why we did this.
JOSH|9|25|We are now in your hands. Do to us whatever seems good and right to you."
JOSH|9|26|So Joshua saved them from the Israelites, and they did not kill them.
JOSH|9|27|That day he made the Gibeonites woodcutters and water carriers for the community and for the altar of the LORD at the place the LORD would choose. And that is what they are to this day.
JOSH|10|1|Now Adoni-Zedek king of Jerusalem heard that Joshua had taken Ai and totally destroyed it, doing to Ai and its king as he had done to Jericho and its king, and that the people of Gibeon had made a treaty of peace with Israel and were living near them.
JOSH|10|2|He and his people were very much alarmed at this, because Gibeon was an important city, like one of the royal cities; it was larger than Ai, and all its men were good fighters.
JOSH|10|3|So Adoni-Zedek king of Jerusalem appealed to Hoham king of Hebron, Piram king of Jarmuth, Japhia king of Lachish and Debir king of Eglon.
JOSH|10|4|"Come up and help me attack Gibeon," he said, "because it has made peace with Joshua and the Israelites."
JOSH|10|5|Then the five kings of the Amorites-the kings of Jerusalem, Hebron, Jarmuth, Lachish and Eglon-joined forces. They moved up with all their troops and took up positions against Gibeon and attacked it.
JOSH|10|6|The Gibeonites then sent word to Joshua in the camp at Gilgal: "Do not abandon your servants. Come up to us quickly and save us! Help us, because all the Amorite kings from the hill country have joined forces against us."
JOSH|10|7|So Joshua marched up from Gilgal with his entire army, including all the best fighting men.
JOSH|10|8|The LORD said to Joshua, "Do not be afraid of them; I have given them into your hand. Not one of them will be able to withstand you."
JOSH|10|9|After an all-night march from Gilgal, Joshua took them by surprise.
JOSH|10|10|The LORD threw them into confusion before Israel, who defeated them in a great victory at Gibeon. Israel pursued them along the road going up to Beth Horon and cut them down all the way to Azekah and Makkedah.
JOSH|10|11|As they fled before Israel on the road down from Beth Horon to Azekah, the LORD hurled large hailstones down on them from the sky, and more of them died from the hailstones than were killed by the swords of the Israelites.
JOSH|10|12|On the day the LORD gave the Amorites over to Israel, Joshua said to the LORD in the presence of Israel: "O sun, stand still over Gibeon, O moon, over the Valley of Aijalon."
JOSH|10|13|So the sun stood still, and the moon stopped, till the nation avenged itself on its enemies, as it is written in the Book of Jashar. The sun stopped in the middle of the sky and delayed going down about a full day.
JOSH|10|14|There has never been a day like it before or since, a day when the LORD listened to a man. Surely the LORD was fighting for Israel!
JOSH|10|15|Then Joshua returned with all Israel to the camp at Gilgal.
JOSH|10|16|Now the five kings had fled and hidden in the cave at Makkedah.
JOSH|10|17|When Joshua was told that the five kings had been found hiding in the cave at Makkedah,
JOSH|10|18|he said, "Roll large rocks up to the mouth of the cave, and post some men there to guard it.
JOSH|10|19|But don't stop! Pursue your enemies, attack them from the rear and don't let them reach their cities, for the LORD your God has given them into your hand."
JOSH|10|20|So Joshua and the Israelites destroyed them completely-almost to a man-but the few who were left reached their fortified cities.
JOSH|10|21|The whole army then returned safely to Joshua in the camp at Makkedah, and no one uttered a word against the Israelites.
JOSH|10|22|Joshua said, "Open the mouth of the cave and bring those five kings out to me."
JOSH|10|23|So they brought the five kings out of the cave-the kings of Jerusalem, Hebron, Jarmuth, Lachish and Eglon.
JOSH|10|24|When they had brought these kings to Joshua, he summoned all the men of Israel and said to the army commanders who had come with him, "Come here and put your feet on the necks of these kings." So they came forward and placed their feet on their necks.
JOSH|10|25|Joshua said to them, "Do not be afraid; do not be discouraged. Be strong and courageous. This is what the LORD will do to all the enemies you are going to fight."
JOSH|10|26|Then Joshua struck and killed the kings and hung them on five trees, and they were left hanging on the trees until evening.
JOSH|10|27|At sunset Joshua gave the order and they took them down from the trees and threw them into the cave where they had been hiding. At the mouth of the cave they placed large rocks, which are there to this day.
JOSH|10|28|That day Joshua took Makkedah. He put the city and its king to the sword and totally destroyed everyone in it. He left no survivors. And he did to the king of Makkedah as he had done to the king of Jericho.
JOSH|10|29|Then Joshua and all Israel with him moved on from Makkedah to Libnah and attacked it.
JOSH|10|30|The LORD also gave that city and its king into Israel's hand. The city and everyone in it Joshua put to the sword. He left no survivors there. And he did to its king as he had done to the king of Jericho.
JOSH|10|31|Then Joshua and all Israel with him moved on from Libnah to Lachish; he took up positions against it and attacked it.
JOSH|10|32|The LORD handed Lachish over to Israel, and Joshua took it on the second day. The city and everyone in it he put to the sword, just as he had done to Libnah.
JOSH|10|33|Meanwhile, Horam king of Gezer had come up to help Lachish, but Joshua defeated him and his army-until no survivors were left.
JOSH|10|34|Then Joshua and all Israel with him moved on from Lachish to Eglon; they took up positions against it and attacked it.
JOSH|10|35|They captured it that same day and put it to the sword and totally destroyed everyone in it, just as they had done to Lachish.
JOSH|10|36|Then Joshua and all Israel with him went up from Eglon to Hebron and attacked it.
JOSH|10|37|They took the city and put it to the sword, together with its king, its villages and everyone in it. They left no survivors. Just as at Eglon, they totally destroyed it and everyone in it.
JOSH|10|38|Then Joshua and all Israel with him turned around and attacked Debir.
JOSH|10|39|They took the city, its king and its villages, and put them to the sword. Everyone in it they totally destroyed. They left no survivors. They did to Debir and its king as they had done to Libnah and its king and to Hebron.
JOSH|10|40|So Joshua subdued the whole region, including the hill country, the Negev, the western foothills and the mountain slopes, together with all their kings. He left no survivors. He totally destroyed all who breathed, just as the LORD, the God of Israel, had commanded.
JOSH|10|41|Joshua subdued them from Kadesh Barnea to Gaza and from the whole region of Goshen to Gibeon.
JOSH|10|42|All these kings and their lands Joshua conquered in one campaign, because the LORD, the God of Israel, fought for Israel.
JOSH|10|43|Then Joshua returned with all Israel to the camp at Gilgal.
JOSH|11|1|When Jabin king of Hazor heard of this, he sent word to Jobab king of Madon, to the kings of Shimron and Acshaph,
JOSH|11|2|and to the northern kings who were in the mountains, in the Arabah south of Kinnereth, in the western foothills and in Naphoth Dor on the west;
JOSH|11|3|to the Canaanites in the east and west; to the Amorites, Hittites, Perizzites and Jebusites in the hill country; and to the Hivites below Hermon in the region of Mizpah.
JOSH|11|4|They came out with all their troops and a large number of horses and chariots-a huge army, as numerous as the sand on the seashore.
JOSH|11|5|All these kings joined forces and made camp together at the Waters of Merom, to fight against Israel.
JOSH|11|6|The LORD said to Joshua, "Do not be afraid of them, because by this time tomorrow I will hand all of them over to Israel, slain. You are to hamstring their horses and burn their chariots."
JOSH|11|7|So Joshua and his whole army came against them suddenly at the Waters of Merom and attacked them,
JOSH|11|8|and the LORD gave them into the hand of Israel. They defeated them and pursued them all the way to Greater Sidon, to Misrephoth Maim, and to the Valley of Mizpah on the east, until no survivors were left.
JOSH|11|9|Joshua did to them as the LORD had directed: He hamstrung their horses and burned their chariots.
JOSH|11|10|At that time Joshua turned back and captured Hazor and put its king to the sword. (Hazor had been the head of all these kingdoms.)
JOSH|11|11|Everyone in it they put to the sword. They totally destroyed them, not sparing anything that breathed, and he burned up Hazor itself.
JOSH|11|12|Joshua took all these royal cities and their kings and put them to the sword. He totally destroyed them, as Moses the servant of the LORD had commanded.
JOSH|11|13|Yet Israel did not burn any of the cities built on their mounds-except Hazor, which Joshua burned.
JOSH|11|14|The Israelites carried off for themselves all the plunder and livestock of these cities, but all the people they put to the sword until they completely destroyed them, not sparing anyone that breathed.
JOSH|11|15|As the LORD commanded his servant Moses, so Moses commanded Joshua, and Joshua did it; he left nothing undone of all that the LORD commanded Moses.
JOSH|11|16|So Joshua took this entire land: the hill country, all the Negev, the whole region of Goshen, the western foothills, the Arabah and the mountains of Israel with their foothills,
JOSH|11|17|from Mount Halak, which rises toward Seir, to Baal Gad in the Valley of Lebanon below Mount Hermon. He captured all their kings and struck them down, putting them to death.
JOSH|11|18|Joshua waged war against all these kings for a long time.
JOSH|11|19|Except for the Hivites living in Gibeon, not one city made a treaty of peace with the Israelites, who took them all in battle.
JOSH|11|20|For it was the LORD himself who hardened their hearts to wage war against Israel, so that he might destroy them totally, exterminating them without mercy, as the LORD had commanded Moses.
JOSH|11|21|At that time Joshua went and destroyed the Anakites from the hill country: from Hebron, Debir and Anab, from all the hill country of Judah, and from all the hill country of Israel. Joshua totally destroyed them and their towns.
JOSH|11|22|No Anakites were left in Israelite territory; only in Gaza, Gath and Ashdod did any survive.
JOSH|11|23|So Joshua took the entire land, just as the LORD had directed Moses, and he gave it as an inheritance to Israel according to their tribal divisions. Then the land had rest from war.
JOSH|12|1|These are the kings of the land whom the Israelites had defeated and whose territory they took over east of the Jordan, from the Arnon Gorge to Mount Hermon, including all the eastern side of the Arabah:
JOSH|12|2|Sihon king of the Amorites, who reigned in Heshbon. He ruled from Aroer on the rim of the Arnon Gorge-from the middle of the gorge-to the Jabbok River, which is the border of the Ammonites. This included half of Gilead.
JOSH|12|3|He also ruled over the eastern Arabah from the Sea of Kinnereth to the Sea of the Arabah (the Salt Sea ), to Beth Jeshimoth, and then southward below the slopes of Pisgah.
JOSH|12|4|And the territory of Og king of Bashan, one of the last of the Rephaites, who reigned in Ashtaroth and Edrei.
JOSH|12|5|He ruled over Mount Hermon, Salecah, all of Bashan to the border of the people of Geshur and Maacah, and half of Gilead to the border of Sihon king of Heshbon.
JOSH|12|6|Moses, the servant of the LORD, and the Israelites conquered them. And Moses the servant of the LORD gave their land to the Reubenites, the Gadites and the half-tribe of Manasseh to be their possession.
JOSH|12|7|These are the kings of the land that Joshua and the Israelites conquered on the west side of the Jordan, from Baal Gad in the Valley of Lebanon to Mount Halak, which rises toward Seir (their lands Joshua gave as an inheritance to the tribes of Israel according to their tribal divisions-
JOSH|12|8|the hill country, the western foothills, the Arabah, the mountain slopes, the desert and the Negev-the lands of the Hittites, Amorites, Canaanites, Perizzites, Hivites and Jebusites):
JOSH|12|9|the king of Jericho one the king of Ai (near Bethel) one
JOSH|12|10|the king of Jerusalem one the king of Hebron one
JOSH|12|11|the king of Jarmuth one the king of Lachish one
JOSH|12|12|the king of Eglon one the king of Gezer one
JOSH|12|13|the king of Debir one the king of Geder one
JOSH|12|14|the king of Hormah one the king of Arad one
JOSH|12|15|the king of Libnah one the king of Adullam one
JOSH|12|16|the king of Makkedah one the king of Bethel one
JOSH|12|17|the king of Tappuah one the king of Hepher one
JOSH|12|18|the king of Aphek one the king of Lasharon one
JOSH|12|19|the king of Madon one the king of Hazor one
JOSH|12|20|the king of Shimron Meron one the king of Acshaph one
JOSH|12|21|the king of Taanach one the king of Megiddo one
JOSH|12|22|the king of Kedesh one the king of Jokneam in Carmel one
JOSH|12|23|the king of Dor (in Naphoth Dor ) one the king of Goyim in Gilgal one
JOSH|12|24|the king of Tirzah one thirty-one kings in all.
JOSH|13|1|When Joshua was old and well advanced in years, the LORD said to him, "You are very old, and there are still very large areas of land to be taken over.
JOSH|13|2|"This is the land that remains: all the regions of the Philistines and Geshurites:
JOSH|13|3|from the Shihor River on the east of Egypt to the territory of Ekron on the north, all of it counted as Canaanite (the territory of the five Philistine rulers in Gaza, Ashdod, Ashkelon, Gath and Ekron-that of the Avvites);
JOSH|13|4|from the south, all the land of the Canaanites, from Arah of the Sidonians as far as Aphek, the region of the Amorites,
JOSH|13|5|the area of the Gebalites; and all Lebanon to the east, from Baal Gad below Mount Hermon to Lebo Hamath.
JOSH|13|6|"As for all the inhabitants of the mountain regions from Lebanon to Misrephoth Maim, that is, all the Sidonians, I myself will drive them out before the Israelites. Be sure to allocate this land to Israel for an inheritance, as I have instructed you,
JOSH|13|7|and divide it as an inheritance among the nine tribes and half of the tribe of Manasseh."
JOSH|13|8|The other half of Manasseh, the Reubenites and the Gadites had received the inheritance that Moses had given them east of the Jordan, as he, the servant of the LORD, had assigned it to them.
JOSH|13|9|It extended from Aroer on the rim of the Arnon Gorge, and from the town in the middle of the gorge, and included the whole plateau of Medeba as far as Dibon,
JOSH|13|10|and all the towns of Sihon king of the Amorites, who ruled in Heshbon, out to the border of the Ammonites.
JOSH|13|11|It also included Gilead, the territory of the people of Geshur and Maacah, all of Mount Hermon and all Bashan as far as Salecah-
JOSH|13|12|that is, the whole kingdom of Og in Bashan, who had reigned in Ashtaroth and Edrei and had survived as one of the last of the Rephaites. Moses had defeated them and taken over their land.
JOSH|13|13|But the Israelites did not drive out the people of Geshur and Maacah, so they continue to live among the Israelites to this day.
JOSH|13|14|But to the tribe of Levi he gave no inheritance, since the offerings made by fire to the LORD, the God of Israel, are their inheritance, as he promised them.
JOSH|13|15|This is what Moses had given to the tribe of Reuben, clan by clan:
JOSH|13|16|The territory from Aroer on the rim of the Arnon Gorge, and from the town in the middle of the gorge, and the whole plateau past Medeba
JOSH|13|17|to Heshbon and all its towns on the plateau, including Dibon, Bamoth Baal, Beth Baal Meon,
JOSH|13|18|Jahaz, Kedemoth, Mephaath,
JOSH|13|19|Kiriathaim, Sibmah, Zereth Shahar on the hill in the valley,
JOSH|13|20|Beth Peor, the slopes of Pisgah, and Beth Jeshimoth
JOSH|13|21|-all the towns on the plateau and the entire realm of Sihon king of the Amorites, who ruled at Heshbon. Moses had defeated him and the Midianite chiefs, Evi, Rekem, Zur, Hur and Reba-princes allied with Sihon-who lived in that country.
JOSH|13|22|In addition to those slain in battle, the Israelites had put to the sword Balaam son of Beor, who practiced divination.
JOSH|13|23|The boundary of the Reubenites was the bank of the Jordan. These towns and their villages were the inheritance of the Reubenites, clan by clan.
JOSH|13|24|This is what Moses had given to the tribe of Gad, clan by clan:
JOSH|13|25|The territory of Jazer, all the towns of Gilead and half the Ammonite country as far as Aroer, near Rabbah;
JOSH|13|26|and from Heshbon to Ramath Mizpah and Betonim, and from Mahanaim to the territory of Debir;
JOSH|13|27|and in the valley, Beth Haram, Beth Nimrah, Succoth and Zaphon with the rest of the realm of Sihon king of Heshbon (the east side of the Jordan, the territory up to the end of the Sea of Kinnereth ).
JOSH|13|28|These towns and their villages were the inheritance of the Gadites, clan by clan.
JOSH|13|29|This is what Moses had given to the half-tribe of Manasseh, that is, to half the family of the descendants of Manasseh, clan by clan:
JOSH|13|30|The territory extending from Mahanaim and including all of Bashan, the entire realm of Og king of Bashan-all the settlements of Jair in Bashan, sixty towns,
JOSH|13|31|half of Gilead, and Ashtaroth and Edrei (the royal cities of Og in Bashan). This was for the descendants of Makir son of Manasseh-for half of the sons of Makir, clan by clan.
JOSH|13|32|This is the inheritance Moses had given when he was in the plains of Moab across the Jordan east of Jericho.
JOSH|13|33|But to the tribe of Levi, Moses had given no inheritance; the LORD, the God of Israel, is their inheritance, as he promised them.
JOSH|14|1|Now these are the areas the Israelites received as an inheritance in the land of Canaan, which Eleazar the priest, Joshua son of Nun and the heads of the tribal clans of Israel allotted to them.
JOSH|14|2|Their inheritances were assigned by lot to the nine-and-a-half tribes, as the LORD had commanded through Moses.
JOSH|14|3|Moses had granted the two-and-a-half tribes their inheritance east of the Jordan but had not granted the Levites an inheritance among the rest,
JOSH|14|4|for the sons of Joseph had become two tribes-Manasseh and Ephraim. The Levites received no share of the land but only towns to live in, with pasturelands for their flocks and herds.
JOSH|14|5|So the Israelites divided the land, just as the LORD had commanded Moses.
JOSH|14|6|Now the men of Judah approached Joshua at Gilgal, and Caleb son of Jephunneh the Kenizzite said to him, "You know what the LORD said to Moses the man of God at Kadesh Barnea about you and me.
JOSH|14|7|I was forty years old when Moses the servant of the LORD sent me from Kadesh Barnea to explore the land. And I brought him back a report according to my convictions,
JOSH|14|8|but my brothers who went up with me made the hearts of the people melt with fear. I, however, followed the LORD my God wholeheartedly.
JOSH|14|9|So on that day Moses swore to me, 'The land on which your feet have walked will be your inheritance and that of your children forever, because you have followed the LORD my God wholeheartedly.'
JOSH|14|10|"Now then, just as the LORD promised, he has kept me alive for forty-five years since the time he said this to Moses, while Israel moved about in the desert. So here I am today, eighty-five years old!
JOSH|14|11|I am still as strong today as the day Moses sent me out; I'm just as vigorous to go out to battle now as I was then.
JOSH|14|12|Now give me this hill country that the LORD promised me that day. You yourself heard then that the Anakites were there and their cities were large and fortified, but, the LORD helping me, I will drive them out just as he said."
JOSH|14|13|Then Joshua blessed Caleb son of Jephunneh and gave him Hebron as his inheritance.
JOSH|14|14|So Hebron has belonged to Caleb son of Jephunneh the Kenizzite ever since, because he followed the LORD, the God of Israel, wholeheartedly.
JOSH|14|15|(Hebron used to be called Kiriath Arba after Arba, who was the greatest man among the Anakites.) Then the land had rest from war.
JOSH|15|1|The allotment for the tribe of Judah, clan by clan, extended down to the territory of Edom, to the Desert of Zin in the extreme south.
JOSH|15|2|Their southern boundary started from the bay at the southern end of the Salt Sea,
JOSH|15|3|crossed south of Scorpion Pass, continued on to Zin and went over to the south of Kadesh Barnea. Then it ran past Hezron up to Addar and curved around to Karka.
JOSH|15|4|It then passed along to Azmon and joined the Wadi of Egypt, ending at the sea. This is their southern boundary.
JOSH|15|5|The eastern boundary is the Salt Sea as far as the mouth of the Jordan. The northern boundary started from the bay of the sea at the mouth of the Jordan,
JOSH|15|6|went up to Beth Hoglah and continued north of Beth Arabah to the Stone of Bohan son of Reuben.
JOSH|15|7|The boundary then went up to Debir from the Valley of Achor and turned north to Gilgal, which faces the Pass of Adummim south of the gorge. It continued along to the waters of En Shemesh and came out at En Rogel.
JOSH|15|8|Then it ran up the Valley of Ben Hinnom along the southern slope of the Jebusite city (that is, Jerusalem). From there it climbed to the top of the hill west of the Hinnom Valley at the northern end of the Valley of Rephaim.
JOSH|15|9|From the hilltop the boundary headed toward the spring of the waters of Nephtoah, came out at the towns of Mount Ephron and went down toward Baalah (that is, Kiriath Jearim).
JOSH|15|10|Then it curved westward from Baalah to Mount Seir, ran along the northern slope of Mount Jearim (that is, Kesalon), continued down to Beth Shemesh and crossed to Timnah.
JOSH|15|11|It went to the northern slope of Ekron, turned toward Shikkeron, passed along to Mount Baalah and reached Jabneel. The boundary ended at the sea.
JOSH|15|12|The western boundary is the coastline of the Great Sea. These are the boundaries around the people of Judah by their clans.
JOSH|15|13|In accordance with the LORD's command to him, Joshua gave to Caleb son of Jephunneh a portion in Judah-Kiriath Arba, that is, Hebron. (Arba was the forefather of Anak.)
JOSH|15|14|From Hebron Caleb drove out the three Anakites-Sheshai, Ahiman and Talmai-descendants of Anak.
JOSH|15|15|From there he marched against the people living in Debir (formerly called Kiriath Sepher).
JOSH|15|16|And Caleb said, "I will give my daughter Acsah in marriage to the man who attacks and captures Kiriath Sepher."
JOSH|15|17|Othniel son of Kenaz, Caleb's brother, took it; so Caleb gave his daughter Acsah to him in marriage.
JOSH|15|18|One day when she came to Othniel, she urged him to ask her father for a field. When she got off her donkey, Caleb asked her, "What can I do for you?"
JOSH|15|19|She replied, "Do me a special favor. Since you have given me land in the Negev, give me also springs of water." So Caleb gave her the upper and lower springs.
JOSH|15|20|This is the inheritance of the tribe of Judah, clan by clan:
JOSH|15|21|The southernmost towns of the tribe of Judah in the Negev toward the boundary of Edom were: Kabzeel, Eder, Jagur,
JOSH|15|22|Kinah, Dimonah, Adadah,
JOSH|15|23|Kedesh, Hazor, Ithnan,
JOSH|15|24|Ziph, Telem, Bealoth,
JOSH|15|25|Hazor Hadattah, Kerioth Hezron (that is, Hazor),
JOSH|15|26|Amam, Shema, Moladah,
JOSH|15|27|Hazar Gaddah, Heshmon, Beth Pelet,
JOSH|15|28|Hazar Shual, Beersheba, Biziothiah,
JOSH|15|29|Baalah, Iim, Ezem,
JOSH|15|30|Eltolad, Kesil, Hormah,
JOSH|15|31|Ziklag, Madmannah, Sansannah,
JOSH|15|32|Lebaoth, Shilhim, Ain and Rimmon-a total of twenty-nine towns and their villages.
JOSH|15|33|In the western foothills: Eshtaol, Zorah, Ashnah,
JOSH|15|34|Zanoah, En Gannim, Tappuah, Enam,
JOSH|15|35|Jarmuth, Adullam, Socoh, Azekah,
JOSH|15|36|Shaaraim, Adithaim and Gederah (or Gederothaim) -fourteen towns and their villages.
JOSH|15|37|Zenan, Hadashah, Migdal Gad,
JOSH|15|38|Dilean, Mizpah, Joktheel,
JOSH|15|39|Lachish, Bozkath, Eglon,
JOSH|15|40|Cabbon, Lahmas, Kitlish,
JOSH|15|41|Gederoth, Beth Dagon, Naamah and Makkedah-sixteen towns and their villages.
JOSH|15|42|Libnah, Ether, Ashan,
JOSH|15|43|Iphtah, Ashnah, Nezib,
JOSH|15|44|Keilah, Aczib and Mareshah-nine towns and their villages.
JOSH|15|45|Ekron, with its surrounding settlements and villages;
JOSH|15|46|west of Ekron, all that were in the vicinity of Ashdod, together with their villages;
JOSH|15|47|Ashdod, its surrounding settlements and villages; and Gaza, its settlements and villages, as far as the Wadi of Egypt and the coastline of the Great Sea.
JOSH|15|48|In the hill country: Shamir, Jattir, Socoh,
JOSH|15|49|Dannah, Kiriath Sannah (that is, Debir),
JOSH|15|50|Anab, Eshtemoh, Anim,
JOSH|15|51|Goshen, Holon and Giloh-eleven towns and their villages.
JOSH|15|52|Arab, Dumah, Eshan,
JOSH|15|53|Janim, Beth Tappuah, Aphekah,
JOSH|15|54|Humtah, Kiriath Arba (that is, Hebron) and Zior-nine towns and their villages.
JOSH|15|55|Maon, Carmel, Ziph, Juttah,
JOSH|15|56|Jezreel, Jokdeam, Zanoah,
JOSH|15|57|Kain, Gibeah and Timnah-ten towns and their villages.
JOSH|15|58|Halhul, Beth Zur, Gedor,
JOSH|15|59|Maarath, Beth Anoth and Eltekon-six towns and their villages.
JOSH|15|60|Kiriath Baal (that is, Kiriath Jearim) and Rabbah-two towns and their villages.
JOSH|15|61|In the desert: Beth Arabah, Middin, Secacah,
JOSH|15|62|Nibshan, the City of Salt and En Gedi-six towns and their villages.
JOSH|15|63|Judah could not dislodge the Jebusites, who were living in Jerusalem; to this day the Jebusites live there with the people of Judah.
JOSH|16|1|The allotment for Joseph began at the Jordan of Jericho, east of the waters of Jericho, and went up from there through the desert into the hill country of Bethel.
JOSH|16|2|It went on from Bethel (that is, Luz), crossed over to the territory of the Arkites in Ataroth,
JOSH|16|3|descended westward to the territory of the Japhletites as far as the region of Lower Beth Horon and on to Gezer, ending at the sea.
JOSH|16|4|So Manasseh and Ephraim, the descendants of Joseph, received their inheritance.
JOSH|16|5|This was the territory of Ephraim, clan by clan: The boundary of their inheritance went from Ataroth Addar in the east to Upper Beth Horon
JOSH|16|6|and continued to the sea. From Micmethath on the north it curved eastward to Taanath Shiloh, passing by it to Janoah on the east.
JOSH|16|7|Then it went down from Janoah to Ataroth and Naarah, touched Jericho and came out at the Jordan.
JOSH|16|8|From Tappuah the border went west to the Kanah Ravine and ended at the sea. This was the inheritance of the tribe of the Ephraimites, clan by clan.
JOSH|16|9|It also included all the towns and their villages that were set aside for the Ephraimites within the inheritance of the Manassites.
JOSH|16|10|They did not dislodge the Canaanites living in Gezer; to this day the Canaanites live among the people of Ephraim but are required to do forced labor.
JOSH|17|1|This was the allotment for the tribe of Manasseh as Joseph's firstborn, that is, for Makir, Manasseh's firstborn. Makir was the ancestor of the Gileadites, who had received Gilead and Bashan because the Makirites were great soldiers.
JOSH|17|2|So this allotment was for the rest of the people of Manasseh-the clans of Abiezer, Helek, Asriel, Shechem, Hepher and Shemida. These are the other male descendants of Manasseh son of Joseph by their clans.
JOSH|17|3|Now Zelophehad son of Hepher, the son of Gilead, the son of Makir, the son of Manasseh, had no sons but only daughters, whose names were Mahlah, Noah, Hoglah, Milcah and Tirzah.
JOSH|17|4|They went to Eleazar the priest, Joshua son of Nun, and the leaders and said, "The LORD commanded Moses to give us an inheritance among our brothers." So Joshua gave them an inheritance along with the brothers of their father, according to the LORD's command.
JOSH|17|5|Manasseh's share consisted of ten tracts of land besides Gilead and Bashan east of the Jordan,
JOSH|17|6|because the daughters of the tribe of Manasseh received an inheritance among the sons. The land of Gilead belonged to the rest of the descendants of Manasseh.
JOSH|17|7|The territory of Manasseh extended from Asher to Micmethath east of Shechem. The boundary ran southward from there to include the people living at En Tappuah.
JOSH|17|8|(Manasseh had the land of Tappuah, but Tappuah itself, on the boundary of Manasseh, belonged to the Ephraimites.)
JOSH|17|9|Then the boundary continued south to the Kanah Ravine. There were towns belonging to Ephraim lying among the towns of Manasseh, but the boundary of Manasseh was the northern side of the ravine and ended at the sea.
JOSH|17|10|On the south the land belonged to Ephraim, on the north to Manasseh. The territory of Manasseh reached the sea and bordered Asher on the north and Issachar on the east.
JOSH|17|11|Within Issachar and Asher, Manasseh also had Beth Shan, Ibleam and the people of Dor, Endor, Taanach and Megiddo, together with their surrounding settlements (the third in the list is Naphoth ).
JOSH|17|12|Yet the Manassites were not able to occupy these towns, for the Canaanites were determined to live in that region.
JOSH|17|13|However, when the Israelites grew stronger, they subjected the Canaanites to forced labor but did not drive them out completely.
JOSH|17|14|The people of Joseph said to Joshua, "Why have you given us only one allotment and one portion for an inheritance? We are a numerous people and the LORD has blessed us abundantly."
JOSH|17|15|"If you are so numerous," Joshua answered, "and if the hill country of Ephraim is too small for you, go up into the forest and clear land for yourselves there in the land of the Perizzites and Rephaites."
JOSH|17|16|The people of Joseph replied, "The hill country is not enough for us, and all the Canaanites who live in the plain have iron chariots, both those in Beth Shan and its settlements and those in the Valley of Jezreel."
JOSH|17|17|But Joshua said to the house of Joseph-to Ephraim and Manasseh-"You are numerous and very powerful. You will have not only one allotment
JOSH|17|18|but the forested hill country as well. Clear it, and its farthest limits will be yours; though the Canaanites have iron chariots and though they are strong, you can drive them out."
JOSH|18|1|The whole assembly of the Israelites gathered at Shiloh and set up the Tent of Meeting there. The country was brought under their control,
JOSH|18|2|but there were still seven Israelite tribes who had not yet received their inheritance.
JOSH|18|3|So Joshua said to the Israelites: "How long will you wait before you begin to take possession of the land that the LORD, the God of your fathers, has given you?
JOSH|18|4|Appoint three men from each tribe. I will send them out to make a survey of the land and to write a description of it, according to the inheritance of each. Then they will return to me.
JOSH|18|5|You are to divide the land into seven parts. Judah is to remain in its territory on the south and the house of Joseph in its territory on the north.
JOSH|18|6|After you have written descriptions of the seven parts of the land, bring them here to me and I will cast lots for you in the presence of the LORD our God.
JOSH|18|7|The Levites, however, do not get a portion among you, because the priestly service of the LORD is their inheritance. And Gad, Reuben and the half-tribe of Manasseh have already received their inheritance on the east side of the Jordan. Moses the servant of the LORD gave it to them."
JOSH|18|8|As the men started on their way to map out the land, Joshua instructed them, "Go and make a survey of the land and write a description of it. Then return to me, and I will cast lots for you here at Shiloh in the presence of the LORD."
JOSH|18|9|So the men left and went through the land. They wrote its description on a scroll, town by town, in seven parts, and returned to Joshua in the camp at Shiloh.
JOSH|18|10|Joshua then cast lots for them in Shiloh in the presence of the LORD, and there he distributed the land to the Israelites according to their tribal divisions.
JOSH|18|11|The lot came up for the tribe of Benjamin, clan by clan. Their allotted territory lay between the tribes of Judah and Joseph:
JOSH|18|12|On the north side their boundary began at the Jordan, passed the northern slope of Jericho and headed west into the hill country, coming out at the desert of Beth Aven.
JOSH|18|13|From there it crossed to the south slope of Luz (that is, Bethel) and went down to Ataroth Addar on the hill south of Lower Beth Horon.
JOSH|18|14|From the hill facing Beth Horon on the south the boundary turned south along the western side and came out at Kiriath Baal (that is, Kiriath Jearim), a town of the people of Judah. This was the western side.
JOSH|18|15|The southern side began at the outskirts of Kiriath Jearim on the west, and the boundary came out at the spring of the waters of Nephtoah.
JOSH|18|16|The boundary went down to the foot of the hill facing the Valley of Ben Hinnom, north of the Valley of Rephaim. It continued down the Hinnom Valley along the southern slope of the Jebusite city and so to En Rogel.
JOSH|18|17|It then curved north, went to En Shemesh, continued to Geliloth, which faces the Pass of Adummim, and ran down to the Stone of Bohan son of Reuben.
JOSH|18|18|It continued to the northern slope of Beth Arabah and on down into the Arabah.
JOSH|18|19|It then went to the northern slope of Beth Hoglah and came out at the northern bay of the Salt Sea, at the mouth of the Jordan in the south. This was the southern boundary.
JOSH|18|20|The Jordan formed the boundary on the eastern side. These were the boundaries that marked out the inheritance of the clans of Benjamin on all sides.
JOSH|18|21|The tribe of Benjamin, clan by clan, had the following cities: Jericho, Beth Hoglah, Emek Keziz,
JOSH|18|22|Beth Arabah, Zemaraim, Bethel,
JOSH|18|23|Avvim, Parah, Ophrah,
JOSH|18|24|Kephar Ammoni, Ophni and Geba-twelve towns and their villages.
JOSH|18|25|Gibeon, Ramah, Beeroth,
JOSH|18|26|Mizpah, Kephirah, Mozah,
JOSH|18|27|Rekem, Irpeel, Taralah,
JOSH|18|28|Zelah, Haeleph, the Jebusite city (that is, Jerusalem), Gibeah and Kiriath-fourteen towns and their villages. This was the inheritance of Benjamin for its clans.
JOSH|19|1|The second lot came out for the tribe of Simeon, clan by clan. Their inheritance lay within the territory of Judah.
JOSH|19|2|It included: Beersheba (or Sheba), Moladah,
JOSH|19|3|Hazar Shual, Balah, Ezem,
JOSH|19|4|Eltolad, Bethul, Hormah,
JOSH|19|5|Ziklag, Beth Marcaboth, Hazar Susah,
JOSH|19|6|Beth Lebaoth and Sharuhen-thirteen towns and their villages;
JOSH|19|7|Ain, Rimmon, Ether and Ashan-four towns and their villages-
JOSH|19|8|and all the villages around these towns as far as Baalath Beer (Ramah in the Negev). This was the inheritance of the tribe of the Simeonites, clan by clan.
JOSH|19|9|The inheritance of the Simeonites was taken from the share of Judah, because Judah's portion was more than they needed. So the Simeonites received their inheritance within the territory of Judah.
JOSH|19|10|The third lot came up for Zebulun, clan by clan: The boundary of their inheritance went as far as Sarid.
JOSH|19|11|Going west it ran to Maralah, touched Dabbesheth, and extended to the ravine near Jokneam.
JOSH|19|12|It turned east from Sarid toward the sunrise to the territory of Kisloth Tabor and went on to Daberath and up to Japhia.
JOSH|19|13|Then it continued eastward to Gath Hepher and Eth Kazin; it came out at Rimmon and turned toward Neah.
JOSH|19|14|There the boundary went around on the north to Hannathon and ended at the Valley of Iphtah El.
JOSH|19|15|Included were Kattath, Nahalal, Shimron, Idalah and Bethlehem. There were twelve towns and their villages.
JOSH|19|16|These towns and their villages were the inheritance of Zebulun, clan by clan.
JOSH|19|17|The fourth lot came out for Issachar, clan by clan.
JOSH|19|18|Their territory included: Jezreel, Kesulloth, Shunem,
JOSH|19|19|Hapharaim, Shion, Anaharath,
JOSH|19|20|Rabbith, Kishion, Ebez,
JOSH|19|21|Remeth, En Gannim, En Haddah and Beth Pazzez.
JOSH|19|22|The boundary touched Tabor, Shahazumah and Beth Shemesh, and ended at the Jordan. There were sixteen towns and their villages.
JOSH|19|23|These towns and their villages were the inheritance of the tribe of Issachar, clan by clan.
JOSH|19|24|The fifth lot came out for the tribe of Asher, clan by clan.
JOSH|19|25|Their territory included: Helkath, Hali, Beten, Acshaph,
JOSH|19|26|Allammelech, Amad and Mishal. On the west the boundary touched Carmel and Shihor Libnath.
JOSH|19|27|It then turned east toward Beth Dagon, touched Zebulun and the Valley of Iphtah El, and went north to Beth Emek and Neiel, passing Cabul on the left.
JOSH|19|28|It went to Abdon, Rehob, Hammon and Kanah, as far as Greater Sidon.
JOSH|19|29|The boundary then turned back toward Ramah and went to the fortified city of Tyre, turned toward Hosah and came out at the sea in the region of Aczib,
JOSH|19|30|Ummah, Aphek and Rehob. There were twenty-two towns and their villages.
JOSH|19|31|These towns and their villages were the inheritance of the tribe of Asher, clan by clan.
JOSH|19|32|The sixth lot came out for Naphtali, clan by clan:
JOSH|19|33|Their boundary went from Heleph and the large tree in Zaanannim, passing Adami Nekeb and Jabneel to Lakkum and ending at the Jordan.
JOSH|19|34|The boundary ran west through Aznoth Tabor and came out at Hukkok. It touched Zebulun on the south, Asher on the west and the Jordan on the east.
JOSH|19|35|The fortified cities were Ziddim, Zer, Hammath, Rakkath, Kinnereth,
JOSH|19|36|Adamah, Ramah, Hazor,
JOSH|19|37|Kedesh, Edrei, En Hazor,
JOSH|19|38|Iron, Migdal El, Horem, Beth Anath and Beth Shemesh. There were nineteen towns and their villages.
JOSH|19|39|These towns and their villages were the inheritance of the tribe of Naphtali, clan by clan.
JOSH|19|40|The seventh lot came out for the tribe of Dan, clan by clan.
JOSH|19|41|The territory of their inheritance included: Zorah, Eshtaol, Ir Shemesh,
JOSH|19|42|Shaalabbin, Aijalon, Ithlah,
JOSH|19|43|Elon, Timnah, Ekron,
JOSH|19|44|Eltekeh, Gibbethon, Baalath,
JOSH|19|45|Jehud, Bene Berak, Gath Rimmon,
JOSH|19|46|Me Jarkon and Rakkon, with the area facing Joppa.
JOSH|19|47|(But the Danites had difficulty taking possession of their territory, so they went up and attacked Leshem, took it, put it to the sword and occupied it. They settled in Leshem and named it Dan after their forefather.)
JOSH|19|48|These towns and their villages were the inheritance of the tribe of Dan, clan by clan.
JOSH|19|49|When they had finished dividing the land into its allotted portions, the Israelites gave Joshua son of Nun an inheritance among them,
JOSH|19|50|as the LORD had commanded. They gave him the town he asked for-Timnath Serah in the hill country of Ephraim. And he built up the town and settled there.
JOSH|19|51|These are the territories that Eleazar the priest, Joshua son of Nun and the heads of the tribal clans of Israel assigned by lot at Shiloh in the presence of the LORD at the entrance to the Tent of Meeting. And so they finished dividing the land.
JOSH|20|1|Then the LORD said to Joshua:
JOSH|20|2|"Tell the Israelites to designate the cities of refuge, as I instructed you through Moses,
JOSH|20|3|so that anyone who kills a person accidentally and unintentionally may flee there and find protection from the avenger of blood.
JOSH|20|4|"When he flees to one of these cities, he is to stand in the entrance of the city gate and state his case before the elders of that city. Then they are to admit him into their city and give him a place to live with them.
JOSH|20|5|If the avenger of blood pursues him, they must not surrender the one accused, because he killed his neighbor unintentionally and without malice aforethought.
JOSH|20|6|He is to stay in that city until he has stood trial before the assembly and until the death of the high priest who is serving at that time. Then he may go back to his own home in the town from which he fled."
JOSH|20|7|So they set apart Kedesh in Galilee in the hill country of Naphtali, Shechem in the hill country of Ephraim, and Kiriath Arba (that is, Hebron) in the hill country of Judah.
JOSH|20|8|On the east side of the Jordan of Jericho they designated Bezer in the desert on the plateau in the tribe of Reuben, Ramoth in Gilead in the tribe of Gad, and Golan in Bashan in the tribe of Manasseh.
JOSH|20|9|Any of the Israelites or any alien living among them who killed someone accidentally could flee to these designated cities and not be killed by the avenger of blood prior to standing trial before the assembly.
JOSH|21|1|Now the family heads of the Levites approached Eleazar the priest, Joshua son of Nun, and the heads of the other tribal families of Israel
JOSH|21|2|at Shiloh in Canaan and said to them, "The LORD commanded through Moses that you give us towns to live in, with pasturelands for our livestock."
JOSH|21|3|So, as the LORD had commanded, the Israelites gave the Levites the following towns and pasturelands out of their own inheritance:
JOSH|21|4|The first lot came out for the Kohathites, clan by clan. The Levites who were descendants of Aaron the priest were allotted thirteen towns from the tribes of Judah, Simeon and Benjamin.
JOSH|21|5|The rest of Kohath's descendants were allotted ten towns from the clans of the tribes of Ephraim, Dan and half of Manasseh.
JOSH|21|6|The descendants of Gershon were allotted thirteen towns from the clans of the tribes of Issachar, Asher, Naphtali and the half-tribe of Manasseh in Bashan.
JOSH|21|7|The descendants of Merari, clan by clan, received twelve towns from the tribes of Reuben, Gad and Zebulun.
JOSH|21|8|So the Israelites allotted to the Levites these towns and their pasturelands, as the LORD had commanded through Moses.
JOSH|21|9|From the tribes of Judah and Simeon they allotted the following towns by name
JOSH|21|10|(these towns were assigned to the descendants of Aaron who were from the Kohathite clans of the Levites, because the first lot fell to them):
JOSH|21|11|They gave them Kiriath Arba (that is, Hebron), with its surrounding pastureland, in the hill country of Judah. (Arba was the forefather of Anak.)
JOSH|21|12|But the fields and villages around the city they had given to Caleb son of Jephunneh as his possession.
JOSH|21|13|So to the descendants of Aaron the priest they gave Hebron (a city of refuge for one accused of murder), Libnah,
JOSH|21|14|Jattir, Eshtemoa,
JOSH|21|15|Holon, Debir,
JOSH|21|16|Ain, Juttah and Beth Shemesh, together with their pasturelands-nine towns from these two tribes.
JOSH|21|17|And from the tribe of Benjamin they gave them Gibeon, Geba,
JOSH|21|18|Anathoth and Almon, together with their pasturelands-four towns.
JOSH|21|19|All the towns for the priests, the descendants of Aaron, were thirteen, together with their pasturelands.
JOSH|21|20|The rest of the Kohathite clans of the Levites were allotted towns from the tribe of Ephraim:
JOSH|21|21|In the hill country of Ephraim they were given Shechem (a city of refuge for one accused of murder) and Gezer,
JOSH|21|22|Kibzaim and Beth Horon, together with their pasturelands-four towns.
JOSH|21|23|Also from the tribe of Dan they received Eltekeh, Gibbethon,
JOSH|21|24|Aijalon and Gath Rimmon, together with their pasturelands-four towns.
JOSH|21|25|From half the tribe of Manasseh they received Taanach and Gath Rimmon, together with their pasturelands-two towns.
JOSH|21|26|All these ten towns and their pasturelands were given to the rest of the Kohathite clans.
JOSH|21|27|The Levite clans of the Gershonites were given: from the half-tribe of Manasseh, Golan in Bashan (a city of refuge for one accused of murder) and Be Eshtarah, together with their pasturelands-two towns;
JOSH|21|28|from the tribe of Issachar, Kishion, Daberath,
JOSH|21|29|Jarmuth and En Gannim, together with their pasturelands-four towns;
JOSH|21|30|from the tribe of Asher, Mishal, Abdon,
JOSH|21|31|Helkath and Rehob, together with their pasturelands-four towns;
JOSH|21|32|from the tribe of Naphtali, Kedesh in Galilee (a city of refuge for one accused of murder), Hammoth Dor and Kartan, together with their pasturelands-three towns.
JOSH|21|33|All the towns of the Gershonite clans were thirteen, together with their pasturelands.
JOSH|21|34|The Merarite clans (the rest of the Levites) were given: from the tribe of Zebulun, Jokneam, Kartah,
JOSH|21|35|Dimnah and Nahalal, together with their pasturelands-four towns;
JOSH|21|36|from the tribe of Reuben, Bezer, Jahaz,
JOSH|21|37|Kedemoth and Mephaath, together with their pasturelands-four towns;
JOSH|21|38|from the tribe of Gad, Ramoth in Gilead (a city of refuge for one accused of murder), Mahanaim,
JOSH|21|39|Heshbon and Jazer, together with their pasturelands-four towns in all.
JOSH|21|40|All the towns allotted to the Merarite clans, who were the rest of the Levites, were twelve.
JOSH|21|41|The towns of the Levites in the territory held by the Israelites were forty-eight in all, together with their pasturelands.
JOSH|21|42|Each of these towns had pasturelands surrounding it; this was true for all these towns.
JOSH|21|43|So the LORD gave Israel all the land he had sworn to give their forefathers, and they took possession of it and settled there.
JOSH|21|44|The LORD gave them rest on every side, just as he had sworn to their forefathers. Not one of their enemies withstood them; the LORD handed all their enemies over to them.
JOSH|21|45|Not one of all the LORD's good promises to the house of Israel failed; every one was fulfilled.
JOSH|22|1|Then Joshua summoned the Reubenites, the Gadites and the half-tribe of Manasseh
JOSH|22|2|and said to them, "You have done all that Moses the servant of the LORD commanded, and you have obeyed me in everything I commanded.
JOSH|22|3|For a long time now-to this very day-you have not deserted your brothers but have carried out the mission the LORD your God gave you.
JOSH|22|4|Now that the LORD your God has given your brothers rest as he promised, return to your homes in the land that Moses the servant of the LORD gave you on the other side of the Jordan.
JOSH|22|5|But be very careful to keep the commandment and the law that Moses the servant of the LORD gave you: to love the LORD your God, to walk in all his ways, to obey his commands, to hold fast to him and to serve him with all your heart and all your soul."
JOSH|22|6|Then Joshua blessed them and sent them away, and they went to their homes.
JOSH|22|7|(To the half-tribe of Manasseh Moses had given land in Bashan, and to the other half of the tribe Joshua gave land on the west side of the Jordan with their brothers.) When Joshua sent them home, he blessed them,
JOSH|22|8|saying, "Return to your homes with your great wealth-with large herds of livestock, with silver, gold, bronze and iron, and a great quantity of clothing-and divide with your brothers the plunder from your enemies."
JOSH|22|9|So the Reubenites, the Gadites and the half-tribe of Manasseh left the Israelites at Shiloh in Canaan to return to Gilead, their own land, which they had acquired in accordance with the command of the LORD through Moses.
JOSH|22|10|When they came to Geliloth near the Jordan in the land of Canaan, the Reubenites, the Gadites and the half-tribe of Manasseh built an imposing altar there by the Jordan.
JOSH|22|11|And when the Israelites heard that they had built the altar on the border of Canaan at Geliloth near the Jordan on the Israelite side,
JOSH|22|12|the whole assembly of Israel gathered at Shiloh to go to war against them.
JOSH|22|13|So the Israelites sent Phinehas son of Eleazar, the priest, to the land of Gilead-to Reuben, Gad and the half-tribe of Manasseh.
JOSH|22|14|With him they sent ten of the chief men, one for each of the tribes of Israel, each the head of a family division among the Israelite clans.
JOSH|22|15|When they went to Gilead-to Reuben, Gad and the half-tribe of Manasseh-they said to them:
JOSH|22|16|"The whole assembly of the LORD says: 'How could you break faith with the God of Israel like this? How could you turn away from the LORD and build yourselves an altar in rebellion against him now?
JOSH|22|17|Was not the sin of Peor enough for us? Up to this very day we have not cleansed ourselves from that sin, even though a plague fell on the community of the LORD!
JOSH|22|18|And are you now turning away from the LORD? "'If you rebel against the LORD today, tomorrow he will be angry with the whole community of Israel.
JOSH|22|19|If the land you possess is defiled, come over to the LORD's land, where the LORD's tabernacle stands, and share the land with us. But do not rebel against the LORD or against us by building an altar for yourselves, other than the altar of the LORD our God.
JOSH|22|20|When Achan son of Zerah acted unfaithfully regarding the devoted things, did not wrath come upon the whole community of Israel? He was not the only one who died for his sin.'"
JOSH|22|21|Then Reuben, Gad and the half-tribe of Manasseh replied to the heads of the clans of Israel:
JOSH|22|22|"The Mighty One, God, the LORD! The Mighty One, God, the LORD! He knows! And let Israel know! If this has been in rebellion or disobedience to the LORD, do not spare us this day.
JOSH|22|23|If we have built our own altar to turn away from the LORD and to offer burnt offerings and grain offerings, or to sacrifice fellowship offerings on it, may the LORD himself call us to account.
JOSH|22|24|"No! We did it for fear that some day your descendants might say to ours, 'What do you have to do with the LORD, the God of Israel?
JOSH|22|25|The LORD has made the Jordan a boundary between us and you-you Reubenites and Gadites! You have no share in the LORD.' So your descendants might cause ours to stop fearing the LORD.
JOSH|22|26|"That is why we said, 'Let us get ready and build an altar-but not for burnt offerings or sacrifices.'
JOSH|22|27|On the contrary, it is to be a witness between us and you and the generations that follow, that we will worship the LORD at his sanctuary with our burnt offerings, sacrifices and fellowship offerings. Then in the future your descendants will not be able to say to ours, 'You have no share in the LORD.'
JOSH|22|28|"And we said, 'If they ever say this to us, or to our descendants, we will answer: Look at the replica of the LORD's altar, which our fathers built, not for burnt offerings and sacrifices, but as a witness between us and you.'
JOSH|22|29|"Far be it from us to rebel against the LORD and turn away from him today by building an altar for burnt offerings, grain offerings and sacrifices, other than the altar of the LORD our God that stands before his tabernacle."
JOSH|22|30|When Phinehas the priest and the leaders of the community-the heads of the clans of the Israelites-heard what Reuben, Gad and Manasseh had to say, they were pleased.
JOSH|22|31|And Phinehas son of Eleazar, the priest, said to Reuben, Gad and Manasseh, "Today we know that the LORD is with us, because you have not acted unfaithfully toward the LORD in this matter. Now you have rescued the Israelites from the LORD's hand."
JOSH|22|32|Then Phinehas son of Eleazar, the priest, and the leaders returned to Canaan from their meeting with the Reubenites and Gadites in Gilead and reported to the Israelites.
JOSH|22|33|They were glad to hear the report and praised God. And they talked no more about going to war against them to devastate the country where the Reubenites and the Gadites lived.
JOSH|22|34|And the Reubenites and the Gadites gave the altar this name: A Witness Between Us that the LORD is God.
JOSH|23|1|After a long time had passed and the LORD had given Israel rest from all their enemies around them, Joshua, by then old and well advanced in years,
JOSH|23|2|summoned all Israel-their elders, leaders, judges and officials-and said to them: "I am old and well advanced in years.
JOSH|23|3|You yourselves have seen everything the LORD your God has done to all these nations for your sake; it was the LORD your God who fought for you.
JOSH|23|4|Remember how I have allotted as an inheritance for your tribes all the land of the nations that remain-the nations I conquered-between the Jordan and the Great Sea in the west.
JOSH|23|5|The LORD your God himself will drive them out of your way. He will push them out before you, and you will take possession of their land, as the LORD your God promised you.
JOSH|23|6|"Be very strong; be careful to obey all that is written in the Book of the Law of Moses, without turning aside to the right or to the left.
JOSH|23|7|Do not associate with these nations that remain among you; do not invoke the names of their gods or swear by them. You must not serve them or bow down to them.
JOSH|23|8|But you are to hold fast to the LORD your God, as you have until now.
JOSH|23|9|"The LORD has driven out before you great and powerful nations; to this day no one has been able to withstand you.
JOSH|23|10|One of you routs a thousand, because the LORD your God fights for you, just as he promised.
JOSH|23|11|So be very careful to love the LORD your God.
JOSH|23|12|"But if you turn away and ally yourselves with the survivors of these nations that remain among you and if you intermarry with them and associate with them,
JOSH|23|13|then you may be sure that the LORD your God will no longer drive out these nations before you. Instead, they will become snares and traps for you, whips on your backs and thorns in your eyes, until you perish from this good land, which the LORD your God has given you.
JOSH|23|14|"Now I am about to go the way of all the earth. You know with all your heart and soul that not one of all the good promises the LORD your God gave you has failed. Every promise has been fulfilled; not one has failed.
JOSH|23|15|But just as every good promise of the LORD your God has come true, so the LORD will bring on you all the evil he has threatened, until he has destroyed you from this good land he has given you.
JOSH|23|16|If you violate the covenant of the LORD your God, which he commanded you, and go and serve other gods and bow down to them, the LORD's anger will burn against you, and you will quickly perish from the good land he has given you."
JOSH|24|1|Then Joshua assembled all the tribes of Israel at Shechem. He summoned the elders, leaders, judges and officials of Israel, and they presented themselves before God.
JOSH|24|2|Joshua said to all the people, "This is what the LORD, the God of Israel, says: 'Long ago your forefathers, including Terah the father of Abraham and Nahor, lived beyond the River and worshiped other gods.
JOSH|24|3|But I took your father Abraham from the land beyond the River and led him throughout Canaan and gave him many descendants. I gave him Isaac,
JOSH|24|4|and to Isaac I gave Jacob and Esau. I assigned the hill country of Seir to Esau, but Jacob and his sons went down to Egypt.
JOSH|24|5|"'Then I sent Moses and Aaron, and I afflicted the Egyptians by what I did there, and I brought you out.
JOSH|24|6|When I brought your fathers out of Egypt, you came to the sea, and the Egyptians pursued them with chariots and horsemen as far as the Red Sea.
JOSH|24|7|But they cried to the LORD for help, and he put darkness between you and the Egyptians; he brought the sea over them and covered them. You saw with your own eyes what I did to the Egyptians. Then you lived in the desert for a long time.
JOSH|24|8|"'I brought you to the land of the Amorites who lived east of the Jordan. They fought against you, but I gave them into your hands. I destroyed them from before you, and you took possession of their land.
JOSH|24|9|When Balak son of Zippor, the king of Moab, prepared to fight against Israel, he sent for Balaam son of Beor to put a curse on you.
JOSH|24|10|But I would not listen to Balaam, so he blessed you again and again, and I delivered you out of his hand.
JOSH|24|11|"'Then you crossed the Jordan and came to Jericho. The citizens of Jericho fought against you, as did also the Amorites, Perizzites, Canaanites, Hittites, Girgashites, Hivites and Jebusites, but I gave them into your hands.
JOSH|24|12|I sent the hornet ahead of you, which drove them out before you-also the two Amorite kings. You did not do it with your own sword and bow.
JOSH|24|13|So I gave you a land on which you did not toil and cities you did not build; and you live in them and eat from vineyards and olive groves that you did not plant.'
JOSH|24|14|"Now fear the LORD and serve him with all faithfulness. Throw away the gods your forefathers worshiped beyond the River and in Egypt, and serve the LORD.
JOSH|24|15|But if serving the LORD seems undesirable to you, then choose for yourselves this day whom you will serve, whether the gods your forefathers served beyond the River, or the gods of the Amorites, in whose land you are living. But as for me and my household, we will serve the LORD."
JOSH|24|16|Then the people answered, "Far be it from us to forsake the LORD to serve other gods!
JOSH|24|17|It was the LORD our God himself who brought us and our fathers up out of Egypt, from that land of slavery, and performed those great signs before our eyes. He protected us on our entire journey and among all the nations through which we traveled.
JOSH|24|18|And the LORD drove out before us all the nations, including the Amorites, who lived in the land. We too will serve the LORD, because he is our God."
JOSH|24|19|Joshua said to the people, "You are not able to serve the LORD. He is a holy God; he is a jealous God. He will not forgive your rebellion and your sins.
JOSH|24|20|If you forsake the LORD and serve foreign gods, he will turn and bring disaster on you and make an end of you, after he has been good to you."
JOSH|24|21|But the people said to Joshua, "No! We will serve the LORD."
JOSH|24|22|Then Joshua said, "You are witnesses against yourselves that you have chosen to serve the LORD.Yes, we are witnesses," they replied.
JOSH|24|23|"Now then," said Joshua, "throw away the foreign gods that are among you and yield your hearts to the LORD, the God of Israel."
JOSH|24|24|And the people said to Joshua, "We will serve the LORD our God and obey him."
JOSH|24|25|On that day Joshua made a covenant for the people, and there at Shechem he drew up for them decrees and laws.
JOSH|24|26|And Joshua recorded these things in the Book of the Law of God. Then he took a large stone and set it up there under the oak near the holy place of the LORD.
JOSH|24|27|"See!" he said to all the people. "This stone will be a witness against us. It has heard all the words the LORD has said to us. It will be a witness against you if you are untrue to your God."
JOSH|24|28|Then Joshua sent the people away, each to his own inheritance.
JOSH|24|29|After these things, Joshua son of Nun, the servant of the LORD, died at the age of a hundred and ten.
JOSH|24|30|And they buried him in the land of his inheritance, at Timnath Serah in the hill country of Ephraim, north of Mount Gaash.
JOSH|24|31|Israel served the LORD throughout the lifetime of Joshua and of the elders who outlived him and who had experienced everything the LORD had done for Israel.
JOSH|24|32|And Joseph's bones, which the Israelites had brought up from Egypt, were buried at Shechem in the tract of land that Jacob bought for a hundred pieces of silver from the sons of Hamor, the father of Shechem. This became the inheritance of Joseph's descendants.
JOSH|24|33|And Eleazar son of Aaron died and was buried at Gibeah, which had been allotted to his son Phinehas in the hill country of Ephraim.
