RUTH|1|1|士師統治的時候，國中有饑荒。在 猶大 的 伯利恆 ，有一個人帶著妻子和兩個兒子往 摩押 地去寄居。
RUTH|1|2|這人名叫 以利米勒 ，他的妻子名叫 拿娥米 ；他兩個兒子，一個名叫 瑪倫 ，一個名叫 基連 ，都是 猶大伯利恆 的 以法他 人。他們到了 摩押 地，就住在那裏。
RUTH|1|3|後來 拿娥米 的丈夫 以利米勒 死了，剩下她和兩個兒子。
RUTH|1|4|兩個兒子娶了 摩押 女子，一個名叫 俄珥巴 ，第二個名叫 路得 ，在那裏住了約有十年。
RUTH|1|5|瑪倫 和 基連 二人也死了，剩下 拿娥米 ，沒有丈夫，也沒有兒子。
RUTH|1|6|拿娥米 與兩個媳婦起身，要從 摩押 地回去，因為她在 摩押 地聽見耶和華眷顧自己的百姓，賜糧食給他們。
RUTH|1|7|她和兩個媳婦就起行，離開所住的地方，上路回 猶大 地去。
RUTH|1|8|拿娥米 對兩個媳婦說：「你們各自回娘家去吧！願耶和華恩待你們，像你們待已故的人和我一樣。
RUTH|1|9|願耶和華使你們各自在新的丈夫家中得歸宿！」於是 拿娥米 與她們親吻，她們就放聲大哭，
RUTH|1|10|對她說：「不，我們要與你一同回你的百姓那裏去。」
RUTH|1|11|拿娥米 說：「我的女兒啊，回去吧！為何要跟我去呢？我還能生兒子作你們的丈夫嗎？
RUTH|1|12|我的女兒啊，回去吧！我年紀老了，不能再有丈夫。就算我還有希望，今夜有丈夫，而且也生了兒子，
RUTH|1|13|你們豈能等著他們長大呢？你們能守住自己不嫁人嗎？我的女兒啊，不要這樣。我比你們更苦，因為耶和華伸手擊打我。」
RUTH|1|14|兩個媳婦又放聲大哭， 俄珥巴 與婆婆吻別，但是 路得 卻緊跟著 拿娥米 。
RUTH|1|15|拿娥米 說：「看哪，你嫂嫂已經回她的百姓和她的神明那裏去了，你也跟你嫂嫂回去吧！」
RUTH|1|16|路得 說： 「不要勸我離開你， 轉去不跟隨你。 你往哪裏去， 我也往哪裏去； 你在哪裏住， 我也在哪裏住； 你的百姓就是我的百姓； 你的上帝就是我的上帝。
RUTH|1|17|你死在哪裏， 我也死在哪裏，葬在哪裏。 只有死能使你我分離； 不然，願耶和華重重懲罰我！」
RUTH|1|18|拿娥米 見 路得 決意要跟自己去，就不再對她說甚麼了。
RUTH|1|19|於是二人同行，來到 伯利恆 。她們到了 伯利恆 ，全城因她們騷動起來。婦女們說：「這是 拿娥米 嗎？」
RUTH|1|20|拿娥米 對她們說： 「不要叫我 拿娥米 ， 要叫我 瑪拉 ， 因為全能者使我受盡了苦。
RUTH|1|21|我滿滿地出去， 耶和華使我空空地回來。 耶和華使我受苦， 全能者降禍於我。 你們為何還叫我 拿娥米 呢？」
RUTH|1|22|拿娥米 從 摩押 地回來了，她的媳婦 摩押 女子 路得 跟她在一起。她們到了 伯利恆 ，正是開始收割大麥的時候。
RUTH|2|1|拿娥米 有一個親戚，是她丈夫 以利米勒 本族的人，名叫 波阿斯 ，是個大財主。
RUTH|2|2|摩押 女子 路得 對 拿娥米 說：「讓我到田裏去拾取麥穗，我在誰的眼中蒙恩，就跟在誰的身後。」 拿娥米 說：「女兒啊，你去吧。」
RUTH|2|3|路得 就去了。她來到田間，在收割的人身後拾取麥穗。她恰巧來到 以利米勒 本族的人 波阿斯 那塊田裏。
RUTH|2|4|看哪， 波阿斯 正從 伯利恆 來，對收割的人說：「願耶和華與你們同在！」他們對他說：「願耶和華賜福給你！」
RUTH|2|5|波阿斯 對監督收割的僕人說：「那是誰家的女子？」
RUTH|2|6|監督收割的僕人回答說：「她是 摩押 女子，跟隨 拿娥米 從 摩押 地回來的。
RUTH|2|7|她說：『請你容許我拾取麥穗，在收割的人身後撿禾捆中掉落的麥穗。』她就來了，從早晨直到如今，除了在屋子裏坐一會兒，她都留在這裏。」
RUTH|2|8|波阿斯 對 路得 說：「女兒啊，聽我說，不要到別人田裏去拾取麥穗，也不要離開這裏，要緊跟著我的女僕們。
RUTH|2|9|你要看好我的僕人正在哪塊田收割，就跟著女僕們去。我已經吩咐僕人不可侵犯你。你渴了，可以到水缸那裏喝僕人打來的水。」　
RUTH|2|10|路得 就臉伏於地叩拜，對他說：「我既是外邦女子，怎麼會在你眼中蒙恩，使你這樣照顧我呢？」
RUTH|2|11|波阿斯 回答她說：「自從你丈夫死後，凡你向婆婆所行的，以及你離開父母和你的出生地，到素不相識的百姓中，這些事人都告訴我了。
RUTH|2|12|願耶和華照你所行的報償你。你來投靠在耶和華－ 以色列 上帝的翅膀下，願你滿得他的報償。」
RUTH|2|13|路得 說：「我主啊，願我在你眼前蒙恩。我雖然不及你的一個婢女，你還安慰我，對你的婢女說關心的話。」
RUTH|2|14|吃飯的時候， 波阿斯 對 路得 說：「你到這裏來吃些餅，把你的一塊蘸在醋裏。」 路得 就在收割的人旁邊坐下。 波阿斯 把烘了的穗子遞給她。她吃飽了，還有剩餘的。
RUTH|2|15|她又起來拾取麥穗， 波阿斯 吩咐僕人說：「她即使在禾捆中拾取麥穗，也不可羞辱她。
RUTH|2|16|你們還要從捆裏抽一些出來，留給她拾取，不可責備她。」
RUTH|2|17|這樣， 路得 在田間拾取麥穗，直到晚上。她把所拾取的麥穗打了約有一伊法的大麥。
RUTH|2|18|路得 把所拾取的帶進城去給婆婆看，又把她吃飽所剩的拿出來，給了婆婆。
RUTH|2|19|婆婆問她說：「你今日在哪裏拾取麥穗？在哪裏做工呢？願那照顧你的得福。」 路得 告訴婆婆，她在誰那裏做工，說：「我今日在一個名叫 波阿斯 的人那裏做工。」
RUTH|2|20|拿娥米 對媳婦說：「願那人蒙耶和華賜福，因為他不斷地恩待活人死人。」 拿娥米 又對她說：「那人是我們本族的人，是一個可以贖我們產業的至親。」
RUTH|2|21|摩押 女子 路得 說：「他還對我說：『你要緊跟著我的僕人拾取麥穗，直到他們把我所有的莊稼收割完畢。』」
RUTH|2|22|拿娥米 對媳婦 路得 說：「女兒啊，你要跟著他的女僕出去，免得你在別人的田間受人騷擾。」
RUTH|2|23|於是 路得 緊跟著 波阿斯 的女僕拾取麥穗，直到大麥和小麥收割完畢。 路得 仍與婆婆同住。
RUTH|3|1|路得 的婆婆 拿娥米 對她說：「女兒啊，我不該為你找個歸宿，使你享福嗎？
RUTH|3|2|你與 波阿斯 的女僕常在一處，現在， 波阿斯 不是我們的親人嗎？看哪，他今夜將在禾場簸大麥。
RUTH|3|3|你要沐浴抹膏，穿上外衣，下到禾場，一直到那人吃喝完了，都不要讓他認出你來。
RUTH|3|4|他躺下的時候，你看準他躺臥的地方，就進去掀露他的腳，躺臥在那裏，他必告訴你所當做的事。」
RUTH|3|5|路得 說：「凡你所吩咐我的，我必遵行。」
RUTH|3|6|路得 就下到禾場，照她婆婆吩咐她的一切去做。
RUTH|3|7|波阿斯 吃喝完了，心情暢快，就去躺臥在麥堆旁邊。 路得 悄悄走來，掀露他的腳，躺臥在那裏。
RUTH|3|8|到了半夜，那人驚醒，翻過身來，看哪，有個女子躺在他的腳旁。
RUTH|3|9|他就說：「你是誰？」 路得 說：「我是你的使女 路得 。請你用你衣服的邊來遮蓋你的使女，因為你是可以贖我產業的至親。」
RUTH|3|10|波阿斯 說：「女兒啊，願你蒙耶和華賜福。你後來的忠誠比先前的更美，因為無論貧富的年輕人，你都沒有跟從。
RUTH|3|11|女兒啊，現在不要懼怕，凡你所說的，我必為你做，因為我城裏的百姓都知道你是個賢德的女子。
RUTH|3|12|現在，我的確是一個可以贖你產業的至親，可是還有一個人比我更親。
RUTH|3|13|你今夜在這裏住宿，明早他若肯為你盡至親的本分，很好，就由他吧！倘若他不肯，我指著永生的耶和華起誓，我必為你盡上至親的本分。你只管躺到早晨。」
RUTH|3|14|路得 就在他腳旁躺到早晨，在人還無法彼此辨認的時候就起來了。 波阿斯 說：「不可讓人知道有女子到禾場來。」　
RUTH|3|15|他又對 路得 說：「把你所披的外衣拿來，握緊它。」她就握緊外衣， 波阿斯 量了六簸箕的大麥，幫 路得 扛上，他就進城去了 。」
RUTH|3|16|路得 回到婆婆那裏，婆婆說：「女兒啊，怎麼樣了 ？」 路得 就把那人向她所做的一切都告訴了婆婆，
RUTH|3|17|又說：「那人給了我這六簸箕的大麥，對我說：『你不可空手回去見婆婆。』」
RUTH|3|18|婆婆說：「女兒啊，等著吧，看這事結果如何，因為那人今日不辦妥這事，必不罷休。」
RUTH|4|1|波阿斯 上到城門，坐在那裏，看哪， 波阿斯 所說那個可以贖產業的至親經過。 波阿斯 說：「某某先生，請你轉回來，坐在這裏。」他就轉回來坐下。
RUTH|4|2|波阿斯 又請了本城的十個長老來，對他們說：「請你們坐在這裏。」他們就都坐下。
RUTH|4|3|波阿斯 對那至親說：「從 摩押 地回來的 拿娥米 ，現在要賣我們弟兄 以利米勒 的那塊地。
RUTH|4|4|我想我應該向你說清楚：你可以買那塊地，當著在座的眾人和我百姓的長老面前，你若要贖就贖吧！倘若你不贖 就告訴我，讓我知道，因為除了你以外，沒有人可以先贖，在你之後才輪到我。」那人說：「我要贖。」
RUTH|4|5|波阿斯 說：「你從 拿娥米 和 摩押 女子 路得 手中買這地的時候，也當買死人的妻子，使死人在產業上留名。」
RUTH|4|6|那至親說：「這樣我就不能贖了，免得對我的產業有損。你儘管去贖我所當贖的吧，我不能贖了！」
RUTH|4|7|從前，在 以色列 中要確認任何交易，無論是贖業或買賣，一方必須脫鞋給另一方。 以色列 中都以此為證。
RUTH|4|8|那至親對 波阿斯 說：「你自己買吧！」於是把鞋脫了下來。
RUTH|4|9|波阿斯 對長老和所有在場的百姓說：「你們今日都是證人；凡屬 以利米勒 ，以及 基連 和 瑪倫 的，我都從 拿娥米 手中買下來了。
RUTH|4|10|我也娶 瑪倫 的妻子 摩押 女子 路得 ，好讓死人可以在產業上留名，免得他的名在本族本鄉的城門中消失了。你們今日都是證人。」
RUTH|4|11|在城門坐著的所有百姓和長老說：「我們都是證人。願耶和華使進你家的這女子，像建立 以色列 家的 拉結 和 利亞 二人一樣。又願你在 以法他 得亨通，在 伯利恆 有名聲。
RUTH|4|12|願耶和華從這年輕女子賜你後裔，使你的家像 她瑪 從 猶大 所生 法勒斯 的家一樣。」
RUTH|4|13|於是， 波阿斯 娶了 路得 為妻，與她同房。耶和華使她懷孕生了一個兒子。
RUTH|4|14|婦女們對 拿娥米 說：「耶和華是應當稱頌的！因為他今日沒有使你斷絕可以贖產業的至親。願這孩子在 以色列 中得名聲。
RUTH|4|15|他必振奮你的精神，奉養你的晚年，因為他是愛慕你的媳婦所生的。有這樣的媳婦，比有七個兒子更好！」
RUTH|4|16|拿娥米 接過孩子來，抱在懷中撫養他。
RUTH|4|17|鄰居的婦人給孩子起名，說：「 拿娥米 得了一個孩子了！」她們就給他起名叫 俄備得 。 俄備得 是 耶西 的父親，是 大衛 的祖父。
RUTH|4|18|這是 法勒斯 的後代： 法勒斯 生 希斯崙 ；
RUTH|4|19|希斯崙 生 蘭 ； 蘭 生 亞米拿達 ；
RUTH|4|20|亞米拿達 生 拿順 ； 拿順 生 撒門 ；
RUTH|4|21|撒門 生 波阿斯 ； 波阿斯 生 俄備得 ；
RUTH|4|22|俄備得 生 耶西 ； 耶西 生 大衛 。
