JOHN|1|1|In the beginning was the Word, and the Word was with God, and the Word was God.
JOHN|1|2|He was with God in the beginning.
JOHN|1|3|Through him all things were made; without him nothing was made that has been made.
JOHN|1|4|In him was life, and that life was the light of men.
JOHN|1|5|The light shines in the darkness, but the darkness has not understood it.
JOHN|1|6|There came a man who was sent from God; his name was John.
JOHN|1|7|He came as a witness to testify concerning that light, so that through him all men might believe.
JOHN|1|8|He himself was not the light; he came only as a witness to the light.
JOHN|1|9|The true light that gives light to every man was coming into the world.
JOHN|1|10|He was in the world, and though the world was made through him, the world did not recognize him.
JOHN|1|11|He came to that which was his own, but his own did not receive him.
JOHN|1|12|Yet to all who received him, to those who believed in his name, he gave the right to become children of God--
JOHN|1|13|children born not of natural descent, nor of human decision or a husband's will, but born of God.
JOHN|1|14|The Word became flesh and made his dwelling among us. We have seen his glory, the glory of the One and Only, who came from the Father, full of grace and truth.
JOHN|1|15|John testifies concerning him. He cries out, saying, "This was he of whom I said, 'He who comes after me has surpassed me because he was before me.'"
JOHN|1|16|From the fullness of his grace we have all received one blessing after another.
JOHN|1|17|For the law was given through Moses; grace and truth came through Jesus Christ.
JOHN|1|18|No one has ever seen God, but God the One and Only,, who is at the Father's side, has made him known.
JOHN|1|19|Now this was John's testimony when the Jews of Jerusalem sent priests and Levites to ask him who he was.
JOHN|1|20|He did not fail to confess, but confessed freely, "I am not the Christ. "
JOHN|1|21|They asked him, "Then who are you? Are you Elijah?" He said, "I am not.Are you the Prophet?" He answered, "No."
JOHN|1|22|Finally they said, "Who are you? Give us an answer to take back to those who sent us. What do you say about yourself?"
JOHN|1|23|John replied in the words of Isaiah the prophet, "I am the voice of one calling in the desert, 'Make straight the way for the Lord.'"
JOHN|1|24|Now some Pharisees who had been sent
JOHN|1|25|questioned him, "Why then do you baptize if you are not the Christ, nor Elijah, nor the Prophet?"
JOHN|1|26|"I baptize with water," John replied, "but among you stands one you do not know.
JOHN|1|27|He is the one who comes after me, the thongs of whose sandals I am not worthy to untie."
JOHN|1|28|This all happened at Bethany on the other side of the Jordan, where John was baptizing.
JOHN|1|29|The next day John saw Jesus coming toward him and said, "Look, the Lamb of God, who takes away the sin of the world!
JOHN|1|30|This is the one I meant when I said, 'A man who comes after me has surpassed me because he was before me.'
JOHN|1|31|I myself did not know him, but the reason I came baptizing with water was that he might be revealed to Israel."
JOHN|1|32|Then John gave this testimony: "I saw the Spirit come down from heaven as a dove and remain on him.
JOHN|1|33|I would not have known him, except that the one who sent me to baptize with water told me, 'The man on whom you see the Spirit come down and remain is he who will baptize with the Holy Spirit.'
JOHN|1|34|I have seen and I testify that this is the Son of God."
JOHN|1|35|The next day John was there again with two of his disciples.
JOHN|1|36|When he saw Jesus passing by, he said, "Look, the Lamb of God!"
JOHN|1|37|When the two disciples heard him say this, they followed Jesus.
JOHN|1|38|Turning around, Jesus saw them following and asked, "What do you want?" They said, "Rabbi" (which means Teacher), "where are you staying?"
JOHN|1|39|"Come," he replied, "and you will see." So they went and saw where he was staying, and spent that day with him. It was about the tenth hour.
JOHN|1|40|Andrew, Simon Peter's brother, was one of the two who heard what John had said and who had followed Jesus.
JOHN|1|41|The first thing Andrew did was to find his brother Simon and tell him, "We have found the Messiah" (that is, the Christ).
JOHN|1|42|And he brought him to Jesus. Jesus looked at him and said, "You are Simon son of John. You will be called Cephas" (which, when translated, is Peter ).
JOHN|1|43|The next day Jesus decided to leave for Galilee. Finding Philip, he said to him, "Follow me."
JOHN|1|44|Philip, like Andrew and Peter, was from the town of Bethsaida.
JOHN|1|45|Philip found Nathanael and told him, "We have found the one Moses wrote about in the Law, and about whom the prophets also wrote--Jesus of Nazareth, the son of Joseph."
JOHN|1|46|"Nazareth! Can anything good come from there?" Nathanael asked. "Come and see," said Philip.
JOHN|1|47|When Jesus saw Nathanael approaching, he said of him, "Here is a true Israelite, in whom there is nothing false."
JOHN|1|48|"How do you know me?" Nathanael asked. Jesus answered, "I saw you while you were still under the fig tree before Philip called you."
JOHN|1|49|Then Nathanael declared, "Rabbi, you are the Son of God; you are the King of Israel."
JOHN|1|50|Jesus said, "You believe because I told you I saw you under the fig tree. You shall see greater things than that."
JOHN|1|51|He then added, "I tell you the truth, you shall see heaven open, and the angels of God ascending and descending on the Son of Man."
JOHN|2|1|On the third day a wedding took place at Cana in Galilee. Jesus' mother was there,
JOHN|2|2|and Jesus and his disciples had also been invited to the wedding.
JOHN|2|3|When the wine was gone, Jesus' mother said to him, "They have no more wine."
JOHN|2|4|"Dear woman, why do you involve me?" Jesus replied, "My time has not yet come."
JOHN|2|5|His mother said to the servants, "Do whatever he tells you."
JOHN|2|6|Nearby stood six stone water jars, the kind used by the Jews for ceremonial washing, each holding from twenty to thirty gallons.
JOHN|2|7|Jesus said to the servants, "Fill the jars with water"; so they filled them to the brim.
JOHN|2|8|Then he told them, "Now draw some out and take it to the master of the banquet."
JOHN|2|9|They did so, and the master of the banquet tasted the water that had been turned into wine. He did not realize where it had come from, though the servants who had drawn the water knew. Then he called the bridegroom aside
JOHN|2|10|and said, "Everyone brings out the choice wine first and then the cheaper wine after the guests have had too much to drink; but you have saved the best till now."
JOHN|2|11|This, the first of his miraculous signs, Jesus performed in Cana of Galilee. He thus revealed his glory, and his disciples put their faith in him.
JOHN|2|12|After this he went down to Capernaum with his mother and brothers and his disciples. There they stayed for a few days.
JOHN|2|13|When it was almost time for the Jewish Passover, Jesus went up to Jerusalem.
JOHN|2|14|In the temple courts he found men selling cattle, sheep and doves, and others sitting at tables exchanging money.
JOHN|2|15|So he made a whip out of cords, and drove all from the temple area, both sheep and cattle; he scattered the coins of the money changers and overturned their tables.
JOHN|2|16|To those who sold doves he said, "Get these out of here! How dare you turn my Father's house into a market!"
JOHN|2|17|His disciples remembered that it is written: "Zeal for your house will consume me."
JOHN|2|18|Then the Jews demanded of him, "What miraculous sign can you show us to prove your authority to do all this?"
JOHN|2|19|Jesus answered them, "Destroy this temple, and I will raise it again in three days."
JOHN|2|20|The Jews replied, "It has taken forty-six years to build this temple, and you are going to raise it in three days?"
JOHN|2|21|But the temple he had spoken of was his body.
JOHN|2|22|After he was raised from the dead, his disciples recalled what he had said. Then they believed the Scripture and the words that Jesus had spoken.
JOHN|2|23|Now while he was in Jerusalem at the Passover Feast, many people saw the miraculous signs he was doing and believed in his name.
JOHN|2|24|But Jesus would not entrust himself to them, for he knew all men.
JOHN|2|25|He did not need man's testimony about man, for he knew what was in a man.
JOHN|3|1|Now there was a man of the Pharisees named Nicodemus, a member of the Jewish ruling council.
JOHN|3|2|He came to Jesus at night and said, "Rabbi, we know you are a teacher who has come from God. For no one could perform the miraculous signs you are doing if God were not with him."
JOHN|3|3|In reply Jesus declared, "I tell you the truth, no one can see the kingdom of God unless he is born again. "
JOHN|3|4|"How can a man be born when he is old?" Nicodemus asked. "Surely he cannot enter a second time into his mother's womb to be born!"
JOHN|3|5|Jesus answered, "I tell you the truth, no one can enter the kingdom of God unless he is born of water and the Spirit.
JOHN|3|6|Flesh gives birth to flesh, but the Spirit gives birth to spirit.
JOHN|3|7|You should not be surprised at my saying, 'You must be born again.'
JOHN|3|8|The wind blows wherever it pleases. You hear its sound, but you cannot tell where it comes from or where it is going. So it is with everyone born of the Spirit."
JOHN|3|9|"How can this be?" Nicodemus asked.
JOHN|3|10|"You are Israel's teacher," said Jesus, "and do you not understand these things?
JOHN|3|11|I tell you the truth, we speak of what we know, and we testify to what we have seen, but still you people do not accept our testimony.
JOHN|3|12|I have spoken to you of earthly things and you do not believe; how then will you believe if I speak of heavenly things?
JOHN|3|13|No one has ever gone into heaven except the one who came from heaven--the Son of Man.
JOHN|3|14|Just as Moses lifted up the snake in the desert, so the Son of Man must be lifted up,
JOHN|3|15|that everyone who believes in him may have eternal life.
JOHN|3|16|"For God so loved the world that he gave his one and only Son, that whoever believes in him shall not perish but have eternal life.
JOHN|3|17|For God did not send his Son into the world to condemn the world, but to save the world through him.
JOHN|3|18|Whoever believes in him is not condemned, but whoever does not believe stands condemned already because he has not believed in the name of God's one and only Son.
JOHN|3|19|This is the verdict: Light has come into the world, but men loved darkness instead of light because their deeds were evil.
JOHN|3|20|Everyone who does evil hates the light, and will not come into the light for fear that his deeds will be exposed.
JOHN|3|21|But whoever lives by the truth comes into the light, so that it may be seen plainly that what he has done has been done through God."
JOHN|3|22|After this, Jesus and his disciples went out into the Judean countryside, where he spent some time with them, and baptized.
JOHN|3|23|Now John also was baptizing at Aenon near Salim, because there was plenty of water, and people were constantly coming to be baptized.
JOHN|3|24|(This was before John was put in prison.)
JOHN|3|25|An argument developed between some of John's disciples and a certain Jew over the matter of ceremonial washing.
JOHN|3|26|They came to John and said to him, "Rabbi, that man who was with you on the other side of the Jordan--the one you testified about--well, he is baptizing, and everyone is going to him."
JOHN|3|27|To this John replied, "A man can receive only what is given him from heaven.
JOHN|3|28|You yourselves can testify that I said, 'I am not the Christ but am sent ahead of him.'
JOHN|3|29|The bride belongs to the bridegroom. The friend who attends the bridegroom waits and listens for him, and is full of joy when he hears the bridegroom's voice. That joy is mine, and it is now complete.
JOHN|3|30|He must become greater; I must become less.
JOHN|3|31|"The one who comes from above is above all; the one who is from the earth belongs to the earth, and speaks as one from the earth. The one who comes from heaven is above all.
JOHN|3|32|He testifies to what he has seen and heard, but no one accepts his testimony.
JOHN|3|33|The man who has accepted it has certified that God is truthful.
JOHN|3|34|For the one whom God has sent speaks the words of God, for God gives the Spirit without limit.
JOHN|3|35|The Father loves the Son and has placed everything in his hands.
JOHN|3|36|Whoever believes in the Son has eternal life, but whoever rejects the Son will not see life, for God's wrath remains on him."
JOHN|4|1|The Pharisees heard that Jesus was gaining and baptizing more disciples than John,
JOHN|4|2|although in fact it was not Jesus who baptized, but his disciples.
JOHN|4|3|When the Lord learned of this, he left Judea and went back once more to Galilee.
JOHN|4|4|Now he had to go through Samaria.
JOHN|4|5|So he came to a town in Samaria called Sychar, near the plot of ground Jacob had given to his son Joseph.
JOHN|4|6|Jacob's well was there, and Jesus, tired as he was from the journey, sat down by the well. It was about the sixth hour.
JOHN|4|7|When a Samaritan woman came to draw water, Jesus said to her, "Will you give me a drink?"
JOHN|4|8|(His disciples had gone into the town to buy food.)
JOHN|4|9|The Samaritan woman said to him, "You are a Jew and I am a Samaritan woman. How can you ask me for a drink?" (For Jews do not associate with Samaritans. )
JOHN|4|10|Jesus answered her, "If you knew the gift of God and who it is that asks you for a drink, you would have asked him and he would have given you living water."
JOHN|4|11|"Sir," the woman said, "you have nothing to draw with and the well is deep. Where can you get this living water?
JOHN|4|12|Are you greater than our father Jacob, who gave us the well and drank from it himself, as did also his sons and his flocks and herds?"
JOHN|4|13|Jesus answered, "Everyone who drinks this water will be thirsty again,
JOHN|4|14|but whoever drinks the water I give him will never thirst. Indeed, the water I give him will become in him a spring of water welling up to eternal life."
JOHN|4|15|The woman said to him, "Sir, give me this water so that I won't get thirsty and have to keep coming here to draw water."
JOHN|4|16|He told her, "Go, call your husband and come back."
JOHN|4|17|"I have no husband," she replied.
JOHN|4|18|Jesus said to her, "You are right when you say you have no husband. The fact is, you have had five husbands, and the man you now have is not your husband. What you have just said is quite true."
JOHN|4|19|"Sir," the woman said, "I can see that you are a prophet.
JOHN|4|20|Our fathers worshiped on this mountain, but you Jews claim that the place where we must worship is in Jerusalem."
JOHN|4|21|Jesus declared, "Believe me, woman, a time is coming when you will worship the Father neither on this mountain nor in Jerusalem.
JOHN|4|22|You Samaritans worship what you do not know; we worship what we do know, for salvation is from the Jews.
JOHN|4|23|Yet a time is coming and has now come when the true worshipers will worship the Father in spirit and truth, for they are the kind of worshipers the Father seeks.
JOHN|4|24|God is spirit, and his worshipers must worship in spirit and in truth."
JOHN|4|25|The woman said, "I know that Messiah" (called Christ) "is coming. When he comes, he will explain everything to us."
JOHN|4|26|Then Jesus declared, "I who speak to you am he."
JOHN|4|27|Just then his disciples returned and were surprised to find him talking with a woman. But no one asked, "What do you want?" or "Why are you talking with her?"
JOHN|4|28|Then, leaving her water jar, the woman went back to the town and said to the people,
JOHN|4|29|"Come, see a man who told me everything I ever did. Could this be the Christ?"
JOHN|4|30|They came out of the town and made their way toward him.
JOHN|4|31|Meanwhile his disciples urged him, "Rabbi, eat something."
JOHN|4|32|But he said to them, "I have food to eat that you know nothing about."
JOHN|4|33|Then his disciples said to each other, "Could someone have brought him food?"
JOHN|4|34|"My food," said Jesus, "is to do the will of him who sent me and to finish his work.
JOHN|4|35|Do you not say, 'Four months more and then the harvest'? I tell you, open your eyes and look at the fields! They are ripe for harvest.
JOHN|4|36|Even now the reaper draws his wages, even now he harvests the crop for eternal life, so that the sower and the reaper may be glad together.
JOHN|4|37|Thus the saying 'One sows and another reaps' is true.
JOHN|4|38|I sent you to reap what you have not worked for. Others have done the hard work, and you have reaped the benefits of their labor."
JOHN|4|39|Many of the Samaritans from that town believed in him because of the woman's testimony, "He told me everything I ever did."
JOHN|4|40|So when the Samaritans came to him, they urged him to stay with them, and he stayed two days.
JOHN|4|41|And because of his words many more became believers.
JOHN|4|42|They said to the woman, "We no longer believe just because of what you said; now we have heard for ourselves, and we know that this man really is the Savior of the world."
JOHN|4|43|After the two days he left for Galilee.
JOHN|4|44|(Now Jesus himself had pointed out that a prophet has no honor in his own country.)
JOHN|4|45|When he arrived in Galilee, the Galileans welcomed him. They had seen all that he had done in Jerusalem at the Passover Feast, for they also had been there.
JOHN|4|46|Once more he visited Cana in Galilee, where he had turned the water into wine. And there was a certain royal official whose son lay sick at Capernaum.
JOHN|4|47|When this man heard that Jesus had arrived in Galilee from Judea, he went to him and begged him to come and heal his son, who was close to death.
JOHN|4|48|"Unless you people see miraculous signs and wonders," Jesus told him, "you will never believe."
JOHN|4|49|The royal official said, "Sir, come down before my child dies."
JOHN|4|50|Jesus replied, "You may go. Your son will live." The man took Jesus at his word and departed.
JOHN|4|51|While he was still on the way, his servants met him with the news that his boy was living.
JOHN|4|52|When he inquired as to the time when his son got better, they said to him, "The fever left him yesterday at the seventh hour."
JOHN|4|53|Then the father realized that this was the exact time at which Jesus had said to him, "Your son will live." So he and all his household believed.
JOHN|4|54|This was the second miraculous sign that Jesus performed, having come from Judea to Galilee.
JOHN|5|1|Some time later, Jesus went up to Jerusalem for a feast of the Jews.
JOHN|5|2|Now there is in Jerusalem near the Sheep Gate a pool, which in Aramaic is called Bethesda and which is surrounded by five covered colonnades.
JOHN|5|3|Here a great number of disabled people used to lie--the blind, the lame, the paralyzed.
JOHN|5|4|See Footnote
JOHN|5|5|One who was there had been an invalid for thirty-eight years.
JOHN|5|6|When Jesus saw him lying there and learned that he had been in this condition for a long time, he asked him, "Do you want to get well?"
JOHN|5|7|"Sir," the invalid replied, "I have no one to help me into the pool when the water is stirred. While I am trying to get in, someone else goes down ahead of me."
JOHN|5|8|Then Jesus said to him, "Get up! Pick up your mat and walk."
JOHN|5|9|At once the man was cured; he picked up his mat and walked. The day on which this took place was a Sabbath,
JOHN|5|10|and so the Jews said to the man who had been healed, "It is the Sabbath; the law forbids you to carry your mat."
JOHN|5|11|But he replied, "The man who made me well said to me, 'Pick up your mat and walk.'"
JOHN|5|12|So they asked him, "Who is this fellow who told you to pick it up and walk?"
JOHN|5|13|The man who was healed had no idea who it was, for Jesus had slipped away into the crowd that was there.
JOHN|5|14|Later Jesus found him at the temple and said to him, "See, you are well again. Stop sinning or something worse may happen to you."
JOHN|5|15|The man went away and told the Jews that it was Jesus who had made him well.
JOHN|5|16|So, because Jesus was doing these things on the Sabbath, the Jews persecuted him.
JOHN|5|17|Jesus said to them, "My Father is always at his work to this very day, and I, too, am working."
JOHN|5|18|For this reason the Jews tried all the harder to kill him; not only was he breaking the Sabbath, but he was even calling God his own Father, making himself equal with God.
JOHN|5|19|Jesus gave them this answer: "I tell you the truth, the Son can do nothing by himself; he can do only what he sees his Father doing, because whatever the Father does the Son also does.
JOHN|5|20|For the Father loves the Son and shows him all he does. Yes, to your amazement he will show him even greater things than these.
JOHN|5|21|For just as the Father raises the dead and gives them life, even so the Son gives life to whom he is pleased to give it.
JOHN|5|22|Moreover, the Father judges no one, but has entrusted all judgment to the Son,
JOHN|5|23|that all may honor the Son just as they honor the Father. He who does not honor the Son does not honor the Father, who sent him.
JOHN|5|24|"I tell you the truth, whoever hears my word and believes him who sent me has eternal life and will not be condemned; he has crossed over from death to life.
JOHN|5|25|I tell you the truth, a time is coming and has now come when the dead will hear the voice of the Son of God and those who hear will live.
JOHN|5|26|For as the Father has life in himself, so he has granted the Son to have life in himself.
JOHN|5|27|And he has given him authority to judge because he is the Son of Man.
JOHN|5|28|"Do not be amazed at this, for a time is coming when all who are in their graves will hear his voice
JOHN|5|29|and come out--those who have done good will rise to live, and those who have done evil will rise to be condemned.
JOHN|5|30|By myself I can do nothing; I judge only as I hear, and my judgment is just, for I seek not to please myself but him who sent me.
JOHN|5|31|"If I testify about myself, my testimony is not valid.
JOHN|5|32|There is another who testifies in my favor, and I know that his testimony about me is valid.
JOHN|5|33|"You have sent to John and he has testified to the truth.
JOHN|5|34|Not that I accept human testimony; but I mention it that you may be saved.
JOHN|5|35|John was a lamp that burned and gave light, and you chose for a time to enjoy his light.
JOHN|5|36|"I have testimony weightier than that of John. For the very work that the Father has given me to finish, and which I am doing, testifies that the Father has sent me.
JOHN|5|37|And the Father who sent me has himself testified concerning me. You have never heard his voice nor seen his form,
JOHN|5|38|nor does his word dwell in you, for you do not believe the one he sent.
JOHN|5|39|You diligently study the Scriptures because you think that by them you possess eternal life. These are the Scriptures that testify about me,
JOHN|5|40|yet you refuse to come to me to have life.
JOHN|5|41|"I do not accept praise from men,
JOHN|5|42|but I know you. I know that you do not have the love of God in your hearts.
JOHN|5|43|I have come in my Father's name, and you do not accept me; but if someone else comes in his own name, you will accept him.
JOHN|5|44|How can you believe if you accept praise from one another, yet make no effort to obtain the praise that comes from the only God?
JOHN|5|45|"But do not think I will accuse you before the Father. Your accuser is Moses, on whom your hopes are set.
JOHN|5|46|If you believed Moses, you would believe me, for he wrote about me.
JOHN|5|47|But since you do not believe what he wrote, how are you going to believe what I say?"
JOHN|6|1|Some time after this, Jesus crossed to the far shore of the Sea of Galilee (that is, the Sea of Tiberias),
JOHN|6|2|and a great crowd of people followed him because they saw the miraculous signs he had performed on the sick.
JOHN|6|3|Then Jesus went up on a mountainside and sat down with his disciples.
JOHN|6|4|The Jewish Passover Feast was near.
JOHN|6|5|When Jesus looked up and saw a great crowd coming toward him, he said to Philip, "Where shall we buy bread for these people to eat?"
JOHN|6|6|He asked this only to test him, for he already had in mind what he was going to do.
JOHN|6|7|Philip answered him, "Eight months' wages would not buy enough bread for each one to have a bite!"
JOHN|6|8|Another of his disciples, Andrew, Simon Peter's brother, spoke up,
JOHN|6|9|"Here is a boy with five small barley loaves and two small fish, but how far will they go among so many?"
JOHN|6|10|Jesus said, "Have the people sit down." There was plenty of grass in that place, and the men sat down, about five thousand of them.
JOHN|6|11|Jesus then took the loaves, gave thanks, and distributed to those who were seated as much as they wanted. He did the same with the fish.
JOHN|6|12|When they had all had enough to eat, he said to his disciples, "Gather the pieces that are left over. Let nothing be wasted."
JOHN|6|13|So they gathered them and filled twelve baskets with the pieces of the five barley loaves left over by those who had eaten.
JOHN|6|14|After the people saw the miraculous sign that Jesus did, they began to say, "Surely this is the Prophet who is to come into the world."
JOHN|6|15|Jesus, knowing that they intended to come and make him king by force, withdrew again to a mountain by himself.
JOHN|6|16|When evening came, his disciples went down to the lake,
JOHN|6|17|where they got into a boat and set off across the lake for Capernaum. By now it was dark, and Jesus had not yet joined them.
JOHN|6|18|A strong wind was blowing and the waters grew rough.
JOHN|6|19|When they had rowed three or three and a half miles, they saw Jesus approaching the boat, walking on the water; and they were terrified.
JOHN|6|20|But he said to them, "It is I; don't be afraid."
JOHN|6|21|Then they were willing to take him into the boat, and immediately the boat reached the shore where they were heading.
JOHN|6|22|The next day the crowd that had stayed on the opposite shore of the lake realized that only one boat had been there, and that Jesus had not entered it with his disciples, but that they had gone away alone.
JOHN|6|23|Then some boats from Tiberias landed near the place where the people had eaten the bread after the Lord had given thanks.
JOHN|6|24|Once the crowd realized that neither Jesus nor his disciples were there, they got into the boats and went to Capernaum in search of Jesus.
JOHN|6|25|When they found him on the other side of the lake, they asked him, "Rabbi, when did you get here?"
JOHN|6|26|Jesus answered, "I tell you the truth, you are looking for me, not because you saw miraculous signs but because you ate the loaves and had your fill.
JOHN|6|27|Do not work for food that spoils, but for food that endures to eternal life, which the Son of Man will give you. On him God the Father has placed his seal of approval."
JOHN|6|28|Then they asked him, "What must we do to do the works God requires?"
JOHN|6|29|Jesus answered, "The work of God is this: to believe in the one he has sent."
JOHN|6|30|So they asked him, "What miraculous sign then will you give that we may see it and believe you? What will you do?
JOHN|6|31|Our forefathers ate the manna in the desert; as it is written: 'He gave them bread from heaven to eat.'"
JOHN|6|32|Jesus said to them, "I tell you the truth, it is not Moses who has given you the bread from heaven, but it is my Father who gives you the true bread from heaven.
JOHN|6|33|For the bread of God is he who comes down from heaven and gives life to the world."
JOHN|6|34|"Sir," they said, "from now on give us this bread."
JOHN|6|35|Then Jesus declared, "I am the bread of life. He who comes to me will never go hungry, and he who believes in me will never be thirsty.
JOHN|6|36|But as I told you, you have seen me and still you do not believe.
JOHN|6|37|All that the Father gives me will come to me, and whoever comes to me I will never drive away.
JOHN|6|38|For I have come down from heaven not to do my will but to do the will of him who sent me.
JOHN|6|39|And this is the will of him who sent me, that I shall lose none of all that he has given me, but raise them up at the last day.
JOHN|6|40|For my Father's will is that everyone who looks to the Son and believes in him shall have eternal life, and I will raise him up at the last day."
JOHN|6|41|At this the Jews began to grumble about him because he said, "I am the bread that came down from heaven."
JOHN|6|42|They said, "Is this not Jesus, the son of Joseph, whose father and mother we know? How can he now say, 'I came down from heaven'?"
JOHN|6|43|"Stop grumbling among yourselves," Jesus answered.
JOHN|6|44|"No one can come to me unless the Father who sent me draws him, and I will raise him up at the last day.
JOHN|6|45|It is written in the Prophets: 'They will all be taught by God.' Everyone who listens to the Father and learns from him comes to me.
JOHN|6|46|No one has seen the Father except the one who is from God; only he has seen the Father.
JOHN|6|47|I tell you the truth, he who believes has everlasting life.
JOHN|6|48|I am the bread of life.
JOHN|6|49|Your forefathers ate the manna in the desert, yet they died.
JOHN|6|50|But here is the bread that comes down from heaven, which a man may eat and not die.
JOHN|6|51|I am the living bread that came down from heaven. If anyone eats of this bread, he will live forever. This bread is my flesh, which I will give for the life of the world."
JOHN|6|52|Then the Jews began to argue sharply among themselves, "How can this man give us his flesh to eat?"
JOHN|6|53|Jesus said to them, "I tell you the truth, unless you eat the flesh of the Son of Man and drink his blood, you have no life in you.
JOHN|6|54|Whoever eats my flesh and drinks my blood has eternal life, and I will raise him up at the last day.
JOHN|6|55|For my flesh is real food and my blood is real drink.
JOHN|6|56|Whoever eats my flesh and drinks my blood remains in me, and I in him.
JOHN|6|57|Just as the living Father sent me and I live because of the Father, so the one who feeds on me will live because of me.
JOHN|6|58|This is the bread that came down from heaven. Your forefathers ate manna and died, but he who feeds on this bread will live forever."
JOHN|6|59|He said this while teaching in the synagogue in Capernaum.
JOHN|6|60|On hearing it, many of his disciples said, "This is a hard teaching. Who can accept it?"
JOHN|6|61|Aware that his disciples were grumbling about this, Jesus said to them, "Does this offend you?
JOHN|6|62|What if you see the Son of Man ascend to where he was before!
JOHN|6|63|The Spirit gives life; the flesh counts for nothing. The words I have spoken to you are spirit and they are life.
JOHN|6|64|Yet there are some of you who do not believe." For Jesus had known from the beginning which of them did not believe and who would betray him.
JOHN|6|65|He went on to say, "This is why I told you that no one can come to me unless the Father has enabled him."
JOHN|6|66|From this time many of his disciples turned back and no longer followed him.
JOHN|6|67|"You do not want to leave too, do you?" Jesus asked the Twelve.
JOHN|6|68|Simon Peter answered him, "Lord, to whom shall we go? You have the words of eternal life.
JOHN|6|69|We believe and know that you are the Holy One of God."
JOHN|6|70|Then Jesus replied, "Have I not chosen you, the Twelve? Yet one of you is a devil!"
JOHN|6|71|(He meant Judas, the son of Simon Iscariot, who, though one of the Twelve, was later to betray him.)
JOHN|7|1|After this, Jesus went around in Galilee, purposely staying away from Judea because the Jews there were waiting to take his life.
JOHN|7|2|But when the Jewish Feast of Tabernacles was near,
JOHN|7|3|Jesus' brothers said to him, "You ought to leave here and go to Judea, so that your disciples may see the miracles you do.
JOHN|7|4|No one who wants to become a public figure acts in secret. Since you are doing these things, show yourself to the world."
JOHN|7|5|For even his own brothers did not believe in him.
JOHN|7|6|Therefore Jesus told them, "The right time for me has not yet come; for you any time is right.
JOHN|7|7|The world cannot hate you, but it hates me because I testify that what it does is evil.
JOHN|7|8|You go to the Feast. I am not yet going up to this Feast, because for me the right time has not yet come."
JOHN|7|9|Having said this, he stayed in Galilee.
JOHN|7|10|However, after his brothers had left for the Feast, he went also, not publicly, but in secret.
JOHN|7|11|Now at the Feast the Jews were watching for him and asking, "Where is that man?"
JOHN|7|12|Among the crowds there was widespread whispering about him. Some said, "He is a good man."
JOHN|7|13|Others replied, "No, he deceives the people." But no one would say anything publicly about him for fear of the Jews.
JOHN|7|14|Not until halfway through the Feast did Jesus go up to the temple courts and begin to teach.
JOHN|7|15|The Jews were amazed and asked, "How did this man get such learning without having studied?"
JOHN|7|16|Jesus answered, "My teaching is not my own. It comes from him who sent me.
JOHN|7|17|If anyone chooses to do God's will, he will find out whether my teaching comes from God or whether I speak on my own.
JOHN|7|18|He who speaks on his own does so to gain honor for himself, but he who works for the honor of the one who sent him is a man of truth; there is nothing false about him.
JOHN|7|19|Has not Moses given you the law? Yet not one of you keeps the law. Why are you trying to kill me?"
JOHN|7|20|"You are demon-possessed," the crowd answered. "Who is trying to kill you?"
JOHN|7|21|Jesus said to them, "I did one miracle, and you are all astonished.
JOHN|7|22|Yet, because Moses gave you circumcision (though actually it did not come from Moses, but from the patriarchs), you circumcise a child on the Sabbath.
JOHN|7|23|Now if a child can be circumcised on the Sabbath so that the law of Moses may not be broken, why are you angry with me for healing the whole man on the Sabbath?
JOHN|7|24|Stop judging by mere appearances, and make a right judgment."
JOHN|7|25|At that point some of the people of Jerusalem began to ask, "Isn't this the man they are trying to kill?
JOHN|7|26|Here he is, speaking publicly, and they are not saying a word to him. Have the authorities really concluded that he is the Christ?
JOHN|7|27|But we know where this man is from; when the Christ comes, no one will know where he is from."
JOHN|7|28|Then Jesus, still teaching in the temple courts, cried out, "Yes, you know me, and you know where I am from. I am not here on my own, but he who sent me is true. You do not know him,
JOHN|7|29|but I know him because I am from him and he sent me."
JOHN|7|30|At this they tried to seize him, but no one laid a hand on him, because his time had not yet come.
JOHN|7|31|Still, many in the crowd put their faith in him. They said, "When the Christ comes, will he do more miraculous signs than this man?"
JOHN|7|32|The Pharisees heard the crowd whispering such things about him. Then the chief priests and the Pharisees sent temple guards to arrest him.
JOHN|7|33|Jesus said, "I am with you for only a short time, and then I go to the one who sent me.
JOHN|7|34|You will look for me, but you will not find me; and where I am, you cannot come."
JOHN|7|35|The Jews said to one another, "Where does this man intend to go that we cannot find him? Will he go where our people live scattered among the Greeks, and teach the Greeks?
JOHN|7|36|What did he mean when he said, 'You will look for me, but you will not find me,' and 'Where I am, you cannot come'?"
JOHN|7|37|On the last and greatest day of the Feast, Jesus stood and said in a loud voice, "If anyone is thirsty, let him come to me and drink.
JOHN|7|38|Whoever believes in me, as the Scripture has said, streams of living water will flow from within him."
JOHN|7|39|By this he meant the Spirit, whom those who believed in him were later to receive. Up to that time the Spirit had not been given, since Jesus had not yet been glorified.
JOHN|7|40|On hearing his words, some of the people said, "Surely this man is the Prophet."
JOHN|7|41|Others said, "He is the Christ."
JOHN|7|42|Still others asked, "How can the Christ come from Galilee? Does not the Scripture say that the Christ will come from David's family and from Bethlehem, the town where David lived?"
JOHN|7|43|Thus the people were divided because of Jesus.
JOHN|7|44|Some wanted to seize him, but no one laid a hand on him.
JOHN|7|45|Finally the temple guards went back to the chief priests and Pharisees, who asked them, "Why didn't you bring him in?"
JOHN|7|46|"No one ever spoke the way this man does," the guards declared.
JOHN|7|47|"You mean he has deceived you also?" the Pharisees retorted.
JOHN|7|48|"Has any of the rulers or of the Pharisees believed in him?
JOHN|7|49|No! But this mob that knows nothing of the law--there is a curse on them."
JOHN|7|50|Nicodemus, who had gone to Jesus earlier and who was one of their own number, asked,
JOHN|7|51|"Does our law condemn anyone without first hearing him to find out what he is doing?"
JOHN|7|52|They replied, "Are you from Galilee, too? Look into it, and you will find that a prophet does not come out of Galilee."
JOHN|7|53|Then each went to his own home.
JOHN|8|1|But Jesus went to the Mount of Olives.
JOHN|8|2|At dawn he appeared again in the temple courts, where all the people gathered around him, and he sat down to teach them.
JOHN|8|3|The teachers of the law and the Pharisees brought in a woman caught in adultery. They made her stand before the group
JOHN|8|4|and said to Jesus, "Teacher, this woman was caught in the act of adultery.
JOHN|8|5|In the Law Moses commanded us to stone such women. Now what do you say?"
JOHN|8|6|They were using this question as a trap, in order to have a basis for accusing him.
JOHN|8|7|But Jesus bent down and started to write on the ground with his finger. When they kept on questioning him, he straightened up and said to them, "If any one of you is without sin, let him be the first to throw a stone at her."
JOHN|8|8|Again he stooped down and wrote on the ground.
JOHN|8|9|At this, those who heard began to go away one at a time, the older ones first, until only Jesus was left, with the woman still standing there.
JOHN|8|10|Jesus straightened up and asked her, "Woman, where are they? Has no one condemned you?"
JOHN|8|11|"No one, sir," she said. "Then neither do I condemn you," Jesus declared. "Go now and leave your life of sin."
JOHN|8|12|When Jesus spoke again to the people, he said, "I am the light of the world. Whoever follows me will never walk in darkness, but will have the light of life."
JOHN|8|13|The Pharisees challenged him, "Here you are, appearing as your own witness; your testimony is not valid."
JOHN|8|14|Jesus answered, "Even if I testify on my own behalf, my testimony is valid, for I know where I came from and where I am going. But you have no idea where I come from or where I am going.
JOHN|8|15|You judge by human standards; I pass judgment on no one.
JOHN|8|16|But if I do judge, my decisions are right, because I am not alone. I stand with the Father, who sent me.
JOHN|8|17|In your own Law it is written that the testimony of two men is valid.
JOHN|8|18|I am one who testifies for myself; my other witness is the Father, who sent me."
JOHN|8|19|Then they asked him, "Where is your father?"
JOHN|8|20|"You do not know me or my Father," Jesus replied. "If you knew me, you would know my Father also." He spoke these words while teaching in the temple area near the place where the offerings were put. Yet no one seized him, because his time had not yet come.
JOHN|8|21|Once more Jesus said to them, "I am going away, and you will look for me, and you will die in your sin. Where I go, you cannot come."
JOHN|8|22|This made the Jews ask, "Will he kill himself? Is that why he says, 'Where I go, you cannot come'?"
JOHN|8|23|But he continued, "You are from below; I am from above. You are of this world; I am not of this world.
JOHN|8|24|I told you that you would die in your sins; if you do not believe that I am the one I claim to be, you will indeed die in your sins."
JOHN|8|25|"Who are you?" they asked.
JOHN|8|26|"Just what I have been claiming all along," Jesus replied. "I have much to say in judgment of you. But he who sent me is reliable, and what I have heard from him I tell the world."
JOHN|8|27|They did not understand that he was telling them about his Father.
JOHN|8|28|So Jesus said, "When you have lifted up the Son of Man, then you will know that I am the one I claim to be and that I do nothing on my own but speak just what the Father has taught me.
JOHN|8|29|The one who sent me is with me; he has not left me alone, for I always do what pleases him."
JOHN|8|30|Even as he spoke, many put their faith in him.
JOHN|8|31|To the Jews who had believed him, Jesus said, "If you hold to my teaching, you are really my disciples.
JOHN|8|32|Then you will know the truth, and the truth will set you free."
JOHN|8|33|They answered him, "We are Abraham's descendants and have never been slaves of anyone. How can you say that we shall be set free?"
JOHN|8|34|Jesus replied, "I tell you the truth, everyone who sins is a slave to sin.
JOHN|8|35|Now a slave has no permanent place in the family, but a son belongs to it forever.
JOHN|8|36|So if the Son sets you free, you will be free indeed.
JOHN|8|37|I know you are Abraham's descendants. Yet you are ready to kill me, because you have no room for my word.
JOHN|8|38|I am telling you what I have seen in the Father's presence, and you do what you have heard from your father. "
JOHN|8|39|"Abraham is our father," they answered. "If you were Abraham's children," said Jesus, "then you would
JOHN|8|40|do the things Abraham did. As it is, you are determined to kill me, a man who has told you the truth that I heard from God. Abraham did not do such things.
JOHN|8|41|You are doing the things your own father does.We are not illegitimate children," they protested. "The only Father we have is God himself."
JOHN|8|42|Jesus said to them, "If God were your Father, you would love me, for I came from God and now am here. I have not come on my own; but he sent me.
JOHN|8|43|Why is my language not clear to you? Because you are unable to hear what I say.
JOHN|8|44|You belong to your father, the devil, and you want to carry out your father's desire. He was a murderer from the beginning, not holding to the truth, for there is no truth in him. When he lies, he speaks his native language, for he is a liar and the father of lies.
JOHN|8|45|Yet because I tell the truth, you do not believe me!
JOHN|8|46|Can any of you prove me guilty of sin? If I am telling the truth, why don't you believe me?
JOHN|8|47|He who belongs to God hears what God says. The reason you do not hear is that you do not belong to God."
JOHN|8|48|The Jews answered him, "Aren't we right in saying that you are a Samaritan and demon-possessed?"
JOHN|8|49|"I am not possessed by a demon," said Jesus, "but I honor my Father and you dishonor me.
JOHN|8|50|I am not seeking glory for myself; but there is one who seeks it, and he is the judge.
JOHN|8|51|I tell you the truth, if anyone keeps my word, he will never see death."
JOHN|8|52|At this the Jews exclaimed, "Now we know that you are demon-possessed! Abraham died and so did the prophets, yet you say that if anyone keeps your word, he will never taste death.
JOHN|8|53|Are you greater than our father Abraham? He died, and so did the prophets. Who do you think you are?"
JOHN|8|54|Jesus replied, "If I glorify myself, my glory means nothing. My Father, whom you claim as your God, is the one who glorifies me.
JOHN|8|55|Though you do not know him, I know him. If I said I did not, I would be a liar like you, but I do know him and keep his word.
JOHN|8|56|Your father Abraham rejoiced at the thought of seeing my day; he saw it and was glad."
JOHN|8|57|"You are not yet fifty years old," the Jews said to him, "and you have seen Abraham!"
JOHN|8|58|"I tell you the truth," Jesus answered, "before Abraham was born, I am!"
JOHN|8|59|At this, they picked up stones to stone him, but Jesus hid himself, slipping away from the temple grounds.
JOHN|9|1|As he went along, he saw a man blind from birth.
JOHN|9|2|His disciples asked him, "Rabbi, who sinned, this man or his parents, that he was born blind?"
JOHN|9|3|"Neither this man nor his parents sinned," said Jesus, "but this happened so that the work of God might be displayed in his life.
JOHN|9|4|As long as it is day, we must do the work of him who sent me. Night is coming, when no one can work.
JOHN|9|5|While I am in the world, I am the light of the world."
JOHN|9|6|Having said this, he spit on the ground, made some mud with the saliva, and put it on the man's eyes.
JOHN|9|7|"Go," he told him, "wash in the Pool of Siloam" (this word means Sent). So the man went and washed, and came home seeing.
JOHN|9|8|His neighbors and those who had formerly seen him begging asked, "Isn't this the same man who used to sit and beg?"
JOHN|9|9|Some claimed that he was. Others said, "No, he only looks like him." But he himself insisted, "I am the man."
JOHN|9|10|"How then were your eyes opened?" they demanded.
JOHN|9|11|He replied, "The man they call Jesus made some mud and put it on my eyes. He told me to go to Siloam and wash. So I went and washed, and then I could see."
JOHN|9|12|"Where is this man?" they asked him. "I don't know," he said.
JOHN|9|13|They brought to the Pharisees the man who had been blind.
JOHN|9|14|Now the day on which Jesus had made the mud and opened the man's eyes was a Sabbath.
JOHN|9|15|Therefore the Pharisees also asked him how he had received his sight. "He put mud on my eyes," the man replied, "and I washed, and now I see."
JOHN|9|16|Some of the Pharisees said, "This man is not from God, for he does not keep the Sabbath." But others asked, "How can a sinner do such miraculous signs?" So they were divided.
JOHN|9|17|Finally they turned again to the blind man, "What have you to say about him? It was your eyes he opened." The man replied, "He is a prophet."
JOHN|9|18|The Jews still did not believe that he had been blind and had received his sight until they sent for the man's parents.
JOHN|9|19|"Is this your son?" they asked. "Is this the one you say was born blind? How is it that now he can see?"
JOHN|9|20|"We know he is our son," the parents answered, "and we know he was born blind.
JOHN|9|21|But how he can see now, or who opened his eyes, we don't know. Ask him. He is of age; he will speak for himself."
JOHN|9|22|His parents said this because they were afraid of the Jews, for already the Jews had decided that anyone who acknowledged that Jesus was the Christ would be put out of the synagogue.
JOHN|9|23|That was why his parents said, "He is of age; ask him."
JOHN|9|24|A second time they summoned the man who had been blind. "Give glory to God, "they said. "We know this man is a sinner."
JOHN|9|25|He replied, "Whether he is a sinner or not, I don't know. One thing I do know. I was blind but now I see!"
JOHN|9|26|Then they asked him, "What did he do to you? How did he open your eyes?"
JOHN|9|27|He answered, "I have told you already and you did not listen. Why do you want to hear it again? Do you want to become his disciples, too?"
JOHN|9|28|Then they hurled insults at him and said, "You are this fellow's disciple! We are disciples of Moses!
JOHN|9|29|We know that God spoke to Moses, but as for this fellow, we don't even know where he comes from."
JOHN|9|30|The man answered, "Now that is remarkable! You don't know where he comes from, yet he opened my eyes.
JOHN|9|31|We know that God does not listen to sinners. He listens to the godly man who does his will.
JOHN|9|32|Nobody has ever heard of opening the eyes of a man born blind.
JOHN|9|33|If this man were not from God, he could do nothing."
JOHN|9|34|To this they replied, "You were steeped in sin at birth; how dare you lecture us!" And they threw him out.
JOHN|9|35|Jesus heard that they had thrown him out, and when he found him, he said, "Do you believe in the Son of Man?"
JOHN|9|36|"Who is he, sir?" the man asked. "Tell me so that I may believe in him."
JOHN|9|37|Jesus said, "You have now seen him; in fact, he is the one speaking with you."
JOHN|9|38|Then the man said, "Lord, I believe," and he worshiped him.
JOHN|9|39|Jesus said, "For judgment I have come into this world, so that the blind will see and those who see will become blind."
JOHN|9|40|Some Pharisees who were with him heard him say this and asked, "What? Are we blind too?"
JOHN|9|41|Jesus said, "If you were blind, you would not be guilty of sin; but now that you claim you can see, your guilt remains.
JOHN|10|1|"I tell you the truth, the man who does not enter the sheep pen by the gate, but climbs in by some other way, is a thief and a robber.
JOHN|10|2|The man who enters by the gate is the shepherd of his sheep.
JOHN|10|3|The watchman opens the gate for him, and the sheep listen to his voice. He calls his own sheep by name and leads them out.
JOHN|10|4|When he has brought out all his own, he goes on ahead of them, and his sheep follow him because they know his voice.
JOHN|10|5|But they will never follow a stranger; in fact, they will run away from him because they do not recognize a stranger's voice."
JOHN|10|6|Jesus used this figure of speech, but they did not understand what he was telling them.
JOHN|10|7|Therefore Jesus said again, "I tell you the truth, I am the gate for the sheep.
JOHN|10|8|All who ever came before me were thieves and robbers, but the sheep did not listen to them.
JOHN|10|9|I am the gate; whoever enters through me will be saved. He will come in and go out, and find pasture.
JOHN|10|10|The thief comes only to steal and kill and destroy; I have come that they may have life, and have it to the full.
JOHN|10|11|"I am the good shepherd. The good shepherd lays down his life for the sheep.
JOHN|10|12|The hired hand is not the shepherd who owns the sheep. So when he sees the wolf coming, he abandons the sheep and runs away. Then the wolf attacks the flock and scatters it.
JOHN|10|13|The man runs away because he is a hired hand and cares nothing for the sheep.
JOHN|10|14|"I am the good shepherd; I know my sheep and my sheep know me--
JOHN|10|15|just as the Father knows me and I know the Father--and I lay down my life for the sheep.
JOHN|10|16|I have other sheep that are not of this sheep pen. I must bring them also. They too will listen to my voice, and there shall be one flock and one shepherd.
JOHN|10|17|The reason my Father loves me is that I lay down my life--only to take it up again.
JOHN|10|18|No one takes it from me, but I lay it down of my own accord. I have authority to lay it down and authority to take it up again. This command I received from my Father."
JOHN|10|19|At these words the Jews were again divided.
JOHN|10|20|Many of them said, "He is demon-possessed and raving mad. Why listen to him?"
JOHN|10|21|But others said, "These are not the sayings of a man possessed by a demon. Can a demon open the eyes of the blind?"
JOHN|10|22|Then came the Feast of Dedication at Jerusalem. It was winter,
JOHN|10|23|and Jesus was in the temple area walking in Solomon's Colonnade.
JOHN|10|24|The Jews gathered around him, saying, "How long will you keep us in suspense? If you are the Christ, tell us plainly."
JOHN|10|25|Jesus answered, "I did tell you, but you do not believe. The miracles I do in my Father's name speak for me,
JOHN|10|26|but you do not believe because you are not my sheep.
JOHN|10|27|My sheep listen to my voice; I know them, and they follow me.
JOHN|10|28|I give them eternal life, and they shall never perish; no one can snatch them out of my hand.
JOHN|10|29|My Father, who has given them to me, is greater than all; no one can snatch them out of my Father's hand.
JOHN|10|30|I and the Father are one."
JOHN|10|31|Again the Jews picked up stones to stone him,
JOHN|10|32|but Jesus said to them, "I have shown you many great miracles from the Father. For which of these do you stone me?"
JOHN|10|33|"We are not stoning you for any of these," replied the Jews, "but for blasphemy, because you, a mere man, claim to be God."
JOHN|10|34|Jesus answered them, "Is it not written in your Law, 'I have said you are gods'?
JOHN|10|35|If he called them 'gods,' to whom the word of God came--and the Scripture cannot be broken--
JOHN|10|36|what about the one whom the Father set apart as his very own and sent into the world? Why then do you accuse me of blasphemy because I said, 'I am God's Son'?
JOHN|10|37|Do not believe me unless I do what my Father does.
JOHN|10|38|But if I do it, even though you do not believe me, believe the miracles, that you may know and understand that the Father is in me, and I in the Father."
JOHN|10|39|Again they tried to seize him, but he escaped their grasp.
JOHN|10|40|Then Jesus went back across the Jordan to the place where John had been baptizing in the early days. Here he stayed
JOHN|10|41|and many people came to him. They said, "Though John never performed a miraculous sign, all that John said about this man was true."
JOHN|10|42|And in that place many believed in Jesus.
JOHN|11|1|Now a man named Lazarus was sick. He was from Bethany, the village of Mary and her sister Martha.
JOHN|11|2|This Mary, whose brother Lazarus now lay sick, was the same one who poured perfume on the Lord and wiped his feet with her hair.
JOHN|11|3|So the sisters sent word to Jesus, "Lord, the one you love is sick."
JOHN|11|4|When he heard this, Jesus said, "This sickness will not end in death. No, it is for God's glory so that God's Son may be glorified through it."
JOHN|11|5|Jesus loved Martha and her sister and Lazarus.
JOHN|11|6|Yet when he heard that Lazarus was sick, he stayed where he was two more days.
JOHN|11|7|Then he said to his disciples, "Let us go back to Judea."
JOHN|11|8|"But Rabbi," they said, "a short while ago the Jews tried to stone you, and yet you are going back there?"
JOHN|11|9|Jesus answered, "Are there not twelve hours of daylight? A man who walks by day will not stumble, for he sees by this world's light.
JOHN|11|10|It is when he walks by night that he stumbles, for he has no light."
JOHN|11|11|After he had said this, he went on to tell them, "Our friend Lazarus has fallen asleep; but I am going there to wake him up."
JOHN|11|12|His disciples replied, "Lord, if he sleeps, he will get better."
JOHN|11|13|Jesus had been speaking of his death, but his disciples thought he meant natural sleep.
JOHN|11|14|So then he told them plainly, "Lazarus is dead,
JOHN|11|15|and for your sake I am glad I was not there, so that you may believe. But let us go to him."
JOHN|11|16|Then Thomas (called Didymus) said to the rest of the disciples, "Let us also go, that we may die with him."
JOHN|11|17|On his arrival, Jesus found that Lazarus had already been in the tomb for four days.
JOHN|11|18|Bethany was less than two miles from Jerusalem,
JOHN|11|19|and many Jews had come to Martha and Mary to comfort them in the loss of their brother.
JOHN|11|20|When Martha heard that Jesus was coming, she went out to meet him, but Mary stayed at home.
JOHN|11|21|"Lord," Martha said to Jesus, "if you had been here, my brother would not have died.
JOHN|11|22|But I know that even now God will give you whatever you ask."
JOHN|11|23|Jesus said to her, "Your brother will rise again."
JOHN|11|24|Martha answered, "I know he will rise again in the resurrection at the last day."
JOHN|11|25|Jesus said to her, "I am the resurrection and the life. He who believes in me will live, even though he dies;
JOHN|11|26|and whoever lives and believes in me will never die. Do you believe this?"
JOHN|11|27|"Yes, Lord," she told him, "I believe that you are the Christ, the Son of God, who was to come into the world."
JOHN|11|28|And after she had said this, she went back and called her sister Mary aside. "The Teacher is here," she said, "and is asking for you."
JOHN|11|29|When Mary heard this, she got up quickly and went to him.
JOHN|11|30|Now Jesus had not yet entered the village, but was still at the place where Martha had met him.
JOHN|11|31|When the Jews who had been with Mary in the house, comforting her, noticed how quickly she got up and went out, they followed her, supposing she was going to the tomb to mourn there.
JOHN|11|32|When Mary reached the place where Jesus was and saw him, she fell at his feet and said, "Lord, if you had been here, my brother would not have died."
JOHN|11|33|When Jesus saw her weeping, and the Jews who had come along with her also weeping, he was deeply moved in spirit and troubled.
JOHN|11|34|"Where have you laid him?" he asked. "Come and see, Lord," they replied.
JOHN|11|35|Jesus wept.
JOHN|11|36|Then the Jews said, "See how he loved him!"
JOHN|11|37|But some of them said, "Could not he who opened the eyes of the blind man have kept this man from dying?"
JOHN|11|38|Jesus, once more deeply moved, came to the tomb. It was a cave with a stone laid across the entrance.
JOHN|11|39|"Take away the stone," he said. "But, Lord," said Martha, the sister of the dead man, "by this time there is a bad odor, for he has been there four days."
JOHN|11|40|Then Jesus said, "Did I not tell you that if you believed, you would see the glory of God?"
JOHN|11|41|So they took away the stone. Then Jesus looked up and said, "Father, I thank you that you have heard me.
JOHN|11|42|I knew that you always hear me, but I said this for the benefit of the people standing here, that they may believe that you sent me."
JOHN|11|43|When he had said this, Jesus called in a loud voice, "Lazarus, come out!"
JOHN|11|44|The dead man came out, his hands and feet wrapped with strips of linen, and a cloth around his face. Jesus said to them, "Take off the grave clothes and let him go."
JOHN|11|45|Therefore many of the Jews who had come to visit Mary, and had seen what Jesus did, put their faith in him.
JOHN|11|46|But some of them went to the Pharisees and told them what Jesus had done.
JOHN|11|47|Then the chief priests and the Pharisees called a meeting of the Sanhedrin.
JOHN|11|48|"What are we accomplishing?" they asked. "Here is this man performing many miraculous signs. If we let him go on like this, everyone will believe in him, and then the Romans will come and take away both our place and our nation."
JOHN|11|49|Then one of them, named Caiaphas, who was high priest that year, spoke up, "You know nothing at all!
JOHN|11|50|You do not realize that it is better for you that one man die for the people than that the whole nation perish."
JOHN|11|51|He did not say this on his own, but as high priest that year he prophesied that Jesus would die for the Jewish nation,
JOHN|11|52|and not only for that nation but also for the scattered children of God, to bring them together and make them one.
JOHN|11|53|So from that day on they plotted to take his life.
JOHN|11|54|Therefore Jesus no longer moved about publicly among the Jews. Instead he withdrew to a region near the desert, to a village called Ephraim, where he stayed with his disciples.
JOHN|11|55|When it was almost time for the Jewish Passover, many went up from the country to Jerusalem for their ceremonial cleansing before the Passover.
JOHN|11|56|They kept looking for Jesus, and as they stood in the temple area they asked one another, "What do you think? Isn't he coming to the Feast at all?"
JOHN|11|57|But the chief priests and Pharisees had given orders that if anyone found out where Jesus was, he should report it so that they might arrest him.
JOHN|12|1|Six days before the Passover, Jesus arrived at Bethany, where Lazarus lived, whom Jesus had raised from the dead.
JOHN|12|2|Here a dinner was given in Jesus' honor. Martha served, while Lazarus was among those reclining at the table with him.
JOHN|12|3|Then Mary took about a pint of pure nard, an expensive perfume; she poured it on Jesus' feet and wiped his feet with her hair. And the house was filled with the fragrance of the perfume.
JOHN|12|4|But one of his disciples, Judas Iscariot, who was later to betray him, objected,
JOHN|12|5|"Why wasn't this perfume sold and the money given to the poor? It was worth a year's wages. "
JOHN|12|6|He did not say this because he cared about the poor but because he was a thief; as keeper of the money bag, he used to help himself to what was put into it.
JOHN|12|7|"Leave her alone," Jesus replied. "It was intended that she should save this perfume for the day of my burial.
JOHN|12|8|You will always have the poor among you, but you will not always have me."
JOHN|12|9|Meanwhile a large crowd of Jews found out that Jesus was there and came, not only because of him but also to see Lazarus, whom he had raised from the dead.
JOHN|12|10|So the chief priests made plans to kill Lazarus as well,
JOHN|12|11|for on account of him many of the Jews were going over to Jesus and putting their faith in him.
JOHN|12|12|The next day the great crowd that had come for the Feast heard that Jesus was on his way to Jerusalem.
JOHN|12|13|They took palm branches and went out to meet him, shouting, "Hosanna! Blessed is he who comes in the name of the Lord!Blessed is the King of Israel!"
JOHN|12|14|Jesus found a young donkey and sat upon it, as it is written,
JOHN|12|15|"Do not be afraid, O Daughter of Zion; see, your king is coming, seated on a donkey's colt."
JOHN|12|16|At first his disciples did not understand all this. Only after Jesus was glorified did they realize that these things had been written about him and that they had done these things to him.
JOHN|12|17|Now the crowd that was with him when he called Lazarus from the tomb and raised him from the dead continued to spread the word.
JOHN|12|18|Many people, because they had heard that he had given this miraculous sign, went out to meet him.
JOHN|12|19|So the Pharisees said to one another, "See, this is getting us nowhere. Look how the whole world has gone after him!"
JOHN|12|20|Now there were some Greeks among those who went up to worship at the Feast.
JOHN|12|21|They came to Philip, who was from Bethsaida in Galilee, with a request. "Sir," they said, "we would like to see Jesus."
JOHN|12|22|Philip went to tell Andrew; Andrew and Philip in turn told Jesus.
JOHN|12|23|Jesus replied, "The hour has come for the Son of Man to be glorified.
JOHN|12|24|I tell you the truth, unless a kernel of wheat falls to the ground and dies, it remains only a single seed. But if it dies, it produces many seeds.
JOHN|12|25|The man who loves his life will lose it, while the man who hates his life in this world will keep it for eternal life.
JOHN|12|26|Whoever serves me must follow me; and where I am, my servant also will be. My Father will honor the one who serves me.
JOHN|12|27|"Now my heart is troubled, and what shall I say? 'Father, save me from this hour'? No, it was for this very reason I came to this hour.
JOHN|12|28|Father, glorify your name!"
JOHN|12|29|Then a voice came from heaven, "I have glorified it, and will glorify it again." The crowd that was there and heard it said it had thundered; others said an angel had spoken to him.
JOHN|12|30|Jesus said, "This voice was for your benefit, not mine.
JOHN|12|31|Now is the time for judgment on this world; now the prince of this world will be driven out.
JOHN|12|32|But I, when I am lifted up from the earth, will draw all men to myself."
JOHN|12|33|He said this to show the kind of death he was going to die.
JOHN|12|34|The crowd spoke up, "We have heard from the Law that the Christ will remain forever, so how can you say, 'The Son of Man must be lifted up'? Who is this 'Son of Man'?"
JOHN|12|35|Then Jesus told them, "You are going to have the light just a little while longer. Walk while you have the light, before darkness overtakes you. The man who walks in the dark does not know where he is going.
JOHN|12|36|Put your trust in the light while you have it, so that you may become sons of light." When he had finished speaking, Jesus left and hid himself from them.
JOHN|12|37|Even after Jesus had done all these miraculous signs in their presence, they still would not believe in him.
JOHN|12|38|This was to fulfill the word of Isaiah the prophet: "Lord, who has believed our message and to whom has the arm of the Lord been revealed?"
JOHN|12|39|For this reason they could not believe, because, as Isaiah says elsewhere:
JOHN|12|40|"He has blinded their eyes and deadened their hearts, so they can neither see with their eyes, nor understand with their hearts, nor turn--and I would heal them."
JOHN|12|41|Isaiah said this because he saw Jesus' glory and spoke about him.
JOHN|12|42|Yet at the same time many even among the leaders believed in him. But because of the Pharisees they would not confess their faith for fear they would be put out of the synagogue;
JOHN|12|43|for they loved praise from men more than praise from God.
JOHN|12|44|Then Jesus cried out, "When a man believes in me, he does not believe in me only, but in the one who sent me.
JOHN|12|45|When he looks at me, he sees the one who sent me.
JOHN|12|46|I have come into the world as a light, so that no one who believes in me should stay in darkness.
JOHN|12|47|"As for the person who hears my words but does not keep them, I do not judge him. For I did not come to judge the world, but to save it.
JOHN|12|48|There is a judge for the one who rejects me and does not accept my words; that very word which I spoke will condemn him at the last day.
JOHN|12|49|For I did not speak of my own accord, but the Father who sent me commanded me what to say and how to say it.
JOHN|12|50|I know that his command leads to eternal life. So whatever I say is just what the Father has told me to say."
JOHN|13|1|It was just before the Passover Feast. Jesus knew that the time had come for him to leave this world and go to the Father. Having loved his own who were in the world, he now showed them the full extent of his love.
JOHN|13|2|The evening meal was being served, and the devil had already prompted Judas Iscariot, son of Simon, to betray Jesus.
JOHN|13|3|Jesus knew that the Father had put all things under his power, and that he had come from God and was returning to God;
JOHN|13|4|so he got up from the meal, took off his outer clothing, and wrapped a towel around his waist.
JOHN|13|5|After that, he poured water into a basin and began to wash his disciples' feet, drying them with the towel that was wrapped around him.
JOHN|13|6|He came to Simon Peter, who said to him, "Lord, are you going to wash my feet?"
JOHN|13|7|Jesus replied, "You do not realize now what I am doing, but later you will understand."
JOHN|13|8|"No," said Peter, "you shall never wash my feet." Jesus answered, "Unless I wash you, you have no part with me."
JOHN|13|9|"Then, Lord," Simon Peter replied, "not just my feet but my hands and my head as well!"
JOHN|13|10|Jesus answered, "A person who has had a bath needs only to wash his feet; his whole body is clean. And you are clean, though not every one of you."
JOHN|13|11|For he knew who was going to betray him, and that was why he said not every one was clean.
JOHN|13|12|When he had finished washing their feet, he put on his clothes and returned to his place. "Do you understand what I have done for you?" he asked them.
JOHN|13|13|"You call me 'Teacher' and 'Lord,' and rightly so, for that is what I am.
JOHN|13|14|Now that I, your Lord and Teacher, have washed your feet, you also should wash one another's feet.
JOHN|13|15|I have set you an example that you should do as I have done for you.
JOHN|13|16|I tell you the truth, no servant is greater than his master, nor is a messenger greater than the one who sent him.
JOHN|13|17|Now that you know these things, you will be blessed if you do them.
JOHN|13|18|"I am not referring to all of you; I know those I have chosen. But this is to fulfill the scripture: 'He who shares my bread has lifted up his heel against me.'
JOHN|13|19|"I am telling you now before it happens, so that when it does happen you will believe that I am He.
JOHN|13|20|I tell you the truth, whoever accepts anyone I send accepts me; and whoever accepts me accepts the one who sent me."
JOHN|13|21|After he had said this, Jesus was troubled in spirit and testified, "I tell you the truth, one of you is going to betray me."
JOHN|13|22|His disciples stared at one another, at a loss to know which of them he meant.
JOHN|13|23|One of them, the disciple whom Jesus loved, was reclining next to him.
JOHN|13|24|Simon Peter motioned to this disciple and said, "Ask him which one he means."
JOHN|13|25|Leaning back against Jesus, he asked him, "Lord, who is it?"
JOHN|13|26|Jesus answered, "It is the one to whom I will give this piece of bread when I have dipped it in the dish." Then, dipping the piece of bread, he gave it to Judas Iscariot, son of Simon.
JOHN|13|27|As soon as Judas took the bread, Satan entered into him.
JOHN|13|28|"What you are about to do, do quickly," Jesus told him, but no one at the meal understood why Jesus said this to him.
JOHN|13|29|Since Judas had charge of the money, some thought Jesus was telling him to buy what was needed for the Feast, or to give something to the poor.
JOHN|13|30|As soon as Judas had taken the bread, he went out. And it was night.
JOHN|13|31|When he was gone, Jesus said, "Now is the Son of Man glorified and God is glorified in him.
JOHN|13|32|If God is glorified in him, God will glorify the Son in himself, and will glorify him at once.
JOHN|13|33|"My children, I will be with you only a little longer. You will look for me, and just as I told the Jews, so I tell you now: Where I am going, you cannot come.
JOHN|13|34|"A new command I give you: Love one another. As I have loved you, so you must love one another.
JOHN|13|35|By this all men will know that you are my disciples, if you love one another."
JOHN|13|36|Simon Peter asked him, "Lord, where are you going?" Jesus replied, "Where I am going, you cannot follow now, but you will follow later."
JOHN|13|37|Peter asked, "Lord, why can't I follow you now? I will lay down my life for you."
JOHN|13|38|Then Jesus answered, "Will you really lay down your life for me? I tell you the truth, before the rooster crows, you will disown me three times!
JOHN|14|1|"Do not let your hearts be troubled. Trust in God; trust also in me.
JOHN|14|2|In my Father's house are many rooms; if it were not so, I would have told you. I am going there to prepare a place for you.
JOHN|14|3|And if I go and prepare a place for you, I will come back and take you to be with me that you also may be where I am.
JOHN|14|4|You know the way to the place where I am going."
JOHN|14|5|Thomas said to him, "Lord, we don't know where you are going, so how can we know the way?"
JOHN|14|6|Jesus answered, "I am the way and the truth and the life. No one comes to the Father except through me.
JOHN|14|7|If you really knew me, you would know my Father as well. From now on, you do know him and have seen him."
JOHN|14|8|Philip said, "Lord, show us the Father and that will be enough for us."
JOHN|14|9|Jesus answered: "Don't you know me, Philip, even after I have been among you such a long time? Anyone who has seen me has seen the Father. How can you say, 'Show us the Father'?
JOHN|14|10|Don't you believe that I am in the Father, and that the Father is in me? The words I say to you are not just my own. Rather, it is the Father, living in me, who is doing his work.
JOHN|14|11|Believe me when I say that I am in the Father and the Father is in me; or at least believe on the evidence of the miracles themselves.
JOHN|14|12|I tell you the truth, anyone who has faith in me will do what I have been doing. He will do even greater things than these, because I am going to the Father.
JOHN|14|13|And I will do whatever you ask in my name, so that the Son may bring glory to the Father.
JOHN|14|14|You may ask me for anything in my name, and I will do it.
JOHN|14|15|"If you love me, you will obey what I command.
JOHN|14|16|And I will ask the Father, and he will give you another Counselor to be with you forever--
JOHN|14|17|the Spirit of truth. The world cannot accept him, because it neither sees him nor knows him. But you know him, for he lives with you and will be in you.
JOHN|14|18|I will not leave you as orphans; I will come to you.
JOHN|14|19|Before long, the world will not see me anymore, but you will see me. Because I live, you also will live.
JOHN|14|20|On that day you will realize that I am in my Father, and you are in me, and I am in you.
JOHN|14|21|Whoever has my commands and obeys them, he is the one who loves me. He who loves me will be loved by my Father, and I too will love him and show myself to him."
JOHN|14|22|Then Judas (not Judas Iscariot) said, "But, Lord, why do you intend to show yourself to us and not to the world?"
JOHN|14|23|Jesus replied, "If anyone loves me, he will obey my teaching. My Father will love him, and we will come to him and make our home with him.
JOHN|14|24|He who does not love me will not obey my teaching. These words you hear are not my own; they belong to the Father who sent me.
JOHN|14|25|"All this I have spoken while still with you.
JOHN|14|26|But the Counselor, the Holy Spirit, whom the Father will send in my name, will teach you all things and will remind you of everything I have said to you.
JOHN|14|27|Peace I leave with you; my peace I give you. I do not give to you as the world gives. Do not let your hearts be troubled and do not be afraid.
JOHN|14|28|"You heard me say, 'I am going away and I am coming back to you.' If you loved me, you would be glad that I am going to the Father, for the Father is greater than I.
JOHN|14|29|I have told you now before it happens, so that when it does happen you will believe.
JOHN|14|30|I will not speak with you much longer, for the prince of this world is coming. He has no hold on me,
JOHN|14|31|but the world must learn that I love the Father and that I do exactly what my Father has commanded me. "Come now; let us leave.
JOHN|15|1|"I am the true vine, and my Father is the gardener.
JOHN|15|2|He cuts off every branch in me that bears no fruit, while every branch that does bear fruit he prunes so that it will be even more fruitful.
JOHN|15|3|You are already clean because of the word I have spoken to you.
JOHN|15|4|Remain in me, and I will remain in you. No branch can bear fruit by itself; it must remain in the vine. Neither can you bear fruit unless you remain in me.
JOHN|15|5|"I am the vine; you are the branches. If a man remains in me and I in him, he will bear much fruit; apart from me you can do nothing.
JOHN|15|6|If anyone does not remain in me, he is like a branch that is thrown away and withers; such branches are picked up, thrown into the fire and burned.
JOHN|15|7|If you remain in me and my words remain in you, ask whatever you wish, and it will be given you.
JOHN|15|8|This is to my Father's glory, that you bear much fruit, showing yourselves to be my disciples.
JOHN|15|9|"As the Father has loved me, so have I loved you. Now remain in my love.
JOHN|15|10|If you obey my commands, you will remain in my love, just as I have obeyed my Father's commands and remain in his love.
JOHN|15|11|I have told you this so that my joy may be in you and that your joy may be complete.
JOHN|15|12|My command is this: Love each other as I have loved you.
JOHN|15|13|Greater love has no one than this, that he lay down his life for his friends.
JOHN|15|14|You are my friends if you do what I command.
JOHN|15|15|I no longer call you servants, because a servant does not know his master's business. Instead, I have called you friends, for everything that I learned from my Father I have made known to you.
JOHN|15|16|You did not choose me, but I chose you and appointed you to go and bear fruit--fruit that will last. Then the Father will give you whatever you ask in my name.
JOHN|15|17|This is my command: Love each other.
JOHN|15|18|"If the world hates you, keep in mind that it hated me first.
JOHN|15|19|If you belonged to the world, it would love you as its own. As it is, you do not belong to the world, but I have chosen you out of the world. That is why the world hates you.
JOHN|15|20|Remember the words I spoke to you: 'No servant is greater than his master.' If they persecuted me, they will persecute you also. If they obeyed my teaching, they will obey yours also.
JOHN|15|21|They will treat you this way because of my name, for they do not know the One who sent me.
JOHN|15|22|If I had not come and spoken to them, they would not be guilty of sin. Now, however, they have no excuse for their sin.
JOHN|15|23|He who hates me hates my Father as well.
JOHN|15|24|If I had not done among them what no one else did, they would not be guilty of sin. But now they have seen these miracles, and yet they have hated both me and my Father.
JOHN|15|25|But this is to fulfill what is written in their Law: 'They hated me without reason.'
JOHN|15|26|"When the Counselor comes, whom I will send to you from the Father, the Spirit of truth who goes out from the Father, he will testify about me.
JOHN|15|27|And you also must testify, for you have been with me from the beginning.
JOHN|16|1|"All this I have told you so that you will not go astray.
JOHN|16|2|They will put you out of the synagogue; in fact, a time is coming when anyone who kills you will think he is offering a service to God.
JOHN|16|3|They will do such things because they have not known the Father or me.
JOHN|16|4|I have told you this, so that when the time comes you will remember that I warned you. I did not tell you this at first because I was with you.
JOHN|16|5|"Now I am going to him who sent me, yet none of you asks me, 'Where are you going?'
JOHN|16|6|Because I have said these things, you are filled with grief.
JOHN|16|7|But I tell you the truth: It is for your good that I am going away. Unless I go away, the Counselor will not come to you; but if I go, I will send him to you.
JOHN|16|8|When he comes, he will convict the world of guilt in regard to sin and righteousness and judgment:
JOHN|16|9|in regard to sin, because men do not believe in me;
JOHN|16|10|in regard to righteousness, because I am going to the Father, where you can see me no longer;
JOHN|16|11|and in regard to judgment, because the prince of this world now stands condemned.
JOHN|16|12|"I have much more to say to you, more than you can now bear.
JOHN|16|13|But when he, the Spirit of truth, comes, he will guide you into all truth. He will not speak on his own; he will speak only what he hears, and he will tell you what is yet to come.
JOHN|16|14|He will bring glory to me by taking from what is mine and making it known to you.
JOHN|16|15|All that belongs to the Father is mine. That is why I said the Spirit will take from what is mine and make it known to you.
JOHN|16|16|"In a little while you will see me no more, and then after a little while you will see me."
JOHN|16|17|Some of his disciples said to one another, "What does he mean by saying, 'In a little while you will see me no more, and then after a little while you will see me,' and 'Because I am going to the Father'?"
JOHN|16|18|They kept asking, "What does he mean by 'a little while'? We don't understand what he is saying."
JOHN|16|19|Jesus saw that they wanted to ask him about this, so he said to them, "Are you asking one another what I meant when I said, 'In a little while you will see me no more, and then after a little while you will see me'?
JOHN|16|20|I tell you the truth, you will weep and mourn while the world rejoices. You will grieve, but your grief will turn to joy.
JOHN|16|21|A woman giving birth to a child has pain because her time has come; but when her baby is born she forgets the anguish because of her joy that a child is born into the world.
JOHN|16|22|So with you: Now is your time of grief, but I will see you again and you will rejoice, and no one will take away your joy.
JOHN|16|23|In that day you will no longer ask me anything. I tell you the truth, my Father will give you whatever you ask in my name.
JOHN|16|24|Until now you have not asked for anything in my name. Ask and you will receive, and your joy will be complete.
JOHN|16|25|"Though I have been speaking figuratively, a time is coming when I will no longer use this kind of language but will tell you plainly about my Father.
JOHN|16|26|In that day you will ask in my name. I am not saying that I will ask the Father on your behalf.
JOHN|16|27|No, the Father himself loves you because you have loved me and have believed that I came from God.
JOHN|16|28|I came from the Father and entered the world; now I am leaving the world and going back to the Father."
JOHN|16|29|Then Jesus' disciples said, "Now you are speaking clearly and without figures of speech.
JOHN|16|30|Now we can see that you know all things and that you do not even need to have anyone ask you questions. This makes us believe that you came from God."
JOHN|16|31|"You believe at last!" Jesus answered.
JOHN|16|32|"But a time is coming, and has come, when you will be scattered, each to his own home. You will leave me all alone. Yet I am not alone, for my Father is with me.
JOHN|16|33|"I have told you these things, so that in me you may have peace. In this world you will have trouble. But take heart! I have overcome the world."
JOHN|17|1|After Jesus said this, he looked toward heaven and prayed:
JOHN|17|2|"Father, the time has come. Glorify your Son, that your Son may glorify you. For you granted him authority over all people that he might give eternal life to all those you have given him.
JOHN|17|3|Now this is eternal life: that they may know you, the only true God, and Jesus Christ, whom you have sent.
JOHN|17|4|I have brought you glory on earth by completing the work you gave me to do.
JOHN|17|5|And now, Father, glorify me in your presence with the glory I had with you before the world began.
JOHN|17|6|"I have revealed you to those whom you gave me out of the world. They were yours; you gave them to me and they have obeyed your word.
JOHN|17|7|Now they know that everything you have given me comes from you.
JOHN|17|8|For I gave them the words you gave me and they accepted them. They knew with certainty that I came from you, and they believed that you sent me.
JOHN|17|9|I pray for them. I am not praying for the world, but for those you have given me, for they are yours.
JOHN|17|10|All I have is yours, and all you have is mine. And glory has come to me through them.
JOHN|17|11|I will remain in the world no longer, but they are still in the world, and I am coming to you. Holy Father, protect them by the power of your name--the name you gave me--so that they may be one as we are one.
JOHN|17|12|While I was with them, I protected them and kept them safe by that name you gave me. None has been lost except the one doomed to destruction so that Scripture would be fulfilled.
JOHN|17|13|"I am coming to you now, but I say these things while I am still in the world, so that they may have the full measure of my joy within them.
JOHN|17|14|I have given them your word and the world has hated them, for they are not of the world any more than I am of the world.
JOHN|17|15|My prayer is not that you take them out of the world but that you protect them from the evil one.
JOHN|17|16|They are not of the world, even as I am not of it.
JOHN|17|17|Sanctify them by the truth; your word is truth.
JOHN|17|18|As you sent me into the world, I have sent them into the world.
JOHN|17|19|For them I sanctify myself, that they too may be truly sanctified.
JOHN|17|20|"My prayer is not for them alone. I pray also for those who will believe in me through their message,
JOHN|17|21|that all of them may be one, Father, just as you are in me and I am in you. May they also be in us so that the world may believe that you have sent me.
JOHN|17|22|I have given them the glory that you gave me, that they may be one as we are one:
JOHN|17|23|I in them and you in me. May they be brought to complete unity to let the world know that you sent me and have loved them even as you have loved me.
JOHN|17|24|"Father, I want those you have given me to be with me where I am, and to see my glory, the glory you have given me because you loved me before the creation of the world.
JOHN|17|25|"Righteous Father, though the world does not know you, I know you, and they know that you have sent me.
JOHN|17|26|I have made you known to them, and will continue to make you known in order that the love you have for me may be in them and that I myself may be in them."
JOHN|18|1|When he had finished praying, Jesus left with his disciples and crossed the Kidron Valley. On the other side there was an olive grove, and he and his disciples went into it.
JOHN|18|2|Now Judas, who betrayed him, knew the place, because Jesus had often met there with his disciples.
JOHN|18|3|So Judas came to the grove, guiding a detachment of soldiers and some officials from the chief priests and Pharisees. They were carrying torches, lanterns and weapons.
JOHN|18|4|Jesus, knowing all that was going to happen to him, went out and asked them, "Who is it you want?"
JOHN|18|5|"Jesus of Nazareth," they replied.
JOHN|18|6|"I am he," Jesus said. (And Judas the traitor was standing there with them.) When Jesus said, "I am he," they drew back and fell to the ground.
JOHN|18|7|Again he asked them, "Who is it you want?" And they said, "Jesus of Nazareth."
JOHN|18|8|"I told you that I am he," Jesus answered. "If you are looking for me, then let these men go."
JOHN|18|9|This happened so that the words he had spoken would be fulfilled: "I have not lost one of those you gave me."
JOHN|18|10|Then Simon Peter, who had a sword, drew it and struck the high priest's servant, cutting off his right ear. (The servant's name was Malchus.)
JOHN|18|11|Jesus commanded Peter, "Put your sword away! Shall I not drink the cup the Father has given me?"
JOHN|18|12|Then the detachment of soldiers with its commander and the Jewish officials arrested Jesus. They bound him
JOHN|18|13|and brought him first to Annas, who was the father-in-law of Caiaphas, the high priest that year.
JOHN|18|14|Caiaphas was the one who had advised the Jews that it would be good if one man died for the people.
JOHN|18|15|Simon Peter and another disciple were following Jesus. Because this disciple was known to the high priest, he went with Jesus into the high priest's courtyard,
JOHN|18|16|but Peter had to wait outside at the door. The other disciple, who was known to the high priest, came back, spoke to the girl on duty there and brought Peter in.
JOHN|18|17|"You are not one of his disciples, are you?" the girl at the door asked Peter. He replied, "I am not."
JOHN|18|18|It was cold, and the servants and officials stood around a fire they had made to keep warm. Peter also was standing with them, warming himself.
JOHN|18|19|Meanwhile, the high priest questioned Jesus about his disciples and his teaching.
JOHN|18|20|"I have spoken openly to the world," Jesus replied. "I always taught in synagogues or at the temple, where all the Jews come together. I said nothing in secret.
JOHN|18|21|Why question me? Ask those who heard me. Surely they know what I said."
JOHN|18|22|When Jesus said this, one of the officials nearby struck him in the face. "Is this the way you answer the high priest?" he demanded.
JOHN|18|23|"If I said something wrong," Jesus replied, "testify as to what is wrong. But if I spoke the truth, why did you strike me?"
JOHN|18|24|Then Annas sent him, still bound, to Caiaphas the high priest.
JOHN|18|25|As Simon Peter stood warming himself, he was asked, "You are not one of his disciples, are you?" He denied it, saying, "I am not."
JOHN|18|26|One of the high priest's servants, a relative of the man whose ear Peter had cut off, challenged him, "Didn't I see you with him in the olive grove?"
JOHN|18|27|Again Peter denied it, and at that moment a rooster began to crow.
JOHN|18|28|Then the Jews led Jesus from Caiaphas to the palace of the Roman governor. By now it was early morning, and to avoid ceremonial uncleanness the Jews did not enter the palace; they wanted to be able to eat the Passover.
JOHN|18|29|So Pilate came out to them and asked, "What charges are you bringing against this man?"
JOHN|18|30|"If he were not a criminal," they replied, "we would not have handed him over to you."
JOHN|18|31|Pilate said, "Take him yourselves and judge him by your own law."
JOHN|18|32|"But we have no right to execute anyone," the Jews objected. This happened so that the words Jesus had spoken indicating the kind of death he was going to die would be fulfilled.
JOHN|18|33|Pilate then went back inside the palace, summoned Jesus and asked him, "Are you the king of the Jews?"
JOHN|18|34|"Is that your own idea," Jesus asked, "or did others talk to you about me?"
JOHN|18|35|"Am I a Jew?" Pilate replied. "It was your people and your chief priests who handed you over to me. What is it you have done?"
JOHN|18|36|Jesus said, "My kingdom is not of this world. If it were, my servants would fight to prevent my arrest by the Jews. But now my kingdom is from another place."
JOHN|18|37|"You are a king, then!" said Pilate. Jesus answered, "You are right in saying I am a king. In fact, for this reason I was born, and for this I came into the world, to testify to the truth. Everyone on the side of truth listens to me."
JOHN|18|38|"What is truth?" Pilate asked. With this he went out again to the Jews and said, "I find no basis for a charge against him.
JOHN|18|39|But it is your custom for me to release to you one prisoner at the time of the Passover. Do you want me to release 'the king of the Jews'?"
JOHN|18|40|They shouted back, "No, not him! Give us Barabbas!" Now Barabbas had taken part in a rebellion.
JOHN|19|1|Then Pilate took Jesus and had him flogged.
JOHN|19|2|The soldiers twisted together a crown of thorns and put it on his head. They clothed him in a purple robe
JOHN|19|3|and went up to him again and again, saying, "Hail, king of the Jews!" And they struck him in the face.
JOHN|19|4|Once more Pilate came out and said to the Jews, "Look, I am bringing him out to you to let you know that I find no basis for a charge against him."
JOHN|19|5|When Jesus came out wearing the crown of thorns and the purple robe, Pilate said to them, "Here is the man!"
JOHN|19|6|As soon as the chief priests and their officials saw him, they shouted, "Crucify! Crucify!" But Pilate answered, "You take him and crucify him. As for me, I find no basis for a charge against him."
JOHN|19|7|The Jews insisted, "We have a law, and according to that law he must die, because he claimed to be the Son of God."
JOHN|19|8|When Pilate heard this, he was even more afraid,
JOHN|19|9|and he went back inside the palace. "Where do you come from?" he asked Jesus, but Jesus gave him no answer.
JOHN|19|10|"Do you refuse to speak to me?" Pilate said. "Don't you realize I have power either to free you or to crucify you?"
JOHN|19|11|Jesus answered, "You would have no power over me if it were not given to you from above. Therefore the one who handed me over to you is guilty of a greater sin."
JOHN|19|12|From then on, Pilate tried to set Jesus free, but the Jews kept shouting, "If you let this man go, you are no friend of Caesar. Anyone who claims to be a king opposes Caesar."
JOHN|19|13|When Pilate heard this, he brought Jesus out and sat down on the judge's seat at a place known as the Stone Pavement (which in Aramaic is Gabbatha).
JOHN|19|14|It was the day of Preparation of Passover Week, about the sixth hour. "Here is your king," Pilate said to the Jews.
JOHN|19|15|But they shouted, "Take him away! Take him away! Crucify him!Shall I crucify your king?" Pilate asked. "We have no king but Caesar," the chief priests answered.
JOHN|19|16|Finally Pilate handed him over to them to be crucified.
JOHN|19|17|So the soldiers took charge of Jesus. Carrying his own cross, he went out to the place of the Skull (which in Aramaic is called Golgotha).
JOHN|19|18|Here they crucified him, and with him two others--one on each side and Jesus in the middle.
JOHN|19|19|Pilate had a notice prepared and fastened to the cross. It read:|sc JESUS OF NAZARETH, THE KING OF THE JEWS.
JOHN|19|20|Many of the Jews read this sign, for the place where Jesus was crucified was near the city, and the sign was written in Aramaic, Latin and Greek.
JOHN|19|21|The chief priests of the Jews protested to Pilate, "Do not write 'The King of the Jews,' but that this man claimed to be king of the Jews."
JOHN|19|22|Pilate answered, "What I have written, I have written."
JOHN|19|23|When the soldiers crucified Jesus, they took his clothes, dividing them into four shares, one for each of them, with the undergarment remaining. This garment was seamless, woven in one piece from top to bottom.
JOHN|19|24|"Let's not tear it," they said to one another. "Let's decide by lot who will get it." This happened that the scripture might be fulfilled which said, "They divided my garments among them and cast lots for my clothing." So this is what the soldiers did.
JOHN|19|25|Near the cross of Jesus stood his mother, his mother's sister, Mary the wife of Clopas, and Mary Magdalene.
JOHN|19|26|When Jesus saw his mother there, and the disciple whom he loved standing nearby, he said to his mother, "Dear woman, here is your son,"
JOHN|19|27|and to the disciple, "Here is your mother." From that time on, this disciple took her into his home.
JOHN|19|28|Later, knowing that all was now completed, and so that the Scripture would be fulfilled, Jesus said, "I am thirsty."
JOHN|19|29|A jar of wine vinegar was there, so they soaked a sponge in it, put the sponge on a stalk of the hyssop plant, and lifted it to Jesus' lips.
JOHN|19|30|When he had received the drink, Jesus said, "It is finished." With that, he bowed his head and gave up his spirit.
JOHN|19|31|Now it was the day of Preparation, and the next day was to be a special Sabbath. Because the Jews did not want the bodies left on the crosses during the Sabbath, they asked Pilate to have the legs broken and the bodies taken down.
JOHN|19|32|The soldiers therefore came and broke the legs of the first man who had been crucified with Jesus, and then those of the other.
JOHN|19|33|But when they came to Jesus and found that he was already dead, they did not break his legs.
JOHN|19|34|Instead, one of the soldiers pierced Jesus' side with a spear, bringing a sudden flow of blood and water.
JOHN|19|35|The man who saw it has given testimony, and his testimony is true. He knows that he tells the truth, and he testifies so that you also may believe.
JOHN|19|36|These things happened so that the scripture would be fulfilled: "Not one of his bones will be broken,"
JOHN|19|37|and, as another scripture says, "They will look on the one they have pierced."
JOHN|19|38|Later, Joseph of Arimathea asked Pilate for the body of Jesus. Now Joseph was a disciple of Jesus, but secretly because he feared the Jews. With Pilate's permission, he came and took the body away.
JOHN|19|39|He was accompanied by Nicodemus, the man who earlier had visited Jesus at night. Nicodemus brought a mixture of myrrh and aloes, about seventy-five pounds.
JOHN|19|40|Taking Jesus' body, the two of them wrapped it, with the spices, in strips of linen. This was in accordance with Jewish burial customs.
JOHN|19|41|At the place where Jesus was crucified, there was a garden, and in the garden a new tomb, in which no one had ever been laid.
JOHN|19|42|Because it was the Jewish day of Preparation and since the tomb was nearby, they laid Jesus there.
JOHN|20|1|Early on the first day of the week, while it was still dark, Mary Magdalene went to the tomb and saw that the stone had been removed from the entrance.
JOHN|20|2|So she came running to Simon Peter and the other disciple, the one Jesus loved, and said, "They have taken the Lord out of the tomb, and we don't know where they have put him!"
JOHN|20|3|So Peter and the other disciple started for the tomb.
JOHN|20|4|Both were running, but the other disciple outran Peter and reached the tomb first.
JOHN|20|5|He bent over and looked in at the strips of linen lying there but did not go in.
JOHN|20|6|Then Simon Peter, who was behind him, arrived and went into the tomb. He saw the strips of linen lying there,
JOHN|20|7|as well as the burial cloth that had been around Jesus' head. The cloth was folded up by itself, separate from the linen.
JOHN|20|8|Finally the other disciple, who had reached the tomb first, also went inside. He saw and believed.
JOHN|20|9|(They still did not understand from Scripture that Jesus had to rise from the dead.)
JOHN|20|10|Then the disciples went back to their homes,
JOHN|20|11|but Mary stood outside the tomb crying. As she wept, she bent over to look into the tomb
JOHN|20|12|and saw two angels in white, seated where Jesus' body had been, one at the head and the other at the foot.
JOHN|20|13|They asked her, "Woman, why are you crying?"
JOHN|20|14|"They have taken my Lord away," she said, "and I don't know where they have put him." At this, she turned around and saw Jesus standing there, but she did not realize that it was Jesus.
JOHN|20|15|"Woman," he said, "why are you crying? Who is it you are looking for?" Thinking he was the gardener, she said, "Sir, if you have carried him away, tell me where you have put him, and I will get him."
JOHN|20|16|Jesus said to her, "Mary." She turned toward him and cried out in Aramaic, "Rabboni!" (which means Teacher).
JOHN|20|17|Jesus said, "Do not hold on to me, for I have not yet returned to the Father. Go instead to my brothers and tell them, 'I am returning to my Father and your Father, to my God and your God.'"
JOHN|20|18|Mary Magdalene went to the disciples with the news: "I have seen the Lord!" And she told them that he had said these things to her.
JOHN|20|19|On the evening of that first day of the week, when the disciples were together, with the doors locked for fear of the Jews, Jesus came and stood among them and said, "Peace be with you!"
JOHN|20|20|After he said this, he showed them his hands and side. The disciples were overjoyed when they saw the Lord.
JOHN|20|21|Again Jesus said, "Peace be with you! As the Father has sent me, I am sending you."
JOHN|20|22|And with that he breathed on them and said, "Receive the Holy Spirit.
JOHN|20|23|If you forgive anyone his sins, they are forgiven; if you do not forgive them, they are not forgiven."
JOHN|20|24|Now Thomas (called Didymus), one of the Twelve, was not with the disciples when Jesus came.
JOHN|20|25|So the other disciples told him, "We have seen the Lord!" But he said to them, "Unless I see the nail marks in his hands and put my finger where the nails were, and put my hand into his side, I will not believe it."
JOHN|20|26|A week later his disciples were in the house again, and Thomas was with them. Though the doors were locked, Jesus came and stood among them and said, "Peace be with you!"
JOHN|20|27|Then he said to Thomas, "Put your finger here; see my hands. Reach out your hand and put it into my side. Stop doubting and believe."
JOHN|20|28|Thomas said to him, "My Lord and my God!"
JOHN|20|29|Then Jesus told him, "Because you have seen me, you have believed; blessed are those who have not seen and yet have believed."
JOHN|20|30|Jesus did many other miraculous signs in the presence of his disciples, which are not recorded in this book.
JOHN|20|31|But these are written that you may believe that Jesus is the Christ, the Son of God, and that by believing you may have life in his name.
JOHN|21|1|Afterward Jesus appeared again to his disciples, by the Sea of Tiberias. It happened this way:
JOHN|21|2|Simon Peter, Thomas (called Didymus), Nathanael from Cana in Galilee, the sons of Zebedee, and two other disciples were together.
JOHN|21|3|"I'm going out to fish," Simon Peter told them, and they said, "We'll go with you." So they went out and got into the boat, but that night they caught nothing.
JOHN|21|4|Early in the morning, Jesus stood on the shore, but the disciples did not realize that it was Jesus.
JOHN|21|5|He called out to them, "Friends, haven't you any fish?No," they answered.
JOHN|21|6|He said, "Throw your net on the right side of the boat and you will find some." When they did, they were unable to haul the net in because of the large number of fish.
JOHN|21|7|Then the disciple whom Jesus loved said to Peter, "It is the Lord!" As soon as Simon Peter heard him say, "It is the Lord," he wrapped his outer garment around him (for he had taken it off) and jumped into the water.
JOHN|21|8|The other disciples followed in the boat, towing the net full of fish, for they were not far from shore, about a hundred yards.
JOHN|21|9|When they landed, they saw a fire of burning coals there with fish on it, and some bread.
JOHN|21|10|Jesus said to them, "Bring some of the fish you have just caught."
JOHN|21|11|Simon Peter climbed aboard and dragged the net ashore. It was full of large fish, 153, but even with so many the net was not torn.
JOHN|21|12|Jesus said to them, "Come and have breakfast." None of the disciples dared ask him, "Who are you?" They knew it was the Lord.
JOHN|21|13|Jesus came, took the bread and gave it to them, and did the same with the fish.
JOHN|21|14|This was now the third time Jesus appeared to his disciples after he was raised from the dead.
JOHN|21|15|When they had finished eating, Jesus said to Simon Peter, "Simon son of John, do you truly love me more than these?Yes, Lord," he said, "you know that I love you." Jesus said, "Feed my lambs."
JOHN|21|16|Again Jesus said, "Simon son of John, do you truly love me?" He answered, "Yes, Lord, you know that I love you." Jesus said, "Take care of my sheep."
JOHN|21|17|The third time he said to him, "Simon son of John, do you love me?" Peter was hurt because Jesus asked him the third time, "Do you love me?" He said, "Lord, you know all things; you know that I love you."
JOHN|21|18|Jesus said, "Feed my sheep. I tell you the truth, when you were younger you dressed yourself and went where you wanted; but when you are old you will stretch out your hands, and someone else will dress you and lead you where you do not want to go."
JOHN|21|19|Jesus said this to indicate the kind of death by which Peter would glorify God. Then he said to him, "Follow me!"
JOHN|21|20|Peter turned and saw that the disciple whom Jesus loved was following them. (This was the one who had leaned back against Jesus at the supper and had said, "Lord, who is going to betray you?")
JOHN|21|21|When Peter saw him, he asked, "Lord, what about him?"
JOHN|21|22|Jesus answered, "If I want him to remain alive until I return, what is that to you? You must follow me."
JOHN|21|23|Because of this, the rumor spread among the brothers that this disciple would not die. But Jesus did not say that he would not die; he only said, "If I want him to remain alive until I return, what is that to you?"
JOHN|21|24|This is the disciple who testifies to these things and who wrote them down. We know that his testimony is true.
JOHN|21|25|Jesus did many other things as well. If every one of them were written down, I suppose that even the whole world would not have room for the books that would be written.
