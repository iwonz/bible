LAM|1|1|ALEPH. Quomodo sedet solacivitas plena populo!Facta est quasi viduadomina gentium;princeps provinciarumfacta est sub tributo.
LAM|1|2|BETH. Plorans plorat in nocte,et lacrimae eius in maxillis eius;non est qui consoletur eamex omnibus caris eius:omnes amici eius spreverunt eamet facti sunt ei inimici.
LAM|1|3|GHIMEL. Migravit Iudas prae afflictioneet multitudine servitutis;habitat inter gentesnec invenit requiem:omnes persecutores eius apprehenderunt eaminter angustias.
LAM|1|4|DALETH. Viae Sion lugent,eo quod non sint qui veniant ad sollemnitatem;omnes portae eius destructae,sacerdotes eius gementes,virgines eius afflictae,et ipsa oppressa amaritudine.
LAM|1|5|HE. Facti sunt hostes eius in caput,inimici eius in securitate,quia Dominus afflixit eampropter multitudinem iniquitatum eius;parvuli eius ducti sunt captiviante faciem tribulantis.
LAM|1|6|VAU. Et egressus est a filia Sionomnis decor eius;facti sunt principes eius velut cervinon invenientes pascuaet abierunt absque fortitudineante faciem persequentis.
LAM|1|7|ZAIN. Recordata est Ierusalemdierum afflictionis suae et peregrinationis,omnium desiderabilium suorum,quae habuerat a diebus antiquis,cum caderet populus eius in manu hostili,et non esset auxiliator;viderunt eam hosteset deriserunt interitum eius.
LAM|1|8|HETH. Peccatum peccavit Ierusalem,propterea abominabilis facta est;omnes, qui glorificabant eam, spreverunt illam,quia viderunt ignominiam eius:ipsa autem gemensconversa est retrorsum.
LAM|1|9|TETH. Sordes eius in fimbriis eius,nec recordata est finis sui;deposita est vehementer,non habens consolatorem. Vide, Domine, afflictionem meam, quoniam erectus est inimicus! ".
LAM|1|10|IOD. Manum suam misit hostisad omnia desiderabilia eius,quia vidit gentesingressas sanctuarium suum,de quibus praeceperas,ne intrarent in ecclesiam tuam.
LAM|1|11|CAPH. Omnis populus eius gemenset quaerens panem;dederunt pretiosa quaeque pro ciboad refocillandam animam. Vide, Domine, et considera,quoniam facta sum vilis!
LAM|1|12|LAMED. O vos omnes, qui transitis per viam,attendite et videte,si est dolor sicut dolor meus,quem paravit mihi,quo afflixit me Dominusin die irae furoris sui.
LAM|1|13|MEM. De excelso misit ignem,in ossa mea immisit eum;expandit rete pedibus meis,convertit me retrorsum:posuit me desolatam,tota die maerore confectam.
LAM|1|14|NUN. Vigilavit super iniquitates meas,in manu eius convolutae suntet impositae collo meo;debilitavit virtutem meam:dedit me Dominus in manu,de qua non potero surgere.
LAM|1|15|SAMECH. Sprevit omnes fortes meosDominus in medio mei;vocavit adversum me conventum,ut contereret iuvenes meos:torcular calcavit Dominusvirgini filiae Iudae.
LAM|1|16|AIN. Idcirco ego plorans,et oculus meus deducens aquas,quia longe factus est a me consolatorreficiens animam meam;facti sunt filii mei desolati,quoniam invaluit inimicus ".
LAM|1|17|PHE. Expandit Sion manus suas,non est qui consoletur eam;mandavit Dominus adversum Iacobin circuitu eius hostes eius:facta est Ierusalemquasi polluta menstruis inter eos.
LAM|1|18|SADE. " Iustus est Dominus,quia contra os eius rebellis fui.Audite, obsecro, universi populi,et videte dolorem meum:virgines meae et iuvenes meiabierunt in captivitatem.
LAM|1|19|COPH. Vocavi amicos meos,et ipsi deceperunt me;sacerdotes mei et senes meiin urbe consumpti sunt,quia quaesierunt cibum sibi,ut refocillarent animam suam.
LAM|1|20|RES. Vide, Domine, quoniam tribulor;efferbuerunt viscera mea,subversum est cor meum in memetipsa,quoniam valde rebellis fui;foris orbavit me gladiuset domi mors.
LAM|1|21|SIN. Audi, quia ingemisco ego,et non est qui consoletur me;omnes inimici mei audierunt malum meum,laetati sunt quoniam tu fecisti.Adduc diem, quem proclamasti,et fient similes mei.
LAM|1|22|THAU. Ingrediatur omne malum eorum coram te,et fac eis,sicut fecisti mihipropter omnes iniquitates meas;multi enim gemitus mei,et cor meum maerens ".
LAM|2|1|ALEPH. Quomodo obtexit caligine in furore suoDominus filiam Sion!Proiecit de caelo in terramgloriam Israelet non est recordatus scabelli pedum suorumin die furoris sui.
LAM|2|2|BETH. Praecipitavit Dominusnec pepercit omnia pascua Iacob;destruxit in furore suomunitiones filiae Iudae;deiecit in terram, polluitregnum et principes eius.
LAM|2|3|GHIMEL. Confregit in ira furoris suiomne cornu Israel;avertit retrorsum dexteram suama facie inimiciet succendit in Iacob quasi ignem flammaedevorantis in gyro.
LAM|2|4|DALETH. Tetendit arcum suum quasi inimicus,firmavit dexteram suam quasi hostiset occidit omne,quod pulchrum erat visu,in tabernaculo filiae Sion;effudit quasi ignem indignationem suam.
LAM|2|5|HE. Factus est Dominus velut inimicus,deglutivit Israel,deglutivit omnia moenia eius,dissipavit munitiones eiuset multiplicavit in filia Iudaemaerorem et maestitiam.
LAM|2|6|VAU. Et dissipavit quasi hortum saepem suam,demolitus est tabernaculum suum; oblivioni tradidit Dominus in Sion festivitatem et sabbatumet despexit in indignatione furoris suiregem et sacerdotem.
LAM|2|7|ZAIN. Reppulit Dominus altare suum,maledixit sanctuario suo;tradidit in manu inimicimuros domorum eius:vocem dederunt in domo Dominisicut in die sollemni.
LAM|2|8|HETH. Cogitavit Dominus dissiparemurum filiae Sion;tetendit funiculum,non avertit manum suam a perditione;et in luctum redegit antemurale et murum:pariter elanguerunt.
LAM|2|9|TETH. Defixae sunt in terra portae eius;perdidit et contrivit vectes eius.Rex eius et principes eius in gentibus;non est lex,et prophetae eius non inveneruntvisionem a Domino.
LAM|2|10|IOD. Sederunt in terra,conticuerunt senes filiae Sion,consperserunt cinere capita sua,accincti sunt ciliciis;abiecerunt in terram capita suavirgines Ierusalem.
LAM|2|11|CAPH. Defecerunt prae lacrimis oculi mei,efferbuerunt viscera mea;effusum est in terra iecur meumsuper contritione filiae populi mei,cum deficeret parvulus et lactansin plateis oppidi.
LAM|2|12|LAMED. Matribus suis dixerunt: Ubi est triticum et vinum? ",cum deficerent quasi vulneratiin plateis civitatis,cum exhalarent animas suasin sinu matrum suarum.
LAM|2|13|MEM. Cui comparabo te vel cui assimilabo te,filia Ierusalem?Cui exaequabo te et consolabor te, virgo filia Sion?Magna est enim velut mare contritio tua;quis medebitur tui?
LAM|2|14|NUN. Prophetae tui viderunt tibi falsa et stultanec aperiebant iniquitatem tuam,ut converterent sortem tuam;viderunt autem tibi oraculamendacii et seductionis.
LAM|2|15|SAMECH. Plauserunt super te manibusomnes transeuntes per viam;sibilaverunt et moverunt caput suumsuper filiam Ierusalem: Haeccine est urbs, quam vocabant perfectum decorem,gaudium universae terrae? ".
LAM|2|16|PHE. Aperuerunt super te os suumomnes inimici tui;sibilaverunt et fremuerunt dentibuset dixerunt: " Devoravimus;en ista est dies, quam exspectabamus:invenimus, vidimus ".
LAM|2|17|AIN. Fecit Dominus, quae cogitavit;complevit sermonem suum,quem praeceperat a diebus antiquis:destruxit et non pepercit.Et laetificavit super te inimicumet exaltavit cornu hostium tuorum.
LAM|2|18|SADE. Clamet cor tuum ad Dominumsuper muros filiae Sion;deduc quasi torrentem lacrimasper diem et noctem.Non des requiem tibi,neque taceat pupilla oculi tui.
LAM|2|19|COPH. Consurge, lamentare in noctein principio vigiliarum,effunde sicut aquam cor tuumante conspectum Domini;leva ad eum manus tuaspro anima parvulorum tuorum,qui defecerunt in famein capite omnium compitorum.
LAM|2|20|RES. " Vide, Domine, et considera,cui feceris ita;ergone comedent mulieres fructum suum,parvulos diligenter fovendos?Num occidetur in sanctuario Dominisacerdos et propheta?
LAM|2|21|SIN. Iacuerunt in terra forispuer et senex;virgines meae et iuvenes meiceciderunt in gladio:interfecisti in die furoris tui,percussisti nec misertus es.
LAM|2|22|THAU. Vocasti quasi ad diem sollemnem,qui terrerent me de circuitu,et non fuit in die furoris Domini,qui effugeret et relinqueretur:quos fovi et enutrivi,inimicus meus consumpsit eos ".
LAM|3|1|ALEPH. Ego vir videns paupertatem meamin virga indignationis eius.
LAM|3|2|ALEPH. Me minavit et adduxitin tenebras et non in lucem.
LAM|3|3|ALEPH. Tantum in me vertit et convertitmanum suam tota die.
LAM|3|4|BETH. Consumpsit pellem meam et carnem meam,contrivit ossa mea.
LAM|3|5|BETH. Aedificavit in gyro meoet circumdedit me felle et labore.
LAM|3|6|BETH. In tenebrosis collocavit mequasi mortuos sempiternos.
LAM|3|7|GHIMEL. Circumaedificavit adversum me, ut non egrediar,aggravavit compedem meum.
LAM|3|8|GHIMEL. Sed et cum clamavero et rogavero,exclusit orationem meam.
LAM|3|9|GHIMEL. Conclusit vias meas lapidibus quadris,semitas meas subvertit.
LAM|3|10|DALETH. Ursus insidians factus est mihi,leo in absconditis.
LAM|3|11|DALETH. Semitas meas subvertit et confregit me,posuit me desolatam.
LAM|3|12|DALETH. Tetendit arcum suum et posuit mequasi signum ad sagittam.
LAM|3|13|HE. Misit in renibus meisfilias pharetrae suae.
LAM|3|14|HE. Factus sum in derisum omni populo meo,canticum eorum tota die.
LAM|3|15|HE. Replevit me amaritudinibus,inebriavit me absinthio.
LAM|3|16|VAU. Et fregit in glarea dentes meos,depressit me cinere.
LAM|3|17|VAU. Et repulsa est a pace anima mea,oblitus sum bonorum.
LAM|3|18|VAU. Et dixi: " Periit splendor meus et spes mea a Domino ".
LAM|3|19|ZAIN. Recordare paupertatis et peregrinationis meae,absinthii et fellis.
LAM|3|20|ZAIN. Memoria memor estet tabescit in me anima mea.
LAM|3|21|ZAIN. Haec recolam in corde meo,ideo sperabo.
LAM|3|22|HETH. Misericordiae Domini, quia non sumus consumpti,quia non defecerunt miserationes eius.
LAM|3|23|HETH. Novae sunt omni mane,magna est fides tua.
LAM|3|24|HETH. " Pars mea Dominus, dixit anima mea;propterea exspectabo eum ".
LAM|3|25|TETH. Bonus est Dominus sperantibus in eum,animae quaerenti illum.
LAM|3|26|TETH. Bonum est praestolari cum silentiosalutare Domini.
LAM|3|27|TETH. Bonum est viro, cum portaveritiugum ab adulescentia sua.
LAM|3|28|IOD. Sedebit solitarius et tacebit,cum istud imponitur ei.
LAM|3|29|IOD. Ponet in pulvere os suum,si forte sit spes.
LAM|3|30|IOD. Dabit percutienti se maxillam,saturabitur opprobriis.
LAM|3|31|CAPH. Quia non repellet in sempiternumDominus.
LAM|3|32|CAPH. Quia si afflixit, et miserebitursecundum multitudinem misericordiarum suarum.
LAM|3|33|CAPH. Non enim humiliat ex corde suoet affligit filios hominum.
LAM|3|34|LAMED. Conterere sub pedibus suisomnes vinctos terrae.
LAM|3|35|LAMED. Declinare iudicium viriin conspectu vultus Altissimi.
LAM|3|36|LAMED. Pervertere hominem in iudicio suo,num Dominus haec ignorat?
LAM|3|37|MEM. Quis est iste, qui dixit, et factum est?Dominus non iussit?
LAM|3|38|MEM. Ex ore Altissimi nonne egrediunturet mala et bona?
LAM|3|39|MEM. Quid murmurabit homo vivens,vir pro peccatis suis?
LAM|3|40|NUN. " Scrutemur vias nostras et quaeramuset revertamur ad Dominum.
LAM|3|41|NUN. Levemus corda nostra cum manibusad Dominum in caelos.
LAM|3|42|NUN. Nos inique egimus et rebelles fuimus;idcirco tu inexorabilis fuisti.
LAM|3|43|SAMECH. Operuisti in furore et percussisti nos;occidisti nec pepercisti.
LAM|3|44|SAMECH. Opposuisti nubem tibi,ne transeat oratio.
LAM|3|45|SAMECH. In eradicationem et abiectionem posuisti nosin medio populorum.
LAM|3|46|PHE. Aperuerunt super nos os suumomnes inimici nostri.
LAM|3|47|PHE. Formido et fovea facta est nobis,vastatio et contritio ".
LAM|3|48|PHE. Rivos aquarum deducit oculus meusin contritione filiae populi mei.
LAM|3|49|AIN. Oculus meus lacrimas effundit nec tacet,eo quod non sit requies.
LAM|3|50|AIN. Donec respiciat et videatDominus de caelis.
LAM|3|51|AIN. Oculus meus affligit animam meamprae cunctis filiabus urbis meae.
LAM|3|52|SADE. Venatione venati sunt me quasi aveminimici mei gratis.
LAM|3|53|SADE. Perdiderunt in lacu vitam meamet iecerunt lapides super me.
LAM|3|54|SADE. Inundaverunt aquae super caput meum,dixi: " Perii ".
LAM|3|55|COPH. Invocavi nomen tuum, Domine,de profunditate lacus.
LAM|3|56|COPH. Vocem meam audisti: " Ne avertasaurem tuam a singultu meo et clamoribus ".
LAM|3|57|COPH. Appropinquasti in die, quando invocavi te,dixisti: " Ne timeas ".
LAM|3|58|RES. Iudicasti, Domine, causam animae meae,redemisti vitam meam.
LAM|3|59|RES. Vidisti, Domine, afflictionem meam;iudica iudicium meum.
LAM|3|60|RES. Vidisti omnem furorem eorum, universas cogitationes eorum adversum me.
LAM|3|61|SIN. Audisti opprobrium eorum, Domine,omnes cogitationes eorum adversum me.
LAM|3|62|SIN. Labia insurgentium mihi et meditationes eorumadversum me tota die.
LAM|3|63|SIN. Sessionem eorum et resurrectionem eorum vide;ego sum psalmus eorum.
LAM|3|64|THAU. Reddes eis vicem, Domine,iuxta opera manuum suarum.
LAM|3|65|THAU. Dabis eis duritiam cordis,exsecrationem tuam.
LAM|3|66|THAU. Persequeris in furore et conteres eossub caelis tuis, Domine.
LAM|4|1|ALEPH. Quomodo obscuratum est aurum,mutatum est obryzum optimum!Dispersi sunt lapides sanctiin capite omnium platearum.
LAM|4|2|BETH. Filii Sion inclitiet ponderati auro primo,quomodo reputati sunt in vasa testea,opus manuum figuli!
LAM|4|3|GHIMEL. Sed et thoes nudaverunt mammam,lactaverunt catulos suos;filia populi mei crudelisquasi struthio in deserto.
LAM|4|4|DALETH. Adhaesit lingua lactantisad palatum eius in siti;parvuli petierunt panem,et non erat qui frangeret eis.
LAM|4|5|HE. Qui vescebantur voluptuose,interierunt in viis;qui nutriebantur in coccinis,amplexati sunt stercora.
LAM|4|6|VAU. Et maior effecta est iniquitas filiae populi meipeccato Sodomae,quae subversa est in momento,et non laborabant in ea manus.
LAM|4|7|ZAIN. Candidiores nazaraei eius nive,nitidiores lacte,rubicundiores in corpore coralliis,sapphirus aspectus eorum.
LAM|4|8|HETH. Denigrata est super carbones facies eorum,et non sunt cogniti in plateis:adhaesit cutis eorum ossibus,aruit et facta est quasi lignum.
LAM|4|9|TETH. Melius fuit occisis gladioquam interfectis fame,quoniam isti extabuerunt consumptia sterilitate terrae.
LAM|4|10|IOD. Manus mulierum misericordiumcoxerunt filios suos:facti sunt cibus earumin contritione filiae populi mei.
LAM|4|11|CAPH. Complevit Dominus furorem suum,effudit iram indignationis suae;et succendit ignem in Sion,qui devoravit fundamenta eius.
LAM|4|12|LAMED. Non crediderunt reges terraeet universi habitatores orbis,quoniam ingrederetur hostis et inimicusper portas Ierusalem.
LAM|4|13|MEM. Propter peccata prophetarum eiuset iniquitates sacerdotum eius,qui effuderunt in medio eiussanguinem iustorum.
LAM|4|14|NUN. Erraverunt caeci in plateis,polluti sunt in sanguine,ita ut nemo posset attingerelacinias eorum.
LAM|4|15|SAMECH. " Recedite! Pollutus est ", clamaverunt eis; Recedite, abite, nolite tangere! ".Cum fugerent et errarent, dixerunt inter gentes: Non addent ultra ut incolant ".
LAM|4|16|PHE. Facies Domini dispersit eos,non addet ut respiciat eos;facies sacerdotum non respexeruntneque senum miserti sunt.
LAM|4|17|AIN. Adhuc deficiunt oculi nostriad auxilium nostrum vanum?In specula nostra respeximusad gentem, quae salvare non potest.
LAM|4|18|SADE. Insidiati sunt vestigiis nostris,ne iremus per plateas nostras. Appropinquavit finis noster, completi sunt dies nostri,quia venit finis noster ".
LAM|4|19|COPH. Velociores fuerunt persecutores nostriaquilis caeli;super montes persecuti sunt nos,in deserto insidiati sunt nobis.
LAM|4|20|RES. Spiritus oris nostri, unctus Domini,captus est in foveis eorum,de quo dicebamus: " Sub umbra suavivemus in gentibus ".
LAM|4|21|SIN. Gaude et laetare, filia Edom,quae habitas in terra Us;ad te quoque perveniet calix,inebriaberis atque nudaberis.
LAM|4|22|THAU. Completa est iniquitas tua, filia Sion,non addet ultra ut transmigret te;visitavit iniquitatem tuam, filia Edom,discooperuit peccata tua.
LAM|5|1|Recordare, Domine, quid acci derit nobis;intuere et respice opprobrium nostrum.
LAM|5|2|Hereditas nostra versa est ad alienos,domus nostrae ad extraneos.
LAM|5|3|Pupilli facti sumus absque patre,matres nostrae quasi viduae.
LAM|5|4|Aquam nostram pecunia bibimus,ligna nostra pretio comparamus.
LAM|5|5|Iugum in cervicibus nostris minamur;lassis non datur requies.
LAM|5|6|Aegyptiis dedimus manum et Assyriis,ut saturaremur pane.
LAM|5|7|Patres nostri peccaverunt et non sunt,et nos iniquitates eorum portamus.
LAM|5|8|Servi dominantur nostri;non est qui redimat de manu eorum.
LAM|5|9|Vitae nostrae periculo afferimus panem nobisa facie gladii in deserto.
LAM|5|10|Pellis nostra quasi clibanus exusta estpropter aestum famis.
LAM|5|11|Mulieres in Sion humiliaveruntet virgines in civitatibus Iudae.
LAM|5|12|Principes manu eorum suspensi sunt;facies senum honorem non habuerunt.
LAM|5|13|Adulescentes molam portaverunt,et pueri sub lignis corruerunt.
LAM|5|14|Senes deficiunt de portis,iuvenes de choro psallentium.
LAM|5|15|Defecit gaudium cordis nostri;versus est in luctum chorus noster.
LAM|5|16|Cecidit corona capitis nostri;vae nobis, quia peccavimus!
LAM|5|17|Propterea maestum factum est cor nostrum,ideo contenebrati sunt oculi nostri,
LAM|5|18|propter montem Sion, quia desolatus est:vulpes ambulant in eo.
LAM|5|19|Tu autem, Domine, in aeternum permanebis,solium tuum in generationem et generationem.
LAM|5|20|Quare in perpetuum oblivisceris nostri,derelinques nos in longitudinem dierum?
LAM|5|21|Converte nos, Domine, ad te, et convertemur;innova dies nostros sicut a principio.
LAM|5|22|Ergone proiciens reppulisti nos,iratus es contra nos vehementer?
