HAB|1|1|Пророцтво, яке бачив пророк Авакум.
HAB|1|2|Аж доки я, Господи, кликати буду, а Ти не почуєш? До тебе я кличу: Насильство! та Ти не спасаєш!
HAB|1|3|Для чого неправість мені Ти показуєш та позираєш на муку? А передо мною грабіж та насильство, і суперечка стається, і носиться сварка.
HAB|1|4|Тому то Закон припиняється, і не виходить до чину назавсіди право, бо несправедливий вигублює праведного, тому правосуддя виходить покривленим.
HAB|1|5|Пригляньтеся ви до народів, і дивіться, і дуже здивуйтесь, бо вчиню Я за ваших днів діло, про яке не повірите ви, коли буде розказане.
HAB|1|6|Бо оце Я поставлю халдеїв, народ лютий та скорий, що ґрасує по широкій землі, щоб захопити оселі, які не його.
HAB|1|7|Страшний та грізний він, від нього самого виходить і право його, і великість його.
HAB|1|8|І від пантер його коні швидші, і від вовків вечерових лютіші.
HAB|1|9|Він приходить увесь на насильство, а ціль їх обличчя вперед, і набере полонених, як того піску.
HAB|1|10|І він глузує з царів, а князі сміх для нього. Він сміється з твердині усякої, бо на вал насипає землі, і її здобуває!
HAB|1|11|Тоді він несеться, як вітер, і перейде, і згрішить, бо зробить за бога свого оцю силу свою.
HAB|1|12|Хіба ж Ти не віддавна, о Господи? Боже Ти мій, мій Святий, не помремо! Господи, Ти для суду поставив його, і, о Скеле, призначив його на карання!
HAB|1|13|Твої очі занадто пречисті, щоб міг Ти дивитись на зло, і на насильство дивитись не можеш. Чому ж дивишся Ти на грабіжників, мовчиш, коли несправедливий винищує справедливішого від себе?
HAB|1|14|Ти ж маєш людей, як у морі тих риб, немов ту черву, що пана над нею нема.
HAB|1|15|Усе це грабіжник витягує вудкою, своїм неводом тягне оце, та збирає оце в свою сітку, тому тішиться він та радіє.
HAB|1|16|Тому жертву приносить він неводові, і кадить для сітки своєї, бо від них ситий уділ його та добірна пожива його!
HAB|1|17|Чи на це випорожнює він свого невода, і завжди готов убивати народи без милости?
HAB|2|1|Нехай я стою на сторожі своїй, і нехай на облозі я стану, і хай виглядаю, щоб бачити, що він буде казати мені, і що відповість на жалобу мою.
HAB|2|2|А Господь відповів та й сказав: Напиши це видіння і поясни на таблицях, щоб читач його легко читав.
HAB|2|3|Бо ще на умовлений час це видіння, і приспішає кінець, і не обмане. Якщо б протягнулось, чекай ти його, бо воно конче прийде, не спізниться.
HAB|2|4|Ось надута, не проста душа його в ньому, а праведний житиме вірою своєю.
HAB|2|5|І що ж, як зрадливе вино, так горда людина спокою не знає: він роззявлює пащу свою, як шеол, і не насичується, як та смерть, і всіх людей він до себе збирає, і всі народи до себе згромаджує.
HAB|2|6|Чи ж усі вони не складуть приповістки на нього та загадки насмішливої йому не прокажуть: Горе тому, хто для себе розмножує те, що не його! Аж доки це буде? Горе тому, хто чинить тяжкою заставу на себе!
HAB|2|7|Хіба нагло не встануть оті, хто тебе буде гризти, і збудяться ті, хто тебе попихає, і за здобич ти станеш для них?
HAB|2|8|За те, що ти грабував був багато народів, вся решта народів тебе пограбує за ту людську кров, і за насильство над краєм, над містом та над усіма, хто мешкає в ньому.
HAB|2|9|Горе тому, хто неправедний зиск побирає для дому свого, щоб покласти гніздо своє на висоті, і тим із рук злого врятованим бути!
HAB|2|10|Нарадив ти сором для дому свого, щоб кінець учинити численним народам, і ти прогрішився за душу свою.
HAB|2|11|Бо камінь з стіни буде кликати, і йому відповість сволок із дерева.
HAB|2|12|Горе тому, хто кров'ю місто будує, хто беззаконням встановлює город!
HAB|2|13|Чи ж оце не від Господа Саваота, що народи трудяться для огню, і мучаться люди на марність?
HAB|2|14|Бо пізнанням Господньої слави наповнена буде земля, як море вода покриває.
HAB|2|15|Горе тому, хто свого ближнього напоює з келіху гніву свого, і поїть, щоб бачити сором його!
HAB|2|16|Ти наситишся ганьбою більше, як славою. Пий також ти, та показуй свій сором! На тебе обернеться келіх правиці Господньої, ганьба ж на славу твою!
HAB|2|17|Бо насилля твоє над Ліваном на тебе спаде, а грабунок худоби зламає тебе за кров людську, та за насилля над краєм, над містом та над усіма, хто мешкає в ньому.
HAB|2|18|Який дасть пожиток бовван, що його вирізьбив творець його, і відлив, і вчитель неправди, що творець його мав охоту чинити богів цих німих?
HAB|2|19|Горе тому, хто дереву каже: Збудись, мовчазливому каменю: Зрушся! Чи він буде навчати? Ось він сріблом та золотом викладений, але жодного духу в ньому нема!
HAB|2|20|А Господь у Своїм храмі святім, мовчи перед обличчям Його, уся земле!
HAB|3|1|Молитва пророка Авакума, для співу на струнному приладі:
HAB|3|2|Господи, звістку Твою я почув та й злякався! Господи, оживи Своє діло в середині років, у середині літ об'яви, у гніві про милість згадай!
HAB|3|3|Бог іде від Теману, і Святий від Парану гори. Села. Велич Його вкрила небо, і слави Його стала повна земля!
HAB|3|4|А сяйво було, наче соняшне світло, проміння при боці у Нього, і там укриття Його потуги.
HAB|3|5|Перед обличчям Його моровиця іде, а по стопах Його пнеться полум'я.
HAB|3|6|Став, і землю Він зміряв, поглянув і народи затряс, і попадали гори довічні, вікові похилились узгір'я. Путі Його вічні.
HAB|3|7|Я бачив намети Кушана під кривдою, тремтять покривала мідіянського краю.
HAB|3|8|Чи на ріки, о Господи, Ти запалав, чи на ріки Твій гнів? Чи Твоє пересердя на море, що їздиш на конях Своїх, на спасенних Своїх колесницях?
HAB|3|9|Лук твій голий, нагий, наповнений стріл сагайдак. Села. Ти річками землю розсік.
HAB|3|10|Тебе вгледівши, гори дрижали, водяна течія потекла, безодня свій голос дала, зняла високо руки свої.
HAB|3|11|Сонце й місяць спинилися в мешканні своєму при світлі Твоїх стріл, що літають при сяйві блискучого списа Твого.
HAB|3|12|У люті ступав Ти землею, у гніві людей молотив.
HAB|3|13|Ти вийшов спасти Свій народ, спасти Помазанця Свого. Ти з дому безбожного голову збив, обнажив Ти основу по шию. Села.
HAB|3|14|Ти пробив його списами голову князя його, як вони піднялись, щоб мене розпорошити; вони тішилися, немов мали пожерти таємно убогого.
HAB|3|15|Ти кіньми Своїми по морю топтав, по водній великій громаді.
HAB|3|16|Я почув і затремтіла утроба моя, задзвеніли на голос цей губи мої, гнилизна ввійшла в мої кості, і тремчу я на місці своїм, бо маю чекати в спокої день утиску, коли прийде народ, який має на вас наступати.
HAB|3|17|Коли б фіґове дерево не зацвіло, і не було б урожаю в виноградниках, обманило зайняття оливкою, а поле їжі не вродило б, позникала отара з кошари і не стало б в оборах худоби,
HAB|3|18|то я Господом тішитись буду й тоді, радітиму Богом спасіння свого!
HAB|3|19|Бог Господь моя сила, і чинить Він ноги мої, як у лані, і водить мене по висотах! Для дириґента хору на моїх струнних знаряддях.
