NAH|1|1|論 尼尼微 的默示， 伊勒歌斯 人 那鴻 所見異象的書。
NAH|1|2|耶和華是忌邪 、報應的上帝。 耶和華施報應，大有憤怒； 耶和華向他的敵人報應， 向他的仇敵懷怒。
NAH|1|3|耶和華不輕易發怒，大有能力， 但耶和華萬不以有罪的為無罪。 他的道路在旋風和暴風之中， 雲彩為他腳下的塵土。
NAH|1|4|他斥責海，使海枯乾， 使一切江河乾涸。 巴珊 和 迦密 衰殘， 黎巴嫩 的花草也衰殘了。
NAH|1|5|大山因他震動， 小山也都融化； 大地在他面前突起， 世界和住在其間的也都如此。
NAH|1|6|他發憤恨，誰能立得住呢？ 他發烈怒，誰能當得起呢？ 他的憤怒如火傾洩而出， 磐石因他崩裂。
NAH|1|7|耶和華本為善， 在患難的日子為人的保障， 並且認識那些投靠他的人；
NAH|1|8|但他必以漲溢的洪水淹沒其地方 ， 又驅逐仇敵進入黑暗。
NAH|1|9|你們籌劃何種計謀攻擊耶和華呢？ 他必終結一切， 仇敵 不會再度興起。
NAH|1|10|你們像雜亂的荊棘， 像喝醉了的人， 又如枯乾的碎秸，全然燒滅。
NAH|1|11|有一人從你那裏出來， 圖謀邪惡，設惡計攻擊耶和華。
NAH|1|12|耶和華如此說： 「他們雖然勢力強大，人數眾多， 也要被剪除，歸於無有。 我雖曾使你受苦， 卻不再使你受苦。
NAH|1|13|現在，我要從你身上折斷他的軛， 解開捆綁你的繩索。」
NAH|1|14|耶和華已經發命令，指著你說： 「你的名下必不再留後； 我要從你神明的廟中除滅雕刻的偶像和鑄造的偶像， 我必因你的卑賤，為你預備墳墓。」
NAH|1|15|看哪，山上有報佳音、傳平安之人的腳蹤。 猶大 啊，守你的節期， 還你的願吧！ 因為惡人不再侵犯你， 他已滅絕淨盡了。
NAH|2|1|那打碎你的人 上到你面前。 要看守堡壘，把守道路， 要挺起腰來，大大使力。
NAH|2|2|耶和華復興 雅各 的榮華， 像復興 以色列 的榮華； 因為蹂躪者曾經蹂躪他們， 毀壞了他們的葡萄枝。
NAH|2|3|他勇士的盾牌是紅的， 精兵都穿朱紅衣服。 在預備打仗的日子， 戰車上的鐵閃爍如火 ， 柏木的槍桿也已舉起 ；
NAH|2|4|戰車在街上疾行， 在廣場上來往奔馳， 形狀如火把， 飛馳如閃電。
NAH|2|5|他 招聚他的貴族； 他們前行時絆跌， 速上城牆， 預備屏障。
NAH|2|6|河閘開放， 宮殿沖沒。
NAH|2|7|這是命定之事： 王后赤身被擄 ， 宮女搥胸， 哀鳴如鴿子。
NAH|2|8|尼尼微 自古以來 如同聚水的池子； 現在居民都在逃跑 。 「站住！站住！」 卻無人回轉。
NAH|2|9|你們搶奪金子吧！ 你們搶奪銀子吧！ 因為所積蓄的無窮， 華美的寶器無數。
NAH|2|10|荒蕪，荒涼，全然荒廢， 人心害怕，雙膝顫抖， 腰部疼痛，臉都變色。
NAH|2|11|獅子的洞， 幼獅餵養之處在哪裏呢？ 公獅、母獅、小獅出入， 無人使牠們驚嚇之地在哪裏呢？
NAH|2|12|公獅撕碎的足夠給幼獅吃， 又為母獅掐死獵物， 把獵物塞滿牠的洞穴， 把撕碎的裝滿牠的窩。
NAH|2|13|看哪，我與你為敵，將它的戰車 焚燒成煙，刀劍必吞滅你的少壯獅子；我必從地上除滅你的獵物，你使者的聲音必不再聽見。這是萬軍之耶和華說的。
NAH|3|1|禍哉！這流人血的城， 欺詐連連，搶奪充斥， 擄掠的事總不止息。
NAH|3|2|鞭聲響亮，車輪轟轟， 馬匹跳躍，戰車奔騰；
NAH|3|3|騎兵爭先，刀劍發光， 槍矛閃爍，被殺的甚多， 屍首成堆，屍骸無數， 人因屍骸而絆跌，
NAH|3|4|都因那美貌的妓女多有淫行， 慣行邪術， 藉淫行誘惑 列國， 用邪術誘惑萬族。
NAH|3|5|看哪，我與你為敵， 掀開你的下襬，蒙在你臉上， 使列邦看見你的赤體， 使列國觀看你的羞辱。 這是萬軍之耶和華說的。
NAH|3|6|我必將可憎污穢之物拋在你身上， 使你被藐視，為眾人所觀看。
NAH|3|7|凡看見你的，都必逃離你，說： 「 尼尼微 荒涼了！有誰為你悲傷呢？ 我何處找到安慰你的人呢？」
NAH|3|8|你能勝過 挪亞們 嗎？ 它坐落在眾河之間， 周圍有水， 海 作它的城郭， 海 作它的城牆。
NAH|3|9|古實 和 埃及 是它的力量， 沒有窮盡， 弗 人和 路比 人是它的幫手。
NAH|3|10|但它被流放，被人擄去， 它的嬰孩也被摔碎在各街頭； 人為它的貴族抽籤， 它的權貴都被鎖鏈鎖住。
NAH|3|11|你也必喝醉，昏迷錯亂， 並因仇敵的緣故尋求庇護。
NAH|3|12|你一切的堡壘必如無花果樹上初熟的果子， 一經搖動，就落在想吃的人口中。
NAH|3|13|看哪，你中間的士兵是婦女， 你國中的關口向仇敵敞開， 你的門閂被火焚燒。
NAH|3|14|你要打水預備受困； 要加強防禦， 取土踹泥， 做成磚模。
NAH|3|15|在那裏，火要吞滅你， 刀必殺戮你， 如蝻子般吞滅你。 你人數增多如蝻子， 增多如蝗蟲吧！
NAH|3|16|你增添商賈，多過天上的星宿； 如蝻子蛻皮飛去。
NAH|3|17|你的領袖多如蝗蟲， 你的將軍彷彿成群的蝗蟲； 天涼時齊落在籬笆上， 太陽一出就飛去， 人不知道落在何處。
NAH|3|18|亞述 王啊， 你的牧人睡覺， 你的貴族躺臥 ， 你的百姓散在山間， 無人招聚。
NAH|3|19|你的損傷並未減輕， 你的傷痕極其重大。 凡聽見這消息的人都因你拍掌。 有誰沒有時常遭受你的暴行呢？
