2PET|1|1|Симеон Петро, раб та апостол Ісуса Христа, до тих, хто одержав із нами рівноцінну віру в правді Бога нашого й Спасителя Ісуса Христа:
2PET|1|2|благодать вам та мир нехай примножиться в пізнанні Бога й Ісуса, Господа нашого!
2PET|1|3|Усе, що потрібне для життя та побожности, подала нам Його Божа сила пізнанням Того, Хто покликав нас славою та чеснотою.
2PET|1|4|Через них даровані нам цінні та великі обітниці, щоб ними ви стали учасниками Божої Істоти, утікаючи від пожадливого світового тління.
2PET|1|5|Тому докладіть до цього всю пильність, і покажіть у вашій вірі чесноту, а в чесноті пізнання,
2PET|1|6|а в пізнанні стримання, а в стриманні терпеливість, а в терпеливості благочестя,
2PET|1|7|а в благочесті братерство, а в братерстві любов.
2PET|1|8|Бо коли це в вас є та примножується, то воно зробить вас нелінивими, ані безплідними для пізнання Господа нашого Ісуса Христа.
2PET|1|9|А хто цього не має, той сліпий, короткозорий, він забув про очищення з своїх давніх гріхів.
2PET|1|10|Тому, браття, тим більше дбайте чинити міцним своє покликання та вибрання, бо, роблячи так, ви ніколи не спіткнетесь.
2PET|1|11|Бо щедро відкриється вам вхід до вічного Царства Господа нашого й Спасителя Ісуса Христа.
2PET|1|12|Тому то ніколи я не занедбую про це вам нагадувати, хоч ви й знаєте, і впевнені в теперішній правді.
2PET|1|13|Бо вважаю я за справедливе, доки я в цій оселі, спонукувати вас нагадуванням,
2PET|1|14|знаючи, що я незабаром повинен покинути оселю свою, як і Господь наш Ісус Христос об'явив був мені.
2PET|1|15|А я пильнуватиму, щоб ви й по моєму відході завжди мали це в пам'яті.
2PET|1|16|Бо ми сповістили вам силу та прихід Господа нашого Ісуса Христа, не йдучи за хитро видуманими байками, але бувши самовидцями Його величі.
2PET|1|17|Бо Він честь та славу прийняв від Бога Отця, як до Нього прийшов від величної слави голос такий: Це Син Мій Улюблений, що Його Я вподобав!
2PET|1|18|І цей голос, що з неба зійшов, ми чули, як із Ним були на святій горі.
2PET|1|19|І ми маємо слово пророче певніше. І ви добре робите, що на нього вважаєте, як на світильника, що світить у темному місці, аж поки зачне розвиднятися, і світова зірниця засяє у ваших серцях,
2PET|1|20|бо ви знаєте перше про те, що жодне пророцтво в Писанні від власного вияснення не залежить.
2PET|1|21|Бо пророцтва ніколи не було з волі людської, а звіщали його святі Божі мужі, проваджені Духом Святим.
2PET|2|1|А між людом були й неправдиві пророки, як і будуть між вас учителі неправдиві, що впровадять згубні єресі, відречуться від Владики, що викупив їх, і стягнуть на себе самі скору погибіль.
2PET|2|2|І багато-хто підуть за пожадливістю їхньою, а через них дорога правдива зневажиться.
2PET|2|3|І в зажерливості вони будуть ловити вас словами облесними. Суд на них віддавна не бариться, а їхня загибіль не дрімає!
2PET|2|4|Бо як Бог Анголів, що згрішили, не помилував був, а в кайданах темряви вкинув до аду, і передав зберігати на суд;
2PET|2|5|і Він не помилував першого світу, а зберіг самовосьмого Ноя, проповідника праведности, і навів потопа на світ безбожних;
2PET|2|6|і міста Содом і Гоморру спопелив, засудивши на знищення, і дав приклада для майбутніх безбожників,
2PET|2|7|а врятував праведного Лота, змученого поводженням розпусних людей,
2PET|2|8|бо цей праведник, живши між ними, день-у-день мучив свою праведну душу, бачачи й чуючи вчинки безбожні,
2PET|2|9|то вміє Господь рятувати побожних від спокуси, а неправедних берегти на день суду для кари,
2PET|2|10|а надто тих, хто ходить за нечистими пожадливостями тіла та погорджує владою; зухвалі свавільці, що не бояться зневажати слави,
2PET|2|11|хоч Анголи, бувши міццю та силою більші за них, не несуть до Господа зневажливого суду на них.
2PET|2|12|Вони, немов звірина нерозумна, зроджена природою на зловлення та загибіль, зневажають те, чого не розуміють, і в тлінні своїм будуть знищені,
2PET|2|13|і приймуть заплату за лихі вчинки. Вони повсякденну розпусту вважають за розкіш; самі бруд та неслава, вони насолоджуються своїми оманами, бенкетуючи з вами.
2PET|2|14|Їхні очі наповнені перелюбом та гріхом безупинним; вони зваблюють душі незміцнені; вони, діти прокляття, мають серце, привчене до зажерливости.
2PET|2|15|Вони покинули просту дорогу та й заблудили, і пішли слідом за Валаамом Беоровим, що полюбив нагороду несправедливости,
2PET|2|16|але був докорений у своїм беззаконні: німа під'яремна ослиця проговорила людським голосом, та й безум пророка спинила.
2PET|2|17|Вони джерела безводні, хмари, бурею гнані; для них приготований морок темряви!
2PET|2|18|Бо, висловлюючи марне базікання, вони зваблюють пожадливістю тіла й розпустою тих, хто ледве втік від тих, хто живе в розпусті.
2PET|2|19|Вони волю обіцюють їм, самі бувши рабами тління. Бо хто ким переможений, той тому й раб.
2PET|2|20|Бо коли хто втече від нечистости світу через пізнання Господа й Спасителя Ісуса Христа, а потому знов заплутуються ними та перемагаються, то останнє буває для них гірше першого.
2PET|2|21|Бо краще було б не пізнати їм дороги праведности, аніж, пізнавши, вернутись назад від переданої їм святої заповіді!
2PET|2|22|Бо їм трапилося за правдивою приказкою: Вертається пес до своєї блювотини, та: Помита свиня йде валятися в калюжу...
2PET|3|1|Це вже другого листа пишу я до вас, улюблені. У них нагадуванням я буджу вашу чисту думку,
2PET|3|2|щоб ви пам'ятали слова, що святі пророки давніше звістили їх вам, і заповідь Господа й Спасителя, що одержали через ваших апостолів.
2PET|3|3|Насамперед знайте оце, що в останні дні прийдуть із насмішками глузії, що ходитимуть за своїми пожадливостями,
2PET|3|4|та й скажуть: Де обітниця Його приходу? Бо від того часу, як позасинали наші батьки, усе залишається так від початку творіння.
2PET|3|5|Бо сховане від тих, хто хоче цього, що небо було напочатку, а земля із води та водою складена словом Божим,
2PET|3|6|тому тодішній світ, водою потоплений, згинув.
2PET|3|7|А теперішні небо й земля заховані тим самим словом, і зберігаються для огню на день суду й загибелі безбожних людей.
2PET|3|8|Нехай же одне це не буде заховане від вас, улюблені, що в Господа один день немов тисяча років, а тисяча років немов один день!
2PET|3|9|Не бариться Господь із обітницею, як деякі вважають це барінням, але вам довготерпить, бо не хоче, щоб хто загинув, але щоб усі навернулися до каяття.
2PET|3|10|День же Господній прибуде, як злодій вночі, коли з гуркотом небо мине, а стихії, розпечені, рунуть, а земля та діла, що на ній, погорять...
2PET|3|11|А коли все оце поруйнується, то якими мусите бути в святому житті та в побожності ви,
2PET|3|12|що чекаєте й прагнете скорого приходу Божого дня, в якім небо, палючися, зникне, а розпалені стихії розтопляться?
2PET|3|13|Але за Його обітницею ми дожидаємо неба нового й нової землі, що правда на них пробуває.
2PET|3|14|Тож, улюблені, чекаючи цього, попильнуйте, щоб ви знайшлися для Нього нескверні та чисті у мирі.
2PET|3|15|А довготерпіння Господа нашого вважайте за спасіння, як і улюблений брат наш Павло написав був до вас за даною йому мудрістю,
2PET|3|16|як і по всіх посланнях, що в них він говорить про це. У них є дещо тяжко зрозуміле, що неуки та незміцнені перекручують, як і інші Писання, на власну загибіль свою.
2PET|3|17|Тож ви, улюблені, знаючи це наперед, стережіться, щоб не були ви зведені блудом безбожних і не відпали від свого вґрунтування,
2PET|3|18|але щоб зростали в благодаті й пізнанні Господа нашого й Спасителя Ісуса Христа. Йому слава і тепер, і дня вічного! Амінь.
