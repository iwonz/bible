2JOHN|1|1|senior electae dominae et natis eius quos ego diligo in veritate et non ego solus sed et omnes qui cognoverunt veritatem
2JOHN|1|2|propter veritatem quae permanet in nobis et nobiscum erit in aeternum
2JOHN|1|3|sit nobiscum gratia misericordia pax a Deo Patre et a Christo Iesu Filio Patris in veritate et caritate
2JOHN|1|4|gavisus sum valde quoniam inveni de filiis tuis ambulantes in veritate sicut mandatum accepimus a Patre
2JOHN|1|5|et nunc rogo te domina non tamquam mandatum novum scribens tibi sed quod habuimus ab initio ut diligamus alterutrum
2JOHN|1|6|et haec est caritas ut ambulemus secundum mandata eius hoc mandatum est ut quemadmodum audistis ab initio in eo ambuletis
2JOHN|1|7|quoniam multi seductores exierunt in mundum qui non confitentur Iesum Christum venientem in carne hic est seductor et antichristus
2JOHN|1|8|videte vosmet ipsos ne perdatis quae operati estis sed ut mercedem plenam accipiatis
2JOHN|1|9|omnis qui praecedit et non manet in doctrina Christi Deum non habet qui permanet in doctrina hic et Filium et Patrem habet
2JOHN|1|10|si quis venit ad vos et hanc doctrinam non adfert nolite recipere eum in domum nec have ei dixeritis
2JOHN|1|11|qui enim dicit illi have communicat operibus illius malignis
2JOHN|1|12|plura habens vobis scribere nolui per cartam et atramentum spero enim me futurum apud vos et os ad os loqui ut gaudium vestrum plenum sit
2JOHN|1|13|salutant te filii sororis tuae electae
