MIC|1|1|当 犹大 王 约坦 、 亚哈斯 、 希西家 在位的时候，耶和华的话临到 摩利沙 人 弥迦 ，他见到有关 撒玛利亚 和 耶路撒冷 的异象。
MIC|1|2|万民哪，你们都要听！ 地和其上所有的，要留心听！ 主耶和华要从他的圣殿 指证你们的不是。
MIC|1|3|看哪，耶和华从他的居所出来， 降临步行地之高处。
MIC|1|4|众山在他底下熔化， 诸谷崩裂， 如蜡熔在火中， 如水冲下山坡。
MIC|1|5|这都是因 雅各 的罪过， 因 以色列 家的罪恶。 雅各 的罪过在哪里呢？ 岂不是在 撒玛利亚 吗？ 犹大 的丘坛在哪里呢？ 岂不是在 耶路撒冷 吗？
MIC|1|6|因此，我必使 撒玛利亚 变为田野的废墟， 用以栽植葡萄； 我必把它的石头倒在山谷， 掀开它的地基。
MIC|1|7|城里一切雕刻的偶像必被打碎， 行淫的赏金全被火烧， 我要毁灭它的一切偶像； 因为从妓女的赏金积聚而来的， 它们仍归为妓女的赏金。
MIC|1|8|为此我要大声哀号， 赤身赤脚行走； 我要呼号如野狗， 哀鸣如鸵鸟。
MIC|1|9|因为 撒玛利亚 的创伤无法医治， 蔓延到 犹大 ， 到了我百姓的城门， 直达 耶路撒冷 。
MIC|1|10|不要在 迦特 宣扬 这事， 千万不要哭泣； 要在 伯．亚弗拉 翻滚于灰尘 中。
MIC|1|11|沙斐 的居民哪，要赤身羞愧地经过， 撒南 的居民不敢出门， 伯．以薛 哀哭，不再支持你们。
MIC|1|12|玛律 的居民心甚忧急，切望得着福气， 因为灾祸已从耶和华那里临到 耶路撒冷 的城门。
MIC|1|13|拉吉 的居民哪，要用快马 套车； 锡安 的罪由你而起， 以色列 的罪过在你那里显出。
MIC|1|14|因此，你要将送别礼送到 摩利设．迦特 ； 亚革悉 的众家族必用诡诈 待 以色列 诸王。
MIC|1|15|玛利沙 的居民哪， 我必使抢夺者来到你这里； 以色列 的贵族 必来到 亚杜兰 。
MIC|1|16|犹大 啊，为了你所喜爱的儿女， 你要剪发，剃光头， 要使你的头光秃，如同秃鹰， 因为他们被掳去离开你了。
MIC|2|1|祸哉，那些在床上图谋罪孽、筹划恶事的人！ 天一亮，他们因手中有能力就去行恶。
MIC|2|2|他们看上田地就占据， 贪图房屋便夺取； 他们欺压户主和他的家庭， 霸占人和他的产业。
MIC|2|3|所以耶和华如此说： 看哪，我筹划灾祸降与这家族； 这灾祸在你们颈项上无法解脱， 你们也不能昂首而行， 因为这是灾祸的时刻。
MIC|2|4|到那日，必有人为你们唱诗歌， 用悲哀的哀歌哀号，说： “我们全然败落， 我百姓的产业易主了！ 耶和华竟然使它离开我， 我们的田地为悖逆的人所瓜分了！”
MIC|2|5|因此，你必无人能在耶和华的会中 抽签拉绳 。
MIC|2|6|他们传讲说：“不可传讲； 人都不可传讲这些事， 羞辱不会临到我们。”
MIC|2|7|雅各 家啊，可这么说吗 ？ 耶和华没有耐心吗？ 这些事是他所行的吗？ 我的言语岂不是与行动正直的人有益吗？
MIC|2|8|然而，近来我的百姓兴起如仇敌。 你们剥去那些安然行路、不愿打仗之人身上的外衣，
MIC|2|9|把我百姓中的妇人从安乐家中赶出， 又将我的荣耀从她们孩子身上永远夺去。
MIC|2|10|起来，走吧！ 这里并非安歇之处； 因为不洁净带来毁坏， 且是大大的毁坏。
MIC|2|11|若有人心存虚假，用谎言说 ： “我向你们传讲可得清酒和烈酒 ”， 那人就必作这百姓的传讲者。
MIC|2|12|雅各 家啊，我定要聚集你们， 定要召集 以色列 的余民， 把他们安置在一处，如 波斯拉 的羊， 又如草场上的羊群， 人数众多，大大喧哗。
MIC|2|13|开路的在他们前面上去， 直闯过城门，从城门出去； 他们的王在前面行， 耶和华在他们的前头。
MIC|3|1|于是我说： 雅各 的领袖， 以色列 家的官长啊， 你们要听！ 你们岂不知道公平吗？
MIC|3|2|你们恶善好恶， 剥我百姓 身上的皮， 从他们的骨头上剔肉，
MIC|3|3|你们吃我百姓的肉， 剥他们的皮， 打断他们的骨头， 如切块 下锅， 如釜中的肉。
MIC|3|4|到了遭灾的时候，这些人要哀求耶和华， 他却不应允他们。 那时，因他们所行的恶， 他必转脸离开他们。
MIC|3|5|论到使我百姓走入歧途的先知， 他们牙齿有所嚼，就呼喊说：“平安！” 谁不给他们吃，就扬言攻击他， 耶和华如此说：
MIC|3|6|你们因此必遭遇黑夜，看不到异象； 遭遇幽暗，无法占卜。 太阳必向先知沉落， 白昼转为黑暗。
MIC|3|7|先见必抱愧， 占卜的必蒙羞， 他们全都捂着胡须， 因为上帝不应允他们。
MIC|3|8|至于我，我藉耶和华的灵， 满有能力、公平和勇气， 可向 雅各 述说他的过犯， 向 以色列 指出他的罪恶。
MIC|3|9|当听这话， 雅各 家的领袖， 以色列 家的官长啊！ 你们厌弃公平， 在一切事上屈枉正直；
MIC|3|10|以血建立 锡安 ， 以罪孽建造 耶路撒冷 。
MIC|3|11|城里的领袖为贿赂行审判， 祭司为酬劳施训诲， 先知为银钱行占卜； 他们却倚赖耶和华，说： “耶和华不是在我们中间吗？ 灾祸必不临到我们。”
MIC|3|12|因此，为你们的缘故， 锡安 要被耕种像一块田地， 耶路撒冷 要变为废墟， 这殿的山必如丛林的高处。
MIC|4|1|末后的日子， 耶和华殿的山必坚立， 超乎诸山，高举过于万岭； 万民都要流归这山。
MIC|4|2|必有许多民族前往，说： “来吧，我们登耶和华的山， 到 雅各 上帝的殿。 他必将他的道指教我们， 我们也要行他的路。” 因为教诲必出于 锡安 ， 耶和华的言语必出于 耶路撒冷 。
MIC|4|3|他必在许多民族中施行审判， 为远方强盛的国断定是非。 他们要将刀打成犁头， 把枪打成镰刀。 这国不举刀攻击那国， 他们也不再学习战事。
MIC|4|4|人人都要坐在自己的葡萄树 和无花果树下， 无人使他们惊吓； 这是万军之耶和华亲口说的。
MIC|4|5|万民都奉自己神明的名行事， 我们却要奉耶和华－我们上帝的名而行， 直到永永远远。
MIC|4|6|耶和华说：在那日， 我必聚集瘸腿的， 召集被赶逐的， 以及我所惩治的人。
MIC|4|7|我要使瘸腿的成为余民， 使被赶到远方的成为强盛之国。 耶和华要在 锡安山 作王治理他们， 从今直到永远。
MIC|4|8|你， 以得台 ， 锡安 的山冈啊， 先前的权柄必归给你， 耶路撒冷 的国权必将归还。
MIC|4|9|现在，你为何大声呼喊呢？ 你中间没有君王， 你的谋士灭绝， 以致疼痛抓住你， 如临产的妇人吗？
MIC|4|10|锡安 哪，你要疼痛生产， 仿佛临产的妇人； 因你必从城里出来，住在田野； 你要到 巴比伦 去， 在那里，你要蒙解救， 在那里，耶和华必救赎你 脱离仇敌的手掌。
MIC|4|11|现在，许多国家聚集攻击你，说： “让 锡安 被玷污！ 让我们亲眼看到！”
MIC|4|12|他们却不知道耶和华的意念， 也不明白他的筹算， 他聚集他们， 像把禾捆聚到禾场。
MIC|4|13|锡安 哪，起来踹谷吧！ 我必使你的角成为铁， 使你的蹄成为铜。 你必打碎许多民族， 将他们的财宝献给耶和华， 将他们的财富献给全地的主。
MIC|5|1|成群的民 哪，现在要聚集成队； 仇敌前来围攻我们， 要用杖击打 以色列 领袖的脸颊。
MIC|5|2|伯利恒 的 以法他 啊， 你在 犹大 诸城中虽小， 将来必有一位从你那里出来， 在 以色列 中为我作掌权者； 他的根源自亘古，从太初就有。
MIC|5|3|因此，耶和华要将 以色列 人交给敌人， 直到临产的妇人生下孩子； 那时，他其余的弟兄 必回到 以色列 人那里。
MIC|5|4|他必倚靠耶和华的大能， 倚靠耶和华－他上帝之名的威严， 站立并牧养， 使他们安然居住； 因为现在他必尊大， 直到地极。
MIC|5|5|这位就是和平 。 当 亚述 侵入我们领土， 践踏我们宫殿时， 我们就立七个牧者， 八个领袖攻击它。
MIC|5|6|他们要用刀剑毁坏 亚述 地 和 宁录 地的关口 。 当 亚述 侵入我们领土， 践踏我们边境时， 他必拯救我们。
MIC|5|7|雅各 的余民 必在许多民族中， 如从耶和华降下的露水， 又如甘霖降在草上； 他们不倚靠人， 也不仰赖世人。
MIC|5|8|雅各 的余民必在列国中， 在许多民族中， 如林间百兽中的狮子， 又如少壮狮子在羊群中； 他若经过就必践踏撕裂， 无人搭救。
MIC|5|9|愿你的手举起，高过敌人！ 愿你的仇敌都被剪除！
MIC|5|10|耶和华说：到那日， 我必从你中间剪除马匹， 毁坏战车；
MIC|5|11|除灭你国中的城镇， 拆毁你一切的堡垒；
MIC|5|12|除掉你手中的邪术， 你那里不再有占卜的人。
MIC|5|13|我必从你中间除灭雕刻的偶像和柱像， 你就不再跪拜自己手所造的；
MIC|5|14|我必从你中间拔除 亚舍拉 ， 毁灭你的城镇；
MIC|5|15|我必在怒气和愤怒中 报应那不听从我的列国。
MIC|6|1|当听耶和华说的话： 起来，向山岭争辩， 使冈陵听见你的声音。
MIC|6|2|山岭啊，要听耶和华的指控！ 大地永久的根基啊，要听！ 因耶和华控告他的百姓， 与 以色列 争辩。
MIC|6|3|“我的百姓啊，我向你做了什么呢？ 我在什么事上使你厌烦？ 你回答我吧！
MIC|6|4|我曾将你从 埃及 地领出来， 从为奴之家救赎你， 我差遣 摩西 、 亚伦 和 米利暗 在你前面带领。
MIC|6|5|我的百姓啊，当记念从前 摩押 王 巴勒 如何筹算， 比珥 的儿子 巴兰 如何回应他， 当记念从 什亭 到 吉甲 所发生的事， 好使你们明白耶和华公义的作为。”
MIC|6|6|“我朝见耶和华， 在至高上帝面前跪拜，当献上什么呢？ 难道献一岁的牛犊为燔祭来朝见他吗？
MIC|6|7|耶和华岂喜悦千千的公羊， 或是万万的油河吗？ 我岂可为自己的过犯献我的长子， 为自己的罪恶献我所亲生的吗？”
MIC|6|8|世人哪，耶和华已指示你何为善。 他向你所要的是什么呢？ 只要你行公义，好怜悯， 存谦卑的心与你的上帝同行。
MIC|6|9|耶和华向这城呼叫 ─看重你的名是真智慧 ─ 你们当听惩罚 和派定惩罚的人 。
MIC|6|10|恶人家中不是仍有不义之财 和惹人生气的变小了的伊法吗？
MIC|6|11|我若用不公道的天平 和袋中诡诈的法码， 岂可算为清白呢？
MIC|6|12|城里的有钱人遍行残暴， 其中的居民说谎话， 口中的舌头尽是诡诈。
MIC|6|13|因此，我也击打你，使你受伤 ， 因你的罪恶使你受惊骇。
MIC|6|14|你要吃，却吃不饱， 你的肚子仍是空空。 你必被挪去，不得逃脱； 如有逃脱的，我必交给刀剑。
MIC|6|15|你撒种，却不得收割； 踹橄榄，却不得油抹身； 有新酒，却不得酒喝。
MIC|6|16|因为你遵守 暗利 的规条， 行 亚哈 家一切所行的， 顺从他们的计谋； 因此，我必使你荒凉， 使你的居民遭人嗤笑， 你们也必担当我百姓的羞辱。
MIC|7|1|我有祸了！我好像夏日收割后的果子， 又如收成之后剩余的葡萄， 没有一挂可吃的， 也没有我心所渴想初熟的无花果。
MIC|7|2|地上的虔诚人灭尽了， 人世间已无正直的人； 他们都埋伏，为要流人的血， 用罗网猎取自己的弟兄。
MIC|7|3|他们双手善于作恶， 君王和审判官都索取贿赂； 位高的人吐出心中的欲望， 彼此勾结 。
MIC|7|4|他们当中最好的，不过像蒺藜； 最正直的，不过如荆棘篱笆。 你守候的日子，惩罚已经来到， 他们必扰乱不安。
MIC|7|5|不可倚赖邻舍， 不可信靠密友； 甚至对躺在你怀中的妻子 也要守住你的口。
MIC|7|6|因为儿子藐视父亲， 女儿抵挡母亲， 媳妇抗拒婆婆， 人的仇敌就是自己家里的人。
MIC|7|7|至于我，我要仰望耶和华， 等候那救我的上帝； 我的上帝必应允我。
MIC|7|8|我的仇敌啊，不要向我夸耀。 我虽跌倒，仍要起来； 虽坐在黑暗里，耶和华却作我的光。
MIC|7|9|我要承受耶和华的恼怒， 直到他为我辩护，为我伸冤， 因我得罪了他； 他要领我进入光明， 我必得见他的公义。
MIC|7|10|那时我的仇敌看见这事就羞愧， 他曾对我说：“耶和华－你的上帝在哪里？” 我必亲眼见他遭报， 现在，他必被践踏，如同街上的泥土。
MIC|7|11|你的城墙重修的日子到了！ 到那日，边界必扩展。
MIC|7|12|到那日，人必从 亚述 ， 从 埃及 的城镇， 从 埃及 到 大河 ， 从这海到那海， 从这山到那山， 都归到你这里。
MIC|7|13|然而，因居民的缘故， 为了他们行事的结果。 这地必然荒凉。
MIC|7|14|求你在 迦密 的树林中， 以你的杖牧放你独居的民， 你产业中的羊群； 愿他们像古时一样， 牧放在 巴珊 和 基列 。
MIC|7|15|我要显奇事给他们看， 好像出 埃及 地的时候一样。
MIC|7|16|列国看见，虽大有势力仍觉惭愧； 他们必用手捂口，掩耳不听。
MIC|7|17|他们要舔土如蛇， 又如地上爬行的动物， 战战兢兢离开他们的营寨； 他们必畏惧耶和华─我们的上帝， 也必因你而害怕。
MIC|7|18|有哪一个神明像你，赦免罪孽， 饶恕他产业中余民的罪过？ 他不永远怀怒，喜爱施恩。
MIC|7|19|他 必转回怜悯我们， 把我们的罪孽踏在脚下。 你必将他们 一切的罪投于深海。
MIC|7|20|你必按古时向我们列祖起誓的话， 以信实待 雅各 ， 向 亚伯拉罕 施慈爱。
