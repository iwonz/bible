1JOHN|1|1|quod fuit ab initio quod audivimus quod vidimus oculis nostris quod perspeximus et manus nostrae temptaverunt de verbo vitae
1JOHN|1|2|et vita manifestata est et vidimus et testamur et adnuntiamus vobis vitam aeternam quae erat apud Patrem et apparuit nobis
1JOHN|1|3|quod vidimus et audivimus adnuntiamus et vobis ut et vos societatem habeatis nobiscum et societas nostra sit cum Patre et cum Filio eius Iesu Christo
1JOHN|1|4|et haec scribimus vobis ut gaudium nostrum sit plenum
1JOHN|1|5|et haec est adnuntiatio quam audivimus ab eo et adnuntiamus vobis quoniam Deus lux est et tenebrae in eo non sunt ullae
1JOHN|1|6|si dixerimus quoniam societatem habemus cum eo et in tenebris ambulamus mentimur et non facimus veritatem
1JOHN|1|7|si autem in luce ambulemus sicut et ipse est in luce societatem habemus ad invicem et sanguis Iesu Filii eius mundat nos ab omni peccato
1JOHN|1|8|si dixerimus quoniam peccatum non habemus ipsi nos seducimus et veritas in nobis non est
1JOHN|1|9|si confiteamur peccata nostra fidelis est et iustus ut remittat nobis peccata et emundet nos ab omni iniquitate
1JOHN|1|10|si dixerimus quoniam non peccavimus mendacem facimus eum et verbum eius non est in nobis
1JOHN|2|1|filioli mei haec scribo vobis ut non peccetis sed et si quis peccaverit advocatum habemus apud Patrem Iesum Christum iustum
1JOHN|2|2|et ipse est propitiatio pro peccatis nostris non pro nostris autem tantum sed etiam pro totius mundi
1JOHN|2|3|et in hoc scimus quoniam cognovimus eum si mandata eius observemus
1JOHN|2|4|qui dicit se nosse eum et mandata eius non custodit mendax est in hoc veritas non est
1JOHN|2|5|qui autem servat verbum eius vere in hoc caritas Dei perfecta est in hoc scimus quoniam in ipso sumus
1JOHN|2|6|qui dicit se in ipso manere debet sicut ille ambulavit et ipse ambulare
1JOHN|2|7|carissimi non mandatum novum scribo vobis sed mandatum vetus quod habuistis ab initio mandatum vetus est verbum quod audistis
1JOHN|2|8|iterum mandatum novum scribo vobis quod est verum et in ipso et in vobis quoniam tenebrae transeunt et lumen verum iam lucet
1JOHN|2|9|qui dicit se in luce esse et fratrem suum odit in tenebris est usque adhuc
1JOHN|2|10|qui diligit fratrem suum in lumine manet et scandalum in eo non est
1JOHN|2|11|qui autem odit fratrem suum in tenebris est et in tenebris ambulat et nescit quo eat quoniam tenebrae obcaecaverunt oculos eius
1JOHN|2|12|scribo vobis filioli quoniam remittuntur vobis peccata propter nomen eius
1JOHN|2|13|scribo vobis patres quoniam cognovistis eum qui ab initio est scribo vobis adulescentes quoniam vicistis malignum
1JOHN|2|14|scripsi vobis infantes quoniam cognovistis Patrem scripsi vobis patres quia cognovistis eum qui ab initio scripsi vobis adulescentes quia fortes estis et verbum Dei in vobis manet et vicistis malignum
1JOHN|2|15|nolite diligere mundum neque ea quae in mundo sunt si quis diligit mundum non est caritas Patris in eo
1JOHN|2|16|quoniam omne quod est in mundo concupiscentia carnis et concupiscentia oculorum est et superbia vitae quae non est ex Patre sed ex mundo est
1JOHN|2|17|et mundus transit et concupiscentia eius qui autem facit voluntatem Dei manet in aeternum
1JOHN|2|18|filioli novissima hora est et sicut audistis quia antichristus venit nunc antichristi multi facti sunt unde scimus quoniam novissima hora est
1JOHN|2|19|ex nobis prodierunt sed non erant ex nobis nam si fuissent ex nobis permansissent utique nobiscum sed ut manifesti sint quoniam non sunt omnes ex nobis
1JOHN|2|20|sed vos unctionem habetis a Sancto et nostis omnia
1JOHN|2|21|non scripsi vobis quasi ignorantibus veritatem sed quasi scientibus eam et quoniam omne mendacium ex veritate non est
1JOHN|2|22|quis est mendax nisi is qui negat quoniam Iesus non est Christus hic est antichristus qui negat Patrem et Filium
1JOHN|2|23|omnis qui negat Filium nec Patrem habet qui confitetur Filium et Patrem habet
1JOHN|2|24|vos quod audistis ab initio in vobis permaneat si in vobis permanserit quod ab initio audistis et vos in Filio et Patre manebitis
1JOHN|2|25|et haec est repromissio quam ipse pollicitus est nobis vitam aeternam
1JOHN|2|26|haec scripsi vobis de eis qui seducunt vos
1JOHN|2|27|et vos unctionem quam accepistis ab eo manet in vobis et non necesse habetis ut aliquis doceat vos sed sicut unctio eius docet vos de omnibus et verum est et non est mendacium et sicut docuit vos manete in eo
1JOHN|2|28|et nunc filioli manete in eo ut cum apparuerit habeamus fiduciam et non confundamur ab eo in adventu eius
1JOHN|2|29|si scitis quoniam iustus est scitote quoniam et omnis qui facit iustitiam ex ipso natus est
1JOHN|3|1|videte qualem caritatem dedit nobis Pater ut filii Dei nominemur et sumus propter hoc mundus non novit nos quia non novit eum
1JOHN|3|2|carissimi nunc filii Dei sumus et nondum apparuit quid erimus scimus quoniam cum apparuerit similes ei erimus quoniam videbimus eum sicuti est
1JOHN|3|3|et omnis qui habet spem hanc in eo sanctificat se sicut et ille sanctus est
1JOHN|3|4|omnis qui facit peccatum et iniquitatem facit et peccatum est iniquitas
1JOHN|3|5|et scitis quoniam ille apparuit ut peccata tolleret et peccatum in eo non est
1JOHN|3|6|omnis qui in eo manet non peccat omnis qui peccat non vidit eum nec cognovit eum
1JOHN|3|7|filioli nemo vos seducat qui facit iustitiam iustus est sicut et ille iustus est
1JOHN|3|8|qui facit peccatum ex diabolo est quoniam ab initio diabolus peccat in hoc apparuit Filius Dei ut dissolvat opera diaboli
1JOHN|3|9|omnis qui natus est ex Deo peccatum non facit quoniam semen ipsius in eo manet et non potest peccare quoniam ex Deo natus est
1JOHN|3|10|in hoc manifesti sunt filii Dei et filii diaboli omnis qui non est iustus non est de Deo et qui non diligit fratrem suum
1JOHN|3|11|quoniam haec est adnuntiatio quam audistis ab initio ut diligamus alterutrum
1JOHN|3|12|non sicut Cain ex maligno erat et occidit fratrem suum et propter quid occidit eum quoniam opera eius maligna erant fratris autem eius iusta
1JOHN|3|13|nolite mirari fratres si odit vos mundus
1JOHN|3|14|nos scimus quoniam translati sumus de morte in vitam quoniam diligimus fratres qui non diligit manet in morte
1JOHN|3|15|omnis qui odit fratrem suum homicida est et scitis quoniam omnis homicida non habet vitam aeternam in se manentem
1JOHN|3|16|in hoc cognovimus caritatem quoniam ille pro nobis animam suam posuit et nos debemus pro fratribus animas ponere
1JOHN|3|17|qui habuerit substantiam mundi et viderit fratrem suum necesse habere et clauserit viscera sua ab eo quomodo caritas Dei manet in eo
1JOHN|3|18|filioli non diligamus verbo nec lingua sed opere et veritate
1JOHN|3|19|in hoc cognoscimus quoniam ex veritate sumus et in conspectu eius suadeamus corda nostra
1JOHN|3|20|quoniam si reprehenderit nos cor maior est Deus corde nostro et novit omnia
1JOHN|3|21|carissimi si cor non reprehenderit nos fiduciam habemus ad Deum
1JOHN|3|22|et quodcumque petierimus accipiemus ab eo quoniam mandata eius custodimus et ea quae sunt placita coram eo facimus
1JOHN|3|23|et hoc est mandatum eius ut credamus in nomine Filii eius Iesu Christi et diligamus alterutrum sicut dedit mandatum nobis
1JOHN|3|24|et qui servat mandata eius in illo manet et ipse in eo et in hoc scimus quoniam manet in nobis de Spiritu quem nobis dedit
1JOHN|4|1|carissimi nolite omni spiritui credere sed probate spiritus si ex Deo sint quoniam multi pseudoprophetae exierunt in mundum
1JOHN|4|2|in hoc cognoscitur Spiritus Dei omnis spiritus qui confitetur Iesum Christum in carne venisse ex Deo est
1JOHN|4|3|et omnis spiritus qui solvit Iesum ex Deo non est et hoc est antichristi quod audistis quoniam venit et nunc iam in mundo est
1JOHN|4|4|vos ex Deo estis filioli et vicistis eos quoniam maior est qui in vobis est quam qui in mundo
1JOHN|4|5|ipsi de mundo sunt ideo de mundo loquuntur et mundus eos audit
1JOHN|4|6|nos ex Deo sumus qui novit Deum audit nos qui non est ex Deo non audit nos in hoc cognoscimus Spiritum veritatis et spiritum erroris
1JOHN|4|7|carissimi diligamus invicem quoniam caritas ex Deo est et omnis qui diligit ex Deo natus est et cognoscit Deum
1JOHN|4|8|qui non diligit non novit Deum quoniam Deus caritas est
1JOHN|4|9|in hoc apparuit caritas Dei in nobis quoniam Filium suum unigenitum misit Deus in mundum ut vivamus per eum
1JOHN|4|10|in hoc est caritas non quasi nos dilexerimus Deum sed quoniam ipse dilexit nos et misit Filium suum propitiationem pro peccatis nostris
1JOHN|4|11|carissimi si sic Deus dilexit nos et nos debemus alterutrum diligere
1JOHN|4|12|Deum nemo vidit umquam si diligamus invicem Deus in nobis manet et caritas eius in nobis perfecta est
1JOHN|4|13|in hoc intellegimus quoniam in eo manemus et ipse in nobis quoniam de Spiritu suo dedit nobis
1JOHN|4|14|et nos vidimus et testificamur quoniam Pater misit Filium salvatorem mundi
1JOHN|4|15|quisque confessus fuerit quoniam Iesus est Filius Dei Deus in eo manet et ipse in Deo
1JOHN|4|16|et nos cognovimus et credidimus caritati quam habet Deus in nobis Deus caritas est et qui manet in caritate in Deo manet et Deus in eo
1JOHN|4|17|in hoc perfecta est caritas nobiscum ut fiduciam habeamus in die iudicii quia sicut ille est et nos sumus in hoc mundo
1JOHN|4|18|timor non est in caritate sed perfecta caritas foras mittit timorem quoniam timor poenam habet qui autem timet non est perfectus in caritate
1JOHN|4|19|nos ergo diligamus quoniam Deus prior dilexit nos
1JOHN|4|20|si quis dixerit quoniam diligo Deum et fratrem suum oderit mendax est qui enim non diligit fratrem suum quem vidit Deum quem non vidit quomodo potest diligere
1JOHN|4|21|et hoc mandatum habemus ab eo ut qui diligit Deum diligat et fratrem suum
1JOHN|5|1|omnis qui credit quoniam Iesus est Christus ex Deo natus est et omnis qui diligit eum qui genuit diligit eum qui natus est ex eo
1JOHN|5|2|in hoc cognoscimus quoniam diligimus natos Dei cum Deum diligamus et mandata eius faciamus
1JOHN|5|3|haec est enim caritas Dei ut mandata eius custodiamus et mandata eius gravia non sunt
1JOHN|5|4|quoniam omne quod natum est ex Deo vincit mundum et haec est victoria quae vincit mundum fides nostra
1JOHN|5|5|quis est qui vincit mundum nisi qui credit quoniam Iesus est Filius Dei
1JOHN|5|6|hic est qui venit per aquam et sanguinem Iesus Christus non in aqua solum sed in aqua et sanguine et Spiritus est qui testificatur quoniam Christus est veritas
1JOHN|5|7|quia tres sunt qui testimonium dant
1JOHN|5|8|Spiritus et aqua et sanguis et tres unum sunt
1JOHN|5|9|si testimonium hominum accipimus testimonium Dei maius est quoniam hoc est testimonium Dei quod maius est quia testificatus est de Filio suo
1JOHN|5|10|qui credit in Filio Dei habet testimonium Dei in se qui non credit Filio mendacem facit eum quoniam non credidit in testimonio quod testificatus est Deus de Filio suo
1JOHN|5|11|et hoc est testimonium quoniam vitam aeternam dedit nobis Deus et haec vita in Filio eius est
1JOHN|5|12|qui habet Filium habet vitam qui non habet Filium Dei vitam non habet
1JOHN|5|13|haec scripsi vobis ut sciatis quoniam vitam habetis aeternam qui creditis in nomine Filii Dei
1JOHN|5|14|et haec est fiducia quam habemus ad eum quia quodcumque petierimus secundum voluntatem eius audit nos
1JOHN|5|15|et scimus quoniam audit nos quicquid petierimus scimus quoniam habemus petitiones quas postulavimus ab eo
1JOHN|5|16|qui scit fratrem suum peccare peccatum non ad mortem petet et dabit ei vitam peccantibus non ad mortem est peccatum ad mortem non pro illo dico ut roget
1JOHN|5|17|omnis iniquitas peccatum est et est peccatum non ad mortem
1JOHN|5|18|scimus quoniam omnis qui natus est ex Deo non peccat sed generatio Dei conservat eum et malignus non tangit eum
1JOHN|5|19|scimus quoniam ex Deo sumus et mundus totus in maligno positus est
1JOHN|5|20|et scimus quoniam Filius Dei venit et dedit nobis sensum ut cognoscamus verum Deum et simus in vero Filio eius hic est verus Deus et vita aeterna
1JOHN|5|21|filioli custodite vos a simulacris
