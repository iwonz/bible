ESTH|1|1|这事发生在 亚哈随鲁 的时代， 亚哈随鲁 从 印度 直到 古实 统治一百二十七个省，
ESTH|1|2|就是 亚哈随鲁 王在 书珊 城堡中坐国度王位的那些日子。
ESTH|1|3|他在位第三年，为所有官员和臣仆摆设宴席，有 波斯 和 玛代 的权贵，各省的贵族与领袖在他面前。
ESTH|1|4|他把他荣耀国度的丰富和他伟大威严的尊贵给他们看了许多日子，共一百八十天。
ESTH|1|5|这些日子满了，王又为所有住 书珊 城堡的百姓，无论大小，在御花园的院子里摆设宴席七日。
ESTH|1|6|院子里有白色棉和蓝色线，用细麻绳、紫色绳系在白玉石柱的银环上，又有金银的床榻摆在红、白、黄、黑大理石镶嵌的地上。
ESTH|1|7|用金器皿盛酒，有很多不同的器皿，照王的厚意提供丰富的御酒。
ESTH|1|8|饮酒有规定，不准勉强人 ，因为王吩咐宫里所有的臣宰，让人各随己意。
ESTH|1|9|瓦实提 王后在 亚哈随鲁 王的宫内也为妇女摆设宴席。
ESTH|1|10|第七日， 亚哈随鲁 王饮酒，心中快乐，就吩咐在他面前侍立的七个太监 米户幔 、 比斯他 、 哈波拿 、 比革他 、 亚拔他 、 西达 、 甲迦 ，
ESTH|1|11|请 瓦实提 王后头戴王后的冠冕到王面前，让各民族和官员观看她的美貌，因为她容貌美丽。
ESTH|1|12|瓦实提 王后却不肯遵照太监所传的王命前来，所以王非常愤怒，怒火中烧。
ESTH|1|13|按王的常规，办事必先询问知例明法的人。那时，王询问通达时务的智慧人，
ESTH|1|14|就是在王左右常见王面、在国中坐高位的 波斯 和 玛代 的七个大臣， 甲示拿 、 示达 、 押玛他 、 他施斯 、 米力 、 玛西拿 、 米慕干 ：
ESTH|1|15|“ 瓦实提 王后不遵照太监所传的王命，照例应当怎样办理呢？”
ESTH|1|16|米慕干 在王和众官长面前回答说：“ 瓦实提 王后这事，不但得罪王，并且有害于 亚哈随鲁 王各省的臣民。
ESTH|1|17|因为王后这事必传到众妇人那里，她们就会藐视自己的丈夫，说：‘ 亚哈随鲁 王吩咐 瓦实提 王后到王面前，她却不来。’
ESTH|1|18|今日 波斯 和 玛代 的众夫人听见王后这事，必向王所有的官长照样说，如此必造成无数的藐视和愤怒。
ESTH|1|19|王若以为好，请降谕旨，写在 波斯 和 玛代 人的条例中，永不更改，不准 瓦实提 再到 亚哈随鲁 王面前，把她王后的位分赐给比她更好的妃子。
ESTH|1|20|王的谕旨一传遍全国，国土纵然辽阔，凡作妻子的，无论丈夫是尊贵或卑贱，都必尊敬他。”
ESTH|1|21|王和众官长都以这话为美，王就照 米慕干 的建议去做。
ESTH|1|22|王下诏书，用各省的文字、各族的语言通知各省，使凡作丈夫的在家中作主，各说本地的语言 。
ESTH|2|1|这些事以后， 亚哈随鲁 王的愤怒平息，就想起 瓦实提 和她所做的，以及自己怎样降旨办她。
ESTH|2|2|于是王的侍臣对王说：“请派人为王寻找美貌的少女；
ESTH|2|3|请王派官员在国中各省招聚所有美貌的少女到 书珊 城堡的女院，交给王所派掌管女子的太监 希该 ，给她们香膏涂抹。
ESTH|2|4|王眼中看为好的女子可以立为王后，代替 瓦实提 。”王以这话为美，就照样做。
ESTH|2|5|书珊 城堡中有一个 犹太 人名叫 末底改 ，是 便雅悯 人 基士 的曾孙， 示每 的孙子， 睚珥 的儿子。
ESTH|2|6|从前 巴比伦 王 尼布甲尼撒 把 犹大 王 耶哥尼雅 和百姓从 耶路撒冷 掳来， 末底改 也在被掳的人当中。
ESTH|2|7|末底改 抚养他叔叔的女儿 哈大沙 ，就是 以斯帖 ，因为她没有父母。这女子容貌美丽；她父母死了， 末底改 收她为自己的女儿。
ESTH|2|8|王的谕旨和敕令传出之后，许多女子被招聚到 书珊 城堡，交给掌管女子的 希该 ； 以斯帖 也被送入王宫，交给 希该 。
ESTH|2|9|希该 眼中宠爱 以斯帖 ，就恩待她，急忙给她涂抹的香膏和当得的份，又从王宫里挑选七个宫女来服事她，使她和她的宫女搬入女院上好的房屋。
ESTH|2|10|以斯帖 未曾将自己的籍贯宗族告诉人，因为 末底改 嘱咐她不可叫人知道。
ESTH|2|11|末底改 天天在女院前徘徊，要知道 以斯帖 是否平安，过得如何。
ESTH|2|12|众女子照例先涂抹身体十二个月：六个月用没药油，六个月用香料和涂抹的香膏。满了日期，每个女子挨次进去朝见 亚哈随鲁 王。
ESTH|2|13|女子进去朝见王是这样：从女院到王宫的时候，凡她所要的都必给她带进去。
ESTH|2|14|晚上她进去，次日回到另一个女院，交给掌管妃嫔的太监 沙甲 。除非王喜爱她，再提名召她，她就不再进去见王。
ESTH|2|15|末底改 的叔叔 亚比孩 的女儿，就是 末底改 收为自己女儿的 以斯帖 ，按次序要进去朝见王的时候，除了掌管女子的太监 希该 所分派给她的，她别无所求。凡看见 以斯帖 的都喜欢她。
ESTH|2|16|亚哈随鲁 王第七年十月，就是提别月， 以斯帖 被引入宫中朝见王。
ESTH|2|17|王爱 以斯帖 过于众女子，她在王面前蒙宠爱胜过众少女。王把王后的冠冕戴在她头上，立她为王后，代替 瓦实提 。
ESTH|2|18|王为所有的官长和臣仆摆设大宴席，称为 以斯帖 的宴席，又豁免各省的租税，并照王的厚意大颁赏赐。
ESTH|2|19|第二次招聚少女的时候， 末底改 坐在朝门。
ESTH|2|20|以斯帖 遵照 末底改 所嘱咐的，没有将籍贯宗族告诉人； 以斯帖 照 末底改 的吩咐去做，正如受他抚养的时候一样。
ESTH|2|21|那时候， 末底改 坐在朝门，王有两个守门的太监， 辟探 和 提列 ，恼恨 亚哈随鲁 王，想要下手害他。
ESTH|2|22|末底改 知道了这件事，就告诉 以斯帖 王后。 以斯帖 以 末底改 的名向王报告。
ESTH|2|23|这事经过查究后发现是真的，二人就被挂在木头上。这事在王面前记录在史籍上。
ESTH|3|1|这些事以后， 亚哈随鲁 王使 亚甲 人 哈米大他 的儿子 哈曼 尊大，提升了他，叫他的爵位超过所有与他同朝的官长。
ESTH|3|2|在朝门，王所有的臣仆都跪拜 哈曼 ，因为王如此吩咐，但 末底改 不跪不拜。
ESTH|3|3|在朝门，王的臣仆对 末底改 说：“你为何违背王的命令呢？”
ESTH|3|4|他们天天劝他，他还是不听，他们就告诉 哈曼 ，要看 末底改 的事是否站得住，因他已经告诉他们自己是 犹太 人。
ESTH|3|5|哈曼 见 末底改 不跪不拜，就非常愤怒。
ESTH|3|6|有人把 末底改 的宗族告诉 哈曼 。 哈曼 看下手只害 末底改 一人是小事，还图谋要灭绝 亚哈随鲁 王全国所有的 犹太 人，就是 末底改 的宗族。
ESTH|3|7|亚哈随鲁 王十二年正月，就是尼散月，人在 哈曼 面前抽普珥，普珥即签，要定何月何日；抽到了十二月，就是亚达月。
ESTH|3|8|哈曼 对 亚哈随鲁 王说：“有一民族散居在王国各省的民族中，与众不同；他们的律例与万民的律例不同，也不守王的律例，所以容留他们对王无益。
ESTH|3|9|王若以为好，请下谕旨灭绝他们，我就捐一万他连得银子交给管财政的人，纳入王的府库。”
ESTH|3|10|于是王从自己手上摘下戒指给 犹太 人的仇敌， 亚甲 人 哈米大他 的儿子 哈曼 。
ESTH|3|11|王对 哈曼 说：“这银子赐给你，这民族也交给你，可以照你眼中看为好的待他们。”
ESTH|3|12|正月十三日，王的一些书记受召而来，照着 哈曼 一切所吩咐的，用各省的文字、各族的语言，奉 亚哈随鲁 王的名写谕旨，又用王的戒指盖印，传给王的总督、各省的省长，以及各族的领袖。
ESTH|3|13|诏书由信差传到王的各省，限令一日之内，就是在十二月，亚达月十三日，把所有的 犹太 人，无论老少妇女孩子，全然剪除，杀戮灭绝，并抢夺他们的财产。
ESTH|3|14|这谕旨的抄本以敕令的方式在各省颁布，通知各族，预备等候那日。
ESTH|3|15|信差奉王的命令急忙起行，敕令传遍了 书珊 城堡。王同 哈曼 坐下饮酒， 书珊 城堡却陷入慌乱中。
ESTH|4|1|末底改 知道所发生的这一切事，就撕裂衣服，披麻蒙灰，在城中行走，痛哭哀号。
ESTH|4|2|他到了朝门前就停住脚步，因为穿麻衣的不可进朝门。
ESTH|4|3|王的谕旨和敕令所到的各省各处， 犹太 人都极其悲哀，禁食哭泣哀号，许多人躺在麻布和炉灰中。
ESTH|4|4|以斯帖 王后的宫女和太监来把这事告诉 以斯帖 ，她非常忧愁，就送衣服给 末底改 穿，要他脱下身上的麻衣，他却不肯接受。
ESTH|4|5|以斯帖 把王所派伺候她的一个太监 哈他革 召来，吩咐他去见 末底改 ，要知道到底发生了什么事，为何如此。
ESTH|4|6|于是 哈他革 出来，到朝门前的广场见 末底改 。
ESTH|4|7|末底改 把自己遭遇的一切，以及 哈曼 为灭绝 犹太 人答应捐入王库的银数都告诉了他；
ESTH|4|8|又把那传遍 书珊 、要灭绝 犹太 人的谕旨抄本交给 哈他革 ，要他给 以斯帖 看，并向她说明，嘱咐她去晋见王，向王恳求，为本族的人在王面前请命。
ESTH|4|9|哈他革 回来，把 末底改 的话告诉 以斯帖 。
ESTH|4|10|以斯帖 吩咐 哈他革 去见 末底改 ，说：
ESTH|4|11|“王所有的臣仆和各省的百姓都知道有一个定例，若未奉召见，擅入内院见王的，无论男女必被处死；除非王向他伸出金杖，不得存活。但我没有被召进去见王已经有三十天了。”
ESTH|4|12|他们把 以斯帖 的话告诉 末底改 。
ESTH|4|13|末底改 托人回覆 以斯帖 说：“你不要自己以为在王宫里强过任何 犹太 人，得以幸免。
ESTH|4|14|此时你若闭口不言， 犹太 人必从别处得解脱，蒙拯救；你和你父家必致灭亡。焉知你得了王后的位分不是为现今的机会吗？”
ESTH|4|15|以斯帖 吩咐人回覆 末底改 说：
ESTH|4|16|“你当去召集 书珊 所有的 犹太 人，为我禁食三昼三夜，不吃不喝；我和我的宫女也要这样禁食。然后我违例去晋见王，我若死就死吧！”
ESTH|4|17|于是 末底改 照 以斯帖 一切所吩咐的去做。
ESTH|5|1|第三日， 以斯帖 穿上朝服，站立在王宫的内院，对着王宫。王在殿里坐在宝座上，对着殿的门。
ESTH|5|2|王见 以斯帖 王后站在院内，她在王的眼中得恩宠，王向她伸出手中的金杖。 以斯帖 往前去摸杖头。
ESTH|5|3|王对她说：“ 以斯帖 王后啊，你要什么？无论你求什么，就是国的一半也必赐给你。”
ESTH|5|4|以斯帖 说：“王若以为好，请王带着 哈曼 今日赴我为王预备的宴席。”
ESTH|5|5|王说：“叫 哈曼 速速照 以斯帖 的话去做。”于是王带着 哈曼 赴 以斯帖 所预备的宴席。
ESTH|5|6|在宴席喝酒的时候，王又对 以斯帖 说：“你要什么，必赐给你；无论你求什么，就是国的一半也必给你。”
ESTH|5|7|以斯帖 回答说：“我所要的、我所求的，嗯......。
ESTH|5|8|我若在王眼前蒙恩，王若愿意赐我所要的，准我所求的，就请王和 哈曼 再赴我为你们预备的宴席。明日我必照王的话去做。”
ESTH|5|9|那日 哈曼 心中快乐，欢欢喜喜地出来。但是当他看见 末底改 在朝门不站起来，也不因他动一下，就满心恼怒 末底改 。
ESTH|5|10|哈曼 忍着气回家，叫人请他的一些朋友和他妻子 细利斯 来。
ESTH|5|11|哈曼 将他的荣华富贵、众多的儿女，和王使他尊大、提升他高过官长和臣仆的事，都述说给他们听。
ESTH|5|12|哈曼 又说：“ 以斯帖 王后预备宴席，除了我之外不许别人随王赴席。明日王后又请我随王赴席。
ESTH|5|13|只是每当我看见 犹太 人 末底改 坐在朝门，这一切对我就都毫无意义了。”
ESTH|5|14|他的妻子 细利斯 和他所有的朋友对他说：“叫人做一个五十肘高的木架，早晨求王把 末底改 挂在其上，然后你可以欢欢喜喜随王赴席。” 哈曼 认为这话很好，就叫人做了木架。
ESTH|6|1|那夜王睡不着觉，吩咐人取历史书，就是史籍，念给他听，
ESTH|6|2|发现书上写着：王有两个守门的太监 辟探 和 提列 ，想要下手害 亚哈随鲁 王， 末底改 告发了这件事。
ESTH|6|3|王说：“ 末底改 做了这事，有没有赐给他什么尊荣或高位呢？”伺候王的臣仆说：“没有赐给他什么。”
ESTH|6|4|王说：“谁在院子里？”那时 哈曼 正进入王宫的外院，要请王把 末底改 挂在他所预备的木架上。
ESTH|6|5|王的臣仆对他说：“看哪， 哈曼 站在院子里。”王说：“叫他进来。”
ESTH|6|6|哈曼 就进去。王对他说：“王所喜爱要赐尊荣的人，当如何待他呢？” 哈曼 心里说：“王所喜爱要赐尊荣的人，除了我，还有谁呢？”
ESTH|6|7|哈曼 就对王说：“王所喜爱要赐尊荣的人，
ESTH|6|8|当把王所穿的王袍拿来，牵了戴冠的御马，
ESTH|6|9|把王袍和御马都交给王一个极尊贵的大臣，吩咐人把王袍给王所喜爱要赐尊荣的人穿上，领他骑着御马走遍城里的广场，在他面前宣告：‘王所喜爱要赐尊荣的人，就是这样待他。’”
ESTH|6|10|王对 哈曼 说：“你速速把这王袍和御马，照你所说的，向坐在朝门的 犹太 人 末底改 去做。凡你所说的，一样都不可缺。”
ESTH|6|11|于是 哈曼 把王袍给 末底改 穿上，领他骑着御马走遍城里的广场，在他面前宣告：“王所喜爱要赐尊荣的人，就是这样待他。”
ESTH|6|12|末底改 仍回到朝门， 哈曼 却忧忧闷闷地蒙着头，急忙回家去了。
ESTH|6|13|哈曼 把所遭遇的一切都说给他妻子 细利斯 和他所有的朋友听。他的智囊团和他的妻子 细利斯 对他说：“你在 末底改 面前开始败落；他既是 犹太 人，你必不能胜过他，终必在他面前败落。”
ESTH|6|14|他们正跟 哈曼 说话的时候，王的几位太监来了，催 哈曼 快去赴 以斯帖 所预备的宴席。
ESTH|7|1|王带着 哈曼 来赴 以斯帖 王后的宴席。
ESTH|7|2|第二天在宴席喝酒的时候，王又对 以斯帖 说：“ 以斯帖 王后啊，你要什么，必赐给你；无论你求什么，就是国的一半也必给你。”
ESTH|7|3|以斯帖 王后回答说：“王啊，我若在你眼前蒙恩，王若以为好，我所要的，是王把我的性命赐给我；我所求的，是求我的本族。
ESTH|7|4|因为我和我的本族被出卖了，要被剪除，杀戮，灭绝。我们若被卖为奴为婢，我就闭口不言；但我们的痛苦比起王的损失，算不得什么 。”
ESTH|7|5|亚哈随鲁 王问 以斯帖 王后说：“擅敢起意如此行的是谁？这人在哪里呢？”
ESTH|7|6|以斯帖 说：“仇人敌人就是这恶人 哈曼 ！” 哈曼 在王和王后面前非常惊惶。
ESTH|7|7|王大怒，起来离开酒席往御花园去了。 哈曼 见王定意要加罪于他，就留下来求 以斯帖 王后救他的命。
ESTH|7|8|王从御花园回到酒席厅，见 哈曼 伏在 以斯帖 所靠的榻上；王说：“他竟敢在宫内、在我面前凌辱王后吗？”这话一出王口， 哈曼 的脸就被蒙住了。
ESTH|7|9|有一个伺候王名叫 哈波拿 的太监说：“看哪， 哈曼 还为那报告给王、救王有功的 末底改 做了一个五十肘高的木架，现今立在 哈曼 的家里。”王说：“把 哈曼 挂在木架上。”
ESTH|7|10|于是 哈曼 被挂在他为 末底改 所预备的木架上；王的愤怒才平息了。
ESTH|8|1|那日， 亚哈随鲁 王把 犹太 人的仇敌 哈曼 的家产赐给 以斯帖 王后。 末底改 也来到王面前，因为 以斯帖 已经告诉王， 末底改 跟她是什么关系。
ESTH|8|2|王摘下自己的戒指，就是从 哈曼 取回的，给了 末底改 。 以斯帖 派 末底改 管理 哈曼 的家产。
ESTH|8|3|以斯帖 又在王面前求情，俯伏在他脚前，流泪哀求他阻止 亚甲 人 哈曼 害 犹太 人的恶谋。
ESTH|8|4|王向 以斯帖 伸出金杖， 以斯帖 就起来，站在王面前，
ESTH|8|5|说：“王若以为好，我若在王面前蒙恩，王若认为合宜，我若在王眼前得喜悦，请王下谕旨，废除 亚甲 人 哈米大他 的儿子 哈曼 设谋，要杀灭王各省的 犹太 人所颁的诏书。
ESTH|8|6|我何忍见我本族的人受害？何忍见我同宗的人被灭呢？”
ESTH|8|7|亚哈随鲁 王对 以斯帖 王后和 犹太 人 末底改 说：“因为 哈曼 要下手害 犹太 人，看哪，我已把他的家产赐给 以斯帖 ，也把 哈曼 挂在木架上了。
ESTH|8|8|你们可以照你们看为好的，奉王的名写谕旨给 犹太 人，用王的戒指盖印；因为奉王的名所写、用王的戒指盖印的谕旨是不能废除的。”
ESTH|8|9|三月，就是西弯月二十三日，当时王的一些书记受召而来，按着 末底改 所吩咐的，用各省的文字、各族的语言，以及 犹太 人的文字语言写谕旨，传给那从 印度 直到 古实 一百二十七省的 犹太 人，以及总督、省长和领袖。
ESTH|8|10|末底改 奉 亚哈随鲁 王的名写谕旨，用王的戒指盖印，交给信差们骑上御用的王室快马去颁布。
ESTH|8|11|王准各城各镇的 犹太 人在一日之内，在十二月，就是亚达月的十三日聚集，在 亚哈随鲁 王的各省保护自己的性命，剪除，杀戮，灭绝那要攻击 犹太 人的各省各族所有的军队，以及他们的妻子儿女，夺取他们的财产为掠物。
ESTH|8|12|
ESTH|8|13|这谕旨的抄本以敕令的方式在各省颁布，通知各族，使 犹太 人预备等候那日，好在仇敌身上报仇。
ESTH|8|14|于是骑御用快马的信差奉王命催促，急忙起行；敕令传遍了 书珊 城堡。
ESTH|8|15|末底改 穿着蓝色白色的朝服，头戴大金冠冕，又穿紫色细麻布的外袍，从王面前出来； 书珊城 充满了欢乐的呼声。
ESTH|8|16|犹太 人有光荣，欢喜快乐，得享尊贵。
ESTH|8|17|王的谕旨和敕令所到的各省各城， 犹太 人都欢喜快乐，摆设宴席，以那日为吉日。国中许多民族的人因惧怕 犹太 人，就自称为 犹太 人。
ESTH|9|1|十二月，就是亚达月十三日，王的谕旨和敕令要执行的那一日， 犹太 人的仇敌盼望制伏他们，但 犹太 人反倒制伏了恨他们的人。
ESTH|9|2|犹太 人在 亚哈随鲁 王各省的城里聚集，下手击杀那些要害他们的人。没有人能在他们面前站立得住，因为各民族都惧怕他们。
ESTH|9|3|各省的领袖、总督、省长，和办理王事务的人，因惧怕 末底改 ，就都帮助 犹太 人。
ESTH|9|4|末底改 在朝中为大，名声传遍各省； 末底改 这人的权势日渐扩大。
ESTH|9|5|犹太 人用刀击杀所有的仇敌，杀灭他们，随意待那些恨他们的人。
ESTH|9|6|在 书珊 城堡中， 犹太 人杀灭了五百人。
ESTH|9|7|他们杀了 巴珊大他 、 达分 、 亚斯帕他 、
ESTH|9|8|破拉他 、 亚大利雅 、 亚利大他 、
ESTH|9|9|帕玛斯他 、 亚利赛 、 亚利代 、 瓦耶撒他 ；
ESTH|9|10|这十人都是 哈米大他 的孙子， 犹太 人的仇敌 哈曼 的儿子。 犹太 人却没有下手夺取财物。
ESTH|9|11|那日， 书珊 城堡中被杀的人数呈报到王面前。
ESTH|9|12|王对 以斯帖 王后说：“ 犹太 人在 书珊 城堡中杀灭了五百人，又杀了 哈曼 的十个儿子，在王其余的各省不知如何。你要什么，必赐给你；你还求什么，也必为你成就。”
ESTH|9|13|以斯帖 说：“王若以为好，求你允准 书珊 的 犹太 人，明日也照今日的谕旨去做，并把 哈曼 十个儿子的尸体挂在木架上。”
ESTH|9|14|王允准这么做。敕令传遍 书珊 ， 哈曼 十个儿子的尸体被挂了起来。
ESTH|9|15|亚达月十四日，在 书珊 的 犹太 人又聚集，在 书珊 杀了三百人，却没有下手夺取财物。
ESTH|9|16|亚达月十三日，在王各省其余的 犹太 人也都聚集，保护自己的性命，摆脱仇敌得享平安。他们杀了七万五千个恨他们的人，却没有下手夺取财物；十四日他们休息，以这日为设宴欢乐的日子。
ESTH|9|17|
ESTH|9|18|但 书珊 的 犹太 人却在十三日、十四日聚集；十五日休息，以这日为设宴欢乐的日子。
ESTH|9|19|所以住在无城墙的乡村的 犹太 人，都以亚达月十四日为设宴欢乐的吉日，彼此馈送礼物。
ESTH|9|20|末底改 记录这些事，写信给 亚哈随鲁 王各省远近所有的 犹太 人，
ESTH|9|21|吩咐他们每年守亚达月十四、十五两日，
ESTH|9|22|以这两日为 犹太 人摆脱仇敌得享平安、转忧为喜、转悲为乐的吉日，并在这两日设宴欢乐，彼此馈送礼物，赒济穷人。
ESTH|9|23|于是， 犹太 人照 末底改 所写给他们的，把开始所做的作为遵守的定例。
ESTH|9|24|因为 犹太 人的仇敌 亚甲 人 哈米大他 的儿子 哈曼 设谋要杀害 犹太 人，抽普珥，普珥即签，为要杀尽灭绝他们；
ESTH|9|25|但这阴谋 到了王面前，王却降旨使 哈曼 谋害 犹太 人的恶事归到他自己的头上，他和他的众子都被挂在木架上。
ESTH|9|26|所以 犹太 人照着普珥这名字称这两日为普珥日。他们因这信上一切的话，又因所看见所遇见的事，
ESTH|9|27|就规定自己与后裔，以及归化他们的人，每年按所写的、按时守这两日，永久不废。
ESTH|9|28|各省各城、世世代代、家家户户都记念并守这两日，使这普珥日在 犹太 人中不可废掉，在他们后裔中也永不遗忘。
ESTH|9|29|亚比孩 的女儿 以斯帖 王后和 犹太 人 末底改 以全权写第二封信，坚立这普珥日，
ESTH|9|30|送信给 亚哈随鲁 王国中一百二十七省所有的 犹太 人，祝他们平安和安稳，
ESTH|9|31|劝他们遵照 犹太 人 末底改 和 以斯帖 王后所规定的，按时守这普珥日，并照着 犹太 人为自己与后裔所规定的，禁食与哀求。
ESTH|9|32|以斯帖 规定了守普珥日的条例，这事也记录在书上。
ESTH|10|1|亚哈随鲁 王向国中和海岛的人征税。
ESTH|10|2|他以权柄能力所做的一切，以及他使 末底改 尊大、提升他的事，岂不都写在 玛代 和 波斯 王的史籍上吗？
ESTH|10|3|犹太 人 末底改 作 亚哈随鲁 王的宰相，在 犹太 人中为大，得许多弟兄的喜悦，为本族的人争取福利，为他所有的后代谋求幸福。
