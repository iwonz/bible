EZRA|1|1|波斯 王 居魯士 元年，耶和華為要應驗藉 耶利米 的口所說的話，就激發 波斯 王 居魯士 的心，使他下詔書通告全國，說：
EZRA|1|2|「 波斯 王 居魯士 如此說：耶和華天上的上帝已將地上萬國賜給我，又委派我在 猶大 的 耶路撒冷 為他建造殿宇。
EZRA|1|3|你們中間凡作他子民的，可以上 猶大 的 耶路撒冷 去，重建耶和華－ 以色列 上帝的殿，他是在 耶路撒冷 的上帝；願上帝與這人同在。
EZRA|1|4|凡存留的人，無論寄居何處，那地的人要用金銀、財物、牲畜幫助他，還要為 耶路撒冷 上帝的殿甘心獻上禮物。」
EZRA|1|5|於是， 猶大 和 便雅憫 的族長、祭司、 利未 人，凡是心被上帝感動的人都起來，要上 耶路撒冷 去建造耶和華的殿。
EZRA|1|6|四圍所有的人都拿銀器 、金子、財物、牲畜、珍寶支持他們 ，此外還有甘心獻的一切禮物 。
EZRA|1|7|居魯士 王也把耶和華殿的器皿拿出來，這些器皿是 尼布甲尼撒 從 耶路撒冷 掠取，放在自己神明廟中的。
EZRA|1|8|波斯 王 居魯士 派 米提利達 司庫把這些器皿拿出來，點交給 猶大 的領袖 設巴薩 。
EZRA|1|9|它們的數目如下：金盤三十個，銀盤一千個，刀二十九把，
EZRA|1|10|金碗三十個，備用銀碗四百一十個，其他器皿一千件。
EZRA|1|11|金銀器皿共有五千四百件。被擄的人從 巴比倫 上 耶路撒冷 的時候， 設巴薩 把這一切都帶了上來。
EZRA|2|1|這些是從被擄之地上來的省民， 巴比倫 王 尼布甲尼撒 把他們擄到 巴比倫 ，他們重返 耶路撒冷 和 猶大 ，各歸本城。
EZRA|2|2|他們是同 所羅巴伯 、 耶書亞 、 尼希米 、 西萊雅 、 利來雅 、 末底改 、 必珊 、 米斯拔 、 比革瓦伊 、 利宏 、 巴拿 一起回來的。 以色列 百姓的人數如下：
EZRA|2|3|巴錄 的子孫二千一百七十二名；
EZRA|2|4|示法提雅 的子孫三百七十二名；
EZRA|2|5|亞拉 的子孫七百七十五名；
EZRA|2|6|巴哈‧摩押 的後裔，就是 耶書亞 和 約押 的子孫二千八百一十二名；
EZRA|2|7|以攔 的子孫一千二百五十四名；
EZRA|2|8|薩土 的子孫九百四十五名；
EZRA|2|9|薩改 的子孫七百六十名；
EZRA|2|10|巴尼 的子孫六百四十二名；
EZRA|2|11|比拜 的子孫六百二十三名；
EZRA|2|12|押甲 的子孫一千二百二十二名；
EZRA|2|13|亞多尼干 的子孫六百六十六名；
EZRA|2|14|比革瓦伊 的子孫二千零五十六名；
EZRA|2|15|亞丁 的子孫四百五十四名；
EZRA|2|16|亞特 的後裔，就是 希西家 的子孫九十八名；
EZRA|2|17|比賽 的子孫三百二十三名；
EZRA|2|18|約拉 的子孫一百一十二名；
EZRA|2|19|哈順 的子孫二百二十三名；
EZRA|2|20|吉罷珥 人九十五名；
EZRA|2|21|伯利恆 人一百二十三名；
EZRA|2|22|尼陀法 人五十六名；
EZRA|2|23|亞拿突 人一百二十八名；
EZRA|2|24|亞斯瑪弗 人四十二名；
EZRA|2|25|基列‧耶琳 人、 基非拉 人、 比錄 人共七百四十三名；
EZRA|2|26|拉瑪 人和 迦巴 人共六百二十一名；
EZRA|2|27|默瑪 人一百二十二名；
EZRA|2|28|伯特利 人和 艾 人共二百二十三名；
EZRA|2|29|尼波 人五十二名；
EZRA|2|30|末必 人一百五十六名；
EZRA|2|31|另一個 以攔 的子孫一千二百五十四名；
EZRA|2|32|哈琳 的子孫三百二十名；
EZRA|2|33|羅德 人、 哈第 人、 阿挪 人共七百二十五名；
EZRA|2|34|耶利哥 人三百四十五名；
EZRA|2|35|西拿 人三千六百三十名。
EZRA|2|36|祭司： 耶書亞 家 耶大雅 的子孫九百七十三名；
EZRA|2|37|音麥 的子孫一千零五十二名；
EZRA|2|38|巴施戶珥 的子孫一千二百四十七名；
EZRA|2|39|哈琳 的子孫一千零一十七名。
EZRA|2|40|利未 人： 何達威雅 的後裔，就是 耶書亞 和 甲篾 的子孫七十四名。
EZRA|2|41|歌唱的： 亞薩 的子孫一百二十八名。
EZRA|2|42|門口的守衛： 沙龍 的子孫、 亞特 的子孫、 達們 的子孫、 亞谷 的子孫、 哈底大 的子孫、 朔拜 的子孫，共一百三十九名。
EZRA|2|43|殿役： 西哈 的子孫、 哈蘇巴 的子孫、 答巴俄 的子孫、
EZRA|2|44|基綠 的子孫、 西亞 的子孫、 巴頓 的子孫、
EZRA|2|45|利巴拿 的子孫、 哈迦巴 的子孫、 亞谷 的子孫、
EZRA|2|46|哈甲 的子孫、 薩買 的子孫、 哈難 的子孫、
EZRA|2|47|吉德 的子孫、 迦哈 的子孫、 利亞雅 的子孫、
EZRA|2|48|利汛 的子孫、 尼哥大 的子孫、 迦散 的子孫、
EZRA|2|49|烏撒 的子孫、 巴西亞 的子孫、 比賽 的子孫、
EZRA|2|50|押拿 的子孫、 米烏寧 的子孫、 尼普心 的子孫、
EZRA|2|51|巴卜 的子孫、 哈古巴 的子孫、 哈忽 的子孫、
EZRA|2|52|巴洗律 的子孫、 米希大 的子孫、 哈沙 的子孫、
EZRA|2|53|巴柯 的子孫、 西西拉 的子孫、 答瑪 的子孫、
EZRA|2|54|尼細亞 的子孫、 哈提法 的子孫。
EZRA|2|55|所羅門 僕人的後裔： 瑣太 的子孫、 瑣斐列 的子孫、 比路大 的子孫、
EZRA|2|56|雅拉 的子孫、 達昆 的子孫、 吉德 的子孫、
EZRA|2|57|示法提雅 的子孫、 哈替 的子孫、 玻黑列‧哈斯巴音 的子孫、 亞米 的子孫。
EZRA|2|58|殿役和 所羅門 僕人的後裔共三百九十二名。
EZRA|2|59|從 特‧米拉 、 特‧哈薩 、 基綠 、 亞頓 、 音麥 上來，不能證明他們的父系家族和後裔是否屬 以色列 的如下：
EZRA|2|60|第萊雅 的子孫、 多比雅 的子孫、 尼哥大 的子孫，共六百五十二名。
EZRA|2|61|祭司中， 哈巴雅 的子孫、 哈哥斯 的子孫、 巴西萊 的子孫， 巴西萊 因為娶了 基列 人 巴西萊 的女兒為妻，所以就以此為名。
EZRA|2|62|這些人在族譜之中尋查自己的譜系，卻尋不著，因此算為不潔，不得作祭司。
EZRA|2|63|省長對他們說，不可吃至聖的物，直到有會用烏陵和土明的祭司興起來。
EZRA|2|64|全會眾共有四萬二千三百六十名。
EZRA|2|65|此外，還有他們的僕婢七千三百三十七名，又有歌唱的男女二百名。
EZRA|2|66|他們有七百三十六匹馬，二百四十五匹騾子，
EZRA|2|67|四百三十五匹駱駝，六千七百二十匹驢。
EZRA|2|68|有些族長到了 耶路撒冷 耶和華的殿，為上帝的殿甘心獻上禮物，要在原有的根基上重新建造。
EZRA|2|69|他們量力捐入工程的庫房，有六萬一千達利克 金子，五千彌那銀子，以及一百件祭司的禮服。
EZRA|2|70|於是祭司、 利未 人、百姓中的一些人、歌唱的、門口的守衛、殿役，各住在自己的城裏； 以色列 眾人都住在自己的城裏。
EZRA|3|1|到了七月， 以色列 人住在自己的城裏；那時他們如同一人，聚集在 耶路撒冷 。
EZRA|3|2|約薩達 的兒子 耶書亞 和他的弟兄眾祭司，以及 撒拉鐵 的兒子 所羅巴伯 和他的弟兄，都起來建築 以色列 上帝的壇，要照神人 摩西 律法書上所寫的，在壇上獻燔祭。
EZRA|3|3|他們在原有的根基上築壇，因為他們懼怕鄰邦民族，又在其上向耶和華早晚獻燔祭，
EZRA|3|4|並照律法書上所寫的守住棚節，按數照例每日獻所當獻的燔祭。
EZRA|3|5|此後，他們獻常獻的燔祭，並在初一和耶和華一切分別為聖的節期獻祭，又向耶和華獻各人的甘心祭。
EZRA|3|6|從七月初一起，雖然耶和華殿的根基尚未立定，他們開始向耶和華獻燔祭。
EZRA|3|7|他們把銀子給石匠、木匠，把糧食、酒、油給 西頓 人、 推羅 人，好將香柏樹從 黎巴嫩 浮海運到 約帕 ，是照 波斯 王 居魯士 所允准他們的。
EZRA|3|8|他們到了 耶路撒冷 上帝殿的第二年，二月的時候， 撒拉鐵 的兒子 所羅巴伯 ， 約薩達 的兒子 耶書亞 和其餘的弟兄，就是祭司和 利未 人，以及所有被擄歸回 耶路撒冷 的人，就開工建造；他們派二十歲以上的 利未 人，監督建造耶和華殿的工作。
EZRA|3|9|於是 何達威雅 的後裔，就是 耶書亞 和他的子孫與弟兄、 甲篾 和他的子孫，他們和 利未 人 希拿達 的子孫與弟兄，都起來如同一人，監督那些在上帝殿裏做工的人。
EZRA|3|10|工匠立耶和華殿根基的時候，祭司穿禮服吹號， 利未 人 亞薩 的子孫敲鈸，都照 以色列 王 大衛 親手所定的，站著讚美耶和華。
EZRA|3|11|他們彼此唱和，讚美稱謝耶和華： 「他本為善， 他向 以色列 永施慈愛。」 他們讚美耶和華的時候，眾百姓大聲呼喊，因為耶和華殿的根基已經立定。
EZRA|3|12|然而有許多祭司、 利未 人和族長，就是見過先前那殿的老年人，現在親眼看見這殿立了根基，就大聲哭號，也有許多人大聲歡呼，
EZRA|3|13|百姓不能分辨歡呼的聲音或哭號的聲音，因為百姓大聲呼喊，聲音連遠處都可聽到。
EZRA|4|1|猶大 和 便雅憫 的敵人聽說被擄歸回的人為耶和華－ 以色列 的上帝建造殿宇，
EZRA|4|2|就去見 所羅巴伯 和族長，對他們說：「請讓我們與你們一同建造，因為我們也與你們一樣尋求你們的上帝。自從 亞述 王 以撒‧哈頓 帶我們上這地的日子以來，我們常向上帝獻祭。」
EZRA|4|3|但 所羅巴伯 、 耶書亞 和其餘 以色列 的族長對他們說：「我們建造上帝的殿與你們無關，因為我們要照 波斯 王 居魯士 所吩咐的，自己為耶和華－ 以色列 的上帝協力建造。」
EZRA|4|4|那地的人就在 猶大 百姓建造的時候，使他們的手發軟，擾亂他們。
EZRA|4|5|從 波斯 王 居魯士 年間，直到 波斯 王 大流士 在位的時候，那些人賄賂謀士，要破壞他們的計劃。
EZRA|4|6|亞哈隨魯 在位，他的國度剛開始的時候，他們上書控告 猶大 和 耶路撒冷 的居民。
EZRA|4|7|亞達薛西 年間， 比施蘭 、 米特利達 、 他別 和他們 的同僚上書奏告 波斯 王 亞達薛西 。奏文是用 亞蘭 文寫的，以 亞蘭 文呈上。
EZRA|4|8|利宏 省長、 伸帥 書記也上奏 亞達薛西 王，控告 耶路撒冷 如下
EZRA|4|9|（那時， 利宏 省長、 伸帥 書記和他們其餘的同僚，法官、官員、軍官、 波斯 官員 、 亞基衛 人、 巴比倫 人，和 書珊迦 人，就是 以攔 人 ，
EZRA|4|10|以及被 亞斯那巴 大人遷移、安置在 撒瑪利亞城 和 大河 西邊一帶地方其餘的人。現在 ，
EZRA|4|11|這是他們上奏 亞達薛西 王奏文的抄本）：「 河西 的臣僕上奏 亞達薛西 王，現在
EZRA|4|12|請王知道，從王那裏上到我們這裏的 猶太 人，已經抵達 耶路撒冷 。他們正在重建這反叛惡劣的城，已經完成了城牆，正要修復根基。
EZRA|4|13|如今請王知道，這城若再建造，城牆完工，他們就不再進貢、納糧、繳稅，王的國庫必受虧損。
EZRA|4|14|如今，我們吃的鹽既然全是宮廷的鹽，就不忍見王吃虧，因此奏告於王，
EZRA|4|15|請王考察先王史籍，必會在史籍上查知這城是反叛的城，對列王和各省有害；自古以來，城中常有悖逆的事，因此這城曾被拆毀。
EZRA|4|16|我們謹奏王知，這城若再建造，城牆完工， 河西 之地王就無份了。」
EZRA|4|17|那時王諭覆 利宏 省長、 伸帥 書記和他們其餘的同僚，就是住 撒瑪利亞 和 河西 一帶地方的人，說：「願你們平安。現在
EZRA|4|18|你們所呈給我們的奏本，已經清楚地在我面前讀了。
EZRA|4|19|我已下令考查，得知這城自古以來果然背叛列王，其中常有反叛悖逆的事。
EZRA|4|20|也曾有強大的君王治理 耶路撒冷 ，統管 河西 全地，人就給他們進貢、納糧、繳稅。
EZRA|4|21|現在你們要下令叫這些人停工，使這城不得建造，等到我再降旨。
EZRA|4|22|你們當謹慎辦這事，不可遲延，何必讓損害加重，使王受虧損呢？」
EZRA|4|23|亞達薛西 王上諭的抄本在 利宏 和 伸帥 書記，以及他們的同僚面前宣讀，他們就急忙往 耶路撒冷 去見 猶太 人，用勢力和強權叫他們停工。
EZRA|4|24|於是，在 耶路撒冷 上帝殿的工程就停止了，直停到 波斯 王 大流士 第二年。
EZRA|5|1|那時， 哈該 先知和 易多 的孫子 撒迦利亞 ，兩個先知奉 以色列 上帝的名向 猶大 和 耶路撒冷 的 猶太 人說預言。
EZRA|5|2|於是 撒拉鐵 的兒子 所羅巴伯 和 約薩達 的兒子 耶書亞 起來，開始建造 耶路撒冷 上帝的殿，有上帝的先知在那裏幫助他們。
EZRA|5|3|當時 河西 的 達乃 總督和 示他‧波斯乃 ，以及他們的同僚來對 猶太 人這樣說：「誰降旨讓你們建造這殿，完成這建築呢？」
EZRA|5|4|於是我們告訴他們建造這建築物的人叫甚麼名字。
EZRA|5|5|但上帝的眼目看顧 猶太 人的長老，以致沒有人叫他們停工，直到奏文上告 大流士 ，得著他對這事的回諭。
EZRA|5|6|這是 河西 的 達乃 總督和 示他‧波斯乃 ，以及他們的同僚，就是住 河西 的官員 ，上書奏告 大流士 王的抄本，
EZRA|5|7|他們上書給王的奏文，其中寫著：「願 大流士 王諸事平安。
EZRA|5|8|請王知道，我們往 猶大 省去，到了至大上帝的殿。這殿是用鑿成的石頭建造的，梁木插入牆內。這項工程進行迅速，在他們手中順利。
EZRA|5|9|於是我們問那些長老，對他們這樣說：『誰降旨讓你們建造這殿，完成這建築呢？』
EZRA|5|10|我們又問他們的名字，要記下他們領袖的名字，奏告於王。
EZRA|5|11|他們這樣回答我們說：『我們是天和地之上帝的僕人，重建多年前所建造的殿，就是 以色列 一位偉大的君王建造完成的。
EZRA|5|12|但因我們祖先惹天上的上帝發怒，上帝把他們交在 迦勒底 人 巴比倫 王 尼布甲尼撒 的手中，他就拆毀這殿，又把百姓擄到 巴比倫 。
EZRA|5|13|然而 巴比倫 王 居魯士 元年，他降旨允准建造上帝的這殿。
EZRA|5|14|上帝殿中的金銀器皿，就是 尼布甲尼撒 從 耶路撒冷 殿中掠取帶到 巴比倫 廟裏的， 居魯士 王從 巴比倫 廟裏取出來，交給派為省長，名叫 設巴薩 的，
EZRA|5|15|對他說：可以將這些器皿帶去，放在 耶路撒冷 的殿中，在原處建造上帝的殿。
EZRA|5|16|於是那位 設巴薩 來建立 耶路撒冷 上帝殿的根基。但從那時直到如今，這殿尚未修建完畢。』
EZRA|5|17|現在，王若以為好，請查閱 巴比倫 王的檔案庫，看 居魯士 王有沒有降旨允准在 耶路撒冷 建造上帝的殿。請降旨指示我們王對這件事的心意。」
EZRA|6|1|於是 大流士 王降旨，要尋察典籍庫，就是在 巴比倫 藏檔案之處；
EZRA|6|2|在 瑪代 省 亞馬他城 的宮內尋得一卷，其中這樣寫著，「紀錄如下：
EZRA|6|3|居魯士 王元年，王降旨論到在 耶路撒冷 上帝的殿，要建造這殿作為獻祭之處，堅固它的根基。殿高六十肘，寬六十肘，
EZRA|6|4|要用三層鑿成的石頭，一層木頭 ，經費可出於王的庫房。
EZRA|6|5|至於上帝殿的金銀器皿，就是 尼布甲尼撒 從 耶路撒冷 的殿中掠取帶到 巴比倫 的，必須歸還，帶回 耶路撒冷 的殿中，各按原處放在上帝的殿裏。」
EZRA|6|6|「現在， 河西 的 達乃 總督和 示他‧波斯乃 ，以及他們的同僚，就是住 河西 的官員，你們當遠離那裏。
EZRA|6|7|不要攔阻這上帝殿的工作，任由 猶太 人的省長和長老在原處建造上帝的這殿。
EZRA|6|8|我又降旨，吩咐你們為建造上帝的殿當向 猶太 人的長老這樣行：從王的財產中，由 河西 所繳納的貢銀，迅速支付這些人，免得工程停頓。
EZRA|6|9|他們向天上的上帝獻燔祭所需用的公牛犢、公綿羊、小綿羊，以及麥子、鹽、酒、油，都要照 耶路撒冷 祭司的話，每日供給他們，不得有誤；
EZRA|6|10|好叫他們獻馨香的祭給天上的上帝，又為王和王眾子的壽命祈禱。
EZRA|6|11|我再降旨，無論誰更改這命令，必從他房屋中拆出一根梁木，把他舉起，懸在其上，又使他的房屋為此成為糞堆。
EZRA|6|12|任何王或百姓若伸手更改這命令，拆毀在 耶路撒冷 上帝的這殿，願那立他名在那裏的上帝將他們滅絕。我 大流士 降這諭旨，你們要速速遵行。」
EZRA|6|13|於是， 河西 的 達乃 總督和 示他‧波斯乃 ，以及他們的同僚，急速遵行 大流士 王所頒的命令。
EZRA|6|14|猶太 人的長老因 哈該 先知和 易多 的孫子 撒迦利亞 的預言，就建造這殿，凡事順利。他們遵照 以色列 上帝的命令和 波斯 王 居魯士 、 大流士 、 亞達薛西 的諭旨，建造完畢。
EZRA|6|15|大流士 王第六年，亞達月初三，這殿完工了。
EZRA|6|16|以色列 人、祭司和 利未 人，以及其餘被擄歸回的人都歡歡喜喜地為上帝的這殿行奉獻禮。
EZRA|6|17|他們為這上帝殿的奉獻禮獻了一百頭公牛，二百隻公綿羊，四百隻小綿羊，又照 以色列 支派的數目獻十二隻公山羊，作 以色列 眾人的贖罪祭。
EZRA|6|18|他們派祭司按著班次， 利未 人也按著班次在 耶路撒冷 事奉上帝，正如 摩西 律法書上所寫的。
EZRA|6|19|正月十四日，被擄歸回的人守逾越節。
EZRA|6|20|祭司和 利未 人一同自潔，他們全都潔淨了。 利未 人為被擄歸回的眾人和他們的弟兄眾祭司，並為自己宰逾越節的羔羊。
EZRA|6|21|從被擄之地歸回的 以色列 人，並所有歸附他們、除掉這地外邦人的污穢、尋求耶和華－ 以色列 上帝的人，都吃這羔羊。
EZRA|6|22|他們歡歡喜喜地守除酵節七日，因為耶和華使他們歡喜。耶和華又使 亞述 王的心轉向他們，堅固他們的手，去做上帝－ 以色列 上帝殿的工。
EZRA|7|1|這些事以後， 波斯 王 亞達薛西 在位的時候，有個人叫 以斯拉 ，他是 西萊雅 的兒子， 西萊雅 是 亞撒利雅 的兒子， 亞撒利雅 是 希勒家 的兒子，
EZRA|7|2|希勒家 是 沙龍 的兒子， 沙龍 是 撒督 的兒子， 撒督 是 亞希突 的兒子，
EZRA|7|3|亞希突 是 亞瑪利雅 的兒子， 亞瑪利雅 是 亞撒利雅 的兒子， 亞撒利雅 是 米拉約 的兒子，
EZRA|7|4|米拉約 是 西拉希雅 的兒子， 西拉希雅 是 烏西 的兒子， 烏西 是 布基 的兒子，
EZRA|7|5|布基 是 亞比書 的兒子， 亞比書 是 非尼哈 的兒子， 非尼哈 是 以利亞撒 的兒子， 以利亞撒 是 亞倫 大祭司的兒子。
EZRA|7|6|這 以斯拉 從 巴比倫 上來，他是一個文士，精通耶和華－ 以色列 上帝所賜 摩西 的律法。王允准他一切所求的，因為耶和華－他上帝的手幫助他。
EZRA|7|7|亞達薛西 王第七年，有些 以色列 人、一些祭司、 利未 人、歌唱的、門口的守衛、殿役，上 耶路撒冷 去。
EZRA|7|8|王第七年五月， 以斯拉 到了 耶路撒冷 。
EZRA|7|9|正月初一，他從 巴比倫 起程，五月初一就到了 耶路撒冷 ，因為他上帝施恩的手幫助他。
EZRA|7|10|以斯拉 立志考究遵行耶和華的律法，又將律例典章教導 以色列 人。
EZRA|7|11|亞達薛西 王賜給精通耶和華誡命和 以色列 律例的文士 以斯拉 祭司的諭旨，抄本如下：
EZRA|7|12|「諸王之王 亞達薛西 ，達於精通天上之上帝律法的 以斯拉 祭司文士等等：現在
EZRA|7|13|住在我國中的 以色列 百姓、祭司、 利未 人，凡願意上 耶路撒冷 去的，我降旨准他們與你同去。
EZRA|7|14|既然王與七個謀士派你去，照你手中上帝的律法視察 猶大 和 耶路撒冷 的景況；
EZRA|7|15|你又帶著王和謀士樂意獻給住 耶路撒冷 、 以色列 上帝的金銀，
EZRA|7|16|和你在 巴比倫 全省所得的一切金銀，以及百姓、祭司甘心獻給 耶路撒冷 他們上帝殿的禮物，
EZRA|7|17|那麼，你就當用這銀子急速買公牛、公綿羊、小綿羊，和同獻的素祭、澆酒祭，獻在 耶路撒冷 你們上帝殿的壇上。
EZRA|7|18|剩下的金銀，你和你的弟兄看怎樣好，就怎樣用，但總要遵照你們上帝的旨意。
EZRA|7|19|你要帶著交託給你、在上帝殿中事奉用的器皿，到 耶路撒冷 上帝面前。
EZRA|7|20|你上帝殿裏若再有需用的經費，是你負責供應的，可以從王的寶庫裏支取。
EZRA|7|21|「我 亞達薛西 王又降旨達於 河西 所有的司庫：『精通天上之上帝律法的 以斯拉 祭司文士無論向你們要甚麼，你們要速速辦理，
EZRA|7|22|直至一百他連得銀子，一百柯珥 麥子，一百罷特酒，一百罷特油，鹽不限其數。
EZRA|7|23|凡天上之上帝所吩咐的，當為天上之上帝的殿切實辦理。何必使憤怒臨到王和王眾子的國呢？
EZRA|7|24|我再吩咐你們：至於任何祭司、 利未 人、歌唱的、門口的守衛和殿役，以及在上帝的這殿事奉的人，不可要求他們進貢，納糧，繳稅。』
EZRA|7|25|「你， 以斯拉 啊，要照著你上帝賜你的智慧，指派所有明白你上帝律法的人作官長、審判官，治理 河西 所有的百姓，教導不明白上帝律法的人。
EZRA|7|26|凡不遵行你上帝律法和王命令的人，當速速定他的罪，或處死，或充軍，或抄家，或囚禁。」
EZRA|7|27|以斯拉 說：「耶和華－我們列祖的上帝是應當稱頌的！因他使王起這心願，使 耶路撒冷 耶和華的殿得榮耀，
EZRA|7|28|他又在王和謀士，以及王所有大能的軍官面前施恩於我。我因耶和華－我上帝的手的幫助，得以堅強，從 以色列 中召集領袖，與我一同上來。」
EZRA|8|1|這些是 亞達薛西 王在位的時候，同我從 巴比倫 上來的族長和他們的家譜：
EZRA|8|2|屬 非尼哈 的子孫有 革順 ；屬 以他瑪 的子孫有 但以理 ；屬 大衛 的子孫有 哈突 ；
EZRA|8|3|屬 示迦尼 的子孫；屬 巴錄 的子孫有 撒迦利亞 ，同著他按家譜計算，男丁一百五十人；
EZRA|8|4|屬 巴哈‧摩押 的子孫有 西拉希雅 的兒子 以利約乃 ，同著他有男丁二百人；
EZRA|8|5|屬 薩土 的子孫有 雅哈悉 的兒子 示迦尼 ，同著他有男丁三百人；
EZRA|8|6|屬 亞丁 的子孫有 約拿單 的兒子 以別 ，同著他有男丁五十人；
EZRA|8|7|屬 以攔 的子孫有 亞他利雅 的兒子 耶篩亞 ，同著他有男丁七十人；
EZRA|8|8|屬 示法提雅 的子孫有 米迦勒 的兒子 西巴第雅 ，同著他有男丁八十人；
EZRA|8|9|屬 約押 的子孫有 耶歇 的兒子 俄巴底亞 ，同著他有男丁二百一十八人；
EZRA|8|10|屬 巴尼 的子孫有 約細斐 的兒子 示羅密 ，同著他有男丁一百六十人；
EZRA|8|11|屬 比拜 的子孫有 比拜 的兒子 撒迦利亞 ，同著他有男丁二十八人；
EZRA|8|12|屬 押甲 的子孫有 哈加坦 的兒子 約哈難 ，同著他有男丁一百一十人；
EZRA|8|13|屬 亞多尼干 的子孫，就是晚到的，他們的名字是 以利法列 、 耶利 、 示瑪雅 ，同著他們有男丁六十人；
EZRA|8|14|屬 比革瓦伊 的子孫有 烏太 和 撒刻 ，同著他們有男丁七十人。
EZRA|8|15|我召集這些人在流入 亞哈瓦 的河旁邊，我們在那裏紮營三日。我查看百姓和祭司，發現並沒有 利未 人在那裏，
EZRA|8|16|就派人到 以利以謝 、 亞列 、 示瑪雅 、 以利拿單 、 雅立 、 以利拿單 、 拿單 、 撒迦利亞 、 米書蘭 等領袖，以及 約雅立 和 以利拿單 教師那裏。
EZRA|8|17|我吩咐他們往 迦西斐雅 地方去見那裏的領袖 易多 ，又告訴他們當向 易多 和他的弟兄，就是 迦西斐雅 那地方的殿役說甚麼話，好為我們上帝的殿帶事奉的人來。
EZRA|8|18|蒙我們上帝施恩的手幫助我們，他們在 以色列 的曾孫， 利未 的孫子， 抹利 的後裔中帶了一個精明的人來，就是 示利比 ，還有他的眾子與兄弟共十八人。
EZRA|8|19|另外，還有 哈沙比雅 ，同著他有 米拉利 的子孫 耶篩亞 ，以及他的眾子和兄弟共二十人。
EZRA|8|20|從前 大衛 和眾領袖派殿役服事 利未 人，現在從這殿役中也帶了二百二十人來，全都是按名指定的。
EZRA|8|21|那時，我在 亞哈瓦河 邊宣告禁食，為要在我們上帝面前刻苦己心，求他使我們和我們的孩子，以及一切所有的，都得平坦的道路。
EZRA|8|22|我以求王撥步兵騎兵幫助我們抵擋路上的仇敵為羞愧，因我們曾對王說：「我們上帝施恩的手必幫助凡尋求他的，但他的能力和憤怒必攻擊凡離棄他的。」
EZRA|8|23|我們為此禁食祈求我們的上帝，他就應允我們。
EZRA|8|24|我分派十二位祭司長，就是 示利比 、 哈沙比雅 和與他們一起的兄弟十人，
EZRA|8|25|把王和謀士、軍官，並在那裏的 以色列 眾人為我們上帝殿所獻的金銀和器皿，都秤了交給他們。
EZRA|8|26|我秤了交在他們手中的有六百五十他連得銀子，一百他連得銀器，一百他連得金子，
EZRA|8|27|二十個金碗，值一千達利克，上等光亮的銅器皿兩個，珍貴如金。
EZRA|8|28|我對他們說：「你們歸耶和華為聖，器皿也歸為聖；金銀是甘心獻給耶和華－你們列祖之上帝的。
EZRA|8|29|你們要警醒看守，直到你們在祭司長和 利未 族長，以及 以色列 的各族長面前，在 耶路撒冷 耶和華殿的庫房內，把這些過了秤。」
EZRA|8|30|於是，祭司和 利未 人把秤過的金銀和器皿接過來，要帶到 耶路撒冷 我們上帝的殿裏。
EZRA|8|31|正月十二日，我們從 亞哈瓦河 邊起行，要往 耶路撒冷 去。我們上帝的手保佑我們，救我們脫離仇敵和路上埋伏之人的手。
EZRA|8|32|我們到了 耶路撒冷 ，在那裏住了三日。
EZRA|8|33|第四日，金銀和器皿都在我們上帝的殿裏過了秤，交在 烏利亞 的兒子 米利末 祭司的手中。同著他的有 非尼哈 的兒子 以利亞撒 ，還有 利未 人 耶書亞 的兒子 約撒拔 和 賓內 的兒子 挪亞底 。
EZRA|8|34|那時，這一切都點過秤過了，重量全寫在冊上。
EZRA|8|35|從被擄之地歸回的人向 以色列 的上帝獻燔祭，為 以色列 眾人獻十二頭公牛，九十六隻公綿羊，七十七隻小綿羊，又獻十二隻公山羊作贖罪祭，這些全都是獻給耶和華的燔祭。
EZRA|8|36|被擄歸回的人把王的諭旨交給王的總督與 河西 的省長，他們就支助百姓和上帝的殿。
EZRA|9|1|這些事完成以後，眾領袖來接近我，說：「 以色列 百姓、祭司和 利未 人沒有棄絕 迦南 人、 赫 人、 比利洗 人、 耶布斯 人、 亞捫 人、 摩押 人、 埃及 人和 亞摩利 人等列邦民族所行可憎的事。
EZRA|9|2|因他們為自己和兒子娶了這些外邦女子，以致聖潔的種籽和列邦民族混雜，而且領袖和官長在這事上是罪魁。」
EZRA|9|3|我一聽見這事，就撕裂衣服和外袍，拔了頭髮和鬍鬚，驚惶地坐著。
EZRA|9|4|凡為 以色列 上帝言語戰兢的人，都因被擄歸回之人所犯的罪，聚集到我這裏來。我驚惶地坐著，直到獻晚祭的時候。
EZRA|9|5|獻晚祭的時候我從愁煩中起來，穿著撕裂的衣服和外袍，雙膝跪下，向耶和華－我的上帝舉手，
EZRA|9|6|說： 「我的上帝啊，我抱愧蒙羞，不敢向你－我的上帝仰面，因為我們的罪孽多到滅頂，我們的罪惡滔天。
EZRA|9|7|從我們祖先的日子直到今日，我們的罪惡深重；因我們的罪孽，我們和君王、祭司都交在鄰國諸王的手中，被殺害，擄掠，搶奪，臉上蒙羞，正如今日的景況。
EZRA|9|8|現在耶和華－我們的上帝暫且向我們施恩，為我們留下一些殘存之民，使我們如釘子釘在他的聖所，讓我們的上帝光照我們的眼目，使我們在受轄制之中稍微復興。
EZRA|9|9|我們是奴僕，然而在受轄制之中，我們的上帝沒有丟棄我們，在 波斯 諸王面前向我們施恩，叫我們復興，能重建我們上帝的殿，修補毀壞之處，使我們在 猶大 和 耶路撒冷 有城牆。
EZRA|9|10|「我們的上帝啊，既然如此，現在我們還有甚麼話可說呢？因為我們離棄了你的誡命，
EZRA|9|11|就是你藉你僕人眾先知所吩咐的，說：『你們要去得為業之地是污穢之地，因列邦民族的污穢和可憎的事，叫這地從這邊到那邊都充滿了污穢。
EZRA|9|12|現在，不可把你們的女兒嫁給他們的兒子，也不可為你們的兒子娶他們的女兒，永不可求他們的平安和他們的利益，這樣你們就可以強盛，吃這地的美物，並把這地留給你們的子孫永遠為業。』
EZRA|9|13|我們因自己的惡行和大罪，遭遇這一切的事，但你－我們的上帝懲罰我們輕於我們罪所當得的，又為我們留下這些殘存之民。
EZRA|9|14|我們豈可再違背你的誡命，與行這些可憎之事的民族結親呢？若我們這樣行，你豈不向我們發怒，將我們滅絕，以致沒有一個餘民或殘存之民嗎？
EZRA|9|15|耶和華－ 以色列 的上帝啊，你是公義的，我們才能剩下這些殘存之民，正如今日的景況。看哪，我們在你面前有罪惡，因此無人能在你面前站立得住。」
EZRA|10|1|以斯拉 禱告，認罪，哭泣，俯伏在上帝殿前的時候，有 以色列 中的男女和孩童聚集到 以斯拉 那裏，成了一個盛大的會，百姓無不痛哭。
EZRA|10|2|以攔 的子孫， 耶歇 的兒子 示迦尼 對 以斯拉 說：「我們娶了這地的外邦女子，干犯了我們的上帝，然而現在 以色列 人在這事上還有指望。
EZRA|10|3|現在，我們要與我們的上帝立約，送走所有的妻子和她們所生的，照著主和那些因我們上帝誡命戰兢之人所議定的，按律法去行。
EZRA|10|4|起來，這是你當辦的事，我們必支持你，你當奮勇而行。」
EZRA|10|5|以斯拉 就起來，叫祭司長和 利未 人，以及 以色列 眾人起誓，要照這話去做；他們就起了誓。
EZRA|10|6|以斯拉 從上帝殿前起來，進入 以利亞實 的兒子 約哈難 的屋裏，到了那裏不吃飯，也不喝水，為被擄歸回之人所犯的罪悲傷。
EZRA|10|7|他們通告 猶大 和 耶路撒冷 ，叫所有被擄歸回的人聚集在 耶路撒冷 。
EZRA|10|8|凡不遵照領袖和長老所議定，三日之內不來的，就必毀壞他所有的財產，把他從被擄歸回之人的會中開除。
EZRA|10|9|於是， 猶大 和 便雅憫 眾人三日之內都聚集在 耶路撒冷 。那時是九月，那月的二十日，眾百姓坐在上帝殿前的廣場，因這事，又因下大雨，就都戰抖。
EZRA|10|10|以斯拉 祭司站起來，對他們說：「你們有罪了，因為你們娶了外邦女子，增添 以色列 的罪惡。
EZRA|10|11|現在當向耶和華－你們列祖的上帝認罪，遵行他的旨意，離開這地的百姓和外邦女子。」
EZRA|10|12|全會眾大聲回答說：「好！我們必照著你的話去做。
EZRA|10|13|只是百姓眾多，又逢大雨的季節，我們沒有氣力站在外面；這也不是一兩天可以辦完的事，因我們在這事上犯了大罪。
EZRA|10|14|讓我們的領袖代表全會眾留在那裏。我們城鎮中凡娶外邦女子的，當按所定的日期，會同本城的長老和審判官前來，直到辦完這事，上帝的烈怒轉離我們 。」
EZRA|10|15|惟有 亞撒黑 的兒子 約拿單 ， 特瓦 的兒子 雅哈謝 反對這事，並有 米書蘭 和 利未 人 沙比太 支持他們。
EZRA|10|16|被擄歸回的人就如此做了。 以斯拉 祭司按著父家指名選派一些族長 。十月初一，他們一同坐下來查辦這事，
EZRA|10|17|到正月初一，才查清所有娶外邦女子的人數。
EZRA|10|18|在祭司中查出娶外邦女子的： 耶書亞 的子孫中，有 約薩達 的兒子，和他兄弟 瑪西雅 、 以利以謝 、 雅立 、 基大利 ，
EZRA|10|19|他們承諾要送走他們的妻子。他們因有罪，就獻羊群中的一隻公綿羊贖罪；
EZRA|10|20|音麥 的子孫中，有 哈拿尼 、 西巴第雅 ；
EZRA|10|21|哈琳 的子孫中，有 瑪西雅 、 以利雅 、 示瑪雅 、 耶歇 、 烏西雅 ；
EZRA|10|22|巴施戶珥 的子孫中，有 以利約乃 、 瑪西雅 、 以實瑪利 、 拿坦業 、 約撒拔 、 以利亞薩 。
EZRA|10|23|利未 人中，有 約撒拔 、 示每 、 基拉雅 ， 基拉雅 就是 基利他 ，還有 毗他希雅 、 猶大 、 以利以謝 。
EZRA|10|24|歌唱的人中有 以利亞實 。門口的守衛中，有 沙龍 、 提聯 、 烏利 。
EZRA|10|25|以色列 人 巴錄 的子孫中，有 拉米 、 耶西雅 、 瑪基雅 、 米雅民 、 以利亞撒 、 瑪基雅 、 比拿雅 。
EZRA|10|26|以攔 的子孫中，有 瑪他尼 、 撒迦利亞 、 耶歇 、 押底 、 耶列末 、 以利雅 。
EZRA|10|27|薩土 的子孫中，有 以利約乃 、 以利亞實 、 瑪他尼 、 耶列末 、 撒拔 、 亞西撒 。
EZRA|10|28|比拜 的子孫中，有 約哈難 、 哈拿尼雅 、 薩拜 、 亞勒 。
EZRA|10|29|巴尼 的子孫中，有 米書蘭 、 瑪鹿 、 亞大雅 、 雅述 、 示押 、 拉末 。
EZRA|10|30|巴哈‧摩押 的子孫中，有 阿底拿 、 基拉 、 比拿雅 、 瑪西雅 、 瑪他尼 、 比撒列 、 賓內 、 瑪拿西 。
EZRA|10|31|哈琳 的子孫中，有 以利以謝 、 伊示雅 、 瑪基雅 、 示瑪雅 、 西緬 、
EZRA|10|32|便雅憫 、 瑪鹿 、 示瑪利雅 。
EZRA|10|33|哈順 的子孫中，有 瑪特乃 、 瑪達他 、 撒拔 、 以利法列 、 耶利買 、 瑪拿西 、 示每 。
EZRA|10|34|巴尼 的子孫中，有 瑪玳 、 暗蘭 、 烏益 、
EZRA|10|35|比拿雅 、 比底雅 、 基祿 、
EZRA|10|36|瓦尼雅 、 米利末 、 以利亞實 、
EZRA|10|37|瑪他尼 、 瑪特乃 、 雅掃 、
EZRA|10|38|巴尼 、 賓內 、 示每 、
EZRA|10|39|示利米雅 、 拿單 、 亞大雅 、
EZRA|10|40|瑪拿底拜 、 沙賽 、 沙賴 、
EZRA|10|41|亞薩利 、 示利米雅 、 示瑪利雅 、
EZRA|10|42|沙龍 、 亞瑪利雅 、 約瑟 。
EZRA|10|43|尼波 的子孫中，有 耶利 、 瑪他提雅 、 撒拔 、 西比拿 、 雅玳 、 約珥 、 比拿雅 。
EZRA|10|44|這些人全都娶了外邦女子，其中也有生了兒女的 。
