HAG|1|1|Во второй год царя Дария, в шестой месяц, в первый день месяца, было слово Господне через Аггея пророка к Зоровавелю, сыну Салафиилеву, правителю Иудеи, и к Иисусу, сыну Иоседекову, великому иерею:
HAG|1|2|так сказал Господь Саваоф: народ сей говорит: "не пришло еще время, не время строить дом Господень".
HAG|1|3|И было слово Господне через Аггея пророка:
HAG|1|4|а вам самим время жить в домах ваших украшенных, тогда как дом сей в запустении?
HAG|1|5|Посему ныне так говорит Господь Саваоф: обратите сердце ваше на пути ваши.
HAG|1|6|Вы сеете много, а собираете мало; едите, но не в сытость; пьете, но не напиваетесь; одеваетесь, а не согреваетесь; зарабатывающий плату зарабатывает для дырявого кошелька.
HAG|1|7|Так говорит Господь Саваоф: обратите сердце ваше на пути ваши.
HAG|1|8|Взойдите на гору и носите дерева, и стройте храм; и Я буду благоволить к нему, и прославлюсь, говорит Господь.
HAG|1|9|Ожидаете многого, а выходит мало; и что принесете домой, то Я развею. – За что? говорит Господь Саваоф: за Мой дом, который в запустении, тогда как вы бежите, каждый к своему дому.
HAG|1|10|Посему–то небо заключилось и не дает вам росы, и земля не дает своих произведений.
HAG|1|11|И Я призвал засуху на землю, на горы, на хлеб, на виноградный сок, на елей и на все, что производит земля, и на человека, и на скот, и на всякий ручной труд.
HAG|1|12|И послушались Зоровавель, сын Салафиилев, и Иисус, сын Иоседеков, и весь прочий народ гласа Господа Бога своего и слов Аггея пророка, как посланного Господом Богом их, и народ убоялся Господа.
HAG|1|13|Тогда Аггей, вестник Господень, посланный от Господа, сказал к народу: Я с вами! говорит Господь.
HAG|1|14|И возбудил Господь дух Зоровавеля, сына Салафиилева, правителя Иудеи, и дух Иисуса, сына Иоседекова, великого иерея, и дух всего остатка народа, и они пришли, и стали производить работы в доме Господа Саваофа, Бога своего,
HAG|1|15|в двадцать четвертый день шестого месяца, во второй год царя Дария.
HAG|2|1|В седьмой месяц, в двадцать первый день месяца, было слово Господне через Аггея пророка:
HAG|2|2|скажи теперь Зоровавелю, сыну Салафиилеву, правителю Иудеи, и Иисусу, сыну Иоседекову, великому иерею, и остатку народа:
HAG|2|3|кто остался между вами, который видел этот дом в прежней его славе, и каким видите вы его теперь? Не есть ли он в глазах ваших как бы ничто?
HAG|2|4|Но ободрись ныне, Зоровавель, говорит Господь, ободрись, Иисус, сын Иоседеков, великий иерей! ободрись, весь народ земли, говорит Господь, и производите работы, ибо Я с вами, говорит Господь Саваоф.
HAG|2|5|Завет Мой, который Я заключил с вами при исшествии вашем из Египта, и дух Мой пребывает среди вас: не бойтесь!
HAG|2|6|Ибо так говорит Господь Саваоф: еще раз, и это будет скоро, Я потрясу небо и землю, море и сушу,
HAG|2|7|и потрясу все народы, и придет Желаемый всеми народами, и наполню дом сей славою, говорит Господь Саваоф.
HAG|2|8|Мое серебро и Мое золото, говорит Господь Саваоф.
HAG|2|9|Слава сего последнего храма будет больше, нежели прежнего, говорит Господь Саваоф; и на месте сем Я дам мир, говорит Господь Саваоф.
HAG|2|10|В двадцать четвертый день девятого месяца, во второй год Дария, было слово Господне через Аггея пророка:
HAG|2|11|так говорит Господь Саваоф: спроси священников о законе и скажи:
HAG|2|12|если бы кто нес освященное мясо в поле одежды своей и полою своею коснулся хлеба, или чего–либо вареного, или вина, или елея, или какой–нибудь пищи: сделается ли это священным? И отвечали священники и сказали: нет.
HAG|2|13|Потом сказал Аггей: а если прикоснется ко всему этому кто–либо, осквернившийся от прикосновения к мертвецу: сделается ли это нечистым? И отвечали священники и сказали: будет нечистым.
HAG|2|14|Тогда отвечал Аггей и сказал: таков этот народ, таково это племя предо Мною, говорит Господь, и таковы все дела рук их! И что они приносят там, все нечисто.
HAG|2|15|Теперь обратите сердце ваше на время от сего дня и назад, когда еще не был положен камень на камень в храме Господнем.
HAG|2|16|Приходили бывало к копне, могущей приносить двадцать мер, и оказывалось только десять; приходили к подточилию, чтобы начерпать пятьдесят мер из подточилия, а оказывалось только двадцать.
HAG|2|17|Поражал Я вас ржавчиною и блеклостью хлеба и градом все труды рук ваших; но вы не обращались ко Мне, говорит Господь.
HAG|2|18|Обратите же сердце ваше на время от сего дня и назад, от двадцать четвертого дня девятого месяца, от того дня, когда основан был храм Господень; обратите сердце ваше:
HAG|2|19|есть ли еще в житницах семена? Доселе ни виноградная лоза, ни смоковница, ни гранатовое дерево, ни маслина не давали плода; а от сего дня Я благословлю их.
HAG|2|20|И было слово Господне к Аггею вторично в двадцать четвертый день месяца, и сказано:
HAG|2|21|скажи Зоровавелю, правителю Иудеи: потрясу Я небо и землю;
HAG|2|22|и ниспровергну престолы царств, и истреблю силу царств языческих, опрокину колесницы и сидящих на них, и низринуты будут кони и всадники их, один мечом другого.
HAG|2|23|В тот день, говорит Господь Саваоф, Я возьму тебя, Зоровавель, сын Салафиилев, раб Мой, говорит Господь, и буду держать тебя как печать, ибо Я избрал тебя, говорит Господь Саваоф.
