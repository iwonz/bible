ISA|1|1|Visio Isaiae filii Amos, quam vidit super Iudam et Ierusalem in diebus Oziae, Ioatham, Achaz, Ezechiae regum Iudae.
ISA|1|2|Audite, caeli, et auribus percipe, terra,quoniam Dominus locutus est: Filios enutrivi et exaltavi,ipsi autem spreverunt me.
ISA|1|3|Cognovit bos possessorem suum,et asinus praesepe domini sui;Israel non cognovit,populus meus non intellexit ".
ISA|1|4|Vae genti peccatrici,populo gravi iniquitate,semini nequam, filiis sceleratis!Dereliquerunt Dominum,blasphemaverunt Sanctum Israel,abalienati sunt retrorsum.
ISA|1|5|Super quo percutiemini vos ultra,addentes praevaricationem?Omne caput languidum,et omne cor maerens.
ISA|1|6|A planta pedis usque ad verticemnon est in eo sanitas;vulnus et livor et plaga tumensnon est circumligatanec curata medicamine neque fota oleo.
ISA|1|7|Terra vestra deserta,civitates vestrae succensae igni;regionem vestram coram vobis alieni devorant,et desolabitur sicut in vastitate hostili.
ISA|1|8|Et derelinquetur filia Sionut umbraculum in vinea,sicut tugurium in cucumerario,sicut civitas, quae obsessa est.
ISA|1|9|Nisi Dominus exercituum reliquisset nobis semen,quasi Sodoma fuissemuset quasi Gomorra similes essemus.
ISA|1|10|Audite verbum Domini,principes Sodomorum;percipite auribus legem Dei nostri, populus Gomorrae.
ISA|1|11|" Quo mihi multitudinem victimarum vestrarum?,dicit Dominus.Plenus sum holocaustis arietumet adipe pinguium;et sanguinem vitulorumet agnorum et hircorum nolui.
ISA|1|12|Cum veneritis ante conspectum meum,quis quaesivit haec de manibus vestris,ut ambularetis in atriis meis?
ISA|1|13|Ne afferatis ultra sacrificium vanum;abominatio mihi incensum,neomenia et sabbatum et conventus;non feram scelus cum coetu sollemni;
ISA|1|14|calendas vestras et sollemnitates vestras odivit anima mea,facta sunt mihi molesta, laboravi sustinens.
ISA|1|15|Et cum extenderitis manus vestras,avertam oculos meos a vobis;et cum multiplicaveritis orationem,non exaudiam:manus enim vestrae sanguine plenae sunt.
ISA|1|16|Lavamini, mundi estote,auferte malum cogitationum vestrarum ab oculis meis;quiescite agere perverse,
ISA|1|17|discite benefacere:quaerite iudicium, subvenite oppresso,iudicate pupillo, defendite viduam.
ISA|1|18|Et venite, et iudicio contendamus,dicit Dominus.Si fuerint peccata vestra ut coccinum,quasi nix dealbabuntur;et, si fuerint rubra quasi vermiculus,velut lana erunt.
ISA|1|19|Si volueritis et audieritis,bona terrae comedetis;
ISA|1|20|quod si nolueritis et me ad iracundiam provocaveritis,gladius devorabit vos,quia os Domini locutum est ".
ISA|1|21|Quomodo facta est meretrixcivitas fidelis, plena iudicii?Iustitia habitavit in ea,nunc autem homicidae.
ISA|1|22|Argentum tuum versum est in scoriam,vinum tuum mixtum est aqua;
ISA|1|23|principes tui infideles, socii furum:omnes diligunt munera, sequuntur retributiones,pupillo non iudicant, et causa viduae non ingreditur ad illos.
ISA|1|24|Propter hoc ait Dominus, Deus exercituum, Fortis Israel: Heu, consolabor super hostibus meiset vindicabor de inimicis meis.
ISA|1|25|Et convertam manum meam ad teet excoquam ad purum scoriam tuamet auferam omne stannum tuum.
ISA|1|26|Et restituam iudices tuos, ut fuerunt prius,et consiliarios tuos sicut antiquitus;post haec vocaberis Civitas iustitiae, Urbs fidelis ".
ISA|1|27|Sion in iudicio redimeturet, qui in ea reversi sunt, in iustitia.
ISA|1|28|Erit autem ruina scelestis et peccatoribus simul;et, qui dereliquerunt Dominum, consumentur.
ISA|1|29|Confundemini enim terebinthis, in quibus delectati estis,et erubescetis super hortis, quos elegistis.
ISA|1|30|Nam eritis velut quercus, defluentibus foliis,et velut hortus absque aqua;
ISA|1|31|et erit fortitudo vestra ut favilla stuppae,et opus eius quasi scintilla,et succendetur utrumque simul, et non erit qui exstinguat.
ISA|2|1|Verbum, quod vidit Isaias filius Amos super Iudam et Ieru salem.
ISA|2|2|Et erit in novissimis diebuspraeparatus mons domus Domini in vertice montium,et elevabitur super colles;et fluent ad eum omnes gentes.
ISA|2|3|Et ibunt populi multi et dicent: Venite, et ascendamus ad montem Domini,ad domum Dei Iacob,ut doceat nos vias suas,et ambulemus in semitis eius ";quia de Sion exibit lex,et verbum Domini de Ierusalem.
ISA|2|4|Et iudicabit genteset arguet populos multos;et conflabunt gladios suos in vomereset lanceas suas in falces;non levabit gens contra gentem gladium,nec exercebuntur ultra ad proelium.
ISA|2|5|Domus Iacob, venite,et ambulemus in lumine Domini.
ISA|2|6|Proiecisti enim populum tuum, domum Iacob,quia repleti sunt hariolis orientalibuset augures habuerunt ut Philisthimet manus alienis porrigunt.
ISA|2|7|Repleta est terra eius argento et auro,et non est finis thesaurorum eius;
ISA|2|8|et repleta est terra eius equis,et innumerabiles quadrigae eius;et repleta est terra eius idolis:opus manuum suarum adoraverunt,quod fecerunt digiti eorum.
ISA|2|9|Et incurvavit se homo,et humiliatus est vir:ne dimittas eis.
ISA|2|10|Ingredere in petram, abscondere in pulverea facie timoris Domini et a gloria maiestatis eius.
ISA|2|11|Oculi sublimes hominis humiliabuntur,et incurvabitur altitudo virorum;exaltabitur autem Dominus solus in die illa.
ISA|2|12|Quia dies Domini exercituumsuper omnem superbum et excelsumet super omnem arrogantem, et humiliabitur;
ISA|2|13|et super omnes cedros Libani sublimes et erectaset super omnes quercus Basan
ISA|2|14|et super omnes montes excelsoset super omnes colles elevatos
ISA|2|15|et super omnem turrim excelsamet super omnem murum munitum
ISA|2|16|et super omnes naves Tharsiset super omnia navigia pulchra.
ISA|2|17|Et incurvabitur sublimitas hominum,et humiliabitur altitudo virorum;et elevabitur Dominus solus in die illa,
ISA|2|18|et idola penitus conterentur.
ISA|2|19|Et introibunt in speluncas petrarumet in voragines terraea facie formidinis Domini et a gloria maiestatis eius,cum surrexerit percutere terram.
ISA|2|20|In die illa proiciet homo idola sua argentea et simulacra sua aurea, quae fecerat sibi, ut adoraret, ad talpas et vespertiliones.
ISA|2|21|Et ingredietur scissuras petrarum et cavernas saxorum a facie formidinis Domini et a gloria maiestatis eius, cum surrexerit percutere terram.
ISA|2|22|Quiescite ergo ab homine, cuius spiritus in naribus eius. Quanti enim aestimabitur ipse?
ISA|3|1|Ecce enim Dominator, Dominus exercituum,aufert a Ierusalem et a Iuda robur et praesidium,omne robur panis et omne robur aquae,
ISA|3|2|fortem et virum bellatorem,iudicem et prophetam et hariolum et senem,
ISA|3|3|principem super quinquaginta et honorabilem vultuet consiliarium et sapientem magumet prudentem incantatorem.
ISA|3|4|Et dabo pueros principes eorum;et infantes dominabuntur eis.
ISA|3|5|Et irruet populus, vir ad virum,unusquisque ad proximum suum:tumultuabitur puer contra senem,et ignobilis contra nobilem.
ISA|3|6|Apprehendet enim vir fratrem suumin domo patris sui: Vestimentum tibi est,princeps esto noster,ruina autem haec sub manu tua ".
ISA|3|7|Clamabit in die illa dicens: Non sum medicus,et in domo mea non est panis neque vestimentum;nolite constituere me principem populi ".
ISA|3|8|Ruit enim Ierusalem, et Iudas concidit,quia lingua eorum et adinventiones eorum contra Dominum,ut provocarent oculos maiestatis eius.
ISA|3|9|Procacitas vultus eorum accusat eos,et peccatum suum quasi Sodomapraedicaverunt nec absconderunt;vae animae eorum,quoniam reddita sunt eis mala!
ISA|3|10|Dicite iusto: " Bene! ",quoniam fructum adinventionum suarum comedet.
ISA|3|11|Vae impio in malum:retributio enim manuum eius fiet ei!
ISA|3|12|Populum meum opprimit infans,et mulieres dominantur ei.Popule meus, qui te beatum dicunt, ipsi te decipiuntet viam gressuum tuorum dissipant.
ISA|3|13|Surgit ad arguendum Dominuset stat ad iudicandos populos.
ISA|3|14|Dominus ad iudicium venietcum senibus populi sui et principibus eius: Vos enim depasti estis vineam,et rapina pauperis in domibus vestris.
ISA|3|15|Quare atteritis populum meumet facies pauperum commolitis? ",dicit Dominus, Deus exercituum.
ISA|3|16|Et dixit Dominus: Pro eo quod elevatae sunt filiae Sionet ambulaverunt extento collo et nutibus oculorum,parvis passibus incedebantet catenulis pedum tinniebant,
ISA|3|17|decalvabit Dominus verticem filiarum Sionet Dominus crinem earum nudabit ".
ISA|3|18|In die illa auferet Dominusornamentum calceamentorum et torques
ISA|3|19|et lunulas et inaureset armillas et mitras,
ISA|3|20|discriminalia et periscelidaset fascias et olfactoriola
ISA|3|21|et anulos et ornamenta narium,
ISA|3|22|mutatoria et palliolaet linteamina et marsupia,
ISA|3|23|specula et sindoneset vittas et pallia.
ISA|3|24|Et erit pro suavi odore foetor,et pro zona funiculus,et pro crispante crine calvitium,et pro fascia pectorali cilicium,stigma pro pulchritudine.
ISA|3|25|Viri tui gladio cadent,et fortes tui in proelio,
ISA|3|26|et maerebunt atque lugebunt portae eius,et desolata in terra sedebit.
ISA|4|1|Et apprehendent septem mulieresvirum unum in die illa dicentes: Panem nostrum comedemuset vestimentis nostris operiemur,tantummodo vocetur nomen tuum super nos:aufer opprobrium nostrum ".
ISA|4|2|In die illa erit germen Domini in splendorem et gloriam,et fructus terrae sublimis et exsultatiohis, qui salvati fuerint de Israel.
ISA|4|3|Et erit: omnis, qui relictus fuerit in Sion,et residuus in Ierusalem, sanctus vocabitur,omnis, qui scriptus est ad vitam in Ierusalem.
ISA|4|4|Cum abluerit Dominus sordem filiarum Sionet sanguinem Ierusalem laverit de medio eiusspiritu iudicii et spiritu ardoris,
ISA|4|5|et creabit Dominus super omnem locum montis Sionet super coetum eiusnubem per diemet fumum et splendorem ignis flammantis in nocte:super omnem enim gloriam protectio,
ISA|4|6|et tabernaculum erit in umbraculum diei ab aestuet in securitatem et absconsionem a turbine et a pluvia.
ISA|5|1|Cantabo dilecto meocanticum amici mei de vinea sua:Vinea facta est dilecto meoin colle pingui;
ISA|5|2|et saepivit eamet lapides elegit ex illaet plantavit in ea vites electaset aedificavit turrim in medio eiuset torcular exstruxit in ea;et exspectavit, ut faceret uvas,et fecit labruscas.
ISA|5|3|Nunc ergo, habitator Ierusalemet vir Iudae,iudicate inter me et vineam meam.
ISA|5|4|Quid est quod debui ultra facere vineae meaeet non feci ei?Cur exspectavi, ut faceret uvas,et fecit labruscas?
ISA|5|5|Et nunc ostendam vobisquid ego faciam vineae meae:auferam saepem eius,et erit in direptionem;diruam maceriam eius,et erit in conculcationem.
ISA|5|6|Et ponam eam desertam:non putabitur et non fodietur,et ascendent vepres et spinae;et nubibus mandabo, ne pluant super eam imbrem.
ISA|5|7|Vinea enim Domini exercituum domus Israel est,et vir Iudae germen eius delectabile;et exspectavi, ut faceret iudicium, et ecce iniquitas,et iustitiam, et ecce nequitia.
ISA|5|8|Vae, qui coniungunt domum ad domumet agrum agro copulant usque ad terminum loci!Numquid habitabitis vos soli in medio terrae?
ISA|5|9|In auribus meis iuravit Dominus exercituum: Certe domus multae desertae erunt,grandes et pulchrae absque habitatore ".
ISA|5|10|Decem enim iugera vinearum facient lagunculam unam,et triginta modii sementis facient modios tres.
ISA|5|11|Vae, qui consurgunt mane ad ebrietatem sectandamet ad potandum usque ad vesperam,ut vinum inflammet eos!
ISA|5|12|Cithara et lyraet tympanum et tibiaet vinum in conviviis eorum,et opus Domini non respiciunt,nec opera manuum eius considerant.
ISA|5|13|Propterea captivus ductus est populus meus,quia non habuit scientiam,et nobiles eius interierunt fame,et multitudo eius siti exaruit.
ISA|5|14|Propterea dilatavit infernus fauces suaset aperuit os suum absque ullo termino;et descendunt fortes Ierusalem, et populus eius,et sublimes et tripudiantes in ea.
ISA|5|15|Et incurvabitur homo, et humiliabitur vir,et oculi sublimium deprimentur;
ISA|5|16|et exaltabitur Dominus exercituum in iudicio,et Deus sanctus sanctificabitur in iustitia,
ISA|5|17|et pascentur agni iuxta ordinem suum velut in prato suo,et alieni comedent in ruinis pinguium.
ISA|5|18|Vae, qui trahunt iniquitatem in funiculis vanitatiset quasi vinculum plaustri peccatum!
ISA|5|19|Qui dicunt: " Festinetet cito veniat opus eius, ut videamus;et appropiet et veniat consilium Sancti Israel,et sciemus illud! ".
ISA|5|20|Vae, qui dicunt malum bonum et bonum malum,ponentes tenebras in lucem et lucem in tenebras,ponentes amarum in dulce et dulce in amarum!
ISA|5|21|Vae, qui sapientes sunt in oculis suiset coram ipsis prudentes!
ISA|5|22|Vae, qui potentes sunt ad bibendum vinum,et viri fortes ad miscendam ebrietatem!
ISA|5|23|Qui absolvunt impium pro muneribuset iustitiam iusti auferunt ab eo!
ISA|5|24|Propter hoc, sicut devorat stipulam lingua ignis,et palea flamma consumitur,sic radix eorum quasi tabes erit,et flos eorum sicut putredo ascendet;abiecerunt enim legem Domini exercituumet eloquium Sancti Israel blasphemaverunt.
ISA|5|25|Ideo exarsit furor Domini in populum suum,et extendit manum suam super eum et percussit eum,et conturbati sunt montes;et facta sunt morticina eorum quasi stercus in medio platearum.In his omnibus non est aversus furor eius,sed adhuc manus eius extenta.
ISA|5|26|Et levabit signum nationibus procul;et sibilabit ad eum de finibus terrae;et ecce festinus velociter veniet.
ISA|5|27|Non est deficiens neque laborans in eo,non dormitabit neque dormiet;neque solvetur cingulum renum eius,nec rumpetur corrigia calceamenti eius.
ISA|5|28|Sagittae eius acutae, et omnes arcus eius extenti;ungulae equorum eius ut silex reputantur,et rotae eius quasi impetus tempestatis.
ISA|5|29|Rugitus eius ut leonis:rugiet ut catuli leonum et frendet;et arripiet praedam et in tuto collocabit,et non erit qui eruat.
ISA|5|30|Et sonabit super eum in die illa sicut sonitus maris.Aspiciet in terram: et ecce tenebrae tribulationis,et lux obtenebrata est in caligine eius.
ISA|6|1|In anno, quo mortuus est rex Ozias, vidi Dominum edentem super solium excelsum et elevatum; et fimbriae eius replebant templum.
ISA|6|2|Seraphim stabant iuxta eum; sex alae uni et sex alae alteri: duabus velabat faciem suam et duabus velabat pedes suos et duabus volabat.
ISA|6|3|Et clamabat alter ad alterum et dicebat: Sanctus, Sanctus, Sanctus Dominus exercituum;plena est omnis terra gloria eius ".
ISA|6|4|Et commota sunt superliminaria cardinum a voce clamantis, et domus repleta est fumo.
ISA|6|5|Et dixi: Vae mihi, quia perii!Quia vir pollutus labiis ego sumet in medio populi polluta labia habentis ego habitoet regem, Dominum exercituum, vidi oculis meis ".
ISA|6|6|Et volavit ad me unus de seraphim, et in manu eius calculus, quem forcipe tulerat de altari,
ISA|6|7|et tetigit os meum et dixit: Ecce tetigit hoc labia tua,et auferetur iniquitas tua,et peccatum tuum mundabitur ".
ISA|6|8|Et audivi vocem Domini dicentis: " Quem mittam? Et quis ibit nobis? ". Et dixi: " Ecce ego, mitte me ".
ISA|6|9|Et dixit: " Vade, et dices populo huic:Audientes audite et nolite intellegere,et videntes videte et nolite cognoscere".
ISA|6|10|Pingue redde cor populi huiuset aures eius aggravaet oculos eius excaeca,ne forte videat oculis suiset auribus suis audiatet corde suo intellegat et convertaturet sanetur ".
ISA|6|11|Et dixi: " Usquequo, Domine? ". Et dixit: Donec desolenturcivitates absque habitatore,et domus sine homine,et terra relinquatur deserta ".
ISA|6|12|Et longe adducet Dominus homines,et magna erit desolatio in medio terrae;
ISA|6|13|et adhuc in ea decimatio,et rursus excisioni tradetursicut terebinthus et sicut quercus,in quibus deiectis manebit aliquid stabile.Semen sanctum erit id quod steterit in ea.
ISA|7|1|Et factum est in diebus Achaz filii Ioatham filii Oziae regis Iu dae, ascendit Rasin rex Syriae et Phacee filius Romeliae rex Israel in Ierusalem ad proeliandum contra eam; et non potuerunt debellare eam.
ISA|7|2|Et nuntiaverunt domui David dicentes: " Requievit Syria super Ephraim ". Et commotum est cor eius et cor populi eius, sicut moventur ligna silvarum a facie venti.
ISA|7|3|Et dixit Dominus ad Isaiam: " Egredere in occursum Achaz, tu et Seariasub (id est Reliquiae revertentur) filius tuus, ad extremum aquaeductus piscinae superioris in viam agri fullonis;
ISA|7|4|et dices ad eum: Vide, ut sileas; noli timere, et cor tuum ne formidet a duabus caudis titionum fumigantium istorum, ob ardorem irae Rasin et Syriae et filii Romeliae,
ISA|7|5|eo quod consilium malum inierit contra te Syria, Ephraim et filius Romeliae dicentes:
ISA|7|6|"Ascendamus ad Iudam et terrorem iniciamus ei et avellamus eum ad nos et ponamus regem in medio eius filium Tabeel" ".
ISA|7|7|Haec dicit Dominus Deus: Non stabit et non erit!
ISA|7|8|Caput enim Syriae Damascus,et caput Damasci Rasin;et adhuc sexaginta et quinque anniet desinet Ephraim esse populus;
ISA|7|9|et caput Ephraim Samaria,et caput Samariae filius Romeliae.Si non credideritis, non permanebitis ".
ISA|7|10|Et adiecit Dominus loqui ad Achaz dicens:
ISA|7|11|" Pete tibi signum a Domino Deo tuo in profundum inferni sive in excelsum supra ".
ISA|7|12|Et dixit Achaz: " Non petam et non tentabo Dominum ".
ISA|7|13|Et dixit: " Audite ergo, domus David; numquid parum vobis est molestos esse hominibus, quia molesti estis et Deo meo?
ISA|7|14|Propter hoc dabit Dominus ipse vobis signum. Ecce, virgo concipiet et pariet filium et vocabit nomen eius Emmanuel;
ISA|7|15|butyrum et mel comedet, ut ipse sciat reprobare malum et eligere bonum.
ISA|7|16|Quia antequam sciat puer reprobare malum et eligere bonum, desolabitur terra, cuius tu formidas duos reges;
ISA|7|17|adducet Dominus super te et super populum tuum et super domum patris tui dies, qui non venerunt a diebus separationis Ephraim a Iuda, regem Assyriorum ".
ISA|7|18|Et erit in die illa:sibilabit Dominus muscae,quae est in extremo fluminum Aegypti,et api, quae est in terra Assur;
ISA|7|19|et venient et requiescent omnesin vallibus praeruptiset in cavernis petrarumet in omnibus frutetiset in omnibus pascuis.
ISA|7|20|In die illa radet Dominusin novacula conducta e regione trans flumenC in rege Assyriorum Ccaput et pilos pedumet barbam quoque abradet.
ISA|7|21|Et erit in die illa:nutriet homo vitulam et duas oves
ISA|7|22|et prae ubertate lactiscomedet butyrum;butyrum enim et mel manducabit omnis,qui relictus fuerit in medio terrae.
ISA|7|23|Et erit in die illa:omnis locus, ubi fuerint mille vites mille argenteis,spinae et vepres erunt.
ISA|7|24|Cum sagittis et arcu ingredientur illuc,vepres enim et spinae erit universa terra.
ISA|7|25|Et in omnes montes, qui in sarculo sarriebantur,nemo veniet prae terrore spinarum et veprium,et erit in pascua bovis et in conculcationem pecoris.
ISA|8|1|Et dixit Dominus ad me: " Sume tibi tabulam grandem et scribe in ea stilo hominis: Maher Salal Has Baz (id est Velociter spolia detrahe, cito praedare).
ISA|8|2|Et adhibui mihi testes fideles, Uriam sacerdotem et Zachariam filium Barachiae;
ISA|8|3|et accessi ad prophetissam, et concepit et peperit filium. Et dixit Dominus ad me: " Voca nomen eius Maher Salal Has Baz,
ISA|8|4|quia antequam sciat puer clamare: "Pater mi" et "Mater mea", afferentur opes Damasci et spolia Samariae coram rege Assyriorum ".
ISA|8|5|Et adiecit Dominus loqui ad me adhuc dicens:
ISA|8|6|" Pro eo quod abiecit populus iste aquas Siloae,quae vadunt cum silentio,et defecit coram Rasin et filio Romeliae,
ISA|8|7|propter hoc ecce Dominus adducet super eosaquas Fluminis fortes et multas,regem Assyriorum et omnem gloriam eius,et ascendet super omnes rivos eiuset fluet super universas ripas eius;
ISA|8|8|et ibit per Iudam inundans et diffluens,usque ad collum veniet.Et erit extensio alarum eiusimplens latitudinem terrae tuae, o Emmanuel ".
ISA|8|9|Clamorem tollite, populi, et consternemini;et audite, universae procul terrae:accingimini et perterremini,accingimini et perterremini.
ISA|8|10|Inite consilium, et dissipabitur;loquimini verbum, et non fiet,quia nobiscum Deus.
ISA|8|11|Haec enim ait Dominus ad me, cum apprehendit me manu et monuit, ne irem in via populi huius, dicens:
ISA|8|12|" Ne vocetis coniurationem,quodcumque populus iste vocat coniurationem,et timorem eius ne timeatis neque paveatis ".
ISA|8|13|Dominum exercituum ipsum sanctificate:ipse pavor vester, et ipse terror vester;
ISA|8|14|et erit in sanctuarium,in lapidem offensionis et in petram scandaliduabus domibus Israel,in laqueum et in insidias habitantibus Ierusalem.
ISA|8|15|Et offendent ex eis plurimiet cadent et conterenturet irretientur et capientur.
ISA|8|16|Liga testimonium, signa legem in discipulis meis.
ISA|8|17|Et exspectabo Dominum, qui abscondit faciem suam a domo Iacob, et praestolabor eum.
ISA|8|18|Ecce ego et pueri, quos dedit mihi Dominus in signum et in portentum Israel a Domino exercituum, qui habitat in monte Sion.
ISA|8|19|Et cum dixerint ad vos: " Quaerite a pythonibus et a divinis, qui susurrant et murmurant; numquid non populus a deo suo requiret, pro vivis a mortuis? ".
ISA|8|20|Ad legem et ad testimonium! Quod si non dixerint iuxta verbum hoc, non erit eis matutina lux.
ISA|8|21|Et transibit per eam afflictus et esuriens;et, cum esurierit, irasceturet maledicet regi suo et deo suoet suspiciet sursum
ISA|8|22|et ad terram intuebitur:et ecce tribulatio et tenebrae,caligo opprimens et obscuritas diffusa.
ISA|8|23|Non erit enim amplius caligo,ubi erat oppressio.Primo tempore contemptibilem reddidit terram Zabulon et terram Nephthali; et novissimo glorificavit viam maris, trans Iordanem, Galilaeam gentium.
ISA|9|1|Populus, qui ambulabat in tenebris,vidit lucem magnam;habitantibus in regione umbrae mortislux orta est eis.
ISA|9|2|Multiplicasti exsultationemet magnificasti laetitiam;laetantur coram tesicut laetantes in messe,sicut exsultant, quando dividunt spolia.
ISA|9|3|Iugum enim oneris eiuset virgam umeri eiuset sceptrum exactoris eiusfregisti, sicut in die Madian.
ISA|9|4|Quia omnis caliga incedentis cum tumultuet vestimentum mixtum sanguineerit in combustionem, cibus ignis.
ISA|9|5|Parvulus enim natus est nobis,filius datus est nobis;et factus est principatus super umerum eius;et vocabitur nomen eiusadmirabilis Consiliarius, Deus fortis,Pater aeternitatis, Princeps pacis.
ISA|9|6|Magnum erit eius imperium,et pacis non erit finissuper solium David et super regnum eius,ut confirmet illud et corroboret in iudicio et iustitiaamodo et usque in sempiternum:zelus Domini exercituum faciet hoc.
ISA|9|7|Verbum misit Dominus in Iacob, et cecidit in Israel.
ISA|9|8|Et sciet omnis populus Ephraim et habitantes Samariamin superbia et magnitudine cordis dicentes:
ISA|9|9|" Lateres ceciderunt, sed quadris lapidibus aedificabimus;sycomori succisae sunt, sed cedris commutabimus ".
ISA|9|10|Et elevavit Dominus hostes super eumet inimicos eius excitavit,
ISA|9|11|Syriam ab oriente et Philisthim ab occidente,qui devoraverunt Israel toto ore.In omnibus his non est aversus furor eius,sed adhuc manus eius extenta.
ISA|9|12|Et populus non est reversus ad percutientem se,et Dominum exercituum non inquisierunt.
ISA|9|13|Et succidit Dominus ab Israel caput et caudam,palmam et arundinem die una:
ISA|9|14|longaevus et honorabilis vultu ipse est caput,et propheta docens mendacium ipse est cauda;
ISA|9|15|rectores populi istius seducenteset, qui regebantur, perierunt.
ISA|9|16|Propter hoc super adulescentulis eius non laetabitur Dominuset pupillorum eius et viduarum non miserebitur,quia omnis impius est et nequam,et universum os loquitur stultitiam.In omnibus his non est aversus furor eius,sed adhuc manus eius extenta.
ISA|9|17|Succensa est enim quasi ignis impietas,veprem et spinam vorat,et succenditur in densitate saltus,et convolvuntur columnae fumi.
ISA|9|18|In ira Domini exercituum incenditur terra;et est populus quasi esca ignis:vir fratri suo non parcit.
ISA|9|19|Et devorat ad dexteram et esuritet comedit ad sinistram et non saturatur;unusquisque carnem proximi sui vorat:
ISA|9|20|Manasses Ephraim, et Ephraim Manassen,simul ipsi contra Iudam.In omnibus his non est aversus furor eius,sed adhuc manus eius extenta.
ISA|10|1|Vae, qui condunt leges iniquaset scribentes iniustitiam scribunt,
ISA|10|2|ut opprimant in iudicio paupereset vim faciant causae humilium populi mei,ut fiant viduae praeda eorum,et pupillos diripiant!
ISA|10|3|Quid facietis in die visitationiset calamitatis de longe venientis?Ad cuius confugietis auxiliumet ubi derelinquetis gloriam vestram?
ISA|10|4|Nam incurvabimini subter captivoset infra occisos cadetis.In omnibus his non est aversus furor eius,sed adhuc manus eius extenta.
ISA|10|5|Vae Assur, virga furoris meiet baculus in manu mea, indignatio mea!
ISA|10|6|Ad gentem impiam mitto eumet contra populum furoris mei mando illi,ut auferat spolia et diripiat praedamet ponat illum in conculcationemquasi lutum platearum.
ISA|10|7|Ipse autem non sic arbitratur,et cor eius non ita existimat;sed in corde suo ad conterendumet ad internecionem gentium non paucarum.
ISA|10|8|Dicet enim: " Numquid non principes mei omnes reges sunt?
ISA|10|9|Numquid non ut Charcamis sic Chalano?Numquid non ut Arphad sic Emath?Numquid non ut Damascus sic Samaria?
ISA|10|10|Quomodo apprehendit manus mea regna idololatra,quorum simulacra plura sunt quam in Ierusalem et in Samaria,
ISA|10|11|numquid non sicut feci Samariae et idolis eius,sic faciam Ierusalem et simulacris eius? ".
ISA|10|12|Et erit: cum impleverit Dominus cuncta opera sua in monte Sion et in Ierusalem, visitabo super fructum superbiae cordis regis Assyriae et super arrogantiam altitudinis oculorum eius.
ISA|10|13|Dixit enim: In fortitudine manus meae feciet in sapientia mea, prudens sum enim;et abstuli terminos populorumet scrinia eorum depraedatus sumet detraxi quasi potens in sublimi sedentes;
ISA|10|14|et apprehendit quasi nidum manus mea fortitudinem populorum;et sicut colliguntur ova derelicta,sic universam terram ego congregavi,et non fuit qui moveret pennam aut aperiret os et ganniret ".
ISA|10|15|Numquid gloriabitur securiscontra eum, qui secat in ea?Aut exaltabitur serracontra eum, qui trahit eam?Quomodo si agitet virga elevantem eam,et exaltet baculus eum, qui non est lignum.
ISA|10|16|Propter hoc mittet Dominator, Dominus exercituum,in pingues eius tenuitatem;et subtus gloriam eiusardor ardebit quasi combustio ignis.
ISA|10|17|Et erit Lumen Israel ignis,et Sanctus eius flamma;et succendetur et devorabit spinas eiuset vepres in die una.
ISA|10|18|Et gloriam saltus eius et horti eiusab anima usque ad carnem consumet,et erit sicut aeger tabescens;
ISA|10|19|et reliquiae ligni saltus eiustam paucae erunt,ut puer scribat ea.
ISA|10|20|Et erit in die illa:non adiciet residuum Israelet, qui effugerint de domo Iacob,inniti super eo, qui percutit eos,sed innitentur super Dominum,Sanctum Israel, in veritate.
ISA|10|21|Reliquiae revertentur,reliquiae, inquam, Iacob, ad Deum fortem.
ISA|10|22|Si enim fuerit populus tuus, Israel, quasi arena maris,reliquiae revertentur ex eo;consummatio decreta redundat in iustitia:
ISA|10|23|interitum enim, qui decretus est,Dominus, Deus exercituum, faciet in medio omnis terrae.
ISA|10|24|Propter hoc haec dicit Dominus, Deus exercituum: " Noli timere, populus meus habitator Sion, ab Assur; in virga percutiet te et baculum suum levabit super te sicut Aegyptus.
ISA|10|25|Adhuc enim paululum modicumque, et consummabitur indignatio et furor meus ad destructionem eorum ".
ISA|10|26|Et suscitabit super eum Dominus exercituum flagellum iuxta plagam Madian in Petra Oreb et virgam suam super mare et levabit eam sicut in Aegypto.
ISA|10|27|Et erit in die illa:auferetur onus eius de umero tuo,et iugum eius de collo tuo.Et vastator ascendit a Remmon.
ISA|10|28|Veniet in Aiath, transibit per Magron,apud Machmas deponit sarcinas suas;
ISA|10|29|transeunt vadum cursim; in Geba pernoctabimus;trepidat Rama, Gabaa Saulis fugit.
ISA|10|30|Hinni voce tua, Bathgallim;attende, Laisa; responde, Anathoth.
ISA|10|31|Migrat Medemena, habitatores Gabim fugiunt;
ISA|10|32|hodie in Nob stabit:agitabit manum suam ad montem filiae Sion,collem Ierusalem.
ISA|10|33|Ecce Dominator, Dominus exercituum,amputat ramos in terrore,et extrema acumina succiduntur,et sublimes humiliantur;
ISA|10|34|et caeduntur condensa saltus ferro,et Libanus cum excelsis suis cadet.
ISA|11|1|Et egredietur virga de stirpe Iesse,et flos de radice eius ascendet;
ISA|11|2|et requiescet super eum spiritus Domini:spiritus sapientiae et intellectus,spiritus consilii et fortitudinis,spiritus scientiae et timoris Domini;
ISA|11|3|et deliciae eius in timore Domini.Non secundum visionem oculorum iudicabitneque secundum auditum aurium decernet;
ISA|11|4|sed iudicabit in iustitia paupereset decernet in aequitate pro mansuetis terrae;et percutiet terram virga oris suiet spiritu labiorum suorum interficiet impium.
ISA|11|5|Et erit iustitia cingulum lumborum eius,et fides cinctorium renum eius.
ISA|11|6|Habitabit lupus cum agno,et pardus cum haedo accubabit;vitulus et leo simul saginabuntur,et puer parvulus minabit eos.
ISA|11|7|Vitula et ursus pascentur,simul accubabunt catuli eorum;et leo sicut bos comedet paleas.
ISA|11|8|Et ludet infans ab uberesuper foramine aspidis;et in cavernam reguli,qui ablactatus fuerit, manum suam mittet.
ISA|11|9|Non nocebunt et non occidentin universo monte sancto meo,quia plena erit terra scientia Domini, sicut aquae mare operiunt.
ISA|11|10|In die illa radix Iessestat in signum populorum;ipsam gentes requirent,et erit sedes eius gloriosa.
ISA|11|11|Et erit in die illa: rursus extendet Dominus manum suamad possidendum residuum populi sui,quod relictum erit ab Assyria et ab Aegyptoet a Phatros et ab Aethiopiaet ab Elam et a Sennaaret ab Emath et ab insulis maris;
ISA|11|12|et levabit signum in nationeset congregabit profugos Israelet dispersos Iudae colliget a quattuor plagis terrae.
ISA|11|13|Et auferetur zelus Ephraim,et hostes Iudae abscindentur;Ephraim non aemulabitur Iudam, et Iudas non pugnabit contra Ephraim.
ISA|11|14|Et volabunt in umeros Philisthim ad mare,simul praedabuntur filios orientis:in Edom et Moab extendent manus suas,et filii Ammon oboedient eis.
ISA|11|15|Et exsiccabit Dominus linguam maris Aegyptiet levabit manum suam super flumen in fortitudine spiritus suiet percutiet illud in septem rivos,ita ut transire faciat eos calceatos.
ISA|11|16|Et erit via residuo populo meo,qui relinquetur ab Assyria,sicut fuit Israeli in die illa,qua ascendit de terra Aegypti.
ISA|12|1|Et dices in die illa: Confitebor tibi, Domine,quoniam cum iratus eras mihi,conversus est furor tuus, et consolatus es me.
ISA|12|2|Ecce Deus salutis meae;fiducialiter agam et non timebo,quia fortitudo mea et laus mea Dominus,et factus est mihi in salutem ".
ISA|12|3|Et haurietis aquas in gaudio de fontibus salutis.
ISA|12|4|Et dicetis in die illa: Confitemini Domino et invocate nomen eius,notas facite in populis adinventiones eius;mementote quoniam excelsum est nomen eius.
ISA|12|5|Cantate Domino, quoniam magnifice fecit;notum sit hoc in universa terra.
ISA|12|6|Exsulta et lauda, quae habitas in Sion,quia magnus in medio tui Sanctus Israel ".
ISA|13|1|Oraculum Babylonis, quod vidit Isaias filius Amos.
ISA|13|2|Super montem decalvatum levate signum,exaltate vocem, levate manum,et ingrediantur portas ducum.
ISA|13|3|Ego mandavi sanctificatis meiset vocavi fortes meos ad iram meam,exsultantes in gloria mea.
ISA|13|4|Vox multitudinis in montibus quasi populi ingentis,vox sonitus regnorum gentium congregatarum.Dominus exercituum recenset militiam belli;
ISA|13|5|veniunt de terra procul a termino caeli,Dominus et vasa furoris eius,ut disperdat omnem terram.
ISA|13|6|Ululate, quia prope est dies Domini;quasi vastitas a Domino veniet.
ISA|13|7|Propter hoc omnes manus dissolventur,et omne cor hominis tabescet.
ISA|13|8|Perterrebuntur.Torsiones et dolores tenebunt eos,quasi parturiens dolebunt;unusquisque ad proximum suum stupebit:facies combustae vultus eorum.
ISA|13|9|Ecce dies Domini venit,crudelis et indignationis plenuset irae furorisque,ad ponendam terram in solitudinem,et peccatores eius conteret de ea.
ISA|13|10|Quoniam stellae caeli et sidera eiusnon expandent lumen suum;obtenebratus est sol in ortu suo,et luna non splendebit in lumine suo.
ISA|13|11|Et visitabo super orbem propter malaet super impios propter iniquitatem eorum;et quiescere faciam superbiam protervorumet arrogantiam fortium humiliabo.
ISA|13|12|Pretiosior erit vir auro,et homo mundo obryzo.
ISA|13|13|Super hoc caelum turbabo,et movebitur terra de loco suoin indignatione Domini exercituumet in die irae furoris eius.
ISA|13|14|Et erit quasi damula fugiens et quasi ovis,et non erit qui congreget;unusquisque ad populum suum convertetur,et singuli ad terram suam fugient.
ISA|13|15|Omnis, qui inventus fuerit, occidetur,et omnis, qui captus fuerit, cadet in gladio;
ISA|13|16|infantes eorum allidentur in oculis eorum,diripientur domus eorum,et uxores eorum violabuntur.
ISA|13|17|Ecce ego suscitabo super eos Medos,qui argentum non quaerant nec aurum velint;
ISA|13|18|sed arcus pueros prosternentet fructui uteri non miserebuntur.
ISA|13|19|Et erit Babylon, splendor regnorum,inclita superbia Chaldaeorum,sicut cum subvertit Dominus Sodomam et Gomorram.
ISA|13|20|Non habitabitur usque in finemet non fundabitur usque ad generationem et generationem,nec ponet ibi tentoria Arabs,nec pastores accubare facient ibi,
ISA|13|21|sed accubabunt ibi bestiae,et replebunt domus eorum ululae,et habitabunt ibi struthiones,et pilosi saltabunt ibi;
ISA|13|22|et respondebunt ibi hyaenae in aedibus eius,et thoes in delubris voluptatis.Prope est ut veniat tempus eius,et dies eius non elongabuntur.
ISA|14|1|Miserebitur enim Dominus Iacobet eliget adhuc de Israelet requiescere eos faciet super humum suam;adiungetur advena ad eoset adhaerebit domui Iacob.
ISA|14|2|Et tenebunt eos populiet adducent eos in locum suum;et possidebit eos domus Israelsuper terram Domini in servos et ancillas;et erunt capientes eos, qui se ceperant,et subicient exactores suos.
ISA|14|3|Et erit in die illa:cum requiem dederit tibi Dominusa labore tuo et a concussione tuaet a servitute dura, qua ante servisti,
ISA|14|4|proferes parabolam istam contra regem Babylonis et dices: Quomodo cessavit exactor, quievit oppressio?
ISA|14|5|Contrivit Dominus baculum impiorum,virgam dominantium,
ISA|14|6|caedentem populos in indignatione plaga sine remissione,subicientem in furore gentes persecutione sine fine.
ISA|14|7|Conquievit et siluit omnis terra,gavisa est, et exsultaverunt.
ISA|14|8|Abietes quoque laetatae sunt super te, et cedri Libani:Ex quo dormisti, non ascendit, qui succidat nos".
ISA|14|9|Infernus subter conturbatus estin occursum adventus tui;suscitat tibi umbras, omnes principes terraesurgere fecit de soliis suis,omnes reges nationum.
ISA|14|10|Universi respondebunt et dicent tibi:Et tu vulneratus es sicut nos,nostri similis effectus es".
ISA|14|11|Detracta est ad inferos superbia tua,sonitus nablorum tuorum;subter te sternitur tinea,et operimentum tuum sunt vermes.
ISA|14|12|Quomodo cecidisti de caelo, lucifer, fili aurorae?Deiectus es in terram, qui deiciebas gentes,
ISA|14|13|qui dicebas in corde tuo:In caelum conscendam,super astra Dei exaltabo solium meum,sedebo in monte conventusin lateribus aquilonis;
ISA|14|14|ascendam super altitudinem nubium,similis ero Altissimo".
ISA|14|15|Verumtamen ad infernum detractus es,in profundum laci.
ISA|14|16|Qui te viderint, te intuenturteque prospicient:Numquid iste est vir, qui conturbavit terram,qui concussit regna,
ISA|14|17|qui posuit orbem desertumet urbes eius destruxit,vinctis eius non aperuit carcerem?
ISA|14|18|Omnes reges gentium universi dormiunt in gloria,vir in domo sua;
ISA|14|19|tu autem proiectus es de sepulcro tuoquasi stirps abominabilis,obvolutus cum his, qui interfecti sunt gladioet descenderunt ad lapides sepulcri,quasi cadaver conculcatum.
ISA|14|20|Non habebis consortium cum eis in sepultura;tu enim terram tuam disperdidisti,tu populum tuum occidisti:non vocabitur in aeternum semen malefactorum.
ISA|14|21|Praeparate filios eius occisioniob iniquitatem patrum suorum;ne consurgant, ut hereditent terram,neque impleant faciem orbis civitatum" ".
ISA|14|22|" Et consurgam contra eos,dicit Dominus exercituum;et perdam Babylonis nomen et reliquiaset germen et progeniem, dicit Dominus;
ISA|14|23|et ponam eam in possessionem ericiiet in paludes aquarum,et scopabo eam in scopa destructionis ",dicit Dominus exercituum.
ISA|14|24|Iuravit Dominus exercituum dicens: Profecto, ut putavi, ita erit;et quomodo mente tractavi, sic eveniet.
ISA|14|25|Conteram Assyrium in terra meaet in montibus meis conculcabo eum;et auferetur ab eis iugum eius,et onus illius ab umero eorum tolletur ".
ISA|14|26|Hoc consilium, quod initum estsuper omnem terram,et haec est manus extentasuper universas gentes.
ISA|14|27|Dominus enim exercituum decrevit,et quis poterit infirmare?Et manus eius extenta,et quis avertet eam?
ISA|14|28|In anno, quo mortuus est rex Achaz, factum est oraculum istud:
ISA|14|29|" Ne laeteris, Philisthaea omnis tu,quoniam comminuta est virga percussoris tui;de radice enim colubri egredietur regulus,et semen eius draco volans.
ISA|14|30|Et pascentur primogeniti egenorum,et pauperes fiducialiter requiescent;et interire faciam in fame radicem tuamet reliquias tuas interficiam.
ISA|14|31|Ulula, porta! Clama, civitas!Contremisce, Philisthaea omnis;ab aquilone enim fumus venit,et non est fugitivus in agminibus eius ".
ISA|14|32|Et quid respondebitur nuntiis gentis? Quia Dominus fundavit Sion,et in ipsam confugiunt pauperes populi eius ".
ISA|15|1|Oraculum Moab.Quia nocte vastata est Ar moab, conticuit;quia nocte vastata est Cirmoab, conticuit.
ISA|15|2|Ascendit filia Dibon ad excelsa in planctum;super Nabo et super Medaba Moab ululavit;in cunctis capitibus eius calvitium, omnis barba rasa.
ISA|15|3|In triviis eius accincti sunt sacco;super tecta eius et in plateis eiusomnes ululant, prorumpunt in fletum.
ISA|15|4|Clamat Hesebon et Eleale,usque Iasa auditur vox eorum;super hoc expediti Moab fremunt,anima eius fremit sibi.
ISA|15|5|Cor meum super Moab clamat,vectes eius usque ad Segor, Eglatselisiam;per ascensum enim Luith flentes ascenduntet in via Oronaim clamorem contritionis levant.
ISA|15|6|Aquae enim Nemrim desertae erunt,quia aruit herba, defecit germen,viror omnis interiit.
ISA|15|7|Ideo supellectiles colligunt, copias divitiarum suastrans torrentem Salicum ducunt.
ISA|15|8|Quoniam circuivit clamor terminum Moab;usque ad Eglaim ululatus eius,et usque ad Beerelim clamor eius.
ISA|15|9|Quia aquae Dimon repletae sunt sanguine;ponam enim super Dimon additamentahis, qui fugerint de Moab leonem, et reliquiis terrae.
ISA|16|1|Emittite agnum dominatori terraede Petra deserti ad montem filiae Sion.
ISA|16|2|Et erit: sicut avis fugiens,et pulli de nido avolantes,sic erunt filiae Moabad vada Arnon.
ISA|16|3|Affer consilium, fac iudicium;pone quasi noctem umbram tuam in meridie,absconde fugientes et vagos ne prodas.
ISA|16|4|Habitent apud te profugi Moab;esto latibulum eorum a facie vastatoris;finitus est enim exactor,consummata est devastatio,defecit calcator a terra.
ISA|16|5|Et firmabitur in misericordia solium;et sedebit super illud in veritate,in tabernaculo David, iudicans et quaerens iudiciumet velociter reddens, quod iustum est.
ISA|16|6|Audivimus superbiam MoabC superbus est valde Csuperbiam eius et arrogantiam eius et indignationem eiuset iactantiam eius non rectam.
ISA|16|7|Idcirco ululabit Moab super Moab,omnes ululabunt;super placentas Cirharesethlamentantur percussi.
ISA|16|8|Quoniam suburbana Hesebon deserta sunt et vinea Sabama;dominos gentium perdiderunt uvae eius;usque ad Iazer pervenerunt,erraverunt in deserto:propagines eius diffusae sunt,transierunt mare.
ISA|16|9|Super hoc plorabo in fletu Iazer vineam Sabama;inebriabo te lacrima mea, Hesebon et Eleale,quoniam super vindemiam tuam et super messem tuamclamor cecidit.
ISA|16|10|Et ablata est laetitia et exsultatio de hortis,et in vineis non exsultant neque iubilant.Vinum in torculari non calcabit, qui calcare consueverat;clamor cessavit.
ISA|16|11|Ideo venter meus super Moab quasi cithara fremit,et viscera mea super Cirhareseth.
ISA|16|12|Et erit: cum apparueritet laboraverit Moab super excelsis,ingredietur ad sancta sua, ut obsecret,et non valebit.
ISA|16|13|Et hoc verbum, quod locutus est Dominus ad Moab ex tunc;
ISA|16|14|nunc autem loquitur Dominus dicens: " In tribus annis, quasi anni mercennarii, auferetur gloria Moab cum omni populo multo, et residuum parvum et modicum nequaquam ingens erit ".
ISA|17|1|Oraculum Damasci. Ecce Damascus desinet esse civitaset erit sicut acervus ruinarum.
ISA|17|2|Derelictae civitates Aroer gregibus erunt;et requiescent ibi, et non erit qui exterreat.
ISA|17|3|Et auferetur munimentum ab Ephraimet regnum a Damasco,et reliquiae Syriae sicut gloria filiorum Israel erunt,dicit Dominus exercituum.
ISA|17|4|Et erit in die illa: attenuabitur gloria Iacob,et pinguedo carnis eius marcescet;
ISA|17|5|et erit, sicut cum messor arripit culmos,et brachium eius spicas legit;et erit, sicut cum quis quaerit spicas in valle Raphaim.
ISA|17|6|Et relinquetur in eo racemus,et sicut cum excutitur olea:duae vel tres olivae in summitate ramisive quattuor aut quinque in cacuminibus arboris fructiferae ",dicit Dominus Deus Israel.
ISA|17|7|In die illa attendet homo ad factorem suum,et oculi eius ad Sanctum Israel respicient;
ISA|17|8|et non attendet ad altaria,quae fecerunt manus eius,et quae operati sunt digiti eius;non respiciet lucos et thymiateria.
ISA|17|9|In die illa erunt civitates fortitudinis eius derelictae,sicut civitates, quas dereliquerunt Hevaei et Amorraeia facie filiorum Israel;et erit desolatio,
ISA|17|10|quia oblita es Dei salutis tuaeet petrae fortitudinis tuae non es recordata:propterea plantabis plantationes iucundaset germen alienum seminabis.
ISA|17|11|In ipso die plantationis tuae saepies easet mane semen tuum florere facies;evanescet messis in die penuriae,et dolor insanabilis erit.
ISA|17|12|Heu!, strepitus populorum multorum;strepunt quasi strepitu maris,et tumultus turbarumquasi sonitu aquarum sonabunt.
ISA|17|13|Sonabunt populi sicut sonitus aquarum inundantium,et increpabit eum, et fugiet procul;et rapietur sicut pulvis montium a facie ventiet sicut turbo coram tempestate.
ISA|17|14|In tempore vespere, et ecce turbatio,ante matutinum non subsistet:haec est pars eorum, qui vastaverunt nos,et sors diripientium nos.
ISA|18|1|Vae terrae alarum strepitantium,quae est trans flumina Aethiopiae!
ISA|18|2|Quae mittit in mari legatoset in vasis papyri super aquas: Ite, nuntii veloces,ad gentem proceram et lucidam,ad populum terribilem,prope et procul,gentem robustam et conculcantem,cuius flumina scindunt terram ".
ISA|18|3|Omnes habitatores orbiset in terra commorantes,cum elevatum fuerit signum in montibus, videbitiset, cum clanguerit tuba, audietis.
ISA|18|4|Quia haec dixit Dominus ad me: Quiescam et considerabo in loco meo,sicut calor torrens orta iam luceet sicut nubes roris in aestu messis ".
ISA|18|5|Etenim ante vindemiam, cum consummatus fuerit flos,et uva germinans maturescens erit,praecidet ramusculos falcibuset propagines abscindet et proiciet;
ISA|18|6|et relinquentur simul avibus montiumet bestiis terrae;et aestate erunt super ea volucres,et omnes bestiae terrae super illa hiemabunt.
ISA|18|7|In tempore illo deferetur munus Domino exercituum a populo procero et lucido, a populo terribili, prope et procul, a gente robusta et conculcante, cuius terram flumina scindunt, ad locum nominis Domini exercituum, montem Sion.
ISA|19|1|Oraculum Aegypti.Ecce Dominus vehitur super nubem levemet ingreditur Aegyptum;et commovebuntur simulacra Aegypti a facie eius,et cor Aegypti tabescet in medio eius.
ISA|19|2|" Et concurrere faciam Aegyptios adversus Aegyptios;et pugnabit vir contra fratrem suum,et vir contra amicum suum,civitas adversus civitatem,regnum adversus regnum.
ISA|19|3|Et dirumpetur spiritus Aegypti in visceribus eius,et consilium eius confundam;et interrogabunt simulacra et divinoset pythones et hariolos.
ISA|19|4|Et tradam Aegyptios in manu domini crudelis,et rex fortis dominabitur eorum ",ait Dominus, Deus exercituum.
ISA|19|5|Et arescet aqua de mari,et fluvius desolabitur atque siccabitur,
ISA|19|6|et putrida fient flumina;attenuabuntur et siccabuntur rivi Aegypti,calamus et iuncus marcescent;
ISA|19|7|nudabuntur ripae Nili,et omnis planta Nili siccabitur;arescet et non erit.
ISA|19|8|Et maerebunt piscatores,et lugebunt omnes mittentes in flumen hamum;et expandentes rete super faciem aquarum languebunt.
ISA|19|9|Confundentur, qui operantur linum,pectentes et texentes byssum.
ISA|19|10|Et opifices eius deprimentur,omnes mercennarii omnino deficient.
ISA|19|11|Quam stulti principes Taneos!Sapientes consiliarii pharaonis dederunt consilium insipiens;quomodo dicetis pharaoni: Filius sapientium ego, filius regum antiquorum "?
ISA|19|12|Ubi nunc sunt sapientes tui?Annuntient tibi et indicentquid cogitaverit Dominus exercituum super Aegyptum.
ISA|19|13|Stulti facti sunt principes Taneos,decepti sunt principes Mempheos,deceperunt Aegyptum anguli tribuum eius.
ISA|19|14|Dominus miscuit in medio eius spiritum vertiginis,et errare fecerunt Aegyptum in omni opere suo,sicut errat ebrius in vomitu suo;
ISA|19|15|et non erit Aegypto opus,quod faciat, caput vel cauda, palma vel arundo.
ISA|19|16|In die illa erunt Aegyptii quasi mulieres et stupebunt et timebunt a facie commotionis manus Domini exercituum, quam ipse movebit super eam.
ISA|19|17|Et erit terra Iudae Aegypto in pavorem: omnis, qui illius fuerit recordatus, pavebit a facie consilii Domini exercituum, quod ipse cogitavit super eam.
ISA|19|18|In die illa erunt quinque civitates in terra Aegypti loquentes lingua Chanaan et iurantes per Dominum exercituum. Civitas Solis vocabitur una.
ISA|19|19|In die illa erit altare Domino in medio terrae Aegypti, et titulus iuxta terminum eius Domino.
ISA|19|20|Et erit in signum et in testimonium Domino exercituum in terra Aegypti. Clamabunt enim ad Dominum a facie tribulantium, et mittet eis salvatorem et propugnatorem, qui liberet eos.
ISA|19|21|Et cognoscetur Dominus ab Aegypto, et cognoscent Aegyptii Dominum in die illa; et colent eum in hostiis et in muneribus et vota vovebunt Domino et solvent.
ISA|19|22|Et percutiet Dominus Aegyptum plaga et sanabit; et revertentur ad Dominum, et placabitur eis et sanabit eos.
ISA|19|23|In die illa erit via de Aegypto in Assyriam; et intrabit Assyrius Aegyptum, et Aegyptius in Assyriam, et servient Aegyptii cum Assyriis.
ISA|19|24|In die illa erit Israel tertius cum Aegypto et Assyria; benedictio in medio terrae,
ISA|19|25|cui benedicet Dominus exercituum dicens: " Benedictus populus meus Aegyptius, et opus manuum mearum Assyrius, et hereditas mea Israel ".
ISA|20|1|In anno quo ingressus est Tharthan in Azotum, cum misisset eum Sargon rex Assyriorum, et pugnasset contra Azotum et cepisset eam,
ISA|20|2|in tempore illo locutus est Dominus in manu Isaiae filii Amos dicens: " Vade et solve saccum de lumbis tuis et calceamenta tua tolle de pedibus tuis ". Et fecit sic, vadens nudus et discalceatus.
ISA|20|3|Et dixit Dominus: " Sicut ambulavit servus meus Isaias nudus et discalceatus tribus annis signum et portentum super Aegyptum et super Aethiopiam,
ISA|20|4|sic minabit rex Assyriorum captivos Aegypti et exsules Aethiopiae, iuvenes et senes, nudos et discalceatos, discoopertis natibus ad ignominiam Aegypti.
ISA|20|5|Et timebunt et confundentur ab Aethiopia spe sua et ab Aegypto gloria sua.
ISA|20|6|Et dicet habitator maritimae regionis huius in die illa: "Ecce, haec erat spes nostra, quo confugimus in auxilium, ut liberaremur a facie regis Assyriorum; et quomodo effugere poterimus nos?" ".
ISA|21|1|Oraculum deserti maris.Sicut turbines per austrum transeuntes,de deserto venit, de terra horribili.
ISA|21|2|Visio dura nuntiata est mihi:praedo praedatur,et vastator vastat.Ascende, Elam;obside, Media;omnem gemitum eius cessare feci.
ISA|21|3|Propterea repleti sunt lumbi mei tremore,angustia possedit me sicut angustia parientis;corrui, cum audirem;conturbatus sum, cum viderem.
ISA|21|4|Vacillat cor meum,pavor invadit me:crepusculum optatumposuit mihi in terrorem.
ISA|21|5|Ponunt mensam,stragulum pandunt, comedunt, bibunt.Surgite, principes,ungite clipeum.
ISA|21|6|Haec enim dixit mihi Dominus: Vade et pone speculatorem;quodcumque viderit, annuntiet.
ISA|21|7|Si viderit currum, bigam equitum,ascensorem asini et ascensorem cameli,intueatur diligenter multo intuitu ".
ISA|21|8|Et clamavit speculator: Super specula, Domine,ego sum stans iugiter per diem,et super custodiam meamego sum stans totis noctibus.
ISA|21|9|Ecce, huc venit agmen virorum,biga equitum ".Et respondit et dixit: Cecidit, cecidit Babylon,et omnia sculptilia deorum eiuscontrita sunt in terram ".
ISA|21|10|Tritura mea et fili areae meae,quae audivi a Domino exercituum, Deo Israel,annuntiavi vobis.
ISA|21|11|Oraculum Duma.Ad me clamat ex Seir: Custos, quid de nocte?Custos, quid de nocte? ".
ISA|21|12|Dixit custos: Venit mane, sed etiam nox;si quaeritis, quaerite,revertimini, venite ".
ISA|21|13|Oraculum in solitudine.In saltu, in solitudine dormietis,turmae Dedanim.
ISA|21|14|Occurrentes sitienti ferte aquam,qui habitatis terram Thema;cum panibus occurrite fugienti:
ISA|21|15|a facie enim gladiorum fugerunt,a facie gladii nudati,a facie arcus extenti,a facie gravis proelii.
ISA|21|16|Quoniam haec dicit Dominus ad me: " Adhuc anno sicut anni mercennarii, et auferetur omnis gloria Cedar;
ISA|21|17|et reliquiae numeri arcuum fortium filiorum Cedar imminuentur; Dominus enim, Deus Israel, locutus est ".
ISA|22|1|Oraculum vallis Visionis.Quidnam tibi est,quia ascendisti omnis in tecta,
ISA|22|2|clamoris plena, urbs tumultuans,civitas exsultans?Interfecti tui non interfecti gladionec mortui in bello;
ISA|22|3|cuncti principes tui fugeruntsimul sine arcu capti;omnes, qui inventi sunt, capti sunt simul,procul fugerunt.
ISA|22|4|Propterea dixi: " Recedite a me,amare flebo;nolite incumbere, ut consolemini mesuper vastitate filiae populi mei ".
ISA|22|5|Dies enim confusioniset conculcationis et fletusDomino, Deo exercituum, in valle Visionis,eversio murorum et vociferatio ad montem.
ISA|22|6|Et Elam sumpsit pharetram,in agmine hominum equitum,et Cir nudavit clipeum.
ISA|22|7|Et electae valles tuaeplenae sunt quadrigarum,et equites ponunt sedes suas in porta.
ISA|22|8|Et revelatum est operimentum Iudae,et respexisti in die illa armamentarium domus Saltus;
ISA|22|9|et scissuras civitatis David vidistis,quia multiplicatae sunt;et congregastis aquas piscinae inferioris.
ISA|22|10|Et domos Ierusalem numerastiset destruxistis domosad muniendum murum;
ISA|22|11|et lacum fecistis inter duos murospro aqua piscinae veteris;sed non suspexistis ad eum, qui fecit haec,et eum, qui haec de longe formavit, non vidistis.
ISA|22|12|Et vocavit Dominus, Deus exercituum, in die illaad fletum et ad planctum,ad calvitium et ad cingendum saccum;
ISA|22|13|et ecce gaudium et laetitia,occidere boves et iugulare pecus,comedere carnes et bibere vinum: Comedamus et bibamus,cras enim moriemur ".
ISA|22|14|Et revelatum est in auribus meisa Domino exercituum: Certe non dimittetur iniquitas haec vobis, donec moriamini! ",dicit Dominus, Deus exercituum.
ISA|22|15|Haec dicit Dominus, Deus exercituum: Vade, ingredere ad procuratorem istum,ad Sobnam praepositum palatii:
ISA|22|16|"Quid tibi hic? Aut quis tibi hic,quia excidisti tibi hic sepulcrum?".Effodiens in excelso sepulcrum suum,excavabat in petra tabernaculum sibi.
ISA|22|17|Ecce Dominus vehementer proiciet te, homo,violenter te apprehendens.
ISA|22|18|In globum te convolvet glomerans;quasi pilam mittet tein terram latam et spatiosam:ibi morieris,et ibi erunt currus gloriae tuae,ignominia domus domini tui.
ISA|22|19|Et expellam te de statione tuaet de ministerio tuo deponam te.
ISA|22|20|Et erit in die illa:vocabo servum meum Eliachim filium Helciae
ISA|22|21|et induam illum tunicam tuamet cingulo tuo cingam eumet potestatem tuam dabo in manu eius;et erit in patrem habitantibus Ierusalemet domui Iudae.
ISA|22|22|Et dabo clavem domus Davidsuper umerum eius;et aperiet, et non erit qui claudat;et claudet, et non erit qui aperiat.
ISA|22|23|Et figam illum paxillum in loco securo,et erit in solium gloriae domui patris sui.
ISA|22|24|Et suspendent super eum omnem gloriam domus patris sui, propagines et stirpes, omne vas parvulum, a pelvibus ad amphoras.
ISA|22|25|In die illa, dicit Dominus exercituum, auferetur paxillus, qui fixus fuerat in loco securo, et frangetur et cadet; et peribit, quod pependerat in eo, quia Dominus locutus est ".
ISA|23|1|Oraculum Tyri.Ululate, naves Tharsis,quia vastatum est refugium vestrum;cum redirent de terra Cetthim, revelatum est eis.
ISA|23|2|Obstupescite, qui habitatis in insula;negotiatores Sidonistransfretantes mare repleverunt te.
ISA|23|3|In aquis multis semen Nili,messis fluminis fruges eius;et facta est negotiatio gentium.
ISA|23|4|Erubesce, Sidon, ait enim mare,fortitudo maris, dicens: Non parturivi et non peperi;et non enutrivi iuvenesnec virgines educavi ".
ISA|23|5|Cum auditum fuerit in Aegypto,dolebunt cum audierint de Tyro.
ISA|23|6|Transite ad Tharsis,ululate, qui habitatis in insula.
ISA|23|7|Estne vestra haec, quae gloriabatur?A diebus pristinis antiquitas eius.Ducebant eam pedes sui longead peregrinandum.
ISA|23|8|Quis cogitavit hocsuper Tyrum quondam coronatam,cuius negotiatores principes,institores eius incliti terrae?
ISA|23|9|Dominus exercituum cogitavit hoc,ut detraheret superbiam omnis gloriaeet viles faceret universos inclitos terrae.
ISA|23|10|Excole terram tuam sicut litus Nili,filia Tharsis, iam non est portus.
ISA|23|11|Manum suam extendit super mare,conturbavit regna.Dominus mandavit adversus Chanaan,ut contereret munimenta eius,
ISA|23|12|et dixit: " Non adicies ultra ut glorieris,violata virgo filia Sidonis;in Cetthim consurgens transfreta:ibi quoque non erit requies tibi ".
ISA|23|13|Ecce terra Chaldaeorum:talis populus non fuit;Assyria fundavit eam pro feris.Erexerunt turres suas;suffoderunt domos eius,posuerunt eam in ruinam.
ISA|23|14|Ululate, naves Tharsis,quia devastatum est praesidium vestrum.
ISA|23|15|Et erit in die illa: in oblivione erit Tyrus septuaginta annis, sicut dies regis unius. Post septuaginta autem annos erit Tyro iuxta canticum meretricis:
ISA|23|16|" Sume citharam, circui civitatem,meretrix oblivioni tradita;bene cane, frequenta canticum,ut memoria tui sit ".
ISA|23|17|Et erit: post septuaginta annos visitabit Dominus Tyrum, et redibit ad mercedes suas et rursum fornicabitur cum universis regnis terrae super faciem terrae.
ISA|23|18|Et erunt negotiatio eius et merces eius sanctificatae Domino; non condentur neque reponentur, quia his, qui habitaverint coram Domino, erit negotiatio eius, ut manducent in saturitate et vestiantur splendide.
ISA|24|1|Ecce Dominus dissipat terram et frangit eamet conturbat faciem eiuset dispergit habitatores eius.
ISA|24|2|Et erit sicut populus sic sacerdos,et sicut servus sic dominus eius,sicut ancilla sic domina eius,sicut emens sic ille qui vendit,sicut fenerator sic is qui mutuum accipit,sicut qui repetit sic qui debet.
ISA|24|3|Dissipatione dissipabitur terraet direptione praedabitur:Dominus enim locutus est verbum hoc.
ISA|24|4|Luget, languet terra,marcescit, languet orbis,marcescit altitudo simul cum terra.
ISA|24|5|Et terra infecta est sub habitatoribus suis,quia transgressi sunt leges,violaverunt mandatum,dissipaverunt foedus sempiternum.
ISA|24|6|Propter hoc maledictio voravit terram,et poenas exsolverunt habitatores eius;ideoque imminuti sunt cultores eius,et relicti sunt homines pauci.
ISA|24|7|Luget mustum,emarcuit vitis,ingemiscunt omnes, qui laetabantur corde.
ISA|24|8|Cessavit gaudium tympanorum,quievit sonitus laetantium,cessavit gaudium citharae;
ISA|24|9|cum cantico non bibent vinum,amara erit potio bibentibus illam.
ISA|24|10|Attrita est civitas inanitatis,clausa est omnis domus, ut nemo introeat;
ISA|24|11|clamor est super vino in plateis,occidit omnis laetitia,translatum est gaudium terrae.
ISA|24|12|Relicta est in urbe solitudo,et in ruinam confracta est porta;
ISA|24|13|quia haec erunt in medio terrae,in medio populorum,quomodo si olivae excutiantur,et finita vindemia colligantur racemi.
ISA|24|14|Hi levabunt vocem suam,laudabunt maiestatem Domini,hinnient de mari.
ISA|24|15|Propter hoc in regionibus lucis glorificate Dominum,in insulis maris nomen Domini, Dei Israel.
ISA|24|16|A finibus terrae laudes audivimus: Gloria iusto ".Et dixi: " Secretum meum mihi,secretum meum mihi.Vae mihi! ".Praevaricantes praevaricati suntet praevaricatione praevaricantium praevaricati sunt.
ISA|24|17|Formido et fovea et laqueus super te,habitator terrae.
ISA|24|18|Et erit: qui fugerit a voce formidinis, cadet in foveam;et, qui ascenderit de fovea,tenebitur laqueo,quia cataractae de excelsis apertae sunt,et concussa sunt fundamenta terrae.
ISA|24|19|Confractione confracta est terra,contritione contrita est terra,commotione commota est terra,
ISA|24|20|agitatione agitabitur terra sicut ebriuset fluctuabit quasi tabernaculum;et gravis erit super eam iniquitas eius,et corruet et non adiciet ut resurgat.
ISA|24|21|Et erit in die illa:visitabit Dominus super militiam caeli in excelsoet super reges terrae super terram;
ISA|24|22|et congregabuntur et vincientur in lacuet claudentur in carcere;et post multos dies visitabuntur.
ISA|24|23|Et erubescet luna, et confundetur sol,quia regnavit Dominus exercituum in monte Sion et in Ierusalemet in conspectu senum suorum glorificabitur.
ISA|25|1|Domine, Deus meus es tu;exaltabo te, confitebor no mini tuo,quoniam fecisti mirabilia,cogitationes antiquas, fideles, veraces.
ISA|25|2|Quia posuisti civitatem in tumulum,urbem munitam in ruinam:arx superborum non amplius est civitas,in sempiternum non reaedificabitur.
ISA|25|3|Super hoc glorificabit te populus fortis,civitas gentium robustarum timebit te;
ISA|25|4|quia factus es fortitudo pauperi,fortitudo egeno in tribulatione sua,protectio a turbine,umbraculum ab aestu:spiritus enim robustorumquasi imber hiemalis.
ISA|25|5|Sicut aestus in aridatumultum superborum humiliabis; sicut aestus in umbra nubiscanticum fortium reprimes.
ISA|25|6|Et faciet Dominus exercituumomnibus populis in monte hocconvivium pinguium,convivium vini meri,pinguium medullatorum,vini deliquati.
ISA|25|7|Et praecipitabit in monte istofaciem vinculi colligati super omnes populoset telam, quam orditus est super omnes nationes.
ISA|25|8|Praecipitabit mortem in sempiternumet absterget Dominus Deus lacrimam ab omni facieet opprobrium populi sui auferet de universa terra,quia Dominus locutus est.
ISA|25|9|Et dicetur in die illa: " Ecce Deus noster iste,exspectavimus eum, ut salvaret nos;iste Dominus, sustinuimus eum:exsultabimus et laetabimur in salutari eius.
ISA|25|10|Quia requiescet manus Domini in monte isto ".Et triturabitur Moab in loco suo,sicuti teruntur paleae in sterquilinio;
ISA|25|11|et extendet manus suas in medio eius,sicut extendit natans ad natandum;et humiliabitur superbia eiuscum allisione manuum eius.
ISA|25|12|Et firmum munimentum murorum tuorum evertit,deiecit, prostravit in terram usque ad pulverem.
ISA|26|1|In die illa cantabitur canticum istud in terra Iudae: Urbs fortis nobis in salutem;posuit muros et antemurale.
ISA|26|2|Aperite portas, et ingrediatur gens iusta,quae servat fidem.
ISA|26|3|Propositum eius est firmum;servabis pacem,quia in te speravit.
ISA|26|4|Sperate in Dominum in saeculis aeternis,Dominus est petra aeterna.
ISA|26|5|Quia evertit habitantes in excelso,civitatem sublimem humiliabit;humiliabit eam usque ad terram,detrahet eam usque ad pulverem.
ISA|26|6|Conculcabit eam pes, pedes pauperis,gressus egenorum.
ISA|26|7|Semita iusti recta est;rectum callem iusti complanas.
ISA|26|8|Et in semita iudiciorum tuorum, Domine, speravimus in te;ad nomen tuum et ad memoriale tuum desiderium animae.
ISA|26|9|Anima mea desiderat te in nocte,sed et spiritu meo in praecordiis meis te quaero.Cum resplenduerint iudicia tua in terra,iustitiam discent habitatores orbis.
ISA|26|10|Fit misericordia impio,non discet iustitiam;in terra probitatis inique geritet non videt maiestatem Domini.
ISA|26|11|Domine, exaltata est manus tua, et non vident;videant confusi zelum tuum in populum,et ignis hostium tuorum devorabit eos.
ISA|26|12|Domine, dabis pacem nobis;omnia enim opera nostra operatus es nobis.
ISA|26|13|Domine Deus noster, possederunt nos domini absque te;tantum in te recordemur nominis tui.
ISA|26|14|Mortui non reviviscent,defuncti non resurgent;propterea visitasti et contrivisti eos et perdidisti omnem memoriam eorum.
ISA|26|15|Auxisti gentem, Domine,auxisti gentem, glorificatus es;elongasti omnes terminos terrae.
ISA|26|16|Domine, in angustia quaesierunt te,fuderunt incantationem, castigatio tua in eis.
ISA|26|17|Sicut quae concipit, cum appropinquaverit ad partumdolens clamat in doloribus suis,sic facti sumus a facie tua, Domine.
ISA|26|18|Concepimus et parturivimus,quasi peperimus ventum.Salutes non fecimus in terra,ideo non nati sunt habitatores terrae.
ISA|26|19|Reviviscent mortui tui, interfecti mei resurgent.Expergiscimini et laudate, qui habitatis in pulvere,quia ros lucis ros tuus,et terra defunctos suos edet in lucem.
ISA|26|20|Vade, populus meus, intra in cubicula tua,claude ostia tua super te,abscondere modicum ad momentum,donec pertranseat indignatio.
ISA|26|21|Ecce enim Dominus egredietur de loco suo,ut visitet iniquitatem habitatoris terrae contra eum;et revelabit terra sanguinem suumet non operiet ultra interfectos suos ".
ISA|27|1|In die illa visitabit Dominusin gladio suo duro et forti et grandisuper Leviathan serpentem fugacemet super Leviathan serpentem tortuosumet occidet draconem, qui in mari est.
ISA|27|2|In die illa vinea erit iucunda;cantate ei.
ISA|27|3|Ego Dominus, qui servo eam;per singula momenta irrigabo eam.Ne forte visitetur contra eam,nocte et die servo eam.
ISA|27|4|Indignatio non est mihi.Quis dabit mihi spinam et veprem?In proelio gradiar super eam,succendam eam pariter,
ISA|27|5|nisi forte protectionem meam apprehendat,faciat pacem mecum,pacem faciat mecum.
ISA|27|6|Diebus futuris radices mittet Iacob,florebit et germinabit Israel,et implebunt faciem orbis fructibus.
ISA|27|7|Numquid iuxta plagam percutientis eum percussit eum?Aut, sicut occiduntur occisi eius, occisus est?
ISA|27|8|In mensura punit eum deiciens eum,impellit in spiritu suo duro, tempore quo spirat eurus.
ISA|27|9|Idcirco super hoc dimittetur iniquitas Iacob,et hic erit omnis fructus ablationis peccati eius:ut scilicet ponat omnes lapides altarissicut lapides calcis comminutos,ne exstent luci et thymiateria.
ISA|27|10|Civitas enim munita desolata est,habitaculum derelictum et dimissum quasi desertum;ibi pascetur vitulus et ibi accubabitet consumet arbusta eius.
ISA|27|11|In siccitate frondes illius conterentur;mulieres venient et comburent eas.Ipse enim non est populus sapiens,propterea non miserebitur eius, qui fecit eum,et, qui formavit eum, non parcet ei.
ISA|27|12|Et erit: in die illa percutiet spicas Dominusa Flumine usque ad torrentem Aegypti;et vos congregabiminiunus et unus, filii Israel.
ISA|27|13|Et erit: in die illa clangetur in tuba magna;et venient, qui perditi fuerant de terra Assyriorum,et qui eiecti erant in terra Aegypti,et adorabunt Dominumin monte sancto in Ierusalem.
ISA|28|1|Vae coronae superbiae ebriorum Ephraimet flori decidenti gloriae maiestatis eius,qui erant in vertice vallis pinguissimae,errantes a vino!
ISA|28|2|Ecce validus et fortis Dominosicut impetus grandinis, turbo confringens,sicut impetus aquarum multarum inundantium,et deiciet in terram violenter.
ISA|28|3|Pedibus conculcabiturcorona superbiae ebriorum Ephraim;
ISA|28|4|et erit flos decidens gloriae maiestatis eius,qui est super verticem vallis pinguium,quasi ficus praecox ante messem,quam quis, ut viderit,manu statim arreptam devorabit.
ISA|28|5|In die illa erit Dominus exercituumcorona gloriaeet sertum maiestatisresiduo populi sui
ISA|28|6|et spiritus iudiciisedenti ad iudicandumet fortitudovertentibus proelium usque ad portam.
ISA|28|7|Verum hi quoque prae vino vacillantet prae ebrietate nutant;sacerdos et propheta vacillant prae ebrietate,absorpti sunt a vino,nutant in ebrietate,vacillant in visione,fluctuant in iudicio.
ISA|28|8|Omnes enim mensae repletae sunt vomitu sordiumque,ita ut non esset ultra locus.
ISA|28|9|Quem docebit scientiam?Et quem intellegere faciet auditum?Ablactatos a lacte,avulsos ab uberibus.
ISA|28|10|Etenim praeceptum ad praeceptum, praeceptum ad praeceptum,regula ad regulam, regula ad regulam,modicum ibi, modicum ibi.
ISA|28|11|Balbis enim labiis et lingua alteraloquetur ad populum istum,
ISA|28|12|cui dixerat: " Haec requies, reficite lassum;et hoc est refrigerium ".Et noluerunt audire.
ISA|28|13|Et erit eis verbum Domini: Praeceptum ad praeceptum, praeceptum ad praeceptum,regula ad regulam, regula ad regulam,modicum ibi, modicum ibi ",ut vadant et cadant retrorsum et conteranturet illaqueentur et capiantur.
ISA|28|14|Propter hoc audite verbum Domini,viri illusores, qui dominamini super populum meum,qui est in Ierusalem.
ISA|28|15|Dixistis enim: " Percussimus foedus cum morteet cum inferno fecimus pactum;flagellum inundans cum transierit,non veniet super nos,quia posuimus mendacium spem nostramet in fallacia absconditi sumus ".
ISA|28|16|Idcirco haec dicit Dominus Deus: Ecce ego fundamentum ponam in Sion, lapidem,lapidem probatum, angularem, pretiosum, fundatum;qui crediderit, non turbabitur.
ISA|28|17|Et ponam iudicium tamquam normamet iustitiam tamquam perpendiculum;et subvertet grando spem mendacii,et latibulum aquae inundabunt.
ISA|28|18|Et delebitur foedus vestrum cum morte,et pactum vestrum cum inferno non stabit;flagellum inundans cum transierit,eritis ei in conculcationem.
ISA|28|19|Quandocumque pertransierit, tollet vos;quoniam mane diluculo pertransibit,in die et in nocte,et erit tantummodo horrendum intellegere auditum ".
ISA|28|20|Coangustatum est enim stratum, ut quis se extendat,et pallium brevius, ut quis se operire possit.
ISA|28|21|Sicut enim in monte Pharasim stabit Dominus,sicut in valle, quae est in Gabaon, irascetur,ut faciat opus suum, novum opus suum,ut operetur operationem suam,peregrinam operationem suam.
ISA|28|22|Et nunc nolite illudere,ne forte constringantur vincula vestra;decretum enim destructionis audivia Domino, Deo exercituum,super universam terram.
ISA|28|23|Auribus percipite et audite vocem meam,attendite et audite eloquium meum.
ISA|28|24|Numquid tota die arat arans, ut serat,proscindit et sarrit humum suam?
ISA|28|25|Nonne, cum adaequaverit faciem eius,spargit nigellam et serit cuminum,ponit triticum et hordeumet far in finibus suis?
ISA|28|26|Erudit enim illum recte,Deus suus docet illum.
ISA|28|27|Non enim in serris trituratur nigella,nec rota plaustri super cuminum circuit;sed in virga excutitur nigella,et cuminum in baculo.
ISA|28|28|Numquid comminuitur triticum?Verum non in perpetuum triturans triturabit illum,neque vexabit eum rota plaustri,nec ungulis suis comminuet eum.
ISA|28|29|Et hoc a Domino, Deo exercituum, exivit;mirabile fecit consilium,magnificavit sapientiam.
ISA|29|1|Vae Ariel, Ariel, civitas,quam circumdedit David!Addite annum ad annum,sollemnitates evolvantur;
ISA|29|2|et circumvallabo Ariel,et erit maeror et maestitia,et erit mihi quasi Ariel.
ISA|29|3|Et circumdabo te quasi sphaeramet iaciam contra te aggeremet munimenta ponam in obsidionem tuam.
ISA|29|4|Humiliaberis, de terra loqueris,et de pulvere vix audietur eloquium tuum,et erit quasi pythonis de terra vox tua,et de humo eloquium tuum mussitabit.
ISA|29|5|Et erit sicut pulvis tenuis multitudo superborum tuorum,et sicut palea volans multitudo fortium.Eritque repente confestim,
ISA|29|6|a Domino exercituum visitaberisin tonitruo et commotione terrae,magno fragore, turbine et tempestateet flamma ignis devorantis.
ISA|29|7|Et erit sicut somnium visionis nocturnaemultitudo omnium gentium, quae dimicant contra Ariel,et omnes, qui pugnant contra eam et contra munimenta eius et oppressores eius;
ISA|29|8|Et sicut somniat esuriens, et ecce comedit,cum autem fuerit expergefactus, vacua est anima eius;et sicut somniat sitiens, et ecce bibitet, postquam fuerit expergefactus, lassus adhuc sitit,et anima eius vacua est,sic erit multitudo omnium gentiumdimicantium contra montem Sion.
ISA|29|9|Obstupescite et admiramini,excaecamini et caeci estote,inebriamini et non a vino,vacillate et non ab ebrietate.
ISA|29|10|Quoniam miscuit vobis Dominus spiritum soporis,clausit oculos vestroset capita vestra operuit.
ISA|29|11|Et erit vobis visio omnis sicut verba libri signati; quem cum dederint scienti litteras dicentes: " Lege istum ", respondebit: " Non possum, signatus est enim ".
ISA|29|12|Et dabitur liber nescienti litteras diceturque ei: " Lege ", et respondebit: " Nescio litteras ".
ISA|29|13|Et dixit Dominus: Eo quod appropinquat populus iste ore suoet labiis suis glorificat me,cor autem eius longe est a me,et est timor eorum erga mevelut mandatum hominum perceptum,
ISA|29|14|ideo ecce ego addam ut admirationem faciampopulo huic miraculo grandi et stupendo:peribit sapientia sapientium eius,et prudentia prudentium eius abscondetur ".
ISA|29|15|Vae, qui profunde a Dominoconsilium abscondunt,quorum sunt in tenebris opera, et dicunt: Quis videt nos, et quis novit nos? ".
ISA|29|16|Perversa cogitatio vestra!Numquid quasi lutum reputabitur figulus,ut dicat opus factori suo: Non fecisti me ";et figmentum dicat fictori suo: Non intellegis "?
ISA|29|17|Nonne adhuc in modico et in brevi convertetur Libanus in hortum,et hortus in saltum reputabitur?
ISA|29|18|Et audient in die illa surdi verba libri,et de tenebris et caligine oculi caecorum videbunt.
ISA|29|19|Et addent mites in Domino laetitiam,et pauperrimi hominum in Sancto Israel exsultabunt;
ISA|29|20|quoniam defecit, qui praevalebat,consummatus est illusor,et succisi sunt omnes, qui vigilabant super iniquitatem,
ISA|29|21|qui peccare faciebant homines in verboet arguentem in porta supplantabantet deiecerunt inanibus verbis iustum.
ISA|29|22|Propter hoc haec dicit Dominusad domum Iacob, qui redemit Abraham: Non modo confundetur Iacob,nec modo vultus eius erubescet;
ISA|29|23|sed, cum viderit opera manuum mearum,in medio sui sanctificabunt nomen meumet sanctificabunt Sanctum Iacobet Deum Israel pavebunt,
ISA|29|24|et scient errantes spiritu sapientiam,et mussitatores discent doctrinam ".
ISA|30|1|" Vae, filii desertores, dicit Dominus,eo quod facitis consilium et non ex me,et pactum statuitis et non per spiritum meum,ut addatis peccatum super peccatum!
ISA|30|2|Qui ambulatis, ut descendatis in Aegyptum,et os meum non interrogastis,sperantes auxilium in fortitudine pharaoniset habentes fiduciam in umbra Aegypti.
ISA|30|3|Et erit vobis fortitudo pharaonis in confusionem,et fiducia sub umbra Aegypti in ignominiam.
ISA|30|4|Cum fuerint enim in Tani principes tui,et nuntii tui usque ad Hanes pervenerint,
ISA|30|5|omnes confundentursuper populo, qui eis prodesse non potest;non erit in auxilium et in utilitatem sed in confusionem et opprobrium ".
ISA|30|6|Oraculum iumentorum Nageb.In terra tribulationis et angustiae,leaenae et leonis rugientis,viperae et draconis volantisportant super umeros iumentorum divitias suaset super gibbum camelorum thesauros suosad populum, qui eis prodesse non poterit.
ISA|30|7|Aegyptus enim frustra et vane auxiliabitur;ideo vocavi Rahab otiosam.
ISA|30|8|Nunc ingredere, scribe coram eis super buxumet in libro diligenter exara illud,et erit in posterumin testimonium usque in aeternum.
ISA|30|9|Populus enim rebellis est,et filii mendaces,filii nolentes audire legem Domini;
ISA|30|10|qui dicunt videntibus: " Nolite videre "et aspicientibus: " Nolite aspicere nobis ea, quae recta sunt;loquimini nobis placentia, aspicite nobis illusiones.
ISA|30|11|Recedite a via, declinate a semita,tollite a facie nostra Sanctum Israel ".
ISA|30|12|Propterea haec dicit Sanctus Israel: Pro eo quod reprobastis verbum hocet sperastis in perversitatem et in perfidiamet innixi estis super eis,
ISA|30|13|propterea erit vobis iniquitas haecsicut interruptio cadens, locus tumens in muro excelso,cuius confractio subito, dum non speratur,venit improviso;
ISA|30|14|et comminuetur, sicut conteritur lagoena figuli,contritione absque misericordia,et non invenietur de fragmentis eius testa,in qua capiatur igniculus de incendio,aut hauriatur aqua de fovea ".
ISA|30|15|Quia haec dixit Dominus Deus, Sanctus Israel: In conversione et quiete salvi eritis;in silentio et in spe erit fortitudo vestra ".Et noluistis
ISA|30|16|et dixistis: Nequaquam, sed super equis fugiemus ",ideo fugietis;et: " Super veloces ascendemus ",ideo veloces erunt, qui persequentur vos.
ISA|30|17|Mille pavebunt a facie terroris unius,et a facie terroris quinque fugietis,donec relinquaminiquasi malus in vertice montiset quasi signum super collem.
ISA|30|18|Propterea exspectat Dominus, ut misereatur vestri,et ideo exaltabitur parcens vobis,quia Deus iudicii Dominus;beati omnes, qui exspectant eum.
ISA|30|19|Nam, popule Sion, qui habitas in Ierusalem,plorans nequaquam plorabis:miserans miserebitur tui ad vocem clamoris tui;statim ut audierit, respondebit tibi.
ISA|30|20|Et dabit vobis Dominuspanem angustiae et aquam afflictionis,sed non amplius avolabit a te doctor tuus;et erunt oculi tui videntes praeceptorem tuum,
ISA|30|21|et aures tuae audient verbum post tergum monentis: Haec via, ambulate in ea ",si declinaveritis ad dexteram vel ad sinistram.
ISA|30|22|Et contaminabis laminas sculptilium argentorum tuorumet vestimentum conflatilis aurei tui;disperges ea sicut immunditiam menstruatae. Egredere " dices ei.
ISA|30|23|Et dabit pluviam semini tuo,quod seminaveris in terra,et panis frugum terrae erit uberrimus et pinguis;pascetur pecus tuum in die illo, agnus in pascuis spatiosis,
ISA|30|24|et boves tui et asini, qui operantur terram,commixtum migma comedentventilatum in pala et ventilabro.
ISA|30|25|Et erunt super omnem montem excelsumet super omnem collem elevatumrivi currentium aquarumin die interfectionis multorum,cum ceciderint turres.
ISA|30|26|Et erit lux lunae sicut lux solis,et lux solis erit septempliciter sicut lux septem dierumin die, qua alligaverit Dominus vulnus populi suiet percussuram plagae eius sanaverit.
ISA|30|27|Ecce nomen Domini venit de longinquo,ardens furor eius, et gravis eius fragor;labia eius repleta sunt indignatione,et lingua eius quasi ignis devorans.
ISA|30|28|Spiritus eius velut torrens inundans,usque ad collum pertingens,ad cribrandas gentes in cribro funesto,et frenum dolosum in maxillis populorum.
ISA|30|29|Canticum erit vobissicut nox sanctificatae sollemnitatis,et laetitia cordissicut eius, qui ad sonum tibiae pergitin montem Domini,ad petram Israel.
ISA|30|30|Et auditam faciet Dominusgloriam vocis suaeet terrorem brachii suiostendet in comminatione furoriset flamma ignis devorantis,in turbine et in imbre et in lapide grandinis.
ISA|30|31|A voce enim Domini pavebitAssyrius virga percussus.
ISA|30|32|Et erit omnis ictus baculi percutientis,quem requiescere faciet Dominussuper eum in tympanis et citharis,et in bellis agitatis expugnabit eos.
ISA|30|33|Praeparata est enim ab heri Topheth,praeparata, profunda et dilatata,in pyra eius ignis et ligna multa;flatus Domini sicut torrens sulphurissuccendit eam.
ISA|31|1|Vae, qui descendunt in Aegyptum ad auxilium,in equis speranteset habentes fiduciam super quadrigis, quia multae sunt,et super equitibus, quia praevalidi nimis,et non intendunt in Sanctum Israelet Dominum non requirunt!
ISA|31|2|Tamen et ipse sapiens adducit malumet verba sua non retractat;et consurget contra domum pessimorumet contra auxilium operantium iniquitatem.
ISA|31|3|Aegyptius homo et non Deus,et equi eorum caro et non spiritus;et Dominus inclinabit manum suam,et corruet auxiliator,et cadet, cui praestatur auxilium,simulque omnes consumentur.
ISA|31|4|Quia haec dicit Dominus ad me: Quomodo si rugit leo et catulus leonis super praedam suam,cum occurrerit ei multitudo pastorum,a voce eorum non formidabit et a multitudine eorum non pavebit,sic descendet Dominus exercituum, ut proelietur super montem Sion et super collem eius.
ISA|31|5|Sicut aves volantes,sic proteget Dominus exercituum Ierusalem,protegens et liberans,parcens et salvans ".
ISA|31|6|Convertimini ad eum, a quo penitus recesseratis,filii Israel.
ISA|31|7|In die enim illa abiciet viridola argentea sua et idola aurea sua,quae fecerunt vobis manus vestrae in peccatum;
ISA|31|8|et cadet Assyria in gladio non viri,et gladius non hominis vorabit eum,et fugiet a facie gladii,et iuvenes eius vectigales erunt.
ISA|31|9|Et fortitudo eius prae terrore transibit,et pavebunt signum principes eius,dixit Dominus, cuius ignis est in Sion,et caminus eius in Ierusalem.
ISA|32|1|Ecce in iustitia regnabit rex,et principes in iudicio praee runt.
ISA|32|2|Et erit vir sicut latibulum a ventoet refugium a tempestate,sicut rivi aquarum in sitiente terraet umbra petrae magnae in terra arida.
ISA|32|3|Non caligabunt oculi videntium,et aures audientium diligenter auscultabunt,
ISA|32|4|et cor stultorum intelleget scientiam,et lingua balborum velociter loquetur et plane.
ISA|32|5|Non vocabitur ultra is, qui insipiens est, nobilis,neque fraudulentus appellabitur maior;
ISA|32|6|stultus enim fatua loquitur,et cor eius cogitat iniquitatem,ut perficiat impietatemet loquatur contra Dominum erroreset vacuam faciat animam esurientemet potum sitienti auferat.
ISA|32|7|Fraudulenti fraudes pessimae sunt;ipse enim cogitationes concinnatad perdendos mites in sermone mendaci,etiam quando pauper iudicium vindicat.
ISA|32|8|Nobilis vero consilia nobilia datet ipse ad nobilia assurget.
ISA|32|9|Mulieres vanae, surgite, audite vocem meam;filiae confidentes, percipite auribus eloquium meum.
ISA|32|10|Post dies enim et annumvos pavebitis confidentes;consummata est enim vindemia,collectio ultra non veniet.
ISA|32|11|Obstupescite, vanae;pavete, confidentes,exuite vos et nudate vos,accingite lumbos vestros.
ISA|32|12|Super ubera plangite,super regione desiderabili,super vinea fertili.
ISA|32|13|Super humum populi meispinae et vepres ascendent,super omnes domos gaudii,super civitatem exsultantem.
ISA|32|14|Domus enim dimissa est;multitudo urbis relicta est,Ophel et Bahan erunt speluncaeusque in aeternum,gaudium onagrorum,pascua gregum,
ISA|32|15|donec effundatur super nosspiritus de excelso.Et erit desertum in hortum,et hortus in saltum reputabitur,
ISA|32|16|et habitabit in solitudine iudicium,et iustitia in horto sedebit;
ISA|32|17|et erit opus iustitiae pax,et cultus iustitiae silentium,et securitas usque in sempiternum.
ISA|32|18|Et sedebit populus meus in habitatione paciset in tabernaculis fiduciaeet in locis securis.
ISA|32|19|Et penitus cadet saltus,et profunde deprimetur civitas.
ISA|32|20|Beati, qui seminatis super omnes aquas,immittentes pedem bovis et asini.
ISA|33|1|Vae, qui praedaris, cum nemo te praedatus sit;qui devastas, cum nemo te devastaverit!Cum consummaveris depraedationem, depraedaberis;cum perfeceris devastationem, te devastabunt.
ISA|33|2|Domine, miserere nostri,te enim exspectavimus;esto brachium nostrum in maneet salus nostra in tempore tribulationis.
ISA|33|3|A voce fragoris fugerunt populi,ab exaltatione tua dispersae sunt gentes.
ISA|33|4|Et congregabuntur spolia, sicut colligitur bruchus;sicut discurrunt locustae, ad ea discurritur.
ISA|33|5|Sublimis est Dominus, quoniam habitat in excelso;implet Sion iudicio et iustitia.
ISA|33|6|Et erit firmitas in temporibus tuis;divitiae salutis sapientia et scientia:timor Domini ipse est thesaurus eius.
ISA|33|7|Ecce praecones clamabunt foris,angeli pacis amare flebunt.
ISA|33|8|Dissipatae sunt viae, cessavit transiens per semitam;irritum fecit pactum,reiecit testes,non reputavit homines.
ISA|33|9|Luget et elanguescit terra,confusus est Libanus et obsorduit,et factus est Saron sicut desertum,et exaruerunt Basan et Carmelus.
ISA|33|10|" Nunc consurgam, dicit Dominus,nunc exaltabor, nunc sublevabor.
ISA|33|11|Concipietis fenum, parietis stipulam;spiritus meus ut ignis vorabit vos.
ISA|33|12|Et erunt populi fornaces calcis:spinae congregatae igne comburentur.
ISA|33|13|Audite, qui longe estis, quae fecerim,et cognoscite, vicini, fortitudinem meam ".
ISA|33|14|Conterriti sunt in Sion peccatores,possedit tremor impios.Quis poterit habitare de vobis cum igne devorante?Quis habitabit ex vobis cum ardoribus sempiternis?
ISA|33|15|Qui ambulat in iustitiis et loquitur aequitates,qui reicit lucra ex rapiniset excutit manus suas, ne munera accipiat,qui obturat aures suas, ne audiat sanguinem,et claudit oculos suos, ne videat malum:
ISA|33|16|iste in excelsis habitabit,munimenta saxorum refugium eius;panis ei datus est, aquae eius fideles sunt.
ISA|33|17|Regem in decore suo videbunt oculi tui,cernent terram longinquam.
ISA|33|18|Cor tuum cum timore inquiret: Ubi est scriba? Ubi ponderator?Ubi computator turrium? ".
ISA|33|19|Populum impudentem non videbis,populum profundi sermonis, ininterpretabilis,linguae barbarae absque intellegentia.
ISA|33|20|Respice Sion civitatem sollemnitatum nostrarum!Oculi tui videbunt Ierusalem,habitationem securam,tabernaculum quod nequaquam transferri poterit;nec auferentur clavi eius in sempiternum,et omnes funiculi eius non rumpentur.
ISA|33|21|Quia ibi potens Dominus pro nobisloco fluviorum, rivorum late patentium;non transibit ibi navis remigum,neque navis magna transgredietur eum.
ISA|33|22|Dominus enim iudex noster, Dominus legifer noster,Dominus rex noster: ipse salvabit nos.
ISA|33|23|Laxati sunt funiculi tuinec sustinent malum suum,ut dilatare velum non queant.Tunc divident caeci praedam multam;claudi diripient rapinam.
ISA|33|24|Nec dicet incola: " Elangui ".Populus, qui habitat in ea,auferetur ab eo iniquitas.
ISA|34|1|Accedite, gentes, ad audien dum;et populi, attendite.Audiat terra et plenitudo eius,orbis et omne germen eius.
ISA|34|2|Quia indignatio Domini super omnes gentes,et furor super universam militiam eorum:ad interitum devovit eos et dedit eos in occisionem.
ISA|34|3|Interfecti eorum proicientur,et de cadaveribus eorum ascendet foetor;dissolventur montes sanguine eorum.
ISA|34|4|Et tabescet omnis militia caelorum,et complicabuntur sicut liber caeli, et omnis militia eorum defluet,sicut defluit folium de vinea et arida frons de ficu.
ISA|34|5|Quoniam inebriatus est in caelo gladius meus:ecce super Edom descendetet super populum interfectionis meae ad iudicium.
ISA|34|6|Gladius Domini repletus est sanguine,incrassatus est adipe,de sanguine agnorum et hircorum, de adipe viscerum arietum;victima enim Domini in Bosra,et interfectio magna in terra Edom.
ISA|34|7|Cadunt bubali cum eis,iuvenci cum tauris;inebriabitur terra eorum sanguine,et humus eorum adipe pinguium,
ISA|34|8|quia dies ultionis Domini,annus retributionum ad vindicandam Sion.
ISA|34|9|Et convertentur torrentes eius in picem,et humus eius in sulphur,et erit terra eius in picem ardentem.
ISA|34|10|Nocte et die non exstinguetur,in sempiternum ascendet fumus eius,a generatione in generationem desolabitur,in saecula saeculorum non erit transiens per eam.
ISA|34|11|Et possidebunt illam onocrotalus et ericius,noctua et corvus habitabunt in ea;et extendet super eam mensuram solitudiniset perpendiculum desolationis.
ISA|34|12|Nobiles eius non erunt,nec regnum proclamabunt;et omnes principes eius erunt in nihilum.
ISA|34|13|Et orientur in domibus eius spinae,urticae et paliurus in munitionibus eius;et erit cubile draconumet pascua struthionum.
ISA|34|14|Et occurrent hyaenae thoibus,et pilosus clamat ad amicum suum;ibi cubat lamiaet invenit sibi requiem.
ISA|34|15|Ibi nidificat serpens ovaque deponitet circumfodit et fovet in umbra eius;illuc congregantur milvi alter ad alterum.
ISA|34|16|Requirite in libro Domini et legite:unum ex eis non deest,alter alterum exspectare non debet;quia os Domini praecepit,et spiritus eius ipse congregavit ea.
ISA|34|17|Et ipse misit eis sortem,et manus eius divisit terram illis in mensura;usque in aeternum possidebunt eam,in generatione et generatione habitabunt in ea.
ISA|35|1|Laetentur deserta et invia,et exsultet solitudo et floreat quasi lilium.
ISA|35|2|Germinet et exsultetlaetabunda et laudans.Gloria Libani data est ei,decor Carmeli et Saron;ipsi videbunt gloriam Domini,maiestatem Dei nostri.
ISA|35|3|Confortate manus dissolutaset genua debilia roborate.
ISA|35|4|Dicite pusillanimis: Confortamini, nolite timere!Ecce Deus vester,ultio veniet, retributio Dei;ipse veniet et salvabit vos ".
ISA|35|5|Tunc aperientur oculi caecorum,et aures surdorum patebunt.
ISA|35|6|Tunc saliet sicut cervus claudus,et exsultabit lingua mutorum,quia erumpent in deserto aquae,et torrentes in solitudine.
ISA|35|7|Et terra arida erit in stagnum,et sitiens in fontes aquarum;in cubilibus, in quibus dracones habitabant,erit locus calami et iunci.
ISA|35|8|Et erit ibi semita et via;et via sancta vocabitur:non transibit per eam pollutus;et erit eis directa via,ita ut stulti non errent per eam.
ISA|35|9|Non erit ibi leo,et rapax bestia non ascendet per eamnec invenietur ibi;et ambulabunt, qui liberati fuerint,
ISA|35|10|et redempti a Domino revertentur.Et venient in Sion cum laude,et laetitia sempiterna super caput eorum:gaudium et laetitiam obtinebunt,et fugiet maeror et gemitus.
ISA|36|1|Et factum est in quarto deci mo anno regis Ezechiae, ascendit Sennacherib rex Assyriorum super omnes civitates Iudae munitas et cepit eas.
ISA|36|2|Et misit rex Assyriorum Rabsacen de Lachis in Ierusalem ad regem Ezechiam in manu gravi, et stetit in aquaeductu piscinae superioris in via agri fullonis.
ISA|36|3|Et egressus est ad eum Eliachim filius Helciae, qui erat super domum, et Sobna scriba et Ioah filius Asaph a commentariis.
ISA|36|4|Et dixit ad eos Rabsaces: " Dicite Ezechiae: Haec dicit rex magnus, rex Assyriorum: Quae est ista fiducia, qua confidis?
ISA|36|5|Dixisti: " Verbum labiorum est consilium et fortitudo ad bellum". Nunc super quem habes fiduciam, quia recessisti a me?
ISA|36|6|Ecce confidis super baculum arundineum confractum istum, super Aegyptum; cui si innixus fuerit homo, intrabit in manum eius et perforabit eam: sic pharao rex Aegypti omnibus, qui confidunt in eo.
ISA|36|7|Quod si responderis mihi: "In Domino Deo nostro confidimus"; nonne ipse est, cuius abstulit Ezechias excelsa et altaria et dixit Iudae et Ierusalem: "Coram altari isto adorabitis"?
ISA|36|8|Et nunc sponde domino meo regi Assyriorum, et dabo tibi duo milia equorum, si poteris ex te praebere ascensores eorum.
ISA|36|9|Et quomodo averteris faciem unius ex servis domini mei minoribus? Et tamen confidis in Aegypto, in quadriga et in equitibus;
ISA|36|10|et nunc, numquid sine Domino ascendi ad terram istam, ut disperderem eam? Dominus dixit ad me: "Ascende super terram istam et disperde eam" ".
ISA|36|11|Et dixit Eliachim et Sobna et Ioah ad Rabsacen: "Loquere ad servos tuos Aramaice; intellegimus enim. Ne loquaris ad nos Iudaice in auribus populi, qui est super murum ".
ISA|36|12|Et dixit Rabsaces: " Numquid ad dominum tuum et ad te misit me dominus meus, ut loquerer omnia verba ista? Et non potius ad viros, qui sedent in muro, ut comedant stercora sua et bibant urinam suam vobiscum? ".
ISA|36|13|Et stetit Rabsaces et clamavit voce magna Iudaice et dixit: " Audite verba regis magni, regis Assyriorum:
ISA|36|14|Haec dicit rex: Non seducat vos Ezechias, quia non poterit eruere vos.
ISA|36|15|Et non vobis tribuat fiduciam Ezechias super Domino dicens: "Eruens liberabit nos Dominus; non dabitur civitas ista in manu regis Assyriorum".
ISA|36|16|Nolite audire Ezechiam. Haec enim dicit rex Assyriorum: Facite mecum benedictionem et egredimini ad me; et comedite unusquisque vineam suam et unusquisque ficum suam, et bibite unusquisque aquam de cisterna sua,
ISA|36|17|donec veniam et tollam vos ad terram, quae est ut terra vestra, terram frumenti et vini, terram panis et vinearum.
ISA|36|18|Ne illudat vos Ezechias dicens: "Dominus liberabit nos". Numquid liberaverunt dii gentium unusquisque terram suam de manu regis Assyriorum?
ISA|36|19|Ubi sunt dii Emath et Arphad? Ubi sunt dii Sepharvaim? Numquid liberaverunt Samariam de manu mea?
ISA|36|20|Quinam ex omnibus diis terrarum istarum eruerunt terram suam de manu mea? Numquid eruet Dominus Ierusalem de manu mea? ".
ISA|36|21|Et siluerunt et non responderunt ei verbum; mandaverat enim rex dicens: Ne respondeatis ei ".
ISA|36|22|Et ingressus est Eliachim filius Helciae, qui erat super domum, et Sobna scriba et Ioah filius Asaph a commentariis ad Ezechiam scissis vestibus; et nuntiaverunt ei verba Rabsacis.
ISA|37|1|Et factum est cum audisset rex Ezechias, scidit vestimen ta sua et obvolutus est sacco et intravit in domum Domini;
ISA|37|2|et misit Eliachim, qui erat super domum, et Sobnam scribam et seniores de sacerdotibus opertos saccis ad Isaiam filium Amos prophetam,
ISA|37|3|et dixerunt ad eum: " Haec dicit Ezechias: Dies tribulationis et correptionis et contumeliae dies haec, quia venerunt filii usque ad partum, et virtus non est pariendi.
ISA|37|4|Forsitan audiet Dominus Deus tuus verba Rabsacis, quem misit rex Assyriorum, dominus suus, ad blasphemandum Deum viventem, et puniet sermones, quos audivit Dominus Deus tuus; leva ergo orationem pro reliquiis, quae repertae sunt ".
ISA|37|5|Et venerunt servi regis Ezechiae ad Isaiam;
ISA|37|6|et dixit ad eos Isaias: "Haec dicetis domino vestro: Haec dicit Dominus: Ne timeas a facie verborum, quae audisti, quibus blasphemaverunt pueri regis Assyriorum me.
ISA|37|7|Ecce ego dabo ei spiritum, et audiet nuntium et revertetur ad terram suam, et corruere eum faciam gladio in terra sua ".
ISA|37|8|Reversus est autem Rabsaces et invenit regem Assyriorum proeliantem adversus Lobnam; audierat enim quia profectus esset de Lachis.
ISA|37|9|Et audivit de Tharaca rege Aethiopiae dicentes: " Egressus est, ut pugnet contra te ".Quod cum audisset, misit nuntios ad Ezechiam dicens:
ISA|37|10|" Haec dicetis Ezechiae regi Iudae loquentes: Non te decipiat Deus tuus, in quo tu confidis, dicens: "Non dabitur Ierusalem in manu regis Assyriorum".
ISA|37|11|Ecce tu audisti omnia, quae fecerunt reges Assyriorum omnibus terris, quas ad interitum devoverunt, et tu poteris liberari?
ISA|37|12|Numquid eruerunt eos dii gentium, quos subverterunt patres mei, Gozan et Charran et Reseph et filios Eden, qui erant in Thelassar?
ISA|37|13|Ubi est rex Emath et rex Arphad et rex urbis Sepharvaim, Ana et Ava? ".
ISA|37|14|Et tulit Ezechias epistulam de manu nuntiorum et legit eam. Et ascendit in domum Domini et expandit eam Ezechias coram Domino.
ISA|37|15|Et oravit Ezechias ad Dominum dicens:
ISA|37|16|" Domine exercituum, Deus Israel, qui sedes super cherubim, tu es Deus solus omnium regnorum terrae, tu fecisti caelum et terram.
ISA|37|17|Inclina, Domine, aurem tuam et audi; aperi, Domine, oculos tuos et vide et audi omnia verba Sennacherib, quae misit ad blasphemandum Deum viventem.
ISA|37|18|Vere enim, Domine, dissipaverunt reges Assyriorum gentes et regiones earum
ISA|37|19|et dederunt deos earum igni: non enim erant dii, sed opera manuum hominum, lignum et lapis; et comminuerunt eos.
ISA|37|20|Et nunc, Domine Deus noster, salva nos de manu eius; et cognoscant omnia regna terrae quia tu, Domine, es solus Deus ".
ISA|37|21|Et misit Isaias filius Amos ad Ezechiam dicens: " Haec dicit Dominus, Deus Israel: Pro quibus rogasti me de Sennacherib rege Assyriorum,
ISA|37|22|hoc est verbum, quod locutus est Dominus super eum:Despexit te, subsannavit te virgo filia Sion;post te caput movit filia Ierusalem.
ISA|37|23|Cui exprobrasti et quem blasphemasti?Et super quem exaltasti vocemet levasti altitudinem oculorum tuorum?Contra Sanctum Israel!
ISA|37|24|In manu servorum tuorum exprobrasti Dominoet dixisti: "In multitudine quadrigarum mearumego ascendi altitudinem montium, iuga Libani;et succidi excelsa cedrorum eiuset electas abietes illiuset introivi altitudinem summitatis eius,silvam condensam.
ISA|37|25|Ego fodi et bibi aquam alienamet exsiccavi vestigio pedis meiomnes rivos Aegypti".
ISA|37|26|Numquid non audisti?A saeculo feci illud; a diebus antiquisego plasmavi illud et nunc adduxi,ut fiat in eradicationem,in lapides eversos civitates munitae.
ISA|37|27|Habitatores earum breviata manucontremuerunt et confusi sunt;facti sunt sicut fenum agriet gramen viride et herba tectorum, quae exaruit a facie austri.
ISA|37|28|Sessionem tuamet egressum tuum et introitum tuum cognoviet insaniam tuam contra me.
ISA|37|29|Cum fureris adversum me,et superbia tua ascenderit in aures meas,ponam circulum in naribus tuiset frenum in labiis tuiset reducam te in viam,per quam venisti.
ISA|37|30|Tibi autem hoc erit signum:Comedantur hoc anno, quae colligi poterunt,et in anno secundo, quae sponte nascuntur;in anno autem tertio seminate et metiteet plantate vineas et comedite fructum earum.
ISA|37|31|Et mittet id, quod salvatum fuerit de domo Iudae,quod reliquum est, radicem deorsumet faciet fructum sursum.
ISA|37|32|Quia de Ierusalem exibit residuum,et, quod salvum fuerit, de monte Sion.Zelus Domini exercituum faciet istud.
ISA|37|33|Propterea haec dicit Dominus de rege Assyriorum:Non introibit civitatem hancet non iaciet ibi sagittamet non opponet ei clipeumet non mittet contra eam aggerem.
ISA|37|34|In via, qua venit, per eam revertetur,et civitatem hanc non ingredietur, dicit Dominus.
ISA|37|35|Et protegam civitatem istam, ut salvem eampropter me et propter David servum meum ".
ISA|37|36|Egressus est autem angelus Domini et percussit in castris Assyriorum centum octoginta quinque milia; et surrexerunt mane, et ecce omnes illi cadavera mortuorum.
ISA|37|37|Et egressus est et abiit; et reversus est Sennacherib rex Assyriorum et habitavit in Nineve.
ISA|37|38|Et factum est, cum adoraret in templo Nesroch dei sui, Adramelech et Sarasar filii eius percusserunt eum gladio fugeruntque in terram Ararat. Et regnavit Asarhaddon filius eius pro eo.
ISA|38|1|In diebus illis aegrotavit Ezechias usque ad mortem. Et introivit ad eum Isaias filius Amos propheta et dixit ei: " Haec dicit Dominus: Dispone domui tuae, quia morieris tu et non vives".
ISA|38|2|Et convertit Ezechias faciem suam ad parietem et oravit ad Dominum
ISA|38|3|et dixit: " Obsecro, Domine; memento, quaeso, quomodo ambulaverim coram te in veritate et in corde perfecto et, quod bonum est in oculis tuis, fecerim ". Et flevit Ezechias fletu magno.
ISA|38|4|Et factum est verbum Domini ad Isaiam dicens:
ISA|38|5|" Vade et dic Ezechiae: "Haec dicit Dominus, Deus David patris tui: Audivi orationem tuam, vidi lacrimas tuas; ecce ego adiciam super dies tuos quindecim annos
ISA|38|6|et de manu regis Assyriorum eruam te et civitatem istam et protegam hanc civitatem".
ISA|38|7|Hoc autem tibi erit signum a Domino quia faciet Dominus verbum hoc, quod locutus est:
ISA|38|8|Ecce ego reverti faciam umbram graduum, per quos descenderat in horologio Achaz in sole retrorsum decem gradibus ". Et reversus est sol decem gradibus per gradus, quos descenderat.
ISA|38|9|Scriptura Ezechiae regis Iudae, cum aegrotasset et convaluisset de infirmitate sua:
ISA|38|10|" Ego dixi: In dimidio dierum meorumvadam ad portas inferi;quaesivi residuum annorum meorum.
ISA|38|11|Dixi: Non videbo Dominum Deum in terra viventium,non aspiciam hominem ultrainter habitatores orbis.
ISA|38|12|Habitaculum meum ablatum est et abductum longe a mequasi tabernaculum pastorum;convolvit sicut textor vitam meam;de stamine succidit me.De mane usque ad vesperam confecisti me.
ISA|38|13|Prostratus sum usque ad mane,quasi leo sic conterit omnia ossa mea;de mane usque ad vesperam confecisti me.
ISA|38|14|Sicut pullus hirundinis, sic mussitabo,meditabor ut columba;attenuati sunt oculi meisuspicientes in excelsum.Domine, vim patior,sponde pro me.
ISA|38|15|Quid dicam, aut quid respondebit mihi?Ipse fecit!Incedam per omnes annos meosin amaritudine animae meae.
ISA|38|16|Domine, in te sperat cor meum;vivat spiritus meus,sana me et vivifica me;
ISA|38|17|ecce in pacem versa est amaritudo mea.Tu autem eruisti animam meama fovea consumptionis,proiecisti enim post tergum tuumomnia peccata mea.
ISA|38|18|Quia non infernus confitebitur tibi,neque mors laudabit te;non exspectabunt, qui descendunt in lacum,veritatem tuam.
ISA|38|19|Vivens, vivens ipse confitebitur tibi,sicut et ego hodie;pater filiis notam faciet veritatem tuam.
ISA|38|20|Domine, salvum me fac,et ad sonum citharae cantabimuscunctis diebus vitae nostraein domo Domini ".
ISA|38|21|Et iussit Isaias, ut tollerent massam de ficis et cataplasmarent super vulnus, et sanaretur.
ISA|38|22|Et dixit Ezechias: " Quod erit signum quia ascendam in domum Domini?".
ISA|39|1|In tempore illo misit Merodachbaladan filius Baladan rex Babylonis litteras et munera ad Ezechiam; audierat enim quod aegrotasset et convaluisset.
ISA|39|2|Laetatus est autem super eis Ezechias et ostendit eis cellam thesauri sui et argentum et aurum et aromata et oleum optimum et omnes apothecas supellectilis suae et universa, quae inventa sunt in thesauris eius. Nihil fuit, quod non ostenderet eis Ezechias in domo sua et in omni potestate sua.
ISA|39|3|Introivit autem Isaias propheta ad Ezechiam regem et dixit ei: " Quid dixerunt viri isti et unde venerunt ad te? ". Et dixit Ezechias: " De terra longinqua venerunt ad me, de Babylone ".
ISA|39|4|Et dixit: "Quid viderunt in domo tua?". Et dixit Ezechias: " Omnia, quae in domo mea sunt, viderunt; non fuit res, quam non ostenderim eis in thesauris meis ".
ISA|39|5|Et dixit Isaias ad Ezechiam: " Audi verbum Domini exercituum:
ISA|39|6|Ecce dies venient, et auferentur omnia, quae in domo tua sunt, et quae thesaurizaverunt patres tui usque ad diem hanc, in Babylonem; non relinquetur quidquam, dicit Dominus.
ISA|39|7|Et de filiis tuis, qui exibunt de te, quos genueris, tollent, et erunt eunuchi in palatio regis Babylonis ".
ISA|39|8|Et dixit Ezechias ad Isaiam: " Bonum verbum Domini, quod locutus est ". Et dixit: " Dummodo fiat pax et securitas in diebus meis ".
ISA|40|1|Consolamini, consolamini populum meum,dicit Deus vester.
ISA|40|2|Loquimini ad cor Ierusalemet clamate ad eam,quoniam completa est militia eius,expiata est iniquitas illius;suscepit de manu Dominiduplicia pro omnibus peccatis suis.
ISA|40|3|Vox clamantis: In deserto parate viam Domini,rectas facite in solitudinesemitas Dei nostri.
ISA|40|4|Omnis vallis exaltetur,et omnis mons et collis humilietur;et fiant prava in directa,et aspera in plana:
ISA|40|5|et revelabitur gloria Domini,et videbit omnis caro pariterquod os Domini locutum est ".
ISA|40|6|Vox dicentis: " Clama! ".Et dixi: " Quid clamabo? ".Omnis caro fenum,et omnis gloria eius quasi flos agri;
ISA|40|7|exsiccatum est fenum, et cecidit flos,quia spiritus Domini sufflavit in eo. Vere fenum est populus.
ISA|40|8|Exsiccatum est fenum, et cecidit flos;verbum autem Dei nostri manet in aeternum.
ISA|40|9|Super montem excelsum ascende,tu, quae evangelizas Sion;exalta in fortitudine vocem tuam,quae evangelizas Ierusalem;exalta, noli timere;dic civitatibus Iudae: Ecce Deus vester,
ISA|40|10|ecce Dominus Deus in virtute venit,et brachium eius dominatur:ecce merces eius cum eo,et praemium illius coram illo.
ISA|40|11|Sicut pastor gregem suum pascit,in brachio suo congregat agnoset in sinu suo levat;fetas ipse portat ".
ISA|40|12|Quis mensus est pugillo aquaset caelos palmo disposuit,modio continuit pulverem terraeet libravit in pondere monteset colles in statera?
ISA|40|13|Quis direxit spiritum Domini?Aut quis consilium suumostendit illi?
ISA|40|14|Cum quo iniit consilium, et instruxit eumet docuit eum semitam iustitiaeet erudivit eum scientiamet viam prudentiae ostendit illi?
ISA|40|15|Ecce gentes quasi stilla situlaeet quasi momentum pulveris in statera reputantur;ecce insulae quasi pulvis exiguus.
ISA|40|16|Et Libanus non sufficiet ad succendendum,et animalia eius non sufficient ad holocaustum.
ISA|40|17|Omnes gentes, quasi non sint, coram eo;quasi nihilum et inane reputantur ab eo.
ISA|40|18|Cui ergo similem facitis Deum?Aut quam imaginem ponitis ei?
ISA|40|19|Sculptile conflat faber,et aurifex auro figurat illud,et laminis argenteis argentarius.
ISA|40|20|Nimis pauper, ut offerat lignum imputribile:exquirit sibi sapientem artificem,ut statuat simulacrum,quod non moveatur.
ISA|40|21|Numquid non scitis? Numquid non audistis?Numquid non annuntiatum est vobis ab initio?Numquid non intellexistis fundamenta terrae?
ISA|40|22|Qui sedet super gyrum terrae,et habitatores eius sunt quasi locustae;qui extendit sicut velum caeloset expandit eos sicut tabernaculum ad inhabitandum;
ISA|40|23|qui redigit in nihilum principes,iudices terrae velut inane facit.
ISA|40|24|Et quidem neque plantatus neque satusneque radicatus in terra truncus eorum;repente flavit in eos, et aruerunt,et turbo quasi stipulam aufert eos.
ISA|40|25|" Et cui assimilabitis me,quasi aequalis ei sim ego? ",dicit Sanctus.
ISA|40|26|Levate in excelsum oculos vestroset videte: Quis creavit haec?Qui educit in numero militiam eorumet omnes ex nomine vocat;prae multitudine fortitudinis et roboris virtutisque eiusneque unum deest.
ISA|40|27|Quare dicis, Iacob,et loqueris, Israel: Abscondita est via mea a Domino,et a Deo meo iudicium meum transit? ".
ISA|40|28|Numquid nescis? Aut non audisti?Deus sempiternus Dominus,qui creavit terminos terrae;non deficiet neque laborabit,nec est investigatio sapientiae eius.
ISA|40|29|Qui dat lasso virtutemet invalido robur multiplicat.
ISA|40|30|Deficient pueri et laborabunt,et iuvenes lapsu labentur;
ISA|40|31|qui autem sperant in Domino,mutabunt fortitudinem,assument pennas sicut aquilae,current et non laborabunt,ambulabunt et non deficient.
ISA|41|1|Taceant ante me insulae,et gentes renovent fortitudinem;accedant et tunc loquantur,simul ad iudicium propinquemus.
ISA|41|2|Quis suscitavit ab oriente eum,cuius gressum sequitur iustitia?Dabit in conspectu eius genteset subiciet ei reges,quos reddet quasi pulverem gladius eius,sicut stipulam vento raptam arcus eius.
ISA|41|3|Persequetur eos, transibit in pace;semita sub pedibus eius non apparebit.
ISA|41|4|Quis operatus est et fecit,vocans generationes ab exordio?Ego Dominus, primuset cum novissimis ego sum.
ISA|41|5|Viderunt insulae et timuerunt,extrema terrae obstupuerunt,appropinquaverunt et accesserunt.
ISA|41|6|Unusquisque proximo suo auxiliabituret fratri suo dicet: " Confortare ".
ISA|41|7|Confortabit faber aurificem,percutiens malleo eum, qui cudit,dicens de glutino: " Bonum est ";et roborat eum clavis,ut non moveatur.
ISA|41|8|Tu autem, Israel, serve meus,Iacob, quem elegi,semen Abraham amici mei,
ISA|41|9|quem apprehendi ab extremis terrae,et a longinquis eius vocavi teet dixi tibi: " Servus meus es tu;elegi te et non abieci te ".
ISA|41|10|Ne timeas, quia ego tecum sum;ne declines, quia ego Deus tuus:confortabo te et auxiliabor tibiet sustentabo te dextera iustitiae meae.
ISA|41|11|Ecce confundentur et erubescentomnes, qui irascuntur adversum te;erunt quasi non sintet peribunt viri, qui contradicunt tibi.
ISA|41|12|Quaeres eos et non inveniesviros, qui rixantur tecum;erunt quasi non sint et veluti nihilum,viri bellantes adversum te.
ISA|41|13|Quia ego Dominus Deus tuusapprehendens manum tuamdicensque tibi: " Ne timeas;ego auxiliabor tibi.
ISA|41|14|Noli timere, vermis Iacob,homines ex Israel.Ego auxiliabor tibi ", dicit Dominuset redemptor tuus, Sanctus Israel.
ISA|41|15|Ecce posui te quasi plaustrum triturans novum,habens rostra serrantia.Triturabis montes et comminueset colles quasi pulverem pones.
ISA|41|16|Ventilabis eos, et ventus tollet eos,et turbo disperget eos;et tu exsultabis in Domino,in Sancto Israel laetaberis.
ISA|41|17|Egeni et pauperes quaerunt aquas, et non sunt,lingua eorum siti aruit.Ego, Dominus, exaudiam eos,Deus Israel non derelinquam eos.
ISA|41|18|Aperiam in decalvatis collibus fluminaet in medio vallium fontes;ponam desertum in stagna aquarumet terram aridam in rivos aquarum.
ISA|41|19|Plantabo in deserto cedrum,acaciam et myrtum et lignum olivae;ponam in solitudine abietem,ulmum et cupressum simul,
ISA|41|20|ut videant et sciantet recogitent et intellegant pariterquia manus Domini fecit hoc,et Sanctus Israel creavit illud.
ISA|41|21|Proferte causam vestram, dicit Dominus;afferte, si quid firmum habetis, dixit Rex Iacob.
ISA|41|22|Accedant et nuntient nobis, quaecumque ventura sunt.Priora, quae fuerunt, nuntiate,ut ponamus cor nostrum et sciamus novissima eorum;et, quae ventura sunt, indicate nobis.
ISA|41|23|Annuntiate, quae ventura sunt in futurum,ut sciamus quia dii estis vos;bene quoque aut male facite,ut inspiciamus et videamus simul.
ISA|41|24|Ecce vos estis nihilum,et opus vestrum nihil valet;abominatio est, qui eligit vos.
ISA|41|25|Suscitavi ab aquilone,et venit ab ortu solis;vocavi eum nomine;et conculcabit potentes quasi lutumet velut plastes calcans humum.
ISA|41|26|Quis annuntiavit ab exordio, ut sciamus,et a principio, ut dicamus: " Iustum est "?Non est neque annuntians neque praedicensneque audiens sermones vestros.
ISA|41|27|Primus ad Sion: Ecce adsunt;et Ierusalem laeta nuntiantem do.
ISA|41|28|Et vidi, et nemo erat,ex istis nullus consiliator,ut, si eos interrogarem,responderent verbum.
ISA|41|29|Ecce omnes iniquitas,vana opera eorum;ventus et inanesimulacra eorum.
ISA|42|1|Ecce servus meus, suscipiam eum;electus meus, complacet sibi in illo anima mea;dedi spiritum meum super eum,iudicium gentibus proferet.
ISA|42|2|Non clamabit neque vociferabitur,nec audietur vox eius foris.
ISA|42|3|Calamum quassatum non conteretet linum fumigans non exstinguet;in veritatem proferet iudicium.
ISA|42|4|Non languebit nec frangetur,donec ponat in terra iudicium;et legem eius insulae exspectant.
ISA|42|5|Haec dicit Dominus Deus,creans caelos et extendens eos,firmans terram et quae germinant ex ea,dans flatum populo, qui est super eam,et spiritum calcantibus eam:
ISA|42|6|" Ego, Dominus, vocavi te in iustitiaet apprehendi manum tuam;et formavi te et dedi tein foedus populi, in lucem gentium,
ISA|42|7|ut aperires oculos caecorumet educeres de conclusione vinctum,de domo carceris sedentes in tenebris.
ISA|42|8|Ego Dominus: hoc est nomen meum;et gloriam meam alteri non daboet laudem meam sculptilibus.
ISA|42|9|Quae prima fuerunt, ecce venerunt;nova quoque ego annuntio:antequam oriantur, audita vobis faciam ".
ISA|42|10|Cantate Domino canticum novum,laus eius ab extremis terrae;qui descenditis in mare, et plenitudo eius,insulae et habitatores earum.
ISA|42|11|Exsultent desertum et civitates eius,vici, quos habitat Cedar.Iubilent habitatores Petrae,de vertice montium clament.
ISA|42|12|Ponant Domino gloriamet laudem eius in insulis nuntient.
ISA|42|13|Dominus sicut fortis egredietur,sicut vir proeliator suscitabit zelum;vociferabitur et conclamabit,super inimicos suos praevalebit.
ISA|42|14|" Tacui semper, silui, patiens fui;sicut parturiens ululabo,gemam et fremam simul.
ISA|42|15|Desertos faciam montes et colleset omne gramen eorum exsiccabo;et ponam flumina in insulaset stagna arefaciam.
ISA|42|16|Et ducam caecos in viam, quam nesciunt,et in semitis, quas ignoraverunt, ambulare eos faciam;ponam tenebras coram eis in lucemet prava in recta.Haec verba faciam eiset non dereliquam eos ".
ISA|42|17|Conversi sunt retrorsum;confundantur confusione, qui confidunt in sculptili,qui dicunt conflatili: Vos dii nostri ".
ISA|42|18|Surdi, audite;et caeci, intuemini ad videndum.
ISA|42|19|Quis caecus sicut servus meus,et surdus sicut nuntius, quem ego mittam?Quis caecus sicut qui restitutus est?Et quis caecus sicut servus Domini?
ISA|42|20|Multa vidisti, sed non servas;aures aperuisti, sed non audis.
ISA|42|21|Dominus voluit propter iustitiam suammagnificare legem et extollere.
ISA|42|22|Ipse autem populus direptus et vastatus;in foveis conclusi omnes,et in domibus carcerum absconditi sunt.Facti sunt in rapinam, nec est qui eruat;in direptionem, nec est qui dicat: " Redde! ".
ISA|42|23|Quis est in vobis, qui audiat hoc,attendat et auscultet futura?
ISA|42|24|Quis dedit in direptionem Iacobet Israel vastantibus?Nonne Dominus ipse, cui peccavimus?Et noluerunt in viis eius ambulareet non audierunt legem eius.
ISA|42|25|Et effudit super eum indignationem furoris suiet forte bellum.Et combussit eum in circuitu, et non cognovit;et succendit eum, et non intellexit.
ISA|43|1|Et nunc haec dicit Dominus,qui creavit te, Iacob, et formavit te, Israel: Noli timere, quia redemi teet vocavi te nomine tuo; meus es tu.
ISA|43|2|Cum transieris per aquas, tecum ero,et flumina non operient te;cum ambulaveris in igne, non combureris,et flamma non ardebit in te,
ISA|43|3|quia ego Dominus Deus tuus,Sanctus Israel, salvator tuus:dedi propitiationem tuam Aegyptum,Aethiopiam et Saba pro te.
ISA|43|4|Quoniam pretiosus factus es in oculis meiset gloriosus, ego diligo teet dabo homines pro teet populos pro anima tua.
ISA|43|5|Noli timere, quoniam ego tecum sum:ab oriente adducam semen tuumet ab occidente congregabo te.
ISA|43|6|Dicam aquiloni: "Da"et austro: "Noli prohibere;affer filios meos de longinquoet filias meas ab extremis terrae.
ISA|43|7|Omnem, qui vocatur nomine meo,in gloriam meam creavi eum,formavi eum et feci eum".
ISA|43|8|Educ foras populum caecum, et oculos habentem,surdos, et aures eis sunt.
ISA|43|9|Omnes gentes congregentur simul,et colligantur nationes:quis in eis annuntiabit istudet priora audire nos faciet?Dent testes suos et iustificenturet audiant et dicant: "Vere".
ISA|43|10|Vos testes mei, dicit Dominus,et servus meus, quem elegi,ut sciatis et credatis mihiet intellegatis quia ego ipse sum;ante me non est formatus Deuset post me non erit.
ISA|43|11|Ego, ego sum Dominus,et non est absque me salvator.
ISA|43|12|Ego, annuntiavi et salvavi;auditum feci, et non fuit in vobis alienus;et vos testes mei, dicit Dominus,et ego Deus,
ISA|43|13|iam ab initio ego ipse.Et non est qui de manu mea eruat; operabor, et quis avertet illud? ".
ISA|43|14|Haec dicit Dominus, redemptor vester,Sanctus Israel: Propter vos misi in Babylonemet detraxi fugitivos universoset Chaldaeos in navibus suis gloriantes.
ISA|43|15|Ego Dominus, Sanctus vester,creans Israel, rex vester ".
ISA|43|16|Haec dicit Dominus,qui dedit in mari viamet in aquis torrentibus semitam;
ISA|43|17|qui eduxit quadrigam et equum,agmen et robustum;simul iacuerunt nec resurgent,contriti sunt quasi linum et exstincti sunt.
ISA|43|18|" Ne memineritis priorumet antiqua ne intueamini:
ISA|43|19|ecce ego facio nova,et nunc orientur: nonne cognoscitis ea?Utique ponam in deserto viamet in invio flumina.
ISA|43|20|Glorificabit me bestia agri,dracones et struthiones,quia dedi in deserto aquas,flumina in invio,ut darem potum populo meo, electo meo.
ISA|43|21|Populum istum formavi mihi;laudem meam narrabunt.
ISA|43|22|Non me invocasti, Iacob;immo taedio mei affectus es, Israel.
ISA|43|23|Non obtulisti mihi agnos holocausti tuiet victimis tuis non glorificasti me;non te gravavi in oblationenec laborem tibi praebui in ture.
ISA|43|24|Non emisti mihi argento calamumet adipe victimarum tuarum non inebriasti me;verumtamen servire me fecisti in peccatis tuis,praebuisti mihi laborem in iniquitatibus tuis.
ISA|43|25|Ego, ego sum ipse, qui deleo iniquitates tuas propter meet peccatorum tuorum non recordabor.
ISA|43|26|Memorem me redde, iudicium agamus simul:narra, ut iustificeris.
ISA|43|27|Pater tuus primus peccavit,et interpretes tui praevaricati sunt in me;
ISA|43|28|et contaminavi principes sanctuarii,dedi ad internecionem Iacobet Israel in opprobrium ".
ISA|44|1|Et nunc audi, Iacob serve meus,et Israel, quem elegi.
ISA|44|2|Haec dicit Dominus, qui fecit teet formavit te ab utero,auxiliator tuus: Noli timere, serve meus Iacob,et dilecte, quem elegi.
ISA|44|3|Effundam enim aquas super terram sitientemet fluenta super aridam;effundam spiritum meum super semen tuumet benedictionem meam super stirpem tuam:
ISA|44|4|et germinabunt inter herbasquasi salices iuxta praeterfluentes aquas.
ISA|44|5|Iste dicet: "Domini ego sum",et ille vocabit se nomine Iacob;et hic scribet manu sua: "Domino", et inscribetur nomine Israel ".
ISA|44|6|Haec dicit Dominus, rex Israelet redemptor eius, Dominus exercituum: Ego primus et ego novissimus,et absque me non est Deus.
ISA|44|7|Quis similis mei? Conclamet et annuntietet exponat mihi,ex quo constitui populum antiquum;ventura et, quae futura sunt, annuntiet nobis.
ISA|44|8|Nolite timere neque conturbemini;nonne ex tunc audire te feci et annuntiavi?Vos estis testes mei.Numquid est Deus absque meaut Petra, quam ego non noverim? ".
ISA|44|9|Plastae idoli omnes nihil sunt, et pretiosa eorum non proderunt eis; testes eorum non vident neque intellegunt, ut confundantur.
ISA|44|10|Quis formavit deum et sculptile conflavit lucrum non quaerens?
ISA|44|11|Ecce omnes participes eius confundentur; fabri enim sunt ex hominibus: conveniant omnes, stent; pavebunt, confundentur simul.
ISA|44|12|Faber ferrarius securim operatur in prunis et in malleis format illam et polit eam in brachio fortitudinis suae; esurit et deficit, non bibit aquam et lassescit.
ISA|44|13|Artifex lignarius extendit normam, describit illud stilo, operatur illud scalpellis et circino describit illud quasi imaginem viri, quasi speciosum hominem, qui resideat in domo.
ISA|44|14|Succidit sibi cedros et arripit ilicem et quercum, quae steterat inter ligna saltus; plantavit pinum, quam pluvia nutrivit.
ISA|44|15|Homini facta sunt ad comburendum; sumit ex eis, ut calefaciat, et succendit et coquit panes. De reliquo autem operatur deum et adorat; facit sculptile et curvatur ante illud.
ISA|44|16|Medium eius comburit igne et medio eius carnes assat, manducat assaturam et saturatur et calefit et dicit: " Vah, calefactus sum, vidi focum ".
ISA|44|17|Reliquum autem eius deum fecit, sculptile sibi; curvatur ante illud et adorat illud et obsecrat dicens: " Libera me, quia deus meus es tu ".
ISA|44|18|Nescierunt neque intellexerunt; nam clausit oculos eorum, ne videant et ne intellegant corde suo.
ISA|44|19|Non recogitant in corde suo, scientia et intellegentia carent, ut dicant: " Medietatem eius combussi igne et coxi super carbones eius panes, coxi carnes et comedi et de reliquo eius abominationem faciam; ante truncum ligni procidam? ".
ISA|44|20|Cinere vescitur; cor insipiens decepit eum, et non liberabit animam suam neque dicet: " Nonne mendacium est in dextera mea? ".
ISA|44|21|Memento horum, Iacob,et Israel, quoniam servus meus es tu;formavi te, servus meus es tu,Israel, non decipies me.
ISA|44|22|Delevi ut nubem iniquitates tuaset quasi nebulam peccata tua;revertere ad me,quoniam redemi te.
ISA|44|23|Exsultate, caeli, quoniam hoc fecit Dominus;iubilate, fundamenta terrae,resonate, montes, laudationem,saltus et omne lignum eius,quoniam redemit Dominus Iacobet in Israel glorificabitur.
ISA|44|24|Haec dicit Dominus, redemptor tuus et formator tuus ex utero: Ego sum Dominus, qui feci omnia,extendi caelos solus,expandi terram; et quis mecum?
ISA|44|25|Qui irrita facio signa divinorumet hariolos stultos reddo;compello sapientes retrorsumet scientiam eorum vanam facio;
ISA|44|26|qui suscito verbum servi meiet consilium nuntiorum meorum compleo.Qui dico Ierusalem: "Habitaberis" et civitatibus Iudae: "Aedificabimini"et deserta eius suscitabo;
ISA|44|27|qui dico profundo: "Desolare,et flumina tua arefaciam";
ISA|44|28|qui dico de Cyro: "Pastor meus estet omnem voluntatem meam complebit";qui dico Ierusalem: "Aedificaberis",et templo: "Fundaberis" ".
ISA|45|1|Haec dicit Dominus de uncto suo Cyro: Apprehendi dexteram eius,ut subiciam ante faciem eius genteset dorsa regum vertamet aperiam coram eo ianuas;et portae non claudentur.
ISA|45|2|Ego ante te iboet montes humiliabo;portas aereas conteramet vectes ferreos confringam.
ISA|45|3|Et dabo tibi thesauros absconditoset divitias occultas,ut scias quia ego Dominus,qui vocavi te nomine tuo, Deus Israel.
ISA|45|4|Propter servum meum Iacobet Israel electum meum,et vocavi te nomine tuo;designavi te, et non cognovisti me.
ISA|45|5|Ego Dominus, et non est amplius:extra me non est Deus.Accinxi te, et non cognovisti me,
ISA|45|6|ut sciant ab ortu solis et ab occidentequoniam absque me nullus est.Ego Dominus, et non est alter,
ISA|45|7|formans lucem et creans tenebras,faciens pacem et creans malum:ego Dominus faciens omnia haec.
ISA|45|8|Rorate, caeli, desuper, et nubes pluant iustitiam;aperiatur terraet germinet salvationem;et iustitia oriatur simul:ego Dominus creavi eam ".
ISA|45|9|Vae, qui contradicit fictori suo,testa de vasis fictilibus terrae!Numquid dicet lutum figulo suo: " Quid facis? "et " Opus tuum absque manibus est "?
ISA|45|10|Vae, qui dicit patri: " Quid generas? "et mulieri: " Quid parturis? ".
ISA|45|11|Haec dicit Dominus,Sanctus Israel, plastes eius: Numquid ventura interrogatis me super filios meoset super opus manuum mearum mandatis mihi?
ISA|45|12|Ego feci terramet hominem super eam creavi ego;manus meae tetenderunt caelos,et omni militiae eorum mandavi.
ISA|45|13|Ego suscitavi eum in iustitiaet omnes vias eius dirigam;ipse aedificabit civitatem meamet captivitatem meam dimittetnon in pretio neque in muneribus ",dicit Dominus exercituum.
ISA|45|14|Haec dicit Dominus: Labor Aegypti et negotiatio Aethiopiaeet Sabaim viri sublimesad te transibunt et tui erunt;post te ambulabunt,vincti manicis pergent et te adorabuntteque deprecabuntur:Tantum in te est Deus,et non est absque te Deus!".
ISA|45|15|Vere tu es Deus absconditus,Deus Israel, salvator.
ISA|45|16|Confusi sunt et erubuerunt omnes,simul abierunt in confusionem fabricatores idolorum.
ISA|45|17|Israel salvatus est in Domino salute aeterna;non confundemini et non erubescetisusque in saeculum saeculi.
ISA|45|18|Quia haec dicit Dominus,qui creavit caelos, ipse Deus,qui formavit terram et fecit eam, ipse fundavit eam;non ut vacua esset, creavit eam,ut habitaretur, formavit eam: Ego Dominus, et non est alius.
ISA|45|19|Non in abscondito locutus sum,in loco terrae tenebroso;non dixi semini Iacob:Frustra quaerite me".Ego Dominus loquens iustitiam,annuntians recta.
ISA|45|20|Congregamini et venite et accedite simul,qui salvati estis ex gentibus.Nescierunt, qui levant lignum sculpturae suaeet rogant deum non salvantem.
ISA|45|21|Annuntiate et venite et consiliamini simul.Quis auditum fecit hoc ab initio,ex tunc praedixit illud?Numquid non ego Dominus,et non est ultra Deus absque me?Deus iustus et salvans non est praeter me.
ISA|45|22|Convertimini ad me et salvi eritis,omnes fines terrae,quia ego Deus, et non est alius.
ISA|45|23|In memetipso iuravi:Egressa est de ore meo iustitia,verbum, quod non revertetur;quia mihi curvabitur omne genu,et iurabit omnis lingua ".
ISA|45|24|" Tantum in Domino " dicent sunt iustitiae et robur! ".Ad eum venient et confundenturomnes, qui repugnant ei;
ISA|45|25|in Domino iustificabitur et laudabituromne semen Israel.
ISA|46|1|Concidit Bel, incurvavit se Nabo;fuerunt simulacra eorum bestiis et iumentis.Statuae vestrae portantur, onera lassis.
ISA|46|2|Se incurvaverunt et conciderunt simul;non potuerunt salvare onuset ipsi in captivitatem ibunt.
ISA|46|3|Audite me, domus Iacobet omne residuum domus Israel,qui portamini ab utero,qui gestamini a vulva.
ISA|46|4|Usque ad senectam ego ipseet usque ad canos ego portabo;et ego feci et ego feram,ego portabo et salvabo.
ISA|46|5|Cui assimilatis me et adaequatiset comparatis me, et erimus similes?
ISA|46|6|Qui effundunt aurum de sacculoet argentum statera ponderant,conducunt aurificem, ut faciat deum,et procidunt et adorant.
ISA|46|7|Portant illum in umeris gestanteset ponentes in loco suo;et stabit ac de loco suo non movebitur;sed et si quis clamat ad eum, non respondet;de tribulatione eius non salvabit eum.
ISA|46|8|Mementote istud et confundamini;redite, praevaricatores, ad cor.
ISA|46|9|Recordamini prioris saeculi,quoniam ego sum Deus,et non est ultra Deus,nec est similis mei.
ISA|46|10|Annuntians ab exordio novissimumet ab initio, quae necdum facta sunt,dicens: " Consilium meum stabit,et omnem voluntatem meam faciam ".
ISA|46|11|Vocans ab oriente avem rapacemet de terra longinqua virum consilii mei;et locutus sum et adducam illud,decrevi et faciam illud.
ISA|46|12|Audite me, duri corde,qui longe estis a iustitia.
ISA|46|13|Prope feci iustitiam meam, non elongabitur;et salus mea non morabitur:et dabo in Sion salutemet Israeli gloriam meam.
ISA|47|1|Descende, sede in pulvere,virgo filia Babylon;sede in terra sine solio,filia Chaldaeorum,quia ultra non vocaberismollis et tenera.
ISA|47|2|Tolle molam et mole farinam;depone velum tuum,subleva stolam, revela crura,transi flumina.
ISA|47|3|Revelabitur ignominia tua,et videbitur opprobrium tuum. Ultionem capiam,nemini parcam ",
ISA|47|4|dicit Redemptor noster, Dominus exercituum nomen illius,Sanctus Israel.
ISA|47|5|Sede tacens et intra in tenebras,filia Chaldaeorum,quia non vocaberis ultraDomina regnorum.
ISA|47|6|Iratus sum super populum meum,contaminavi hereditatem meamet dedi eos in manu tua;non posuisti eis misericordias,super senem aggravasti iugum tuum valde
ISA|47|7|et dixisti: " In sempiternum ero domina ".Non posuisti haec super cor tuumneque recordata es novissimi tui.
ISA|47|8|Et nunc audi haec, delicata,quae habitas confidenteret dicis in corde tuo: Ego, et praeter me non est altera, non sedebo vidua et orbitatem ignorabo ".
ISA|47|9|Venient tibi duo haecsubito in die una,orbitas et viduitas;repente venerunt super tepropter multitudinem maleficiorum tuorum,propter abundantiam incantationum tuarum.
ISA|47|10|Et fiduciam habuisti in malitia tuaet dixisti: " Non est qui videat me ".Sapientia tua et scientia tua,haec decepit te.Et dixisti in corde tuo: Ego, et praeter me non est altera ".
ISA|47|11|Veniet super te malum,et nescies avertere;et irruet super te calamitas,quam non poteris expiare;veniet super te repentemiseria, quam nescies.
ISA|47|12|Sta cum incantationibus tuiset cum multitudine maleficiorum tuorum,in quibus laborasti ab adulescentia tua:forte poteris iuvari, forte terrebis.
ISA|47|13|Defecisti in multitudine consiliorum tuorum;stent et salvent te, qui metiuntur caelum,qui contemplantur sideraet annuntiant singulis noviluniisventura tibi.
ISA|47|14|Ecce facti sunt quasi stipula,ignis combussit eos.Non liberabunt seipsosde manu flammae;non sunt prunae, quibus calefiant,nec focus, ut sedeant ad eum.
ISA|47|15|Sic fiunt tibi incantatores tui,in quibuscumque laborasti ab adulescentia tua;unusquisque in via sua errat,non est qui salvet te.
ISA|48|1|Audite hoc, domus Iacob,qui vocamini nomine Israelet de aquis Iudae existis,qui iuratis in nomine Dominiet Deum Israel invocatisnon in veritate neque in iustitia.
ISA|48|2|De civitate enim sancta vocati suntet super Deum Israel constabiliti sunt;Dominus exercituum nomen eius.
ISA|48|3|Priora ex tunc annuntiavi,et ex ore meo exierunt,et audita feci ea;repente operatus sum, et venerunt.
ISA|48|4|Scivi enim quia durus es tu,et nervus ferreus cervix tua,et frons tua aerea.
ISA|48|5|Praedixi tibi ex tunc;antequam venirent, indicavi tibi,ne forte diceres: "Idolum meum operatum est haec,et sculptile meum et conflatile mandaverunt ista ".
ISA|48|6|Quae audisti, vide omnia;vos autem num annuntiabitis?Audita facio tibi nova ex nuncet occulta, quae nescis.
ISA|48|7|Nunc creata sunt et non ex tunc,et ante eorum diem, et non audisti ea,ne forte diceres: "Ecce ego cognovi ea ".
ISA|48|8|Neque audisti neque cognovisti,neque ex tunc aperta est auris tua;scio enim quia praevaricans praevaricariset transgressor ex utero vocaris.
ISA|48|9|Propter nomen meum longe faciam furorem meumet propter laudem meam infrenabo me super te,ne perdam te.
ISA|48|10|Ecce excoxi te, sed non quasi argentum;probavi te in camino paupertatis.
ISA|48|11|Propter me, propter me faciam,ut non blasphemer;et gloriam meam alteri non dabo.
ISA|48|12|Audi me, Iacob,et Israel, quem ego vocavi;ego, ego primuset ego novissimus.
ISA|48|13|Manus mea fundavit terram,et dextera mea expandit caelos;ego voco eos, et stant simul.
ISA|48|14|Congregamini, omnes vos, et audite:Quis de eis annuntiavit haec?Dominus dilexit eum;faciet voluntatem suam in Babyloneet brachium suum in Chaldaeis.
ISA|48|15|Ego, ego locutus sum et vocavi eum;adduxi eum, et prospera fuit via eius.
ISA|48|16|Accedite ad me et audite hoc:Non a principio in abscondito locutus sum;ex tempore, antequam fieret, ibi eram;et nunc Dominus Deus misit me cum spiritu suo.
ISA|48|17|Haec dicit Dominus,redemptor tuus, Sanctus Israel:Ego Dominus Deus tuus docens te utilia,gubernans te in via, qua ambulas.
ISA|48|18|Utinam attendisses mandata mea!Facta fuisset sicut flumen pax tua,et iustitia tua sicut gurgites maris;
ISA|48|19|et fuisset quasi arena semen tuum,et stirps uteri tui ut lapilli eius;non interisset et non fuisset attritumnomen eius a facie mea.
ISA|48|20|Egredimini de Babylone, fugite a Chaldaeis,in voce exsultationis annuntiate;auditum facite hoc, efferte illud usque ad extrema terrae,dicite: " Redemit Dominus servum suum Iacob ".
ISA|48|21|Non sitierunt, cum per desertum duceret eos;aquam de petra produxit eiset scidit petram, et fluxerunt aquae.
ISA|48|22|Non est pax impiis, dicit Dominus.
ISA|49|1|Audite me, insulae, et attendite, populi de longe;Dominus ab utero vocavit me,de ventre matris meae recordatus est nominis mei;
ISA|49|2|et posuit os meum quasi gladium acutum,in umbra manus suae protexit meet posuit me sicut sagittam electam,in pharetra sua abscondit me
ISA|49|3|et dixit mihi: " Servus meus es tu,Israel, in quo gloriabor ".
ISA|49|4|Et ego dixi: " In vacuum laboravi,sine causa et vane fortitudinem meam consumpsi;verumtamen iudicium meum cum Domino,et merces mea cum Deo meo ".
ISA|49|5|Et nunc dicit Dominus,qui formavit me ex utero servum sibi,ut reducerem Iacob ad eum,et Israel ei congregaretur;et glorificatus sum in oculis Domini,et Deus meus factus est fortitudo mea.
ISA|49|6|Et dixit: " Parum est ut sis mihi servusad suscitandas tribus Iacobet reliquias Israel reducendas:dabo te in lucem gentium,ut sit salus mea usque ad extremum terrae ".
ISA|49|7|Haec dicit Dominus,redemptor Israel, Sanctus eius,ad contemptum in anima,ad abominatum in gente,ad servum dominorum: Reges videbunt et consurgent,principes quoque et adorabunt,propter Dominum, quia fidelis est,Sanctum Israel, qui elegit te ".
ISA|49|8|Haec dicit Dominus: In tempore beneplaciti exaudivi teet in die salutis auxiliatus sum tui;et servavi te et dedi te in foedus populi,ut suscitares terramet distribueres hereditates dissipatas;
ISA|49|9|ut diceres his, qui vincti sunt: "Exite",et his, qui in tenebris: "Revelamini".Super vias pascentur,et in omnibus collibus decalvatis pascua eorum;
ISA|49|10|non esurient neque sitient,et non percutiet eos aestus vel sol,quia miserator eorum reget eoset ad fontes aquarum adducet eos.
ISA|49|11|Et ponam omnes montes meos in viam,et semitae meae exaltabuntur.
ISA|49|12|Ecce isti de longe venient,et ecce illi ab aquilone et mari,et isti de terra Sinim ".
ISA|49|13|Laudate, caeli, et exsulta, terra;iubilate, montes, laudem,quia consolatur Dominus populum suumet pauperum suorum miseretur.
ISA|49|14|Et dixit Sion: " Dereliquit me Dominus,et Dominus oblitus est mei ".
ISA|49|15|Numquid oblivisci potest mulier infantem suum,ut non misereatur filio uteri sui?Et si illa oblita fuerit,ego tamen non obliviscar tui.
ISA|49|16|Ecce in manibus meis descripsi te;muri tui coram me semper.
ISA|49|17|Festinant structores tui;destruentes te et dissipantes a te exibunt.
ISA|49|18|Leva in circuitu oculos tuos et vide:omnes isti congregati sunt, venerunt tibi. Vivo ego, dicit Dominus,quia omnibus his velut ornamento vestieriset circumdabis tibi eos quasi sponsa ".
ISA|49|19|Quia ruinae tuae et solitudines tuaeet terra eversa:nunc angusta eris prae habitatoribus;et longe erunt, qui devorabant te.
ISA|49|20|Adhuc dicent in auribus tuisfilii orbitatis tuae: Angustus est mihi locus;fac spatium mihi, ut habitem ".
ISA|49|21|Et dices in corde tuo: Quis genuit mihi istos?Ego orbata et non pariens,transmigrata et captiva;et istos quis enutrivit?Ecce ego relicta eram sola;et isti ubi erant? ".
ISA|49|22|Haec dicit Dominus Deus: Ecce levabo ad gentes manum meamet ad populos exaltabo signum meum;et afferent filios tuos in ulnis,et filiae tuae super umeros portabuntur.
ISA|49|23|Et erunt reges nutricii tui,et reginae nutrices tuae;vultu in terram demisso adorabunt teet pulverem pedum tuorum lingent.Et scies quia ego Dominus:non confundentur, qui sperant in me ".
ISA|49|24|Numquid tolletur a forti praeda,aut, quod captum fuerit, a robusto salvari poterit?
ISA|49|25|Quia haec dicit Dominus: Equidem et captivus a forti tolletur,et, quod ablatum fuerit a robusto, salvabitur;cum his, qui contendebant tecum, ego contendamet filios tuos ego salvabo.
ISA|49|26|Et cibabo hostes tuos carnibus suis,et quasi musto sanguine suo inebriabuntur;et sciet omnis caro quia ego Dominus salvator tuus,et redemptor tuus Fortis Iacob ".
ISA|50|1|Haec dicit Dominus: Ubinam est liber repudii matris vestrae,quo dimisi eam?Aut quis est creditor meus,cui vendidi vos?Ecce in iniquitatibus vestris venditi estis,et in sceleribus vestris dimissa est mater vestra.
ISA|50|2|Cur veni, et non erat vir,vocavi, et non erat qui responderet?Numquid abbreviata est manus mea,ut non possim redimere?Aut non est in me virtus ad liberandum?Ecce in increpatione mea exsiccabo mare,ponam flumina in siccum;computrescent pisces sine aquaet morientur in siti.
ISA|50|3|Induam caelos luctuet saccum ponam operimentum eorum ".
ISA|50|4|Dominus Deus dedit mihi linguam eruditam,ut sciam sustentare eum, qui lassus est, verbo;excitat mane, mane excitat mihi aurem,ut audiam quasi discipulus.
ISA|50|5|Dominus Deus aperuit mihi aurem;ego autem non rebellavi, retrorsum non abii.
ISA|50|6|Dorsum meum dedi percutientibuset genas meas vellentibus:faciem meam non avertiab increpationibus et sputis.
ISA|50|7|Dominus Deus auxiliator meus;ideo non sum confusus,ideo posui faciem meam ut petram durissimamet scio quoniam non confundar.
ISA|50|8|Iuxta est qui iustificat me;quis contradicet mihi? Stemus simul.Quis est adversarius meus? Accedat ad me.
ISA|50|9|Ecce Dominus Deus auxiliator meus;quis est qui condemnet me?Ecce omnes quasi vestimentum conterentur,tinea comedet eos.
ISA|50|10|Quis ex vobis timet Dominum,audiens vocem servi sui?Qui ambulavit in tenebris,et non est lumen ei,speret in nomine Dominiet innitatur super Deum suum.
ISA|50|11|Ecce vos omnes, qui accenditis ignem,accincti sagittis,ambulate in lumine ignis vestriet in sagittis, quas succendistis.De manu mea factum est hoc vobis;in doloribus recumbetis.
ISA|51|1|Audite me, qui sequimini iustitiam,qui quaeritis Dominum;attendite ad petram, unde excisi estis,et ad cavernam laci, de qua praecisi estis.
ISA|51|2|Attendite ad Abraham patrem vestrumet ad Saram, quae peperit vos;quia unum vocavi eumet benedixi ei et multiplicavi eum.
ISA|51|3|Consolatur enim Dominus Sion,consolatur omnes ruinas eius;et ponit desertum eius quasi Edenet solitudinem eius quasi hortum Domini.Gaudium et laetitia invenietur in ea,gratiarum actio et vox laudis.
ISA|51|4|Attendite ad me, popule meus;et nationes, me audite,quia lex a me exiet,et iudicium meum in lucem populorum statuam.
ISA|51|5|Prope est iustitia mea,egressa est salus mea,et brachia mea populos iudicabunt;in me insulae sperabuntet ad brachium meum attendent.
ISA|51|6|Levate in caelum oculos vestroset inspicite in terram deorsum,quia caeli sicut fumus liquescent,et terra sicut vestimentum atteretur,et habitatores eius sicut haec interibunt.Salus autem mea in sempiternum erit,et iustitia mea non deficiet.
ISA|51|7|Audite me, qui scitis iustitiam,popule, in cuius corde est lex mea:nolite timere opprobrium hominumet blasphemias eorum ne metuatis.
ISA|51|8|Sicut enim vestimentum sic comedet eos vermis,et sicut lanam sic devorabit eos tinea;iustitia autem mea in sempiternum erit,et salus mea in generationes generationum.
ISA|51|9|Consurge, consurge, induere fortitudinem,brachium Domini;consurge sicut in diebus antiquis,in generationibus saeculorum.Numquid non tu percussisti Rahab,vulnerasti draconem?
ISA|51|10|Numquid non tu siccasti mare,aquam abyssi vehementis,qui posuisti profundum maris viam,ut transirent liberati?
ISA|51|11|Et redempti a Domino revertenturet venient in Sion laudantes;et laetitia sempiterna super capita eorum,gaudium et laetitiam obtinebunt;fugiet dolor et gemitus.
ISA|51|12|Ego, ego ipse consolator vester.Quis tu, ut timeas ab homine mortaliet a filio hominis, qui quasi fenum ita arescet?
ISA|51|13|Et oblitus es Domini factoris tui,qui tetendit caelos et fundavit terram;et formidasti iugiter tota diea facie furoris eius, qui te tribulabat,cum parabat ad perdendum.Ubi nunc est furor tribulantis?
ISA|51|14|Cito captivus liberabituret non morietur in fovea,nec deficiet panis eius.
ISA|51|15|Ego enim sum Dominus Deus tuus,qui conturbo mare,et intumescunt fluctus eius;Dominus exercituum nomen eius.
ISA|51|16|Posui verba mea in ore tuoet in umbra manus meae protexi te,cum extendebam caelos et fundabam terramet dicebam ad Sion: "Populus meus es tu ".
ISA|51|17|Elevare, elevare, consurge, Ierusalem,quae bibisti de manu Domini calicem irae eius;poculum soporis bibisti,epotasti.
ISA|51|18|Non est qui sustentet eamex omnibus filiis, quos genuit;et non est qui apprehendat manum eiusex omnibus filiis, quos enutrivit.
ISA|51|19|Duo sunt quae occurrerunt tibi;quis contristabitur super te?Vastitas et contritio et fames et gladius;quis consolabitur te?
ISA|51|20|Filii tui defecerunt,iacent in capite omnium viarumsicut oryx illaqueatus,pleni indignatione Domini,increpatione Dei tui.
ISA|51|21|Idcirco audi hoc, pauperculaet ebria, sed non a vino.
ISA|51|22|Haec dicit dominator tuus,Dominus et Deus tuus, qui contendit pro populo suo: Ecce tuli de manu tua calicem soporis,poculum indignationis meae;non adicies, ut bibas illum ultra.
ISA|51|23|Et ponam illum in manu eorum, qui te humiliaveruntet dixerunt tibi: "Incurvare, ut transeamus";et ponebas ut terram dorsum tuumet quasi viam transeuntibus ".
ISA|52|1|Consurge, consurge,induere fortitudine tua, Sion;induere vestimentis gloriae tuae,Ierusalem, civitas sanctitatis,quia non adiciet ultra, ut pertranseat per teincircumcisus et immundus.
ISA|52|2|Excutere de pulvere, consurge,captiva Ierusalem;solve vincula colli tui,captiva filia Sion.
ISA|52|3|Quia haec dicit Dominus: " Gratis venumdati estis et sine argento redimemini ".
ISA|52|4|Quia haec dicit Dominus Deus: " In Aegyptum descendit populus meus in principio, ut colonus esset ibi; et Assur sine causa oppressit eum.
ISA|52|5|Et nunc quid mihi est hic, dicit Dominus, quoniam ablatus est populus meus gratis? Dominatores eius ululant, dicit Dominus, et iugiter tota die nomen meum blasphematur.
ISA|52|6|Propter hoc sciet populus meus nomen meum in die illa, quia ego ipse, qui loquebar: "Ecce adsum" ".
ISA|52|7|Quam pulchri super montespedes annuntiantis, praedicantis pacem,annuntiantis bonum, praedicantis salutem,dicentis Sion: "Regnavit Deus tuus!".
ISA|52|8|Vox speculatorum tuorum: levaverunt vocem,simul exsultabunt,quia oculo ad oculum videbunt,cum redierit Dominus ad Sion.
ISA|52|9|Gaudete et exsultate simul,deserta Ierusalem,quia consolatus est Dominus populum suum,redemit Ierusalem.
ISA|52|10|Nudavit Dominus brachium sanctum suumin oculis omnium gentium;et videbunt omnes fines terraesalutare Dei nostri.
ISA|52|11|Recedite, recedite, exite inde,pollutum nolite tangere;exite de medio eius, mundamini,qui fertis vasa Domini.
ISA|52|12|Quoniam non in festinatione exibitisnec in fuga properabitis;praecedet enim vos Dominus,et colliget vos Deus Israel.
ISA|52|13|Ecce prospere aget servus meus;exaltabitur et elevabitur et sublimis erit valde.
ISA|52|14|Sicut obstupuerunt super eum multi,sic deformis erat, quasi non esset hominis species eius,filiorum hominis aspectus eius,
ISA|52|15|sic disperget gentes multas.Super ipsum continebunt reges os suum,quia, quae non sunt narrata eis, videruntet, quae non audierunt, contemplati sunt.
ISA|53|1|" Quis credidit auditui nostro,et brachium Domini cui revelatum est?
ISA|53|2|Et ascendit sicut virgultum coram eoet sicut radix de terra sitienti.Non erat species ei neque decor, ut aspiceremus eum,et non erat aspectus, ut desideraremus eum.
ISA|53|3|Despectus erat et novissimus virorum,vir dolorum et sciens infirmitatem,et quasi abscondebamus vultum coram eo;despectus, unde nec reputabamus eum.
ISA|53|4|Vere languores nostros ipse tulitet dolores nostros ipse portavit;et nos putavimus eum quasi plagatum,percussum a Deo et humiliatum.
ISA|53|5|Ipse autem vulneratus est propter iniquitates nostras,attritus est propter scelera nostra;disciplina pacis nostrae super eum,et livore eius sanati sumus.
ISA|53|6|Omnes nos quasi oves erravimus,unusquisque in viam suam declinavit;et posuit Dominus in eoiniquitatem omnium nostrum ".
ISA|53|7|Afflictus est et ipse subiecit seet non aperuit os suum;sicut agnus, qui ad occisionem ducitur,et quasi ovis, quae coram tondentibus se obmutuitet non aperuit os suum.
ISA|53|8|Angustia et iudicio sublatus est.De generatione eius quis curabit?Quia abscissus est de terra viventium;propter scelus populi mei percussus est ad mortem.
ISA|53|9|Et posuerunt sepulcrum eius cum impiis,cum divitibus tumulum eius,eo quod iniquitatem non fecerit,neque dolus fuerit in ore eius.
ISA|53|10|Et Dominus voluit conterere eum infirmitate.Si posuerit in piaculum animam suam,videbit semen longaevum,et voluntas Domini in manu eius prosperabitur.
ISA|53|11|Propter laborem animae eiusvidebit lucem, saturabitur in scientia sua.Iustificabit iustus servus meus multoset iniquitates eorum ipse portabit.
ISA|53|12|Ideo dispertiam ei multos,et cum fortibus dividet spolia,pro eo quod tradidit in mortem animam suamet cum sceleratis reputatus est;et ipse peccatum multorum tulitet pro transgressoribus rogat.
ISA|54|1|Exsulta, sterilis, quae non peperisti,laetare, gaude, quae non parturisti,quoniam multi sunt filii desertaemagis quam filii nuptae, dicit Dominus.
ISA|54|2|Dilata locum tentorii tuiet pelles tabernaculorum tuorum extende, ne parcas;longos fac funiculos tuoset clavos tuos consolida.
ISA|54|3|Ad dexteram enim et ad laevam penetrabis,et semen tuum hereditabit gentes,quae civitates desertas inhabitabunt.
ISA|54|4|Noli timere, quia non confunderis,neque erubescas, quia non te pudebit;nam confusionis adulescentiae tuae oblivisceriset opprobrii viduitatis tuae non recordaberis amplius.
ISA|54|5|Qui enim fecit te, erit sponsus tuus,Dominus exercituum nomen eius;et redemptor tuus Sanctus Israel,Deus omnis terrae vocabitur.
ISA|54|6|Quia ut mulierem derelictam et maerentem spirituvocavit te Dominus,et uxorem ab adulescentia abiectamdixit Deus tuus.
ISA|54|7|Ad punctum in modico dereliqui teet in miserationibus magnis congregabo te.
ISA|54|8|In momento indignationisabscondi faciem meam parumper a teet in misericordia sempiterna misertus sum tui,dixit redemptor tuus Dominus.
ISA|54|9|Sicut in diebus Noe istud mihi est,cui iuravi, ne inducerem aquas Noe ultra supra terram;sic iuravi, ut non irascar tibiet non increpem te.
ISA|54|10|Montes enim recedent,et colles movebuntur,misericordia autem mea non recedet a te,et foedus pacis meae non movebitur,dixit miserator tuus Dominus.
ISA|54|11|Paupercula, tempestate convulsa absque ulla consolatione,ecce ego sternam super carbunculos lapides tuoset fundabo te in sapphiris;
ISA|54|12|et ponam iaspidem propugnacula tuaet portas tuas in lapides pretiososet omnes terminos tuos in lapides desiderabiles.
ISA|54|13|Universi filii tui erunt discipuli Domini,et magna erit pax filiis tuis;
ISA|54|14|in iustitia fundaberis.Procul eris ab oppressione, quia non timebis,et a pavore, quia non appropinquabit tibi.
ISA|54|15|Ecce, si impetus fiet, non erit ex me; qui impetum fecerit in te, cadet contra te.
ISA|54|16|Ecce, ego creavi fabrumsufflantem in igne prunaset proferentem vas in opus suum;et ego creavi etiam vastatorem ad disperdendum.
ISA|54|17|Omne vas, quod fictum est contra te, frustra erit.Et omnem linguam insurgentem tibi in iudicio confutabis:haec est hereditas servorum Dominiet iustitia eorum ex me, dicit Dominus.
ISA|55|1|Heu! Omnes sitientes, venite ad aquas;et, qui non habetis argentum, properate,emite et comedite, venite, emite absque argentoet absque ulla commutatione vinum et lac.
ISA|55|2|Quare appenditis argentum non in panibuset laborem vestrum non in saturitate?Audite, audientes me, et comedite bonum,ut delectetur in crassitudine anima vestra.
ISA|55|3|Inclinate aurem vestram et venite ad me;audite, ut vivat anima vestra,et feriam vobiscum pactum sempiternum,misericordias David fideles.
ISA|55|4|Ecce testem populis dedi eum,ducem ac praeceptorem gentibus.
ISA|55|5|Ecce gentem, quam nesciebas, vocabis,et gentes, quae te non cognoverunt, ad te current,propter Dominum Deum tuumet Sanctum Israel, quia glorificavit te.
ISA|55|6|Quaerite Dominum, dum inveniri potest;invocate eum, dum prope est.
ISA|55|7|Derelinquat impius viam suam,et vir iniquus cogitationes suas;et revertatur ad Dominum, et miserebitur eius,et ad Deum nostrum, quoniam multus est ad ignoscendum.
ISA|55|8|Non enim cogitationes meae cogitationes vestrae,neque viae vestrae viae meae, dicit Dominus.
ISA|55|9|Quia sicut exaltantur caeli a terra,sic exaltatae sunt viae meae a viis vestris,et cogitationes meae a cogitationibus vestris.
ISA|55|10|Et quomodo descendit imber et nix de caeloet illuc ultra non revertitur,sed inebriat terram et infundit eamet germinare eam facitet dat semen serenti et panem comedenti,
ISA|55|11|sic erit verbum meum, quod egredietur de ore meo:non revertetur ad me vacuum,sed faciet, quaecumque volui,et prosperabitur in his, ad quae misi illud.
ISA|55|12|Quia in laetitia egredieminiet in pace deducemini;montes et colles cantabunt coram vobis laudem,et omnia ligna regionis plaudent manu.
ISA|55|13|Pro vepribus ascendet cupressus,et pro urtica crescet myrtus;et erit Domino in gloriam,in signum aeternum, quod non auferetur.
ISA|56|1|Haec dicit Dominus: Custodite iudicium et faciteiustitiam,quia iuxta est salus mea, ut veniat,et iustitia mea, ut reveletur ".
ISA|56|2|Beatus vir, qui facit hoc,et filius hominis, qui apprehendit istud,custodiens sabbatum, ne polluat illud,custodiens manum suam, ne faciat omne malum.
ISA|56|3|Et non dicat filius advenae, qui adhaeret Domino,dicens: " Separatione dividet me Dominus a populo suo ".Et non dicat eunuchus: Ecce, ego lignum aridum ".
ISA|56|4|Quia haec dicit Dominus eunuchis: Qui custodierint sabbata meaet elegerint, quae ego volui,et tenuerint foedus meum,
ISA|56|5|dabo eis in domo mea et in muris meislocum et nomen melius a filiis et filiabus:nomen sempiternum dabo eis,quod non peribit.
ISA|56|6|Et filios advenae, qui adhaerent Domino,ut colant eum,ut diligant nomen Domini,ut sint ei in servos,omnes custodientes sabbatum, ne polluant illud,et tenentes foedus meum,
ISA|56|7|adducam eos in montem sanctum meumet laetificabo eos in domo orationis meae:holocausta eorum et victimae eorumplacebunt mihi super altari meo,quia domus mea domus orationisvocabitur cunctis populis ".
ISA|56|8|Ait Dominus Deus, qui congregat dispersos Israel: Adhuc congregabo ad eum praeter congregatos eius ".
ISA|56|9|Omnes bestiae agri, venite ad devorandum,universae bestiae saltus.
ISA|56|10|Speculatores eius caeci, omnes nescierunt;universi sunt canes muti non valentes latrare,insanientes, cubantes, amantes soporem;
ISA|56|11|et canes voraces nescierunt saturitatem,ipsi pastores ignoraverunt intellegentiam:omnes in viam suam declinaverunt,unusquisque ad avaritiam suam,a summo usque ad novissimum.
ISA|56|12|" Venite, sumam vinum, et impleamur ebrietate;et cras erit sicut hodieet multo amplius ".
ISA|57|1|Iustus perit, et non est qui recogitet in corde suo;et viri misericordiae colliguntur,tamen non est qui intellegat:a facie enim malitiae collectus est iustus.
ISA|57|2|In pacem ingreditur, requiescit in cubili suo,qui ambulat in directione sua.
ISA|57|3|Vos autem accedite huc, filii auguratricis,semen adulteri et fornicariae.
ISA|57|4|Super quem luditis?Super quem dilatatis os et eicitis linguam?Numquid non vos filii scelesti, semen mendax,
ISA|57|5|qui exardescitis in terebinthissubter omne lignum frondosum,immolantes parvulos in vallibussubter scissuras petrarum?
ISA|57|6|In partibus vallis pars tua,hae sunt sors tua;et ipsis effundisti libamen, obtulisti sacrificium.Numquid super his consolabor?
ISA|57|7|Super montem excelsum et sublimem posuisti cubile tuum,et illuc ascendisti, ut immolares hostias.
ISA|57|8|Et post ostium et postem posuisti memoriale tuum;nam longe a me discooperuisti et ascendisti,dilatasti cubile tuum,et pepigisti cum eis foedus;dilexisti stratum eorum, manum respexisti.
ISA|57|9|Et ingressa es ad regem cum unguentoet multiplicasti pigmenta tua;misisti legatos tuos proculet humiliata es usque ad inferos.
ISA|57|10|In multitudine viae tuae laborasti;non dixisti: " Vanum est! ".Vitam manus tuae invenisti,propterea non aegrotasti.
ISA|57|11|Pro quo sollicita timuisti,quia mentita es et mei non es recordataneque cogitasti in corde tuo?Nonne, quia ego tacui et longo tempore,me non times?
ISA|57|12|Ego annuntiabo iustitiam tuamet opera tua, quae non proderunt tibi.
ISA|57|13|Cum clamaveris, liberent te lucra tua;et omnia illa auferet ventus, tollet aura.Qui autem fiduciam habet in me, hereditabit terramet possidebit montem sanctum meum.
ISA|57|14|Et dicent: " Sternite, sternite,parate viam, auferte offendicula de via populi mei ".
ISA|57|15|Quia haec dicit Excelsus et Sublimis,habitans aeternitatem, et sanctum nomen eius: Excelsus et sanctus habitoet cum contrito et humili spiritu,ut vivificem spiritum humiliumet vivificem cor contritorum.
ISA|57|16|Non enim in sempiternum litigaboneque usque ad finem irascar,quia spiritus a facie mea deficeret,halitus, quem ego feci.
ISA|57|17|Propter iniquitatem avaritiae eius iratus sum et percussi eum,abscondi faciem meam et indignatus sum;et abiit vagus in via cordis sui.
ISA|57|18|Vias eius vidi et sanabo eum et reducam eumet reddam consolationes ipsi et lugentibus eius.
ISA|57|19|Creo fructum labiorum pacem;pacem ei, qui longe est et qui prope, dixit Dominus,et sanabo eum ".
ISA|57|20|Impii autem quasi mare fervens,quod quiescere non potest,et redundant fluctus eius in limum et lutum.
ISA|57|21|Non est pax impiis, dicit Deus meus.
ISA|58|1|Clama fortiter, ne cesses;quasi tuba exalta vocem tuamet annuntia populo meo scelera eorumet domui Iacob peccata eorum.
ISA|58|2|Me etenim de die in diem quaerunt et scire vias meas volunt,quasi gens, quae iustitiam feceritet iudicium Dei sui non dereliquerit.Rogant me iudicia iustitiae,appropinquare Deum volunt.
ISA|58|3|" Quare ieiunavimus, et non aspexisti,humiliavimus animam nostram, et nescisti? ".Ecce, in die ieiunii vestri agitis negotiaet omnes operarios vestros opprimitis.
ISA|58|4|Ecce, ad lites et contentiones ieiunatiset percutitis pugno impie.Nolite ieiunare sicut hodie,ut audiatur in excelso clamor vester.
ISA|58|5|Numquid tale est ieiunium, quod elegi,dies, quo homo affligit animam suam?Numquid contorquere quasi iuncum caput suumet saccum et cinerem sternere?Numquid istud vocabis ieiuniumet diem acceptabilem Domino?
ISA|58|6|Nonne hoc est ieiunium, quod elegi:dissolvere vincula iniqua,solvere funes iugi,dimittere eos, qui confracti sunt, liberos,et omne iugum dirumpere?
ISA|58|7|Nonne frangere esurienti panem tuum,et egenos, vagos inducere in domum?Cum videris nudum, operi eumet carnem tuam ne despexeris.
ISA|58|8|Tunc erumpet quasi aurora lumen tuum,et sanatio tua citius orietur;et anteibit faciem tuam iustitia tua,et gloria Domini colliget te.
ISA|58|9|Tunc invocabis, et Dominus exaudiet;clamabis, et dicet: " Ecce adsum ".Si abstuleris de medio tui iugumet desieris extendere digitumet loqui iniquitatem;
ISA|58|10|si effuderis esurienti animam tuamet animam afflictam satiaveris,orietur in tenebris lux tua,et caligo tua erit sicut meridies.
ISA|58|11|Et te ducet Dominus semper,et satiabit in locis aridis animam tuamet ossa tua firmabit;et eris quasi hortus irriguuset sicut fons aquarum,cuius non deficient aquae.
ISA|58|12|Et reaedificabit gens tua ruinas antiquas;fundamenta generationis et generationis suscitabis:et vocaberis restitutor ruinarum,instaurator viarum, ut habitentur.
ISA|58|13|Si averteris a sabbato pedem tuum,facere negotia tua in die sancto meo,et vocaveris sabbatum deliciaset diem Domino sacrum gloriosum;et glorificaveris eum relinquens vias tuaset negotia tua et sermones tuos,
ISA|58|14|tunc delectaberis super Domino;et vehi te faciam super altitudines terraeet cibabo te hereditate Iacob patris tui.Os enim Domini locutum est.
ISA|59|1|Ecce non est abbreviata manus Domini,ut salvare nequeat,neque aggravata est auris eius,ut non exaudiat;
ISA|59|2|sed iniquitates vestrae diviseruntinter vos et Deum vestrum,et peccata vestra absconderunt faciem eiusa vobis, ne exaudiret.
ISA|59|3|Manus enim vestrae pollutae sunt sanguine,et digiti vestri iniquitate;labia vestra locuta sunt mendacium,et lingua vestra iniquitatem fatur.
ISA|59|4|Non est qui invocet iustitiam,neque est qui iudicet vere;confidunt in nihilo et loquuntur vanitates:conceperunt laborem et pepererunt iniquitatem.
ISA|59|5|Ova aspidum rumpuntet telas araneae texunt;qui comederit de ovis eorum, morietur,et, quod fractum est, erumpet in regulum.
ISA|59|6|Telae eorum non erunt in vestimentum,neque operientur operibus suis;opera eorum opera iniquitatis,et facinora violentiae in manibus eorum.
ISA|59|7|Pedes eorum ad malum curruntet festinant, ut effundant sanguinem innocentem;cogitationes eorum cogitationes iniquitatis,vastitas et contritio in viis eorum.
ISA|59|8|Viam pacis nescierunt,et non est iudicium in gressibus eorum;semitae eorum incurvatae sunt eis:omnis, qui calcat in eis, ignorat pacem.
ISA|59|9|Propter hoc elongatum est iudicium a nobis,et non apprehendit nos iustitia;exspectamus lucem, et ecce tenebrae,splendorem, et in caligine ambulamus.
ISA|59|10|Palpamus sicut caeci parietemet quasi absque oculis attrectamus;impegimus meridie quasi in crepusculo,inter sanos quasi mortui.
ISA|59|11|Rugimus quasi ursi omneset quasi columbae gementes gemimus;exspectamus iudicium, et non est,salutem, et elongata est a nobis.
ISA|59|12|Multiplicatae sunt enim iniquitates nostrae coram te,et peccata nostra respondent nobis;quia scelera nostra nobiscum,et iniquitates nostras cognovimus:
ISA|59|13|peccare et mentiri contra Dominumet recedere a Deo nostro,loqui violentiam et transgressionem,concipere et murmurare de corde verba mendacii.
ISA|59|14|Et conversum est retrorsum iudicium,et iustitia longe stat,quia corruit in platea veritas,et aequitas non potuit ingredi.
ISA|59|15|Et facta est veritas in oblivionem,et, qui recedit a malo, spoliatur.Et vidit Dominus, et malum apparuit in oculis eius,quia non est iudicium.
ISA|59|16|Et vidit quia non est vir,et aporiatus est, quia non est qui occurrat;et salvavit sibi brachium suum,et iustitia eius ipsa confirmavit eum.
ISA|59|17|Indutus est iustitia ut lorica,et galea salutis in capite eius;indutus est vestimentis ultioniset operuit se zelo quasi pallio.
ISA|59|18|Secundum opera sic retribuet:iram hostibus suis,retributionem inimicis suis,insulis vicem reddet.
ISA|59|19|Et timebunt, qui ab occidente, nomen Domini,et, qui ab ortu solis, gloriam eius,cum venerit quasi fluvius violentus,quem spiritus Domini cogit.
ISA|59|20|Et veniet pro Sion redemptoret eis, qui redeunt ab iniquitate in Iacob,dixit Dominus.
ISA|59|21|Hoc foedus meum cum eis,dixit Dominus: Spiritus meus, qui est super te,et verba mea, quae posui in ore tuo,non recedent de ore tuoet de ore seminis tuiet de ore seminis seminis tui,dixit Dominus, amodo et usque in sempiternum ".
ISA|60|1|Surge, illuminare, quia venit lumen tuum,et gloria Domini super te orta est.
ISA|60|2|Quia ecce tenebrae operient terramet caligo populos;super te autem orietur Dominus,et gloria eius in te videbitur.
ISA|60|3|Et ambulabunt gentes in lumine tuo,et reges in splendore ortus tui.
ISA|60|4|Leva in circuitu oculos tuos et vide:omnes isti congregati sunt, venerunt tibi;filii tui de longe veniunt,et filiae tuae in ulnis gestantur.
ISA|60|5|Tunc videbis et illuminaberis,et palpitabit et dilatabitur cor tuum,quia confluet ad te multitudo maris,fortitudo gentium veniet tibi;
ISA|60|6|inundatio camelorum operiet te,dromedarii Madian et Epha;omnes de Saba venient,aurum et tus deferenteset laudem Domini annuntiantes.
ISA|60|7|Omne pecus Cedar congregabitur tibi,arietes Nabaioth ministrabunt tibi;offerentur super placabili altari meo,et domum gloriae meae glorificabo.
ISA|60|8|Quae sunt istae, quae ut nubes volant,et quasi columbae ad fenestras suas?
ISA|60|9|Me enim insulae exspectabunt,et in principio naves Tharsis,ut adducant filios tuos de longe,argentum eorum et aurum eorum cum eis,nomini Domini Dei tui et Sancto Israel,quia glorificavit te.
ISA|60|10|Et aedificabunt filii peregrinorum muros tuos,et reges eorum ministrabunt tibi;in indignatione enim mea percussi te,sed in beneplacito meo misertus sum tui.
ISA|60|11|Et aperientur portae tuae iugiter,die ac nocte non claudentur,ut afferatur ad te fortitudo gentium,et reges earum adducantur.
ISA|60|12|Gens enim et regnum, quae non servierint tibi, peribunt,et gentes vastitate vastabuntur.
ISA|60|13|Gloria Libani ad te veniet,cupressus, ulmus et abies simul,ad ornandum locum sanctuarii mei;et locum pedum meorum glorificabo.
ISA|60|14|Et venient ad te curvi filii eorum, qui humiliaverunt te,et adorabunt vestigia pedum tuorum omnes, qui detrahebant tibi, et vocabunt te Civitatem Domini,Sion Sancti Israel.
ISA|60|15|Pro eo quod fuisti derelicta et odio habita,et non erat qui per te transiret,ponam te in superbiam saeculorum,gaudium in generationem et generationem;
ISA|60|16|et suges lac gentiumet mamilla regum lactaberiset scies quia ego Dominus salvator tuus,et redemptor tuus Fortis Iacob.
ISA|60|17|Pro aere afferam aurumet pro ferro afferam argentumet pro lignis aeset pro lapidibus ferrum;et ponam custodes tuos pacemet praepositos tuos iustitiam.
ISA|60|18|Non audietur ultra violentia in terra tua,vastitas et contritio in terminis tuis;et vocabis Salutem muros tuoset portas tuas Laudem.
ISA|60|19|Non erit tibi amplius sol ad lucendum per diem,nec splendor lunae illuminabit te,sed erit tibi Dominus in lucem sempiternam,et Deus tuus in gloriam tuam.
ISA|60|20|Non occidet ultra sol tuus,et luna tua non minuetur,quia erit tibi Dominus in lucem sempiternam,et complebuntur dies luctus tui.
ISA|60|21|Populus autem tuus omnes iusti;in perpetuum hereditabunt terram,germen plantationis meae,opus manus meae ad glorificandum.
ISA|60|22|Minimus erit in mille,et parvulus in gentem fortem.Ego Dominus in tempore eius subito faciam istud.
ISA|61|1|Spiritus Domini Dei super me,eo quod unxerit Dominus me;ad annuntiandum laeta mansuetis misit me,ut mederer contritis cordeet praedicarem captivis liberationemet clausis apertionem;
ISA|61|2|ut praedicarem annum placabilem Dominoet diem ultionis Deo nostro;ut consolarer omnes lugentes,
ISA|61|3|ut ponerem lugentibus Sionet darem eis coronam pro cinere,oleum gaudii pro luctu,pallium laudis pro spiritu maeroris.Et vocabuntur Terebinthi iustitiae,plantatio Domini ad glorificandum.
ISA|61|4|Et aedificabunt deserta a saeculoet ruinas antiquas erigentet instaurabunt civitates desertas,dissipatas in generatione et generatione.
ISA|61|5|Et stabunt alieni et pascent pecora vestra,et filii peregrinorum agricolae et vinitores vestri erunt;
ISA|61|6|vos autem Sacerdotes Domini vocabimini,Ministri Dei nostri dicetur vobis;fortitudinem gentium comedetiset in gloria earum superbietis.
ISA|61|7|Pro confusione eorum dupliciet ignominia laudabunt partem suam;propterea in terra sua duplicia possidebunt,laetitia sempiterna erit eis.
ISA|61|8|Quia ego Dominus diligens iudicium,odio habens rapinam et iniquitatem;et dabo opus eorum in veritateet foedus perpetuum feriam eis.
ISA|61|9|Et scietur in gentibus semen eorum,et germen eorum in medio populorum;omnes, qui viderint eos, cognoscent illos,quia isti sunt semen, cui benedixit Dominus.
ISA|61|10|Gaudens gaudebo in Domino,et exsultabit anima mea in Deo meo,quia induit me vestimentis salutiset indumento iustitiae circumdedit me,quasi sponsum decoratum coronaet quasi sponsam ornatam monilibus suis.
ISA|61|11|Sicut enim terra profert germen suum,et sicut hortus semen suum germinat,sic Dominus Deus germinabit iustitiamet laudem coram universis gentibus.
ISA|62|1|Propter Sion non taceboet propter Ierusalem nonquiescam,donec egrediatur ut splendor iustitia eius,et salus eius ut lampas accendatur.
ISA|62|2|Et videbunt gentes iustitiam tuam,et cuncti reges gloriam tuam;et vocaberis nomine novo,quod os Domini nominabit.
ISA|62|3|Et eris corona gloriae in manu Domini,et diadema regni in manu Dei tui.
ISA|62|4|Non vocaberis ultra Derelicta,et terra tua non vocabitur amplius Desolata;sed vocaberis Beneplacitum meum in ea,et terra tua Nupta,quia complacuit Domino in te,et terra tua erit nupta.
ISA|62|5|Nam ut iuvenis uxorem ducit virginem,ita ducent te filii tui;ut gaudet sponsus super sponsam,ita gaudebit super te Deus tuus.
ISA|62|6|Super muros tuos, Ierusalem, constitui custodes;tota die et tota nocte, in perpetuo non tacebunt.Qui commonetis Dominum, ne taceatis
ISA|62|7|et ne detis silentium ei,donec stabiliat et donec ponat Ierusalemlaudem in terra.
ISA|62|8|Iuravit Dominus in dextera suaet in brachio fortitudinis suae: Non dabo triticum tuum ultracibum inimicis tuis,neque bibent filii alienivinum tuum, in quo laborasti.
ISA|62|9|Quia, qui collegerint illud, comedentet laudabunt Dominum;et, qui vindemiam fecerint,illud bibent in atriis sanctuarii mei.
ISA|62|10|Transite, transite per portas,parate viam populo.Sternite, sternite semitam, eligite lapides,elevate signum ad populos ".
ISA|62|11|Ecce Dominus auditum fecit in extremis terrae: Dicite filiae Sion:Ecce salus tua venit,ecce merces eius cum eo,et praemium eius coram illo.
ISA|62|12|Et vocabunt eos Populus sanctus,Redempti a Domino;tu autem vocaberis Quaesita,Civitas non derelicta ".
ISA|63|1|" Quis est iste, qui venit de Edom,tinctis vestibus de Bosra?Iste formosus in stola sua,gradiens in multitudine fortitudinis suae ". Sum ego, qui loquor iustitiam,potens ad salvandum ".
ISA|63|2|" Quare ergo rubrum est indumentum tuum,et vestimenta tua sicut calcantis in torculari? ".
ISA|63|3|" Torcular calcavi solus,et de gentibus non erat vir mecum;calcavi eos in furore meoet conculcavi eos in ira mea.Et aspersus est sanguis eorum super vestimenta mea,et omnia indumenta mea inquinavi.
ISA|63|4|Dies enim ultionis in corde meo,annus redemptionis meae venit.
ISA|63|5|Circumspexi, et non erat auxiliator,miratus sum, et non fuit qui adiuvaret;et salvavit mihi brachium meum,et indignatio mea ipsa auxiliata est mihi.
ISA|63|6|Et conculcavi populos in furore meoet contrivi eos in indignatione meaet effudi in terram sanguinem eorum ".
ISA|63|7|Miserationum Domini recordabor,laudum Dominisuper omnibus, quae reddidit nobis Dominus,et super multitudinem bonorum domui Israel,quae largitus est eis secundum misericordias suaset secundum multitudinem miserationum suarum.
ISA|63|8|Et dixit: " Verumtamen populus meus est,filii, qui non deludent ";et factus est eis salvator.
ISA|63|9|In omni tribulatione eorum non legatus neque angelus,sed ipse salvavit eos.In dilectione sua et in indulgentia suaipse redemit eoset sustulit eos et portavit eoscunctis diebus saeculi.
ISA|63|10|Ipsi autem ad iracundiam provocaveruntet afflixerunt spiritum sanctitatis eius;et conversus est eis in inimicumet ipse debellavit eos.
ISA|63|11|Et recordatus est dierum antiquorum,Moysi et populi sui.Ubi est qui eduxit eos de maricum pastore gregis sui?Ubi est qui posuit in medio eiusspiritum sanctitatis suae?
ISA|63|12|Qui adduxit ad dexteram Moysibrachium maiestatis suae,qui scidit aquas ante eos,ut faceret sibi nomen sempiternum,
ISA|63|13|qui deduxit eos per abyssosquasi equum per desertum, et non impingebant?
ISA|63|14|Sicut armentum, quod descendit per vallem,spiritus Domini fecit eos quiescere;sic conduxisti populum tuum,ut faceres tibi nomen gloriae.
ISA|63|15|Attende de caelo et videde habitaculo sancto tuo et gloriae tuae;ubi est zelus tuus et fortitudo tua?Commotio viscerum tuorum et misericordiae tuaesuper me continuerunt se.
ISA|63|16|Tu enim pater noster.Abraham enim nescit nos,et Israel ignorat nos;tu, Domine, pater noster,redemptor noster: a saeculo nomen tuum.
ISA|63|17|Quare errare nos fecisti, Domine, de viis tuis,indurasti cor nostrum, ne timeremus te?Convertere propter servos tuos,tribus hereditatis tuae.
ISA|63|18|Brevi tempore hereditaverunt populum sanctum tuum,hostes nostri conculcaverunt sanctuarium tuum.
ISA|63|19|Facti sumus a saeculo,cum non dominareris nostri,neque invocaretur nomen tuum super nos.Utinam dirumperes caelos et descenderes!A facie tua montes defluerent.
ISA|64|1|Sicut ignis succendit sarmenta,aquam ebullire facit ignis,ut notum facias nomen tuum inimicis tuis,a facie tua gentes turbentur,
ISA|64|2|cum feceris mirabilia,quae non sperabamus.Descendisti, et a facie tua montes defluxerunt.
ISA|64|3|A saeculo non audierunt, neque aures perceperunt;oculus non vidit Deum, absque te,qui operaretur pro sperantibus in eum.
ISA|64|4|Occurris laetanti, facienti iustitiamet his, qui in viis tuis recordantur tui.Ecce tu iratus es, et peccavimus;in ipsis a saeculo nos salvabimur.
ISA|64|5|Et facti sumus ut immundus omnes nos,et quasi pannus inquinatus universae iustitiae nostrae;et marcuimus quasi folium universi,et iniquitates nostrae quasi ventus abstulerunt nos.
ISA|64|6|Non est qui invocet nomen tuum,qui consurgat et adhaereat tibi,quia abscondisti faciem tuam a nobiset dissolvisti nos in manu iniquitatis nostrae.
ISA|64|7|Et nunc, Domine, pater noster es tu,nos vero lutum; et fictor noster tu,et opera manuum tuarum omnes nos.
ISA|64|8|Ne irascaris, Domine, nimiset ne ultra memineris iniquitatis;ecce, respice: populus tuus omnes nos.
ISA|64|9|Urbes sanctitatis tuae factae sunt in desertum,Sion deserta facta est,Ierusalem desolata est.
ISA|64|10|Domus sanctitatis nostrae et gloriae nostrae,ubi laudaverunt te patres nostri,facta est in exustionem ignis,et omnia desiderabilia nostra versa sunt in ruinas.
ISA|64|11|Numquid super his continebis te, Domine,tacebis et affliges nos vehementer?
ISA|65|1|" Quaesitus sum ab his, qui non consulebant me,inventus sum ab his, qui non quaerebant me.Dixi: "Ecce ego, ecce ego!"ad gentem, quae non invocabat nomen meum.
ISA|65|2|Expandi manus meas tota diead populum rebellem,qui graditur in via non bonapost cogitationes suas;
ISA|65|3|populus, qui ad iracundiam provocat meante faciem meam semper,qui immolant in hortiset sacrificant super lateres,
ISA|65|4|qui morantur in sepulcriset in locis occultis pernoctant,qui comedunt carnem suillamet ius abominabile in vasis eorum,
ISA|65|5|qui dicunt: "Recede!Non appropinques mihi, quia sanctificarem te".Isti fumus sunt in naribus meis,ignis ardens tota die.
ISA|65|6|Ecce scriptum est coram me;non tacebo, sed retribuam,et retribuam in sinum eorum
ISA|65|7|iniquitates vestras et iniquitates patrum vestrorumsimul, dicit Dominus,qui sacrificaverunt super monteset super colles exprobraverunt mihi;et remetiar opus eorum primoin sinu eorum ".
ISA|65|8|Haec dicit Dominus: Quomodo si inveniatur mustum in botroet dicatur: "Ne dissipes illud,quoniam benedictio est in eo",sic faciam propter servos meos,ut non disperdam totum.
ISA|65|9|Et educam de Iacob semenet de Iuda possidentem montes meos;et hereditabunt terram electi mei,et servi mei habitabunt ibi.
ISA|65|10|Et erit Saron in pascua gregum,et vallis Achor in cubile armentorumpopulo meo, qui quaesierunt me.
ISA|65|11|Vos autem, qui derelinquitis Dominum,qui obliviscimini montem sanctum meum,qui ponitis Gad mensamet amphoram impletis Meni,
ISA|65|12|numerabo vos in gladio,et omnes in caede corruetis;pro eo quod vocavi, et non respondistis,locutus sum, et non audistis,sed fecistis malum in oculis meiset, quod displicet mihi, elegistis ".
ISA|65|13|Propter hoc haec dicit Dominus Deus: Ecce servi mei comedent,et vos esurietis;ecce servi mei bibent,et vos sitietis;ecce servi mei laetabuntur,et vos confundemini;
ISA|65|14|ecce servi mei laudabunt in exsultatione cordis,et vos clamabitis prae dolore cordiset prae contritione spiritus ululabitis.
ISA|65|15|Et relinquetis nomen vestrumin iuramentum electis meis:Interficiat te Dominus Deus";et servos suos vocabit nomine alio.
ISA|65|16|Quicumque benedicit sibi in terra,benedicet sibi in Deo Amen;et, quicumque iurat in terra,iurabit in Deo Amen;quia oblivioni tradentur angustiae priores,et quia abscondentur ab oculis meis.
ISA|65|17|Ecce enim ego creocaelos novos et terram novam,et non erunt in memoria prioraet non ascendent super cor.
ISA|65|18|Sed gaudebunt et exsultabunt usque in sempiternumin his, quae ego creo,quia ecce ego creo Ierusalem exsultationemet populum eius gaudium.
ISA|65|19|Et exsultabo in Ierusalemet gaudebo in populo meo,et non audietur in ea ultravox fletus et vox clamoris.
ISA|65|20|Non erit ibi amplius infans dierumet senex, qui non impleat dies suos.Quoniam puer erit,qui centenarius moriatur;et, qui non attingat centum annos,maledictus erit.
ISA|65|21|Et aedificabunt domos et habitabuntet plantabunt vineas et comedent fructus earum.
ISA|65|22|Non aedificabunt, ut alius habitet,non plantabunt, ut alius comedat:secundum enim dies ligni erunt dies populi mei,et operibus manuum suarum diu fruentur electi mei.
ISA|65|23|Non laborabunt frustraneque generabunt in interitum repentinum,quia semen benedictorum erunt Domini,et nepotes eorum cum eis.
ISA|65|24|Eritque: antequam clament, ego respondebo;adhuc illis loquentibus, ego exaudiam.
ISA|65|25|Lupus et agnus pascentur simul,et leo sicut bos comedet paleas,et serpenti pulvis panis eius.Non nocebunt neque occidentin omni monte sancto meo ",dicit Dominus.
ISA|66|1|Haec dicit Dominus: Caelum thronus meus,terra autem scabellum pedum meorum.Quae ista domus, quam aedificabitis mihi,et quis iste locus quietis meae?
ISA|66|2|Omnia haec manus mea fecit,et mea sunt universa ista,dicit Dominus.Ad hunc autem respiciam,ad pauperculum et contritum spirituet trementem sermones meos.
ISA|66|3|Qui immolat bovem, interficit virum;qui sacrificat ovem, excerebrat canem;qui offert oblationem, idemque sanguinem suillum;qui adolet incensum, benedicit idolo.Sicut isti elegerunt vias suas,et in abominationibus suis anima eorum delectatur,
ISA|66|4|sic ego eligam malam sortem eorumet, quae timebant, adducam eis;quia vocavi, et non erat qui responderet,locutus sum, et non audieruntfeceruntque malum in oculis meiset, quod displicet mihi, elegerunt ".
ISA|66|5|Audite verbum Domini,qui tremitis ad verbum eius.Dixerunt fratres vestri odientes voset abicientes vos propter nomen meum: Gloriam suam manifestet Dominus,ut videamus laetitiam vestram";ipsi autem confundentur.
ISA|66|6|Vox clamoris de civitate,vox de templo,vox Dominireddentis retributionem inimicis suis.
ISA|66|7|Antequam parturiret, peperit;antequam veniret partus eius, peperit masculum.
ISA|66|8|Quis audivit umquam tale?Et quis vidit huic simile?Numquid oritur terra in die una,aut parietur gens in momento?Quia parturivit, iam peperit Sion filios suos.
ISA|66|9|" Numquid aperiam uterum et parere non faciam? ",dicit Dominus. Aut ego, qui parere facio, uterum claudam? ",ait Deus tuus.
ISA|66|10|Laetamini cum Ierusalem et exsultate in ea,omnes, qui diligitis eam;gaudete cum ea gaudio,universi, qui lugebatis super eam,
ISA|66|11|ut sugatis et repleaminiab ubere consolationis eius,ut mulgeatis et deliciis affluatisex uberibus gloriae eius.
ISA|66|12|Quia haec dicit Dominus: Ecce ego dirigam ad eam quasi fluvium pacemet quasi torrentem inundantem gloriam gentium.Sugetis, in ulnis portabimini,et super genua blandientur vobis.
ISA|66|13|Quomodo si quem mater consolatur,ita ego consolabor vos;et in Ierusalem consolabimini.
ISA|66|14|Videbitis, et gaudebit cor vestrum,et ossa vestra quasi herba germinabunt,et manifestabitur manus Domini in servis eius,et indignabitur inimicis suis.
ISA|66|15|Quia ecce Dominus in igne veniet,et quasi turbo quadrigae eius,reddere in indignatione furorem suumet increpationem suam in flamma ignis;
ISA|66|16|quia in igne Dominus diiudicabitet in gladio suo omnem carnem,et multiplicabuntur interfecti a Domino.
ISA|66|17|Qui sanctificantur et purificantur, ut ingredianturin hortos post aliquem stantem in medio,qui comedunt carnem suillamet abominationem et murem,simul consumentur,dicit Dominus.
ISA|66|18|Ego autem cognoscens opera eorum et cogitationes eorum veniam, ut congregem omnes gentes et linguas; et venient et videbunt gloriam meam.
ISA|66|19|Et ponam in eis signum et mittam ex eis, qui salvati fuerint, ad gentes in Tharsis, Phut, Lud, Mosoch, Ros, Thubal et Iavan, ad insulas longinquas, ad eos, qui non audierunt de me et non viderunt gloriam meam, et annuntiabunt gloriam meam gentibus;
ISA|66|20|et adducent omnes fratres vestros de cunctis gentibus oblationem Domino, in equis et in quadrigis et in lecticis et in mulis et in dromedariis, ad montem sanctum meum Ierusalem, dicit Dominus: quomodo si inferant filii Israel oblationem in vase mundo in domum Domini.
ISA|66|21|Et assumam ex eis in sacerdotes et Levitas, dicit Dominus.
ISA|66|22|Quia sicut caeli noviet terra nova, quae ego faciam,stabunt coram me,dicit Dominus,sic stabit semen vestrum et nomen vestrum.
ISA|66|23|Et erit: unoquoque novilunioet quovis sabbatoveniet omnis caro, ut adoret coram facie mea,dicit Dominus.
ISA|66|24|Et egredientur et videbunt cadavera virorum,qui praevaricati sunt in me;nam vermis eorum non morietur,et ignis eorum non exstinguetur,et erunt abominationi omni carni ".
