2THESS|1|1|保罗 、 西拉 和 提摩太 写信给 帖撒罗尼迦 、在我们的父上帝与主耶稣基督里的教会。
2THESS|1|2|愿恩惠、平安 从我们的 父上帝和主耶稣基督归给你们！
2THESS|1|3|弟兄们，我们该常常为你们感谢上帝，这本是合宜的；因为你们的信心格外增长，你们众人彼此相爱的心也都增加。
2THESS|1|4|所以，我们在上帝的各教会里为你们夸耀，因为你们在所受的一切压迫患难中仍牢守着耐心和信心。
2THESS|1|5|这正是上帝公义判断的明证，使你们配得上他的国，你们就是为这国受苦。
2THESS|1|6|既然上帝是公义的，他必以患难报复那加患难给你们的人，
2THESS|1|7|也必使你们这受患难的人与我们同得平安。那时，主耶稣同他有权能的天使从天上在火焰中显现，要报应那些不认识上帝和不听从我们的主耶稣福音的人。
2THESS|1|8|
2THESS|1|9|他们要受惩罚，永远沉沦，与主的面和他权能的荣光隔绝。
2THESS|1|10|这正是主再来，要在他圣徒的身上得荣耀，就是要使一切信的人感到惊讶的那日子，因为你们信了我们对你们作的见证。
2THESS|1|11|为此，我们常为你们祷告，愿我们的上帝看你们与他的呼召相配，又用大能成就你们一切良善的美意和因信心所做的工作，
2THESS|1|12|使我们主耶稣的名，照着我们的上帝和主耶稣基督的恩，在你们身上得荣耀，你们也在他身上得荣耀。
2THESS|2|1|弟兄们，关于我们主耶稣基督的来临和我们到他那里聚集，我劝你们：
2THESS|2|2|无论藉着灵，藉着言语，藉着冒我的名写的书信，说主的日子已经到了，不要轻易动心，也不要惊慌。
2THESS|2|3|不要让任何人用什么法子欺骗你们，因为那日子以前必有叛教的事，并有那不法的人，那沉沦之子出现。
2THESS|2|4|那抵挡者高抬自己超过一切称为神明的，和一切受人敬拜的，甚至坐在上帝的殿里，自称为上帝。
2THESS|2|5|我还在你们那里的时候曾把这些事告诉你们，你们不记得吗？
2THESS|2|6|现在你们也知道那拦阻他的是什么，为要使他到了时机才出现。
2THESS|2|7|因为那不法的隐秘已经运作，只是现在有一个阻挡的，要等到那阻挡的被除去才会发作，
2THESS|2|8|那时这不法的人必出现，主耶稣 要用口中的气灭绝他，以自己来临的光辉摧毁他。
2THESS|2|9|这不法的人来，是靠撒但的运作，行各样的异能、神迹和一切虚假的奇事，
2THESS|2|10|并且在那沉沦的人身上行各样不义的诡诈，因为他们不领受爱真理的心，好让他们得救。
2THESS|2|11|故此，上帝就给他们一个引发错误的心，叫他们信从虚谎，
2THESS|2|12|使一切不信真理、倒喜爱不义的人都被定罪。
2THESS|2|13|主所爱的弟兄们哪，我们本该常为你们感谢上帝，因为他拣选你们为初熟的果子 ，使你们因信真道，又蒙圣灵感化成圣，得到拯救。
2THESS|2|14|为此，上帝藉着我们所传的福音呼召你们，好得着我们主耶稣基督的荣光。
2THESS|2|15|所以，弟兄们，你们要站立得稳，凡所领受的教导，无论是我们口传的，是信上写的，都要坚守。
2THESS|2|16|愿我们主耶稣基督自己，和那爱我们、开恩将永远的安慰及美好的盼望赐给我们的父上帝，
2THESS|2|17|安慰你们的心，并且在一切善行善言上坚固你们！
2THESS|3|1|末了，弟兄们，请你们为我们祷告，好让主的道快快传开，得着荣耀，正如在你们中间一样，
2THESS|3|2|也让我们能脱离无理和邪恶人的手，因为不是人人都有信仰。
2THESS|3|3|但主是信实的，他要坚固你们，保护你们脱离那邪恶者。
2THESS|3|4|我们靠主对你们有信心，你们现在遵行，以后也必遵行我们所吩咐的。
2THESS|3|5|愿主引导你们的心去爱上帝，并学基督的忍耐！
2THESS|3|6|弟兄们，我们奉主耶稣基督的名吩咐你们，凡有弟兄懒散，不遵守我们所传授的教导，要远离他。
2THESS|3|7|你们自己知道该怎样效法我们。因为我们在你们当中从未懒散过，
2THESS|3|8|也从未白吃人的饭，倒是辛苦劳碌，昼夜做工，免得使你们中间有人受累。
2THESS|3|9|这并不是因我们没有权柄，而是要给你们作榜样，好让你们效法我们。
2THESS|3|10|我们在你们那里的时候曾吩咐你们，说若有人不肯做工，就不可吃饭。
2THESS|3|11|因为我们听说，在你们中间有人懒散，什么工都不做，反倒专管闲事。
2THESS|3|12|我们靠主耶稣基督吩咐并劝戒这样的人，要安分做工，自食其力。
2THESS|3|13|弟兄们，你们行善不可丧志。
2THESS|3|14|若有人不听从我们这信上的话，要把他记下，不和他交往，使他自觉羞愧；
2THESS|3|15|但不要把他当仇人，要劝他如劝弟兄。
2THESS|3|16|愿赐平安 的主随时随事亲自赐给你们平安！愿主与你们众人同在！
2THESS|3|17|我— 保罗 亲笔向你们问安。凡我的信都以此为记，我的笔迹就是这样。
2THESS|3|18|愿我们主耶稣基督的恩惠与你们众人同在！
