NAH|1|1|onus Nineve liber visionis Naum Helcesei
NAH|1|2|Deus aemulator et ulciscens Dominus ulciscens Dominus et habens furorem ulciscens Dominus in hostes suos et irascens ipse inimicis suis
NAH|1|3|Dominus patiens et magnus fortitudine et mundans non faciet innocentem Dominus in tempestate et turbine viae eius et nebulae pulvis pedum eius
NAH|1|4|increpans mare et exsiccans illud et omnia flumina ad desertum deducens infirmatus est Basan et Carmelus et flos Libani elanguit
NAH|1|5|montes commoti sunt ab eo et colles adsolati sunt et contremuit terra a facie eius et orbis et omnes habitantes in eo
NAH|1|6|ante faciem indignationis eius quis stabit et quis resistet in ira furoris eius indignatio eius effusa est ut ignis et petrae dissolutae sunt ab eo
NAH|1|7|bonus Dominus et confortans in die tribulationis et sciens sperantes in se
NAH|1|8|et in diluvio praetereunte consummationem faciet loci eius et inimicos eius persequentur tenebrae
NAH|1|9|quid cogitatis contra Dominum consummationem ipse faciet non consurget duplex tribulatio
NAH|1|10|quia sicut spinae se invicem conplectuntur sic convivium eorum pariter potantium consumentur quasi stipula ariditate plena
NAH|1|11|ex te exivit cogitans contra Dominum malitiam mente pertractans praevaricationem
NAH|1|12|haec dicit Dominus si perfecti fuerint et ita plures sic quoque adtondentur et pertransibit adflixi te et non adfligam te ultra
NAH|1|13|et nunc conteram virgam eius de dorso tuo et vincula tua disrumpam
NAH|1|14|et praecipiet super te Dominus non seminabitur ex nomine tuo amplius de domo Dei tui interficiam sculptile et conflatile ponam sepulchrum tuum quia inhonoratus es
NAH|1|15|ecce super montes pedes evangelizantis et adnuntiantis pacem celebra Iuda festivitates tuas et redde vota tua quia non adiciet ultra ut pertranseat in te Belial universus interiit
NAH|2|1|ascendit qui dispergat coram te qui custodit obsidionem contemplare viam conforta lumbos robora virtutem valde
NAH|2|2|quia reddidit Dominus superbiam Iacob sicut superbiam Israhel quia vastatores dissipaverunt eos et propagines eorum corruperunt
NAH|2|3|clypeus fortium eius ignitus viri exercitus in coccineis igneae habenae currus in die praeparationis eius et agitatores consopiti sunt
NAH|2|4|in itineribus conturbati sunt quadrigae conlisae sunt in plateis aspectus eorum quasi lampades quasi fulgura discurrentia
NAH|2|5|recordabitur fortium suorum ruent in itineribus suis velociter ascendent muros eius et praeparabitur umbraculum
NAH|2|6|portae fluviorum apertae sunt et templum ad solum dirutum
NAH|2|7|et miles captivus abductus est et ancillae eius minabantur gementes ut columbae murmurantes in cordibus suis
NAH|2|8|et Nineve quasi piscina aquarum aquae eius ipsi vero fugerunt state state et non est qui revertatur
NAH|2|9|diripite argentum diripite aurum et non est finis divitiarum ex omnibus vasis desiderabilibus
NAH|2|10|dissipata et scissa et dilacerata et cor tabescens et dissolutio geniculorum et defectio in cunctis renibus et facies omnium sicut nigredo ollae
NAH|2|11|ubi est habitaculum leonum et pascua catulorum leonum ad quam ivit leo ut ingrederetur illuc catulus leonis et non est qui exterreat
NAH|2|12|leo cepit sufficienter catulis suis et necavit leaenis suis et implevit praeda speluncas suas et cubile suum rapina
NAH|2|13|ecce ego ad te dicit Dominus exercituum et succendam usque ad fumum quadrigas eius et leunculos tuos comedet gladius et exterminabo de terra praedam tuam et non audietur ultra vox nuntiorum tuorum
NAH|3|1|vae civitas sanguinum universa mendacii dilaceratione plena non recedet a te rapina
NAH|3|2|vox flagelli et vox impetus rotae et equi frementis et quadrigae ferventis equitis ascendentis
NAH|3|3|et micantis gladii et fulgurantis hastae et multitudinis interfectae et gravis ruinae nec est finis cadaverum et corruent in corporibus suis
NAH|3|4|propter multitudinem fornicationum meretricis speciosae et gratae et habentis maleficia quae vendidit gentes in fornicationibus suis et familias in maleficiis suis
NAH|3|5|ecce ego ad te dicit Dominus exercituum et revelabo pudenda tua in facie tua et ostendam gentibus nuditatem tuam et regnis ignominiam tuam
NAH|3|6|et proiciam super te abominationes et contumeliis te adficiam et ponam te in exemplum
NAH|3|7|et erit omnis qui viderit te resiliet a te et dicet vastata est Nineve quis commovebit super te caput unde quaeram consolatorem tibi
NAH|3|8|numquid melior es ab Alexandria populorum quae habitat in fluminibus aqua in circuitu eius cuius divitiae mare aquae muri eius
NAH|3|9|Aethiopia fortitudo et Aegyptus et non est finis Africa et Lybies fuerunt in auxilio tuo
NAH|3|10|sed et ipsa in transmigrationem ducta est in captivitatem parvuli eius elisi sunt in capite omnium viarum et super inclitos eius miserunt sortem et omnes optimates eius confixi sunt in conpedibus
NAH|3|11|et tu ergo inebriaberis eris despecta et tu quaeres auxilium ab inimico
NAH|3|12|omnes munitiones tuae sicuti ficus cum grossis suis si concussae fuerint cadent in os comedentis
NAH|3|13|ecce populus tuus mulieres in medio tui inimicis tuis adapertione pandentur portae terrae tuae devorabit ignis vectes tuos
NAH|3|14|aquam propter obsidionem hauri tibi extrue munitiones tuas intra in lutum et calca subigens tene laterem
NAH|3|15|ibi comedet te ignis peribis gladio devorabit te ut bruchus congregare ut bruchus multiplicare ut lucusta
NAH|3|16|plures fecisti negotiationes tuas quam stellae sunt caeli bruchus expansus est et avolavit
NAH|3|17|custodes tui quasi lucustae et parvuli tui quasi lucustae lucustarum quae considunt in sepibus in die frigoris sol ortus est et avolaverunt et non est cognitus locus earum ubi fuerint
NAH|3|18|dormitaverunt pastores tui rex Assur sepelientur principes tui latitavit populus tuus in montibus et non est qui congreget
NAH|3|19|non est obscura contritio tua pessima est plaga tua omnes qui audierunt auditionem tuam conpresserunt manum super te quia super quem non transiit malitia tua semper
