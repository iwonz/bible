ZEPH|1|1|Verbum Domini, quod factum est ad Sophoniam filium Chusi filii Godoliae filii Amariae filii Ezechiae, in diebus Iosiae filii Amon regis Iudae.
ZEPH|1|2|" Auferens auferam omniaa facie terrae,dicit Dominus,
ZEPH|1|3|auferam hominem et pecus,auferam volatile caeliet pisces maris.Et ruinae impiorum erunt;et disperdam homines a facie terrae,dicit Dominus.
ZEPH|1|4|Et extendam manum meam super Iudamet super omnes habitantes Ierusalem;et disperdam de loco hoc reliquias Baalet nomina aedituorum cum sacerdotibus
ZEPH|1|5|et eos, qui adorant super tectamilitiam caeliet adorant et iurant in Dominoet iurant in Melchom,
ZEPH|1|6|et qui avertuntur de post tergum Domini,et qui non quaerunt Dominum nec investigant eum ".
ZEPH|1|7|Silete a facie Domini Dei,quia iuxta est dies Domini;quia praeparavit Dominus hostiam,sanctificavit vocatos suos.
ZEPH|1|8|" Et erit in die hostiae Domini:visitabo super principeset super filios regiset super omnes, qui induti suntveste peregrina;
ZEPH|1|9|et visitabo super omnem,qui arroganter ingreditur super limen in die illa,qui complent domum domini suiiniquitate et dolo.
ZEPH|1|10|Et erit in die illa,dicit Dominus,vox clamoris a porta Piscium,et ululatus ab urbe Nova,et contritio magna a collibus.
ZEPH|1|11|Ululate, habitatores Pilae,quia interiit omnis populus Chanaan,disperierunt omnes involuti argento.
ZEPH|1|12|Et erit in tempore illo:scrutabor Ierusalem in lucerniset visitabo super virosdefixos in faecibus suis,qui dicunt in cordibus suis:Non faciet bene Dominuset non faciet male".
ZEPH|1|13|Et erunt opes eorum in direptionem,et domus eorum in desertum;et aedificabunt domoset non habitabunt,et plantabunt vineaset non bibent vinum earum ".
ZEPH|1|14|Iuxta est dies Domini magnus,iuxta et velox nimis;vox diei Domini amara,tribulabitur ibi fortis.
ZEPH|1|15|Dies irae dies illa,dies tribulationis et angustiae,dies vastitatis et desolationis,dies tenebrarum et caliginis,dies nebulae et turbinis,
ZEPH|1|16|dies tubae et clangorissuper civitates munitaset super angulos excelsos.
ZEPH|1|17|Et tribulabo homines,et ambulabunt ut caeci,quia Domino peccaverunt;et effundetur sanguis eorum sicut humus,et viscera eorum sicut stercora.
ZEPH|1|18|Sed et argentum eorum et aurum eorumnon poterit liberare eosin die irae Domini;in igne zeli eiusdevorabitur omnis terra,quia consummationem cum festinatione facietcunctis habitantibus terram.
ZEPH|2|1|Convenite, congregamini,gens non amabilis,
ZEPH|2|2|priusquam dispergaminiquasi pulvis transeuntes,antequam veniat super vosira furoris Domini,antequam veniat super vosdies furoris Domini.
ZEPH|2|3|Quaerite Dominum,omnes mansueti terrae,qui iudicium eius estis operati;quaerite iustitiam, quaerite mansuetudinem,si quomodo abscondaminiin die furoris Domini.
ZEPH|2|4|Quia Gaza deserta erit,et Ascalon desolata,Azotum in meridie eicient,et Accaron eradicabitur.
ZEPH|2|5|Vae, qui habitatis funiculum maris, gens Cretensium!Verbum Domini super vos,Chanaan, terra Philisthinorum: Disperdam te,ita ut non sit inhabitator ".
ZEPH|2|6|Et erit funiculus marisrequies pastorum et caulae pecorum.
ZEPH|2|7|Et erit funiculus marisreliquiis domus Iudae:ibi pascentur,in domibus Ascalonis ad vesperam requiescent,quia visitabit eos Dominus Deus eorumet convertet sortem eorum.
ZEPH|2|8|" Audivi opprobrium Moabet blasphemias filiorum Ammon, qui exprobraverunt populo meoet magnificati sunt super terminos eorum.
ZEPH|2|9|Propterea vivo ego,dicit Dominus exercituum, Deus Israel,quia Moab ut Sodoma erit,et filii Ammon quasi Gomorra,possessio spinarum et acervi saliset desertum usque in aeternum;reliquiae populi mei diripient eos,et residui gentis meae possidebunt illos ".
ZEPH|2|10|Hoc eis eveniet pro superbia sua, quia blasphemaverunt et magnificati suntsuper populum Domini exercituum.
ZEPH|2|11|Horribilis Dominus super eos,quia attenuabit omnes deos terrae;et adorabunt eum, singuli de loco suo,omnes insulae gentium.
ZEPH|2|12|" Sed et vos, Aethiopes,interfecti gladio meo eritis ".
ZEPH|2|13|Et extendet manum suam super aquilonemet perdet Assyriam;et ponet Nineven in solitudinemet in aridam, quasi desertum.
ZEPH|2|14|Et accubabunt in medio eius greges,omne genus animalium.Et onocrotalus et ululain capitellis eius morabuntur;vox cantat in fenestra,corvus in limine,quoniam tabulatum cedrinum sublatum est.
ZEPH|2|15|Haec est civitas exsultans,habitans in confidentia,quae dicebat in corde suo: Ego sum, et extra me non est alia amplius! ".Quomodo facta est in desertum,cubile bestiae?Omnis, qui transit per eam,sibilabit et movebit manum suam.
ZEPH|3|1|Vae, provocatrix et inquinata,civitas violenta!
ZEPH|3|2|Non audivit vocem,non suscepit disciplinam;in Domino non est confisa,ad Deum suum non appropiavit.
ZEPH|3|3|Principes eius in medio eiusleones rugientes;iudices eius lupi deserti,ossa non relinquunt in mane.
ZEPH|3|4|Prophetae eius vaniloqui,viri fallaces;sacerdotes eius polluerunt sanctum, iniuste egerunt contra legem.
ZEPH|3|5|Dominus iustus in medio eiusnon faciet iniquitatem;mane, mane iudicium suum dabit, sicut lucem, quae non deficit;nescivit autem iniquus confusionem.
ZEPH|3|6|" Disperdidi gentes,dissipati sunt anguli earum;desertas feci vias eorum,dum non est qui transeat;desolatae sunt civitates eorum,non remanente viro nec ullo habitatore.
ZEPH|3|7|Dixi: Nunc timebis me,suscipies disciplinam!Et non evanescent ab oculis eius omnia, in quibus visitavi eam.Verumtamen acceleraverunt corrumpereomnes actiones suas.
ZEPH|3|8|Quapropter exspecta me,dicit Dominus,in die qua surgam ut testis;quia iudicium meum, ut congregem genteset colligam regna,ut effundam super eas indignationem meam,omnem iram furoris mei;in igne enim zeli meidevorabitur omnis terra.
ZEPH|3|9|Quia tunc reddam populislabium purum,ut invocent omnes in nomine Dominiet serviant ei umero uno.
ZEPH|3|10|Ultra flumina Aethiopiae,inde supplices mei,filii dispersorum meorumdeferent munus mihi.
ZEPH|3|11|In die illa non confunderissuper cunctis actionibus tuis,quibus praevaricata es in me;quia tunc auferam de medio tuimagniloquos superbos tuos,et non adicies exaltari ampliusin monte sancto meo.
ZEPH|3|12|Et derelinquam in medio tuipopulum pauperem et egenum ".Et sperabunt in nomine Dominireliquiae Israel.
ZEPH|3|13|Non facient iniquitatemnec loquentur mendacium;et non invenietur in ore eorumlingua dolosa,quoniam ipsi pascentur et accubabunt,et non erit qui exterreat.
ZEPH|3|14|Lauda, filia Sion;iubilate, Israel!Laetare et exsulta in omni corde,filia Ierusalem!
ZEPH|3|15|Abstulit Dominus iudicium tuum,avertit inimicos tuos;rex Israel, Dominus, in medio tui,non timebis malum ultra.
ZEPH|3|16|In die illa dicetur Ierusalem: Noli timere, Sion;ne dissolvantur manus tuae!
ZEPH|3|17|Dominus Deus tuus in medio tui,fortis ipse salvabit;gaudebit super te in laetitia,commotus in dilectione sua;exsultabit super te in laude
ZEPH|3|18|sicut in die conventus ". Auferam a te calamitatem,ut non ultra habeas super ea opprobrium.
ZEPH|3|19|Ecce ego interficiamomnes, qui afflixerunt tein tempore illo;et salvabo claudicantemet eam, quae eiecta fuerat, congregabo;et ponam eos in laudem et in nomen in omni terra confusionis eorum,
ZEPH|3|20|in tempore illo, quo adducam vos,et in tempore, quo congregabo vos. Dabo enim vos in nomen et in laudemomnibus populis terrae,cum convertero sortem vestramcoram oculis vestris ",dicit Dominus.
