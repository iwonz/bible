HAB|1|1|The burden which Habakkuk the prophet did see.
HAB|1|2|O LORD, how long shall I cry, and thou wilt not hear! even cry out unto thee of violence, and thou wilt not save!
HAB|1|3|Why dost thou shew me iniquity, and cause me to behold grievance? for spoiling and violence are before me: and there are that raise up strife and contention.
HAB|1|4|Therefore the law is slacked, and judgment doth never go forth: for the wicked doth compass about the righteous; therefore wrong judgment proceedeth.
HAB|1|5|Behold ye among the heathen, and regard, and wonder marvelously: for I will work a work in your days which ye will not believe, though it be told you.
HAB|1|6|For, lo, I raise up the Chaldeans, that bitter and hasty nation, which shall march through the breadth of the land, to possess the dwellingplaces that are not their's.
HAB|1|7|They are terrible and dreadful: their judgment and their dignity shall proceed of themselves.
HAB|1|8|Their horses also are swifter than the leopards, and are more fierce than the evening wolves: and their horsemen shall spread themselves, and their horsemen shall come from far; they shall fly as the eagle that hasteth to eat.
HAB|1|9|They shall come all for violence: their faces shall sup up as the east wind, and they shall gather the captivity as the sand.
HAB|1|10|And they shall scoff at the kings, and the princes shall be a scorn unto them: they shall deride every strong hold; for they shall heap dust, and take it.
HAB|1|11|Then shall his mind change, and he shall pass over, and offend, imputing this his power unto his god.
HAB|1|12|Art thou not from everlasting, O LORD my God, mine Holy One? we shall not die. O LORD, thou hast ordained them for judgment; and, O mighty God, thou hast established them for correction.
HAB|1|13|Thou art of purer eyes than to behold evil, and canst not look on iniquity: wherefore lookest thou upon them that deal treacherously, and holdest thy tongue when the wicked devoureth the man that is more righteous than he?
HAB|1|14|And makest men as the fishes of the sea, as the creeping things, that have no ruler over them?
HAB|1|15|They take up all of them with the angle, they catch them in their net, and gather them in their drag: therefore they rejoice and are glad.
HAB|1|16|Therefore they sacrifice unto their net, and burn incense unto their drag; because by them their portion is fat, and their meat plenteous.
HAB|1|17|Shall they therefore empty their net, and not spare continually to slay the nations?
HAB|2|1|I will stand upon my watch, and set me upon the tower, and will watch to see what he will say unto me, and what I shall answer when I am reproved.
HAB|2|2|And the LORD answered me, and said, Write the vision, and make it plain upon tables, that he may run that readeth it.
HAB|2|3|For the vision is yet for an appointed time, but at the end it shall speak, and not lie: though it tarry, wait for it; because it will surely come, it will not tarry.
HAB|2|4|Behold, his soul which is lifted up is not upright in him: but the just shall live by his faith.
HAB|2|5|Yea also, because he transgresseth by wine, he is a proud man, neither keepeth at home, who enlargeth his desire as hell, and is as death, and cannot be satisfied, but gathereth unto him all nations, and heapeth unto him all people:
HAB|2|6|Shall not all these take up a parable against him, and a taunting proverb against him, and say, Woe to him that increaseth that which is not his! how long? and to him that ladeth himself with thick clay!
HAB|2|7|Shall they not rise up suddenly that shall bite thee, and awake that shall vex thee, and thou shalt be for booties unto them?
HAB|2|8|Because thou hast spoiled many nations, all the remnant of the people shall spoil thee; because of men's blood, and for the violence of the land, of the city, and of all that dwell therein.
HAB|2|9|Woe to him that coveteth an evil covetousness to his house, that he may set his nest on high, that he may be delivered from the power of evil!
HAB|2|10|Thou hast consulted shame to thy house by cutting off many people, and hast sinned against thy soul.
HAB|2|11|For the stone shall cry out of the wall, and the beam out of the timber shall answer it.
HAB|2|12|Woe to him that buildeth a town with blood, and stablisheth a city by iniquity!
HAB|2|13|Behold, is it not of the LORD of hosts that the people shall labour in the very fire, and the people shall weary themselves for very vanity?
HAB|2|14|For the earth shall be filled with the knowledge of the glory of the LORD, as the waters cover the sea.
HAB|2|15|Woe unto him that giveth his neighbour drink, that puttest thy bottle to him, and makest him drunken also, that thou mayest look on their nakedness!
HAB|2|16|Thou art filled with shame for glory: drink thou also, and let thy foreskin be uncovered: the cup of the LORD's right hand shall be turned unto thee, and shameful spewing shall be on thy glory.
HAB|2|17|For the violence of Lebanon shall cover thee, and the spoil of beasts, which made them afraid, because of men's blood, and for the violence of the land, of the city, and of all that dwell therein.
HAB|2|18|What profiteth the graven image that the maker thereof hath graven it; the molten image, and a teacher of lies, that the maker of his work trusteth therein, to make dumb idols?
HAB|2|19|Woe unto him that saith to the wood, Awake; to the dumb stone, Arise, it shall teach! Behold, it is laid over with gold and silver, and there is no breath at all in the midst of it.
HAB|2|20|But the LORD is in his holy temple: let all the earth keep silence before him.
HAB|3|1|A prayer of Habakkuk the prophet upon Shigionoth.
HAB|3|2|O LORD, I have heard thy speech, and was afraid: O LORD, revive thy work in the midst of the years, in the midst of the years make known; in wrath remember mercy.
HAB|3|3|God came from Teman, and the Holy One from mount Paran. Selah. His glory covered the heavens, and the earth was full of his praise.
HAB|3|4|And his brightness was as the light; he had horns coming out of his hand: and there was the hiding of his power.
HAB|3|5|Before him went the pestilence, and burning coals went forth at his feet.
HAB|3|6|He stood, and measured the earth: he beheld, and drove asunder the nations; and the everlasting mountains were scattered, the perpetual hills did bow: his ways are everlasting.
HAB|3|7|I saw the tents of Cushan in affliction: and the curtains of the land of Midian did tremble.
HAB|3|8|Was the LORD displeased against the rivers? was thine anger against the rivers? was thy wrath against the sea, that thou didst ride upon thine horses and thy chariots of salvation?
HAB|3|9|Thy bow was made quite naked, according to the oaths of the tribes, even thy word. Selah. Thou didst cleave the earth with rivers.
HAB|3|10|The mountains saw thee, and they trembled: the overflowing of the water passed by: the deep uttered his voice, and lifted up his hands on high.
HAB|3|11|The sun and moon stood still in their habitation: at the light of thine arrows they went, and at the shining of thy glittering spear.
HAB|3|12|Thou didst march through the land in indignation, thou didst thresh the heathen in anger.
HAB|3|13|Thou wentest forth for the salvation of thy people, even for salvation with thine anointed; thou woundedst the head out of the house of the wicked, by discovering the foundation unto the neck. Selah.
HAB|3|14|Thou didst strike through with his staves the head of his villages: they came out as a whirlwind to scatter me: their rejoicing was as to devour the poor secretly.
HAB|3|15|Thou didst walk through the sea with thine horses, through the heap of great waters.
HAB|3|16|When I heard, my belly trembled; my lips quivered at the voice: rottenness entered into my bones, and I trembled in myself, that I might rest in the day of trouble: when he cometh up unto the people, he will invade them with his troops.
HAB|3|17|Although the fig tree shall not blossom, neither shall fruit be in the vines; the labour of the olive shall fail, and the fields shall yield no meat; the flock shall be cut off from the fold, and there shall be no herd in the stalls:
HAB|3|18|Yet I will rejoice in the LORD, I will joy in the God of my salvation.
HAB|3|19|The LORD God is my strength, and he will make my feet like hinds' feet, and he will make me to walk upon mine high places. To the chief singer on my stringed instruments.
