ZECH|1|1|In the eighth month, in the second year of Darius, the word of the LORD came to the prophet Zechariah, the son of Berechiah, son of Iddo, saying,
ZECH|1|2|"The LORD was very angry with your fathers.
ZECH|1|3|Therefore say to them, Thus declares the LORD of hosts: Return to me, says the LORD of hosts, and I will return to you, says the LORD of hosts.
ZECH|1|4|Do not be like your fathers, to whom the former prophets cried out, 'Thus says the LORD of hosts, Return from your evil ways and from your evil deeds.' But they did not hear or pay attention to me, declares the LORD.
ZECH|1|5|Your fathers, where are they? And the prophets, do they live forever?
ZECH|1|6|But my words and my statutes, which I commanded my servants the prophets, did they not overtake your fathers? So they repented and said, As the LORD of hosts purposed to deal with us for our ways and deeds, so has he dealt with us."
ZECH|1|7|On the twenty-fourth day of the eleventh month, which is the month of Shebat, in the second year of Darius, the word of the LORD came to the prophet Zechariah, the son of Berechiah, son of Iddo, saying,
ZECH|1|8|"I saw in the night, and behold, a man riding on a red horse! He was standing among the myrtle trees in the glen, and behind him were red, sorrel, and white horses.
ZECH|1|9|Then I said, 'What are these, my lord?' The angel who talked with me said to me, 'I will show you what they are.'
ZECH|1|10|So the man who was standing among the myrtle trees answered, 'These are they whom the LORD has sent to patrol the earth.'
ZECH|1|11|And they answered the angel of the LORD who was standing among the myrtle trees, and said, 'We have patrolled the earth, and behold, all the earth remains at rest.'
ZECH|1|12|Then the angel of the LORD said, 'O LORD of hosts, how long will you have no mercy on Jerusalem and the cities of Judah, against which you have been angry these seventy years?'
ZECH|1|13|And the LORD answered gracious and comforting words to the angel who talked with me.
ZECH|1|14|So the angel who talked with me said to me, 'Cry out, Thus says the LORD of hosts: I am exceedingly jealous for Jerusalem and for Zion.
ZECH|1|15|And I am exceedingly angry with the nations that are at ease; for while I was angry but a little, they furthered the disaster.
ZECH|1|16|Therefore, thus says the LORD, I have returned to Jerusalem with mercy; my house shall be built in it, declares the LORD of hosts, and the measuring line shall be stretched out over Jerusalem.
ZECH|1|17|Cry out again, Thus says the LORD of hosts: My cities shall again overflow with prosperity, and the LORD will again comfort Zion and again choose Jerusalem.'"
ZECH|1|18|And I lifted my eyes and saw, and behold, four horns!
ZECH|1|19|And I said to the angel who talked with me, "What are these?" And he said to me, "These are the horns that have scattered Judah, Israel, and Jerusalem."
ZECH|1|20|Then the LORD showed me four craftsmen.
ZECH|1|21|And I said, "What are these coming to do?" He said, "These are the horns that scattered Judah, so that no one raised his head. And these have come to terrify them, to cast down the horns of the nations who lifted up their horns against the land of Judah to scatter it."
ZECH|2|1|And I lifted my eyes and saw, and behold, a man with a measuring line in his hand!
ZECH|2|2|Then I said, "Where are you going?" And he said to me, "To measure Jerusalem, to see what is its width and what is its length."
ZECH|2|3|And behold, the angel who talked with me came forward, and another angel came forward to meet him
ZECH|2|4|and said to him, "Run, say to that young man, 'Jerusalem shall be inhabited as villages without walls, because of the multitude of people and livestock in it.
ZECH|2|5|And I will be to her a wall of fire all around, declares the LORD, and I will be the glory in her midst.'"
ZECH|2|6|Up! Up! Flee from the land of the north, declares the LORD. For I have spread you abroad as the four winds of the heavens, declares the LORD.
ZECH|2|7|Up! Escape to Zion, you who dwell with the daughter of Babylon.
ZECH|2|8|For thus said the LORD of hosts, after his glory sent me to the nations who plundered you, for he who touches you touches the apple of his eye:
ZECH|2|9|"Behold, I will shake my hand over them, and they shall become plunder for those who served them. Then you will know that the LORD of hosts has sent me.
ZECH|2|10|Sing and rejoice, O daughter of Zion, for behold, I come and I will dwell in your midst, declares the LORD.
ZECH|2|11|And many nations shall join themselves to the LORD in that day, and shall be my people. And I will dwell in your midst, and you shall know that the LORD of hosts has sent me to you.
ZECH|2|12|And the LORD will inherit Judah as his portion in the holy land, and will again choose Jerusalem."
ZECH|2|13|Be silent, all flesh, before the LORD, for he has roused himself from his holy dwelling.
ZECH|3|1|Then he showed me Joshua the high priest standing before the angel of the LORD, and Satan standing at his right hand to accuse him.
ZECH|3|2|And the LORD said to Satan, "The LORD rebuke you, O Satan! The LORD who has chosen Jerusalem rebuke you! Is not this a brand plucked from the fire?"
ZECH|3|3|Now Joshua was standing before the angel, clothed with filthy garments.
ZECH|3|4|And the angel said to those who were standing before him, "Remove the filthy garments from him." And to him he said, "Behold, I have taken your iniquity away from you, and I will clothe you with pure vestments."
ZECH|3|5|And I said, "Let them put a clean turban on his head." So they put a clean turban on his head and clothed him with garments. And the angel of the LORD was standing by.
ZECH|3|6|And the angel of the LORD solemnly assured Joshua,
ZECH|3|7|"Thus says the LORD of hosts: If you will walk in my ways and keep my charge, then you shall rule my house and have charge of my courts, and I will give you the right of access among those who are standing here.
ZECH|3|8|Hear now, O Joshua the high priest, you and your friends who sit before you, for they are men who are a sign: behold, I will bring my servant the Branch.
ZECH|3|9|For behold, on the stone that I have set before Joshua, on a single stone with seven eyes, I will engrave its inscription, declares the LORD of hosts, and I will remove the iniquity of this land in a single day.
ZECH|3|10|In that day, declares the LORD of hosts, every one of you will invite his neighbor to come under his vine and under his fig tree."
ZECH|4|1|And the angel who talked with me came again and woke me, like a man who is awakened out of his sleep.
ZECH|4|2|And he said to me, "What do you see?" I said, "I see, and behold, a lampstand all of gold, with a bowl on the top of it, and seven lamps on it, with seven lips on each of the lamps that are on the top of it.
ZECH|4|3|And there are two olive trees by it, one on the right of the bowl and the other on its left."
ZECH|4|4|And I said to the angel who talked with me, "What are these, my lord?"
ZECH|4|5|Then the angel who talked with me answered and said to me, "Do you not know what these are?" I said, "No, my lord."
ZECH|4|6|Then he said to me, "This is the word of the LORD to Zerubbabel: Not by might, nor by power, but by my Spirit, says the LORD of hosts.
ZECH|4|7|Who are you, O great mountain? Before Zerubbabel you shall become a plain. And he shall bring forward the top stone amid shouts of 'Grace, grace to it!'"
ZECH|4|8|Then the word of the LORD came to me, saying,
ZECH|4|9|"The hands of Zerubbabel have laid the foundation of this house; his hands shall also complete it. Then you will know that the LORD of hosts has sent me to you.
ZECH|4|10|For whoever has despised the day of small things shall rejoice, and shall see the plumb line in the hand of Zerubbabel. "These seven are the eyes of the LORD, which range through the whole earth."
ZECH|4|11|Then I said to him, "What are these two olive trees on the right and the left of the lampstand?"
ZECH|4|12|And a second time I answered and said to him, "What are these two branches of the olive trees, which are beside the two golden pipes from which the golden oil is poured out?"
ZECH|4|13|He said to me, "Do you not know what these are?" I said, "No, my lord."
ZECH|4|14|Then he said, "These are the two anointed ones who stand by the Lord of the whole earth."
ZECH|5|1|Again I lifted my eyes and saw, and behold, a flying scroll!
ZECH|5|2|And he said to me, "What do you see?" I answered, "I see a flying scroll. Its length is twenty cubits, and its width ten cubits."
ZECH|5|3|Then he said to me, "This is the curse that goes out over the face of the whole land. For everyone who steals shall be cleaned out according to what is on one side, and everyone who swears falsely shall be cleaned out according to what is on the other side.
ZECH|5|4|I will send it out, declares the LORD of hosts, and it shall enter the house of the thief, and the house of him who swears falsely by my name. And it shall remain in his house and consume it, both timber and stones."
ZECH|5|5|Then the angel who talked with me came forward and said to me, "Lift your eyes and see what this is that is going out."
ZECH|5|6|And I said, "What is it?" He said, "This is the basket that is going out." And he said, "This is their iniquity in all the land."
ZECH|5|7|And behold, the leaden cover was lifted, and there was a woman sitting in the basket!
ZECH|5|8|And he said, "This is Wickedness." And he thrust her back into the basket, and thrust down the leaden weight on its opening.
ZECH|5|9|Then I lifted my eyes and saw, and behold, two women coming forward! The wind was in their wings. They had wings like the wings of a stork, and they lifted up the basket between earth and heaven.
ZECH|5|10|Then I said to the angel who talked with me, "Where are they taking the basket?"
ZECH|5|11|He said to me, "To the land of Shinar, to build a house for it. And when this is prepared, they will set the basket down there on its base."
ZECH|6|1|Again I lifted my eyes and saw, and behold, four chariots came out from between two mountains. And the mountains were mountains of bronze.
ZECH|6|2|The first chariot had red horses, the second black horses,
ZECH|6|3|the third white horses, and the fourth chariot dappled horses- all of them strong.
ZECH|6|4|Then I answered and said to the angel who talked with me, "What are these, my lord?"
ZECH|6|5|And the angel answered and said to me, "These are going out to the four winds of heaven, after presenting themselves before the LORD of all the earth.
ZECH|6|6|The chariot with the black horses goes toward the north country, the white ones go after them, and the dappled ones go toward the south country."
ZECH|6|7|When the strong horses came out, they were impatient to go and patrol the earth. And he said, "Go, patrol the earth." So they patrolled the earth.
ZECH|6|8|Then he cried to me, "Behold, those who go toward the north country have set my Spirit at rest in the north country."
ZECH|6|9|And the word of the LORD came to me:
ZECH|6|10|"Take from the exiles Heldai, Tobijah, and Jedaiah, who have arrived from Babylon, and go the same day to the house of Josiah, the son of Zephaniah.
ZECH|6|11|Take from them silver and gold, and make a crown, and set it on the head of Joshua, the son of Jehozadak, the high priest.
ZECH|6|12|And say to him, 'Thus says the LORD of hosts, "Behold, the man whose name is the Branch: for he shall branch out from his place, and he shall build the temple of the LORD.
ZECH|6|13|It is he who shall build the temple of the LORD and shall bear royal honor, and shall sit and rule on his throne. And there shall be a priest on his throne, and the counsel of peace shall be between them both."'
ZECH|6|14|And the crown shall be in the temple of the LORD as a reminder to Helem, Tobijah, Jedaiah, and Hen the son of Zephaniah.
ZECH|6|15|"And those who are far off shall come and help to build the temple of the LORD. And you shall know that the LORD of hosts has sent me to you. And this shall come to pass, if you will diligently obey the voice of the LORD your God."
ZECH|7|1|In the fourth year of King Darius, the word of the LORD came to Zechariah on the fourth day of the ninth month, which is Chislev.
ZECH|7|2|Now the people of Bethel had sent Sharezer and Regem-melech and their men to entreat the favor of the LORD,
ZECH|7|3|saying to the priests of the house of the LORD of hosts and the prophets, "Should I weep and abstain in the fifth month, as I have done for so many years?"
ZECH|7|4|Then the word of the LORD of hosts came to me:
ZECH|7|5|"Say to all the people of the land and the priests, When you fasted and mourned in the fifth month and in the seventh, for these seventy years, was it for me that you fasted?
ZECH|7|6|And when you eat and when you drink, do you not eat for yourselves and drink for yourselves?
ZECH|7|7|Were not these the words that the LORD proclaimed by the former prophets, when Jerusalem was inhabited and prosperous, with her cities around her, and the South and the lowland were inhabited?"
ZECH|7|8|And the word of the LORD came to Zechariah, saying,
ZECH|7|9|"Thus says the LORD of hosts, Render true judgments, show kindness and mercy to one another,
ZECH|7|10|do not oppress the widow, the fatherless, the sojourner, or the poor, and let none of you devise evil against another in your heart."
ZECH|7|11|But they refused to pay attention and turned a stubborn shoulder and stopped their ears that they might not hear.
ZECH|7|12|They made their hearts diamond-hard lest they should hear the law and the words that the LORD of hosts had sent by his Spirit through the former prophets. Therefore great anger came from the LORD of hosts.
ZECH|7|13|"As I called, and they would not hear, so they called, and I would not hear," says the LORD of hosts,
ZECH|7|14|"and I scattered them with a whirlwind among all the nations that they had not known. Thus the land they left was desolate, so that no one went to and fro, and the pleasant land was made desolate."
ZECH|8|1|And the word of the LORD of hosts came, saying,
ZECH|8|2|"Thus says the LORD of hosts: I am jealous for Zion with great jealousy, and I am jealous for her with great wrath.
ZECH|8|3|Thus says the LORD: I have returned to Zion and will dwell in the midst of Jerusalem, and Jerusalem shall be called the faithful city, and the mountain of the LORD of hosts, the holy mountain.
ZECH|8|4|Thus says the LORD of hosts: Old men and old women shall again sit in the streets of Jerusalem, each with staff in hand because of great age.
ZECH|8|5|And the streets of the city shall be full of boys and girls playing in its streets.
ZECH|8|6|Thus says the LORD of hosts: If it is marvelous in the sight of the remnant of this people in those days, should it also be marvelous in my sight, declares the LORD of hosts?
ZECH|8|7|Thus says the LORD of hosts: behold, I will save my people from the east country and from the west country,
ZECH|8|8|and I will bring them to dwell in the midst of Jerusalem. And they shall be my people, and I will be their God, in faithfulness and in righteousness."
ZECH|8|9|Thus says the LORD of hosts: "Let your hands be strong, you who in these days have been hearing these words from the mouth of the prophets who were present on the day that the foundation of the house of the LORD of hosts was laid, that the temple might be built.
ZECH|8|10|For before those days there was no wage for man or any wage for beast, neither was there any safety from the foe for him who went out or came in, for I set every man against his neighbor.
ZECH|8|11|But now I will not deal with the remnant of this people as in the former days, declares the LORD of hosts.
ZECH|8|12|For there shall be a sowing of peace. The vine shall give its fruit, and the ground shall give its produce, and the heavens shall give their dew. And I will cause the remnant of this people to possess all these things.
ZECH|8|13|And as you have been a byword of cursing among the nations, O house of Judah and house of Israel, so will I save you, and you shall be a blessing. Fear not, but let your hands be strong."
ZECH|8|14|For thus says the LORD of hosts: "As I purposed to bring disaster to you when your fathers provoked me to wrath, and I did not relent, says the LORD of hosts,
ZECH|8|15|so again have I purposed in these days to bring good to Jerusalem and to the house of Judah; fear not.
ZECH|8|16|These are the things that you shall do: Speak the truth to one another; render in your gates judgments that are true and make for peace;
ZECH|8|17|do not devise evil in your hearts against one another, and love no false oath, for all these things I hate, declares the LORD."
ZECH|8|18|And the word of the LORD of hosts came to me, saying,
ZECH|8|19|"Thus says the LORD of hosts: The fast of the fourth month and the fast of the fifth and the fast of the seventh and the fast of the tenth shall be to the house of Judah seasons of joy and gladness and cheerful feasts. Therefore love truth and peace.
ZECH|8|20|"Thus says the LORD of hosts: Peoples shall yet come, even the inhabitants of many cities.
ZECH|8|21|The inhabitants of one city shall go to another, saying, 'Let us go at once to entreat the favor of the LORD and to seek the LORD of hosts; I myself am going.'
ZECH|8|22|Many peoples and strong nations shall come to seek the LORD of hosts in Jerusalem and to entreat the favor of the LORD.
ZECH|8|23|Thus says the LORD of hosts: In those days ten men from the nations of every tongue shall take hold of the robe of a Jew, saying, 'Let us go with you, for we have heard that God is with you.'"
ZECH|9|1|The burden of the word of the LORD is against the land of Hadrach and Damascus is its resting place. For the LORD has an eye on mankind and on all the tribes of Israel,
ZECH|9|2|and on Hamath also, which borders on it, Tyre and Sidon, though they are very wise.
ZECH|9|3|Tyre has built herself a rampart and heaped up silver like dust, and fine gold like the mud of the streets.
ZECH|9|4|But behold, the Lord will strip her of her possessions and strike down her power on the sea, and she shall be devoured by fire.
ZECH|9|5|Ashkelon shall see it, and be afraid; Gaza too, and shall writhe in anguish; Ekron also, because its hopes are confounded. The king shall perish from Gaza; Ashkelon shall be uninhabited;
ZECH|9|6|a mixed people shall dwell in Ashdod, and I will cut off the pride of Philistia.
ZECH|9|7|I will take away its blood from its mouth, and its abominations from between its teeth; it too shall be a remnant for our God; it shall be like a clan in Judah, and Ekron shall be like the Jebusites.
ZECH|9|8|Then I will encamp at my house as a guard, so that none shall march to and fro; no oppressor shall again march over them, for now I see with my own eyes.
ZECH|9|9|Rejoice greatly, O daughter of Zion! Shout aloud, O daughter of Jerusalem! behold, your king is coming to you; righteous and having salvation is he, humble and mounted on a donkey, on a colt, the foal of a donkey.
ZECH|9|10|I will cut off the chariot from Ephraim and the war horse from Jerusalem; and the battle bow shall be cut off, and he shall speak peace to the nations; his rule shall be from sea to sea, and from the River to the ends of the earth.
ZECH|9|11|As for you also, because of the blood of my covenant with you, I will set your prisoners free from the waterless pit.
ZECH|9|12|Return to your stronghold, O prisoners of hope; today I declare that I will restore to you double.
ZECH|9|13|For I have bent Judah as my bow; I have made Ephraim its arrow. I will stir up your sons, O Zion, against your sons, O Greece, and wield you like a warrior's sword.
ZECH|9|14|Then the LORD will appear over them, and his arrow will go forth like lightning; the Lord GOD will sound the trumpet and will march forth in the whirlwinds of the south.
ZECH|9|15|The LORD of hosts will protect them, and they shall devour, and tread down the sling stones, and they shall drink and roar as if drunk with wine, and be full like a bowl, drenched like the corners of the altar.
ZECH|9|16|On that day the LORD their God will save them, as the flock of his people; for like the jewels of a crown they shall shine on his land.
ZECH|9|17|For how great is his goodness, and how great his beauty! Grain shall make the young men flourish, and new wine the young women.
ZECH|10|1|Ask rain from the LORD in the season of the spring rain, from the LORD who makes the storm clouds, and he will give them showers of rain, to everyone the vegetation in the field.
ZECH|10|2|For the household gods utter nonsense, and the diviners see lies; they tell false dreams and give empty consolation. Therefore the people wander like sheep; they are afflicted for lack of a shepherd.
ZECH|10|3|"My anger is hot against the shepherds, and I will punish the leaders; for the LORD of hosts cares for his flock, the house of Judah, and will make them like his majestic steed in battle.
ZECH|10|4|From him shall come the cornerstone, from him the tent peg, from him the battle bow, from him every ruler- all of them together.
ZECH|10|5|They shall be like mighty men in battle, trampling the foe in the mud of the streets; they shall fight because the LORD is with them, and they shall put to shame the riders on horses.
ZECH|10|6|"I will strengthen the house of Judah, and I will save the house of Joseph. I will bring them back because I have compassion on them, and they shall be as though I had not rejected them, for I am the LORD their God and I will answer them.
ZECH|10|7|Then Ephraim shall become like a mighty warrior, and their hearts shall be glad as with wine. Their children shall see it and be glad; their hearts shall rejoice in the LORD.
ZECH|10|8|"I will whistle for them and gather them in, for I have redeemed them, and they shall be as many as they were before.
ZECH|10|9|Though I scattered them among the nations, yet in far countries they shall remember me, and with their children they shall live and return.
ZECH|10|10|I will bring them home from the land of Egypt, and gather them from Assyria, and I will bring them to the land of Gilead and to Lebanon, till there is no room for them.
ZECH|10|11|He shall pass through the sea of troubles and strike down the waves of the sea, and all the depths of the Nile shall be dried up. The pride of Assyria shall be laid low, and the scepter of Egypt shall depart.
ZECH|10|12|I will make them strong in the LORD, and they shall walk in his name," declares the LORD.
ZECH|11|1|Open your doors, O Lebanon, that the fire may devour your cedars!
ZECH|11|2|Wail, O cypress, for the cedar has fallen, for the glorious trees are ruined! Wail, oaks of Bashan, for the thick forest has been felled!
ZECH|11|3|The sound of the wail of the shepherds, for their glory is ruined! The sound of the roar of the lions, for the thicket of the Jordan is ruined!
ZECH|11|4|Thus said the LORD my God: "Become shepherd of the flock doomed to slaughter.
ZECH|11|5|Those who buy them slaughter them and go unpunished, and those who sell them say, 'Blessed be the LORD, I have become rich,' and their own shepherds have no pity on them.
ZECH|11|6|For I will no longer have pity on the inhabitants of this land, declares the LORD. Behold, I will cause each of them to fall into the hand of his neighbor, and each into the hand of his king, and they shall crush the land, and I will deliver none from their hand."
ZECH|11|7|So I became the shepherd of the flock doomed to be slaughtered by the sheep traders. And I took two staffs, one I named Favor, the other I named Union. And I tended the sheep.
ZECH|11|8|In one month I destroyed the three shepherds. But I became impatient with them, and they also detested me.
ZECH|11|9|So I said, "I will not be your shepherd. What is to die, let it die. What is to be destroyed, let it be destroyed. And let those who are left devour the flesh of one another."
ZECH|11|10|And I took my staff Favor, and I broke it, annulling the covenant that I had made with all the peoples.
ZECH|11|11|So it was annulled on that day, and the sheep traders, who were watching me, knew that it was the word of the LORD.
ZECH|11|12|Then I said to them, "If it seems good to you, give me my wages; but if not, keep them." And they weighed out as my wages thirty pieces of silver.
ZECH|11|13|Then the LORD said to me, "Throw it to the potter"- the lordly price at which I was priced by them. So I took the thirty pieces of silver and threw them into the house of the LORD, to the potter.
ZECH|11|14|Then I broke my second staff Union, annulling the brotherhood between Judah and Israel.
ZECH|11|15|Then the LORD said to me, "Take once more the equipment of a foolish shepherd.
ZECH|11|16|For behold, I am raising up in the land a shepherd who does not care for those being destroyed, or seek the young or heal the maimed or nourish the healthy, but devours the flesh of the fat ones, tearing off even their hoofs.
ZECH|11|17|"Woe to my worthless shepherd, who deserts the flock! May the sword strike his arm and his right eye! Let his arm be wholly withered, his right eye utterly blinded!"
ZECH|12|1|The burden of the word of the LORD concerning Israel: Thus declares the LORD, who stretched out the heavens and founded the earth and formed the spirit of man within him:
ZECH|12|2|"Behold, I am about to make Jerusalem a cup of staggering to all the surrounding peoples. The siege of Jerusalem will also be against Judah.
ZECH|12|3|On that day I will make Jerusalem a heavy stone for all the peoples. All who lift it will surely hurt themselves. And all the nations of the earth will gather against it.
ZECH|12|4|On that day, declares the LORD, I will strike every horse with panic, and its rider with madness. But for the sake of the house of Judah I will keep my eyes open, when I strike every horse of the peoples with blindness.
ZECH|12|5|Then the clans of Judah shall say to themselves, 'The inhabitants of Jerusalem have strength through the LORD of hosts, their God.'
ZECH|12|6|"On that day I will make the clans of Judah like a blazing pot in the midst of wood, like a flaming torch among sheaves. And they shall devour to the right and to the left all the surrounding peoples, while Jerusalem shall again be inhabited in its place, in Jerusalem.
ZECH|12|7|"And the LORD will give salvation to the tents of Judah first, that the glory of the house of David and the glory of the inhabitants of Jerusalem may not surpass that of Judah.
ZECH|12|8|On that day the LORD will protect the inhabitants of Jerusalem, so that the feeblest among them on that day shall be like David, and the house of David shall be like God, like the angel of the LORD, going before them.
ZECH|12|9|And on that day I will seek to destroy all the nations that come against Jerusalem.
ZECH|12|10|"And I will pour out on the house of David and the inhabitants of Jerusalem a spirit of grace and pleas for mercy, so that, when they look on me, on him whom they have pierced, they shall mourn for him, as one mourns for an only child, and weep bitterly over him, as one weeps over a firstborn.
ZECH|12|11|On that day the mourning in Jerusalem will be as great as the mourning for Hadad-rimmon in the plain of Megiddo.
ZECH|12|12|The land shall mourn, each family by itself: the family of the house of David by itself, and their wives by themselves; the family of the house of Nathan by itself, and their wives by themselves;
ZECH|12|13|the family of the house of Levi by itself, and their wives by themselves; the family of the Shimeites by itself, and their wives by themselves;
ZECH|12|14|and all the families that are left, each by itself, and their wives by themselves.
ZECH|13|1|"On that day there shall be a fountain opened for the house of David and the inhabitants of Jerusalem, to cleanse them from sin and uncleanness.
ZECH|13|2|"And on that day, declares the LORD of hosts, I will cut off the names of the idols from the land, so that they shall be remembered no more. And also I will remove from the land the prophets and the spirit of uncleanness.
ZECH|13|3|And if anyone again prophesies, his father and mother who bore him will say to him, 'You shall not live, for you speak lies in the name of the LORD.' And his father and mother who bore him shall pierce him through when he prophesies.
ZECH|13|4|"On that day every prophet will be ashamed of his vision when he prophesies. He will not put on a hairy cloak in order to deceive,
ZECH|13|5|but he will say, 'I am no prophet, I am a worker of the soil, for a man sold me in my youth.'
ZECH|13|6|And if one asks him, 'What are these wounds on your back?' he will say, 'The wounds I received in the house of my friends.'
ZECH|13|7|"Awake, O sword, against my shepherd, against the man who stands next to me," declares the LORD of hosts. "Strike the shepherd, and the sheep will be scattered; I will turn my hand against the little ones.
ZECH|13|8|In the whole land, declares the LORD, two thirds shall be cut off and perish, and one third shall be left alive.
ZECH|13|9|And I will put this third into the fire, and refine them as one refines silver, and test them as gold is tested. They will call upon my name, and I will answer them. I will say, 'They are my people'; and they will say, 'The LORD is my God.'"
ZECH|14|1|Behold, a day is coming for the LORD, when the spoil taken from you will be divided in your midst.
ZECH|14|2|For I will gather all the nations against Jerusalem to battle, and the city shall be taken and the houses plundered and the women raped. Half of the city shall go out into exile, but the rest of the people shall not be cut off from the city.
ZECH|14|3|Then the LORD will go out and fight against those nations as when he fights on a day of battle.
ZECH|14|4|On that day his feet shall stand on the Mount of Olives that lies before Jerusalem on the east, and the Mount of Olives shall be split in two from east to west by a very wide valley, so that one half of the Mount shall move northward, and the other half southward.
ZECH|14|5|And you shall flee to the valley of my mountains, for the valley of the mountains shall reach to Azal. And you shall flee as you fled from the earthquake in the days of Uzziah king of Judah. Then the LORD my God will come, and all the holy ones with him.
ZECH|14|6|On that day there shall be no light, cold, or frost.
ZECH|14|7|And there shall be a unique day, which is known to the LORD, neither day nor night, but at evening time there shall be light.
ZECH|14|8|On that day living waters shall flow out from Jerusalem, half of them to the eastern sea and half of them to the western sea. It shall continue in summer as in winter.
ZECH|14|9|And the LORD will be king over all the earth. On that day the LORD will be one and his name one.
ZECH|14|10|The whole land shall be turned into a plain from Geba to Rimmon south of Jerusalem. But Jerusalem shall remain aloft on its site from the Gate of Benjamin to the place of the former gate, to the Corner Gate, and from the Tower of Hananel to the king's winepresses.
ZECH|14|11|And it shall be inhabited, for there shall never again be a decree of utter destruction. Jerusalem shall dwell in security.
ZECH|14|12|And this shall be the plague with which the LORD will strike all the peoples that wage war against Jerusalem: their flesh will rot while they are still standing on their feet, their eyes will rot in their sockets, and their tongues will rot in their mouths.
ZECH|14|13|And on that day a great panic from the LORD shall fall on them, so that each will seize the hand of another, and the hand of the one will be raised against the hand of the other.
ZECH|14|14|Even Judah will fight against Jerusalem. And the wealth of all the surrounding nations shall be collected, gold, silver, and garments in great abundance.
ZECH|14|15|And a plague like this plague shall fall on the horses, the mules, the camels, the donkeys, and whatever beasts may be in those camps.
ZECH|14|16|Then everyone who survives of all the nations that have come against Jerusalem shall go up year after year to worship the King, the LORD of hosts, and to keep the Feast of Booths.
ZECH|14|17|And if any of the families of the earth do not go up to Jerusalem to worship the King, the LORD of hosts, there will be no rain on them.
ZECH|14|18|And if the family of Egypt does not go up and present themselves, then on them there shall be no rain; there shall be the plague with which the LORD afflicts the nations that do not go up to keep the Feast of Booths.
ZECH|14|19|This shall be the punishment to Egypt and the punishment to all the nations that do not go up to keep the Feast of Booths.
ZECH|14|20|And on that day there shall be inscribed on the bells of the horses, "Holy to the LORD." And the pots in the house of the LORD shall be as the bowls before the altar.
ZECH|14|21|And every pot in Jerusalem and Judah shall be holy to the LORD of hosts, so that all who sacrifice may come and take of them and boil the meat of the sacrifice in them. And there shall no longer be a trader in the house of the LORD of hosts on that day.
