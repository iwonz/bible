COL|1|1|Paul, an apostle of Christ Jesus by the will of God, and Timothy our brother,
COL|1|2|To the saints and faithful brothers in Christ at Colossae: Grace to you and peace from God our Father.
COL|1|3|We always thank God, the Father of our Lord Jesus Christ, when we pray for you,
COL|1|4|since we heard of your faith in Christ Jesus and of the love that you have for all the saints,
COL|1|5|because of the hope laid up for you in heaven. Of this you have heard before in the word of the truth, the gospel,
COL|1|6|which has come to you, as indeed in the whole world it is bearing fruit and growing- as it also does among you, since the day you heard it and understood the grace of God in truth,
COL|1|7|just as you learned it from Epaphras our beloved fellow servant. He is a faithful minister of Christ on your behalf
COL|1|8|and has made known to us your love in the Spirit.
COL|1|9|And so, from the day we heard, we have not ceased to pray for you, asking that you may be filled with the knowledge of his will in all spiritual wisdom and understanding,
COL|1|10|so as to walk in a manner worthy of the Lord, fully pleasing to him, bearing fruit in every good work and increasing in the knowledge of God.
COL|1|11|May you be strengthened with all power, according to his glorious might, for all endurance and patience with joy,
COL|1|12|giving thanks to the Father, who has qualified you to share in the inheritance of the saints in light.
COL|1|13|He has delivered us from the domain of darkness and transferred us to the kingdom of his beloved Son,
COL|1|14|in whom we have redemption, the forgiveness of sins.
COL|1|15|He is the image of the invisible God, the firstborn of all creation.
COL|1|16|For by him all things were created, in heaven and on earth, visible and invisible, whether thrones or dominions or rulers or authorities- all things were created through him and for him.
COL|1|17|And he is before all things, and in him all things hold together.
COL|1|18|And he is the head of the body, the church. He is the beginning, the firstborn from the dead, that in everything he might be preeminent.
COL|1|19|For in him all the fullness of God was pleased to dwell,
COL|1|20|and through him to reconcile to himself all things, whether on earth or in heaven, making peace by the blood of his cross.
COL|1|21|And you, who once were alienated and hostile in mind, doing evil deeds,
COL|1|22|he has now reconciled in his body of flesh by his death, in order to present you holy and blameless and above reproach before him,
COL|1|23|if indeed you continue in the faith, stable and steadfast, not shifting from the hope of the gospel that you heard, which has been proclaimed in all creation under heaven, and of which I, Paul, became a minister.
COL|1|24|Now I rejoice in my sufferings for your sake, and in my flesh I am filling up what is lacking in Christ's afflictions for the sake of his body, that is, the church,
COL|1|25|of which I became a minister according to the stewardship from God that was given to me for you, to make the word of God fully known,
COL|1|26|the mystery hidden for ages and generations but now revealed to his saints.
COL|1|27|To them God chose to make known how great among the Gentiles are the riches of the glory of this mystery, which is Christ in you, the hope of glory.
COL|1|28|Him we proclaim, warning everyone and teaching everyone with all wisdom, that we may present everyone mature in Christ.
COL|1|29|For this I toil, struggling with all his energy that he powerfully works within me.
COL|2|1|For I want you to know how great a struggle I have for you and for those at Laodicea and for all who have not seen me face to face,
COL|2|2|that their hearts may be encouraged, being knit together in love, to reach all the riches of full assurance of understanding and the knowledge of God's mystery, which is Christ,
COL|2|3|in whom are hidden all the treasures of wisdom and knowledge.
COL|2|4|I say this in order that no one may delude you with plausible arguments.
COL|2|5|For though I am absent in body, yet I am with you in spirit, rejoicing to see your good order and the firmness of your faith in Christ.
COL|2|6|Therefore, as you received Christ Jesus the Lord, so walk in him,
COL|2|7|rooted and built up in him and established in the faith, just as you were taught, abounding in thanksgiving.
COL|2|8|See to it that no one takes you captive by philosophy and empty deceit, according to human tradition, according to the elemental spirits of the world, and not according to Christ.
COL|2|9|For in him the whole fullness of deity dwells bodily,
COL|2|10|and you have been filled in him, who is the head of all rule and authority.
COL|2|11|In him also you were circumcised with a circumcision made without hands, by putting off the body of the flesh, by the circumcision of Christ,
COL|2|12|having been buried with him in baptism, in which you were also raised with him through faith in the powerful working of God, who raised him from the dead.
COL|2|13|And you, who were dead in your trespasses and the uncircumcision of your flesh, God made alive together with him, having forgiven us all our trespasses,
COL|2|14|by canceling the record of debt that stood against us with its legal demands. This he set aside, nailing it to the cross.
COL|2|15|He disarmed the rulers and authorities and put them to open shame, by triumphing over them in him.
COL|2|16|Therefore let no one pass judgment on you in questions of food and drink, or with regard to a festival or a new moon or a Sabbath.
COL|2|17|These are a shadow of the things to come, but the substance belongs to Christ.
COL|2|18|Let no one disqualify you, insisting on asceticism and worship of angels, going on in detail about visions, puffed up without reason by his sensuous mind,
COL|2|19|and not holding fast to the Head, from whom the whole body, nourished and knit together through its joints and ligaments, grows with a growth that is from God.
COL|2|20|If with Christ you died to the elemental spirits of the world, why, as if you were still alive in the world, do you submit to regulations-
COL|2|21|"Do not handle, Do not taste, Do not touch"
COL|2|22|(referring to things that all perish as they are used)- according to human precepts and teachings?
COL|2|23|These have indeed an appearance of wisdom in promoting self-made religion and asceticism and severity to the body, but they are of no value in stopping the indulgence of the flesh.
COL|3|1|If then you have been raised with Christ, seek the things that are above, where Christ is, seated at the right hand of God.
COL|3|2|Set your minds on things that are above, not on things that are on earth.
COL|3|3|For you have died, and your life is hidden with Christ in God.
COL|3|4|When Christ who is your life appears, then you also will appear with him in glory.
COL|3|5|Put to death therefore what is earthly in you: sexual immorality, impurity, passion, evil desire, and covetousness, which is idolatry.
COL|3|6|On account of these the wrath of God is coming.
COL|3|7|In these you too once walked, when you were living in them.
COL|3|8|But now you must put them all away: anger, wrath, malice, slander, and obscene talk from your mouth.
COL|3|9|Do not lie to one another, seeing that you have put off the old self with its practices
COL|3|10|and have put on the new self, which is being renewed in knowledge after the image of its creator.
COL|3|11|Here there is not Greek and Jew, circumcised and uncircumcised, barbarian, Scythian, slave, free; but Christ is all, and in all.
COL|3|12|Put on then, as God's chosen ones, holy and beloved, compassion, kindness, humility, meekness, and patience,
COL|3|13|bearing with one another and, if one has a complaint against another, forgiving each other; as the Lord has forgiven you, so you also must forgive.
COL|3|14|And above all these put on love, which binds everything together in perfect harmony.
COL|3|15|And let the peace of Christ rule in your hearts, to which indeed you were called in one body. And be thankful.
COL|3|16|Let the word of Christ dwell in you richly, teaching and admonishing one another in all wisdom, singing psalms and hymns and spiritual songs, with thankfulness in your hearts to God.
COL|3|17|And whatever you do, in word or deed, do everything in the name of the Lord Jesus, giving thanks to God the Father through him.
COL|3|18|Wives, submit to your husbands, as is fitting in the Lord.
COL|3|19|Husbands, love your wives, and do not be harsh with them.
COL|3|20|Children, obey your parents in everything, for this pleases the Lord.
COL|3|21|Fathers, do not provoke your children, lest they become discouraged.
COL|3|22|Slaves, obey in everything those who are your earthly masters, not by way of eye-service, as people-pleasers, but with sincerity of heart, fearing the Lord.
COL|3|23|Whatever you do, work heartily, as for the Lord and not for men,
COL|3|24|knowing that from the Lord you will receive the inheritance as your reward. You are serving the Lord Christ.
COL|3|25|For the wrongdoer will be paid back for the wrong he has done, and there is no partiality.
COL|4|1|Masters, treat your slaves justly and fairly, knowing that you also have a Master in heaven.
COL|4|2|Continue steadfastly in prayer, being watchful in it with thanksgiving.
COL|4|3|At the same time, pray also for us, that God may open to us a door for the word, to declare the mystery of Christ, on account of which I am in prison-
COL|4|4|that I may make it clear, which is how I ought to speak.
COL|4|5|Conduct yourselves wisely toward outsiders, making the best use of the time.
COL|4|6|Let your speech always be gracious, seasoned with salt, so that you may know how you ought to answer each person.
COL|4|7|Tychicus will tell you all about my activities. He is a beloved brother and faithful minister and fellow servant in the Lord.
COL|4|8|I have sent him to you for this very purpose, that you may know how we are and that he may encourage your hearts,
COL|4|9|and with him Onesimus, our faithful and beloved brother, who is one of you. They will tell you of everything that has taken place here.
COL|4|10|Aristarchus my fellow prisoner greets you, and Mark the cousin of Barnabas (concerning whom you have received instructions- if he comes to you, welcome him),
COL|4|11|and Jesus who is called Justus. These are the only men of the circumcision among my fellow workers for the kingdom of God, and they have been a comfort to me.
COL|4|12|Epaphras, who is one of you, a servant of Christ Jesus, greets you, always struggling on your behalf in his prayers, that you may stand mature and fully assured in all the will of God.
COL|4|13|For I bear him witness that he has worked hard for you and for those in Laodicea and in Hierapolis.
COL|4|14|Luke the beloved physician greets you, as does Demas.
COL|4|15|Give my greetings to the brothers at Laodicea, and to Nympha and the church in her house.
COL|4|16|And when this letter has been read among you, have it also read in the church of the Laodiceans; and see that you also read the letter from Laodicea.
COL|4|17|And say to Archippus, "See that you fulfill the ministry that you have received in the Lord."
COL|4|18|I, Paul, write this greeting with my own hand. Remember my chains. Grace be with you.
